module top( mc_cke_pad_o__pad , mc_vpen_pad_o_pad , \mem_ack_r_reg/P0001  , \poc_o[0]_pad  , \poc_o[10]_pad  , \poc_o[11]_pad  , \poc_o[12]_pad  , \poc_o[13]_pad  , \poc_o[14]_pad  , \poc_o[15]_pad  , \poc_o[16]_pad  , \poc_o[17]_pad  , \poc_o[18]_pad  , \poc_o[19]_pad  , \poc_o[1]_pad  , \poc_o[20]_pad  , \poc_o[21]_pad  , \poc_o[22]_pad  , \poc_o[23]_pad  , \poc_o[24]_pad  , \poc_o[25]_pad  , \poc_o[26]_pad  , \poc_o[27]_pad  , \poc_o[28]_pad  , \poc_o[29]_pad  , \poc_o[2]_pad  , \poc_o[30]_pad  , \poc_o[31]_pad  , \poc_o[3]_pad  , \poc_o[4]_pad  , \poc_o[5]_pad  , \poc_o[6]_pad  , \poc_o[7]_pad  , \poc_o[8]_pad  , \poc_o[9]_pad  , suspended_o_pad , \u0_cs_reg[0]/NET0131  , \u0_cs_reg[1]/NET0131  , \u0_csc_mask_r_reg[0]/NET0131  , \u0_csc_mask_r_reg[10]/NET0131  , \u0_csc_mask_r_reg[1]/NET0131  , \u0_csc_mask_r_reg[2]/NET0131  , \u0_csc_mask_r_reg[3]/NET0131  , \u0_csc_mask_r_reg[4]/NET0131  , \u0_csc_mask_r_reg[5]/NET0131  , \u0_csc_mask_r_reg[6]/NET0131  , \u0_csc_mask_r_reg[7]/NET0131  , \u0_csc_mask_r_reg[8]/NET0131  , \u0_csc_mask_r_reg[9]/NET0131  , \u0_csc_reg[10]/NET0131  , \u0_csc_reg[11]/NET0131  , \u0_csc_reg[1]/NET0131  , \u0_csc_reg[2]/NET0131  , \u0_csc_reg[3]/NET0131  , \u0_csc_reg[4]/NET0131  , \u0_csc_reg[5]/NET0131  , \u0_csc_reg[6]/NET0131  , \u0_csc_reg[7]/NET0131  , \u0_csc_reg[9]/NET0131  , \u0_csr_r2_reg[0]/NET0131  , \u0_csr_r2_reg[1]/NET0131  , \u0_csr_r2_reg[2]/NET0131  , \u0_csr_r2_reg[3]/NET0131  , \u0_csr_r2_reg[4]/NET0131  , \u0_csr_r2_reg[5]/NET0131  , \u0_csr_r2_reg[6]/NET0131  , \u0_csr_r2_reg[7]/NET0131  , \u0_csr_r_reg[0]/P0001  , \u0_csr_r_reg[10]/NET0131  , \u0_csr_r_reg[2]/NET0131  , \u0_csr_r_reg[3]/NET0131  , \u0_csr_r_reg[4]/NET0131  , \u0_csr_r_reg[5]/NET0131  , \u0_csr_r_reg[6]/NET0131  , \u0_csr_r_reg[7]/NET0131  , \u0_csr_r_reg[8]/NET0131  , \u0_csr_r_reg[9]/NET0131  , \u0_init_ack_r_reg/P0001  , \u0_init_req_reg/NET0131  , \u0_lmr_ack_r_reg/P0001  , \u0_lmr_req_reg/NET0131  , \u0_rf_we_reg/NET0131  , \u0_rst_r2_reg/NET0131  , \u0_sp_csc_reg[10]/NET0131  , \u0_sp_csc_reg[1]/NET0131  , \u0_sp_csc_reg[2]/NET0131  , \u0_sp_csc_reg[3]/NET0131  , \u0_sp_csc_reg[4]/NET0131  , \u0_sp_csc_reg[5]/NET0131  , \u0_sp_csc_reg[6]/NET0131  , \u0_sp_csc_reg[7]/NET0131  , \u0_sp_csc_reg[9]/NET0131  , \u0_sp_tms_reg[0]/NET0131  , \u0_sp_tms_reg[10]/NET0131  , \u0_sp_tms_reg[11]/NET0131  , \u0_sp_tms_reg[12]/NET0131  , \u0_sp_tms_reg[13]/NET0131  , \u0_sp_tms_reg[14]/NET0131  , \u0_sp_tms_reg[15]/NET0131  , \u0_sp_tms_reg[16]/NET0131  , \u0_sp_tms_reg[17]/NET0131  , \u0_sp_tms_reg[18]/NET0131  , \u0_sp_tms_reg[19]/NET0131  , \u0_sp_tms_reg[1]/NET0131  , \u0_sp_tms_reg[20]/NET0131  , \u0_sp_tms_reg[21]/NET0131  , \u0_sp_tms_reg[22]/NET0131  , \u0_sp_tms_reg[23]/NET0131  , \u0_sp_tms_reg[24]/NET0131  , \u0_sp_tms_reg[25]/NET0131  , \u0_sp_tms_reg[26]/NET0131  , \u0_sp_tms_reg[27]/NET0131  , \u0_sp_tms_reg[2]/NET0131  , \u0_sp_tms_reg[3]/NET0131  , \u0_sp_tms_reg[4]/NET0131  , \u0_sp_tms_reg[5]/NET0131  , \u0_sp_tms_reg[6]/NET0131  , \u0_sp_tms_reg[7]/NET0131  , \u0_sp_tms_reg[8]/NET0131  , \u0_sp_tms_reg[9]/NET0131  , \u0_spec_req_cs_reg[0]/NET0131  , \u0_spec_req_cs_reg[1]/NET0131  , \u0_sreq_cs_le_reg/NET0131  , \u0_tms_reg[0]/NET0131  , \u0_tms_reg[10]/NET0131  , \u0_tms_reg[11]/NET0131  , \u0_tms_reg[12]/NET0131  , \u0_tms_reg[13]/NET0131  , \u0_tms_reg[14]/NET0131  , \u0_tms_reg[15]/NET0131  , \u0_tms_reg[16]/NET0131  , \u0_tms_reg[17]/NET0131  , \u0_tms_reg[18]/NET0131  , \u0_tms_reg[19]/NET0131  , \u0_tms_reg[1]/NET0131  , \u0_tms_reg[20]/NET0131  , \u0_tms_reg[21]/NET0131  , \u0_tms_reg[22]/NET0131  , \u0_tms_reg[23]/NET0131  , \u0_tms_reg[24]/NET0131  , \u0_tms_reg[25]/NET0131  , \u0_tms_reg[26]/NET0131  , \u0_tms_reg[27]/NET0131  , \u0_tms_reg[2]/NET0131  , \u0_tms_reg[3]/NET0131  , \u0_tms_reg[4]/NET0131  , \u0_tms_reg[5]/NET0131  , \u0_tms_reg[6]/NET0131  , \u0_tms_reg[7]/NET0131  , \u0_tms_reg[8]/NET0131  , \u0_tms_reg[9]/NET0131  , \u0_u0_addr_r_reg[2]/P0001  , \u0_u0_addr_r_reg[3]/P0001  , \u0_u0_addr_r_reg[4]/P0001  , \u0_u0_addr_r_reg[5]/P0001  , \u0_u0_addr_r_reg[6]/P0001  , \u0_u0_csc_reg[0]/NET0131  , \u0_u0_csc_reg[10]/P0001  , \u0_u0_csc_reg[11]/P0001  , \u0_u0_csc_reg[12]/P0001  , \u0_u0_csc_reg[13]/P0001  , \u0_u0_csc_reg[14]/P0001  , \u0_u0_csc_reg[15]/P0001  , \u0_u0_csc_reg[16]/P0001  , \u0_u0_csc_reg[17]/P0001  , \u0_u0_csc_reg[18]/P0001  , \u0_u0_csc_reg[19]/P0001  , \u0_u0_csc_reg[1]/NET0131  , \u0_u0_csc_reg[20]/P0001  , \u0_u0_csc_reg[21]/P0001  , \u0_u0_csc_reg[22]/P0001  , \u0_u0_csc_reg[23]/P0001  , \u0_u0_csc_reg[24]/P0001  , \u0_u0_csc_reg[25]/P0001  , \u0_u0_csc_reg[26]/P0001  , \u0_u0_csc_reg[27]/P0001  , \u0_u0_csc_reg[28]/P0001  , \u0_u0_csc_reg[29]/P0001  , \u0_u0_csc_reg[2]/NET0131  , \u0_u0_csc_reg[30]/P0001  , \u0_u0_csc_reg[31]/P0001  , \u0_u0_csc_reg[3]/NET0131  , \u0_u0_csc_reg[4]/P0001  , \u0_u0_csc_reg[5]/P0001  , \u0_u0_csc_reg[6]/P0001  , \u0_u0_csc_reg[7]/P0001  , \u0_u0_csc_reg[8]/P0001  , \u0_u0_csc_reg[9]/P0001  , \u0_u0_init_req_reg/NET0131  , \u0_u0_init_req_we_reg/NET0131  , \u0_u0_inited_reg/NET0131  , \u0_u0_lmr_req_reg/NET0131  , \u0_u0_lmr_req_we_reg/NET0131  , \u0_u0_tms_reg[0]/P0001  , \u0_u0_tms_reg[10]/P0001  , \u0_u0_tms_reg[11]/P0001  , \u0_u0_tms_reg[12]/P0001  , \u0_u0_tms_reg[13]/P0001  , \u0_u0_tms_reg[14]/P0001  , \u0_u0_tms_reg[15]/P0001  , \u0_u0_tms_reg[16]/P0001  , \u0_u0_tms_reg[17]/P0001  , \u0_u0_tms_reg[18]/P0001  , \u0_u0_tms_reg[19]/P0001  , \u0_u0_tms_reg[1]/P0001  , \u0_u0_tms_reg[20]/P0001  , \u0_u0_tms_reg[21]/P0001  , \u0_u0_tms_reg[22]/P0001  , \u0_u0_tms_reg[23]/P0001  , \u0_u0_tms_reg[24]/P0001  , \u0_u0_tms_reg[25]/P0001  , \u0_u0_tms_reg[26]/P0001  , \u0_u0_tms_reg[27]/P0001  , \u0_u0_tms_reg[28]/P0001  , \u0_u0_tms_reg[29]/P0001  , \u0_u0_tms_reg[2]/P0001  , \u0_u0_tms_reg[30]/P0001  , \u0_u0_tms_reg[31]/P0001  , \u0_u0_tms_reg[3]/P0001  , \u0_u0_tms_reg[4]/P0001  , \u0_u0_tms_reg[5]/P0001  , \u0_u0_tms_reg[6]/P0001  , \u0_u0_tms_reg[7]/P0001  , \u0_u0_tms_reg[8]/P0001  , \u0_u0_tms_reg[9]/P0001  , \u0_u1_csc_reg[0]/NET0131  , \u0_u1_csc_reg[10]/P0001  , \u0_u1_csc_reg[11]/P0001  , \u0_u1_csc_reg[12]/P0001  , \u0_u1_csc_reg[13]/P0001  , \u0_u1_csc_reg[14]/P0001  , \u0_u1_csc_reg[15]/P0001  , \u0_u1_csc_reg[16]/P0001  , \u0_u1_csc_reg[17]/P0001  , \u0_u1_csc_reg[18]/P0001  , \u0_u1_csc_reg[19]/P0001  , \u0_u1_csc_reg[1]/NET0131  , \u0_u1_csc_reg[20]/P0001  , \u0_u1_csc_reg[21]/P0001  , \u0_u1_csc_reg[22]/P0001  , \u0_u1_csc_reg[23]/P0001  , \u0_u1_csc_reg[24]/P0001  , \u0_u1_csc_reg[25]/P0001  , \u0_u1_csc_reg[26]/P0001  , \u0_u1_csc_reg[27]/P0001  , \u0_u1_csc_reg[28]/P0001  , \u0_u1_csc_reg[29]/P0001  , \u0_u1_csc_reg[2]/NET0131  , \u0_u1_csc_reg[30]/P0001  , \u0_u1_csc_reg[31]/P0001  , \u0_u1_csc_reg[3]/NET0131  , \u0_u1_csc_reg[4]/P0001  , \u0_u1_csc_reg[5]/P0001  , \u0_u1_csc_reg[6]/P0001  , \u0_u1_csc_reg[7]/P0001  , \u0_u1_csc_reg[8]/P0001  , \u0_u1_csc_reg[9]/P0001  , \u0_u1_init_req_reg/NET0131  , \u0_u1_init_req_we_reg/NET0131  , \u0_u1_inited_reg/NET0131  , \u0_u1_lmr_req_reg/NET0131  , \u0_u1_lmr_req_we_reg/NET0131  , \u0_u1_tms_reg[0]/P0001  , \u0_u1_tms_reg[10]/P0001  , \u0_u1_tms_reg[11]/P0001  , \u0_u1_tms_reg[12]/P0001  , \u0_u1_tms_reg[13]/P0001  , \u0_u1_tms_reg[14]/P0001  , \u0_u1_tms_reg[15]/P0001  , \u0_u1_tms_reg[16]/P0001  , \u0_u1_tms_reg[17]/P0001  , \u0_u1_tms_reg[18]/P0001  , \u0_u1_tms_reg[19]/P0001  , \u0_u1_tms_reg[1]/P0001  , \u0_u1_tms_reg[20]/P0001  , \u0_u1_tms_reg[21]/P0001  , \u0_u1_tms_reg[22]/P0001  , \u0_u1_tms_reg[23]/P0001  , \u0_u1_tms_reg[24]/P0001  , \u0_u1_tms_reg[25]/P0001  , \u0_u1_tms_reg[26]/P0001  , \u0_u1_tms_reg[27]/P0001  , \u0_u1_tms_reg[28]/P0001  , \u0_u1_tms_reg[29]/P0001  , \u0_u1_tms_reg[2]/P0001  , \u0_u1_tms_reg[30]/P0001  , \u0_u1_tms_reg[31]/P0001  , \u0_u1_tms_reg[3]/P0001  , \u0_u1_tms_reg[4]/P0001  , \u0_u1_tms_reg[5]/P0001  , \u0_u1_tms_reg[6]/P0001  , \u0_u1_tms_reg[7]/P0001  , \u0_u1_tms_reg[8]/P0001  , \u0_u1_tms_reg[9]/P0001  , \u0_wp_err_reg/NET0131  , \u1_acs_addr_reg[0]/P0001  , \u1_acs_addr_reg[10]/P0001  , \u1_acs_addr_reg[11]/P0001  , \u1_acs_addr_reg[12]/P0001  , \u1_acs_addr_reg[13]/P0001  , \u1_acs_addr_reg[14]/P0001  , \u1_acs_addr_reg[15]/P0001  , \u1_acs_addr_reg[16]/P0001  , \u1_acs_addr_reg[17]/P0001  , \u1_acs_addr_reg[18]/P0001  , \u1_acs_addr_reg[19]/P0001  , \u1_acs_addr_reg[1]/P0001  , \u1_acs_addr_reg[20]/P0001  , \u1_acs_addr_reg[21]/P0001  , \u1_acs_addr_reg[22]/P0001  , \u1_acs_addr_reg[23]/P0001  , \u1_acs_addr_reg[2]/P0001  , \u1_acs_addr_reg[3]/P0001  , \u1_acs_addr_reg[4]/P0001  , \u1_acs_addr_reg[5]/P0001  , \u1_acs_addr_reg[6]/P0001  , \u1_acs_addr_reg[7]/P0001  , \u1_acs_addr_reg[8]/P0001  , \u1_acs_addr_reg[9]/P0001  , \u1_bank_adr_reg[0]/P0001  , \u1_bank_adr_reg[1]/P0001  , \u1_col_adr_reg[0]/P0001  , \u1_col_adr_reg[1]/P0001  , \u1_col_adr_reg[2]/P0001  , \u1_col_adr_reg[3]/P0001  , \u1_col_adr_reg[4]/P0001  , \u1_col_adr_reg[5]/P0001  , \u1_col_adr_reg[6]/P0001  , \u1_col_adr_reg[7]/P0001  , \u1_col_adr_reg[8]/P0001  , \u1_col_adr_reg[9]/P0001  , \u1_row_adr_reg[0]/P0001  , \u1_row_adr_reg[10]/P0001  , \u1_row_adr_reg[11]/P0001  , \u1_row_adr_reg[12]/P0001  , \u1_row_adr_reg[1]/P0001  , \u1_row_adr_reg[2]/P0001  , \u1_row_adr_reg[3]/P0001  , \u1_row_adr_reg[4]/P0001  , \u1_row_adr_reg[5]/P0001  , \u1_row_adr_reg[6]/P0001  , \u1_row_adr_reg[7]/P0001  , \u1_row_adr_reg[8]/P0001  , \u1_row_adr_reg[9]/P0001  , \u1_sram_addr_reg[0]/P0001  , \u1_sram_addr_reg[10]/P0001  , \u1_sram_addr_reg[11]/P0001  , \u1_sram_addr_reg[12]/P0001  , \u1_sram_addr_reg[13]/P0001  , \u1_sram_addr_reg[14]/P0001  , \u1_sram_addr_reg[15]/P0001  , \u1_sram_addr_reg[16]/P0001  , \u1_sram_addr_reg[17]/P0001  , \u1_sram_addr_reg[18]/P0001  , \u1_sram_addr_reg[19]/P0001  , \u1_sram_addr_reg[1]/P0001  , \u1_sram_addr_reg[20]/P0001  , \u1_sram_addr_reg[21]/P0001  , \u1_sram_addr_reg[22]/P0001  , \u1_sram_addr_reg[23]/P0001  , \u1_sram_addr_reg[2]/P0001  , \u1_sram_addr_reg[3]/P0001  , \u1_sram_addr_reg[4]/P0001  , \u1_sram_addr_reg[5]/P0001  , \u1_sram_addr_reg[6]/P0001  , \u1_sram_addr_reg[7]/P0001  , \u1_sram_addr_reg[8]/P0001  , \u1_sram_addr_reg[9]/P0001  , \u1_u0_out_r_reg[0]/P0001  , \u1_u0_out_r_reg[10]/P0001  , \u1_u0_out_r_reg[11]/P0001  , \u1_u0_out_r_reg[12]/P0001  , \u1_u0_out_r_reg[1]/P0001  , \u1_u0_out_r_reg[2]/P0001  , \u1_u0_out_r_reg[3]/P0001  , \u1_u0_out_r_reg[4]/P0001  , \u1_u0_out_r_reg[5]/P0001  , \u1_u0_out_r_reg[6]/P0001  , \u1_u0_out_r_reg[7]/P0001  , \u1_u0_out_r_reg[8]/P0001  , \u1_u0_out_r_reg[9]/P0001  , \u2_bank_open_reg/P0001  , \u2_row_same_reg/P0001  , \u2_u0_b0_last_row_reg[0]/P0001  , \u2_u0_b0_last_row_reg[10]/P0001  , \u2_u0_b0_last_row_reg[11]/P0001  , \u2_u0_b0_last_row_reg[12]/P0001  , \u2_u0_b0_last_row_reg[1]/P0001  , \u2_u0_b0_last_row_reg[2]/P0001  , \u2_u0_b0_last_row_reg[3]/P0001  , \u2_u0_b0_last_row_reg[4]/P0001  , \u2_u0_b0_last_row_reg[5]/P0001  , \u2_u0_b0_last_row_reg[6]/P0001  , \u2_u0_b0_last_row_reg[7]/P0001  , \u2_u0_b0_last_row_reg[8]/P0001  , \u2_u0_b0_last_row_reg[9]/P0001  , \u2_u0_b1_last_row_reg[0]/P0001  , \u2_u0_b1_last_row_reg[10]/P0001  , \u2_u0_b1_last_row_reg[11]/P0001  , \u2_u0_b1_last_row_reg[12]/P0001  , \u2_u0_b1_last_row_reg[1]/P0001  , \u2_u0_b1_last_row_reg[2]/P0001  , \u2_u0_b1_last_row_reg[3]/P0001  , \u2_u0_b1_last_row_reg[4]/P0001  , \u2_u0_b1_last_row_reg[5]/P0001  , \u2_u0_b1_last_row_reg[6]/P0001  , \u2_u0_b1_last_row_reg[7]/P0001  , \u2_u0_b1_last_row_reg[8]/P0001  , \u2_u0_b1_last_row_reg[9]/P0001  , \u2_u0_b2_last_row_reg[0]/P0001  , \u2_u0_b2_last_row_reg[10]/P0001  , \u2_u0_b2_last_row_reg[11]/P0001  , \u2_u0_b2_last_row_reg[12]/P0001  , \u2_u0_b2_last_row_reg[1]/P0001  , \u2_u0_b2_last_row_reg[2]/P0001  , \u2_u0_b2_last_row_reg[3]/P0001  , \u2_u0_b2_last_row_reg[4]/P0001  , \u2_u0_b2_last_row_reg[5]/P0001  , \u2_u0_b2_last_row_reg[6]/P0001  , \u2_u0_b2_last_row_reg[7]/P0001  , \u2_u0_b2_last_row_reg[8]/P0001  , \u2_u0_b2_last_row_reg[9]/P0001  , \u2_u0_b3_last_row_reg[0]/P0001  , \u2_u0_b3_last_row_reg[10]/P0001  , \u2_u0_b3_last_row_reg[11]/P0001  , \u2_u0_b3_last_row_reg[12]/P0001  , \u2_u0_b3_last_row_reg[1]/P0001  , \u2_u0_b3_last_row_reg[2]/P0001  , \u2_u0_b3_last_row_reg[3]/P0001  , \u2_u0_b3_last_row_reg[4]/P0001  , \u2_u0_b3_last_row_reg[5]/P0001  , \u2_u0_b3_last_row_reg[6]/P0001  , \u2_u0_b3_last_row_reg[7]/P0001  , \u2_u0_b3_last_row_reg[8]/P0001  , \u2_u0_b3_last_row_reg[9]/P0001  , \u2_u0_bank0_open_reg/NET0131  , \u2_u0_bank1_open_reg/NET0131  , \u2_u0_bank2_open_reg/NET0131  , \u2_u0_bank3_open_reg/NET0131  , \u2_u1_b0_last_row_reg[0]/P0001  , \u2_u1_b0_last_row_reg[10]/P0001  , \u2_u1_b0_last_row_reg[11]/P0001  , \u2_u1_b0_last_row_reg[12]/P0001  , \u2_u1_b0_last_row_reg[1]/P0001  , \u2_u1_b0_last_row_reg[2]/P0001  , \u2_u1_b0_last_row_reg[3]/P0001  , \u2_u1_b0_last_row_reg[4]/P0001  , \u2_u1_b0_last_row_reg[5]/P0001  , \u2_u1_b0_last_row_reg[6]/P0001  , \u2_u1_b0_last_row_reg[7]/P0001  , \u2_u1_b0_last_row_reg[8]/P0001  , \u2_u1_b0_last_row_reg[9]/P0001  , \u2_u1_b1_last_row_reg[0]/P0001  , \u2_u1_b1_last_row_reg[10]/P0001  , \u2_u1_b1_last_row_reg[11]/P0001  , \u2_u1_b1_last_row_reg[12]/P0001  , \u2_u1_b1_last_row_reg[1]/P0001  , \u2_u1_b1_last_row_reg[2]/P0001  , \u2_u1_b1_last_row_reg[3]/P0001  , \u2_u1_b1_last_row_reg[4]/P0001  , \u2_u1_b1_last_row_reg[5]/P0001  , \u2_u1_b1_last_row_reg[6]/P0001  , \u2_u1_b1_last_row_reg[7]/P0001  , \u2_u1_b1_last_row_reg[8]/P0001  , \u2_u1_b1_last_row_reg[9]/P0001  , \u2_u1_b2_last_row_reg[0]/P0001  , \u2_u1_b2_last_row_reg[10]/P0001  , \u2_u1_b2_last_row_reg[11]/P0001  , \u2_u1_b2_last_row_reg[12]/P0001  , \u2_u1_b2_last_row_reg[1]/P0001  , \u2_u1_b2_last_row_reg[2]/P0001  , \u2_u1_b2_last_row_reg[3]/P0001  , \u2_u1_b2_last_row_reg[4]/P0001  , \u2_u1_b2_last_row_reg[5]/P0001  , \u2_u1_b2_last_row_reg[6]/P0001  , \u2_u1_b2_last_row_reg[7]/P0001  , \u2_u1_b2_last_row_reg[8]/P0001  , \u2_u1_b2_last_row_reg[9]/P0001  , \u2_u1_b3_last_row_reg[0]/P0001  , \u2_u1_b3_last_row_reg[10]/P0001  , \u2_u1_b3_last_row_reg[11]/P0001  , \u2_u1_b3_last_row_reg[12]/P0001  , \u2_u1_b3_last_row_reg[1]/P0001  , \u2_u1_b3_last_row_reg[2]/P0001  , \u2_u1_b3_last_row_reg[3]/P0001  , \u2_u1_b3_last_row_reg[4]/P0001  , \u2_u1_b3_last_row_reg[5]/P0001  , \u2_u1_b3_last_row_reg[6]/P0001  , \u2_u1_b3_last_row_reg[7]/P0001  , \u2_u1_b3_last_row_reg[8]/P0001  , \u2_u1_b3_last_row_reg[9]/P0001  , \u2_u1_bank0_open_reg/NET0131  , \u2_u1_bank1_open_reg/NET0131  , \u2_u1_bank2_open_reg/NET0131  , \u2_u1_bank3_open_reg/NET0131  , \u3_byte0_reg[0]/P0001  , \u3_byte0_reg[1]/P0001  , \u3_byte0_reg[2]/P0001  , \u3_byte0_reg[3]/P0001  , \u3_byte0_reg[4]/P0001  , \u3_byte0_reg[5]/P0001  , \u3_byte0_reg[6]/P0001  , \u3_byte0_reg[7]/P0001  , \u3_byte1_reg[0]/P0001  , \u3_byte1_reg[1]/P0001  , \u3_byte1_reg[2]/P0001  , \u3_byte1_reg[3]/P0001  , \u3_byte1_reg[4]/P0001  , \u3_byte1_reg[5]/P0001  , \u3_byte1_reg[6]/P0001  , \u3_byte1_reg[7]/P0001  , \u3_byte2_reg[0]/P0001  , \u3_byte2_reg[1]/P0001  , \u3_byte2_reg[2]/P0001  , \u3_byte2_reg[3]/P0001  , \u3_byte2_reg[4]/P0001  , \u3_byte2_reg[5]/P0001  , \u3_byte2_reg[6]/P0001  , \u3_byte2_reg[7]/P0001  , \u3_u0_r0_reg[0]/P0001  , \u3_u0_r0_reg[10]/P0001  , \u3_u0_r0_reg[11]/P0001  , \u3_u0_r0_reg[12]/P0001  , \u3_u0_r0_reg[13]/P0001  , \u3_u0_r0_reg[14]/P0001  , \u3_u0_r0_reg[15]/P0001  , \u3_u0_r0_reg[16]/P0001  , \u3_u0_r0_reg[17]/P0001  , \u3_u0_r0_reg[18]/P0001  , \u3_u0_r0_reg[19]/P0001  , \u3_u0_r0_reg[1]/P0001  , \u3_u0_r0_reg[20]/P0001  , \u3_u0_r0_reg[21]/P0001  , \u3_u0_r0_reg[22]/P0001  , \u3_u0_r0_reg[23]/P0001  , \u3_u0_r0_reg[24]/P0001  , \u3_u0_r0_reg[25]/P0001  , \u3_u0_r0_reg[26]/P0001  , \u3_u0_r0_reg[27]/P0001  , \u3_u0_r0_reg[28]/P0001  , \u3_u0_r0_reg[29]/P0001  , \u3_u0_r0_reg[2]/P0001  , \u3_u0_r0_reg[30]/P0001  , \u3_u0_r0_reg[31]/P0001  , \u3_u0_r0_reg[32]/P0001  , \u3_u0_r0_reg[33]/P0001  , \u3_u0_r0_reg[34]/P0001  , \u3_u0_r0_reg[35]/P0001  , \u3_u0_r0_reg[3]/P0001  , \u3_u0_r0_reg[4]/P0001  , \u3_u0_r0_reg[5]/P0001  , \u3_u0_r0_reg[6]/P0001  , \u3_u0_r0_reg[7]/P0001  , \u3_u0_r0_reg[8]/P0001  , \u3_u0_r0_reg[9]/P0001  , \u3_u0_r1_reg[0]/P0001  , \u3_u0_r1_reg[10]/P0001  , \u3_u0_r1_reg[11]/P0001  , \u3_u0_r1_reg[12]/P0001  , \u3_u0_r1_reg[13]/P0001  , \u3_u0_r1_reg[14]/P0001  , \u3_u0_r1_reg[15]/P0001  , \u3_u0_r1_reg[16]/P0001  , \u3_u0_r1_reg[17]/P0001  , \u3_u0_r1_reg[18]/P0001  , \u3_u0_r1_reg[19]/P0001  , \u3_u0_r1_reg[1]/P0001  , \u3_u0_r1_reg[20]/P0001  , \u3_u0_r1_reg[21]/P0001  , \u3_u0_r1_reg[22]/P0001  , \u3_u0_r1_reg[23]/P0001  , \u3_u0_r1_reg[24]/P0001  , \u3_u0_r1_reg[25]/P0001  , \u3_u0_r1_reg[26]/P0001  , \u3_u0_r1_reg[27]/P0001  , \u3_u0_r1_reg[28]/P0001  , \u3_u0_r1_reg[29]/P0001  , \u3_u0_r1_reg[2]/P0001  , \u3_u0_r1_reg[30]/P0001  , \u3_u0_r1_reg[31]/P0001  , \u3_u0_r1_reg[32]/P0001  , \u3_u0_r1_reg[33]/P0001  , \u3_u0_r1_reg[34]/P0001  , \u3_u0_r1_reg[35]/P0001  , \u3_u0_r1_reg[3]/P0001  , \u3_u0_r1_reg[4]/P0001  , \u3_u0_r1_reg[5]/P0001  , \u3_u0_r1_reg[6]/P0001  , \u3_u0_r1_reg[7]/P0001  , \u3_u0_r1_reg[8]/P0001  , \u3_u0_r1_reg[9]/P0001  , \u3_u0_r2_reg[0]/P0001  , \u3_u0_r2_reg[10]/P0001  , \u3_u0_r2_reg[11]/P0001  , \u3_u0_r2_reg[12]/P0001  , \u3_u0_r2_reg[13]/P0001  , \u3_u0_r2_reg[14]/P0001  , \u3_u0_r2_reg[15]/P0001  , \u3_u0_r2_reg[16]/P0001  , \u3_u0_r2_reg[17]/P0001  , \u3_u0_r2_reg[18]/P0001  , \u3_u0_r2_reg[19]/P0001  , \u3_u0_r2_reg[1]/P0001  , \u3_u0_r2_reg[20]/P0001  , \u3_u0_r2_reg[21]/P0001  , \u3_u0_r2_reg[22]/P0001  , \u3_u0_r2_reg[23]/P0001  , \u3_u0_r2_reg[24]/P0001  , \u3_u0_r2_reg[25]/P0001  , \u3_u0_r2_reg[26]/P0001  , \u3_u0_r2_reg[27]/P0001  , \u3_u0_r2_reg[28]/P0001  , \u3_u0_r2_reg[29]/P0001  , \u3_u0_r2_reg[2]/P0001  , \u3_u0_r2_reg[30]/P0001  , \u3_u0_r2_reg[31]/P0001  , \u3_u0_r2_reg[32]/P0001  , \u3_u0_r2_reg[33]/P0001  , \u3_u0_r2_reg[34]/P0001  , \u3_u0_r2_reg[35]/P0001  , \u3_u0_r2_reg[3]/P0001  , \u3_u0_r2_reg[4]/P0001  , \u3_u0_r2_reg[5]/P0001  , \u3_u0_r2_reg[6]/P0001  , \u3_u0_r2_reg[7]/P0001  , \u3_u0_r2_reg[8]/P0001  , \u3_u0_r2_reg[9]/P0001  , \u3_u0_r3_reg[0]/P0001  , \u3_u0_r3_reg[10]/P0001  , \u3_u0_r3_reg[11]/P0001  , \u3_u0_r3_reg[12]/P0001  , \u3_u0_r3_reg[13]/P0001  , \u3_u0_r3_reg[14]/P0001  , \u3_u0_r3_reg[15]/P0001  , \u3_u0_r3_reg[16]/P0001  , \u3_u0_r3_reg[17]/P0001  , \u3_u0_r3_reg[18]/P0001  , \u3_u0_r3_reg[19]/P0001  , \u3_u0_r3_reg[1]/P0001  , \u3_u0_r3_reg[20]/P0001  , \u3_u0_r3_reg[21]/P0001  , \u3_u0_r3_reg[22]/P0001  , \u3_u0_r3_reg[23]/P0001  , \u3_u0_r3_reg[24]/P0001  , \u3_u0_r3_reg[25]/P0001  , \u3_u0_r3_reg[26]/P0001  , \u3_u0_r3_reg[27]/P0001  , \u3_u0_r3_reg[28]/P0001  , \u3_u0_r3_reg[29]/P0001  , \u3_u0_r3_reg[2]/P0001  , \u3_u0_r3_reg[30]/P0001  , \u3_u0_r3_reg[31]/P0001  , \u3_u0_r3_reg[32]/P0001  , \u3_u0_r3_reg[33]/P0001  , \u3_u0_r3_reg[34]/P0001  , \u3_u0_r3_reg[35]/P0001  , \u3_u0_r3_reg[3]/P0001  , \u3_u0_r3_reg[4]/P0001  , \u3_u0_r3_reg[5]/P0001  , \u3_u0_r3_reg[6]/P0001  , \u3_u0_r3_reg[7]/P0001  , \u3_u0_r3_reg[8]/P0001  , \u3_u0_r3_reg[9]/P0001  , \u3_u0_rd_adr_reg[0]/NET0131  , \u3_u0_rd_adr_reg[1]/NET0131  , \u3_u0_rd_adr_reg[2]/NET0131  , \u3_u0_rd_adr_reg[3]/NET0131  , \u3_u0_wr_adr_reg[0]/NET0131  , \u3_u0_wr_adr_reg[1]/NET0131  , \u3_u0_wr_adr_reg[2]/NET0131  , \u3_u0_wr_adr_reg[3]/NET0131  , \u4_ps_cnt_reg[0]/NET0131  , \u4_ps_cnt_reg[1]/NET0131  , \u4_ps_cnt_reg[2]/NET0131  , \u4_ps_cnt_reg[3]/NET0131  , \u4_ps_cnt_reg[4]/NET0131  , \u4_ps_cnt_reg[5]/NET0131  , \u4_ps_cnt_reg[6]/NET0131  , \u4_ps_cnt_reg[7]/NET0131  , \u4_rfr_ce_reg/NET0131  , \u4_rfr_clr_reg/P0001  , \u4_rfr_cnt_reg[0]/NET0131  , \u4_rfr_cnt_reg[1]/NET0131  , \u4_rfr_cnt_reg[2]/NET0131  , \u4_rfr_cnt_reg[3]/NET0131  , \u4_rfr_cnt_reg[4]/NET0131  , \u4_rfr_cnt_reg[5]/NET0131  , \u4_rfr_cnt_reg[6]/NET0131  , \u4_rfr_cnt_reg[7]/NET0131  , \u4_rfr_early_reg/NET0131  , \u4_rfr_en_reg/NET0131  , \u4_rfr_req_reg/NET0131  , \u5_ack_cnt_reg[0]/NET0131  , \u5_ack_cnt_reg[1]/NET0131  , \u5_ack_cnt_reg[2]/NET0131  , \u5_ack_cnt_reg[3]/NET0131  , \u5_ap_en_reg/NET0131  , \u5_burst_act_rd_reg/P0001  , \u5_burst_cnt_reg[0]/NET0131  , \u5_burst_cnt_reg[10]/NET0131  , \u5_burst_cnt_reg[1]/NET0131  , \u5_burst_cnt_reg[2]/NET0131  , \u5_burst_cnt_reg[3]/NET0131  , \u5_burst_cnt_reg[4]/NET0131  , \u5_burst_cnt_reg[5]/NET0131  , \u5_burst_cnt_reg[6]/NET0131  , \u5_burst_cnt_reg[7]/NET0131  , \u5_burst_cnt_reg[8]/NET0131  , \u5_burst_cnt_reg[9]/NET0131  , \u5_cke_o_del_reg/P0001  , \u5_cke_r_reg/NET0131  , \u5_cmd_a10_r_reg/P0001  , \u5_cmd_asserted2_reg/NET0131  , \u5_cmd_asserted_reg/NET0131  , \u5_cmd_del_reg[0]/NET0131  , \u5_cmd_del_reg[1]/NET0131  , \u5_cmd_del_reg[2]/NET0131  , \u5_cmd_del_reg[3]/NET0131  , \u5_cnt_reg/NET0131  , \u5_cs_le_r_reg/P0001  , \u5_cs_le_reg/P0001  , \u5_data_oe_r2_reg/NET0131  , \u5_data_oe_reg/NET0131  , \u5_dv_r_reg/NET0131  , \u5_ir_cnt_done_reg/P0001  , \u5_ir_cnt_reg[0]/P0001  , \u5_ir_cnt_reg[1]/P0001  , \u5_ir_cnt_reg[2]/P0001  , \u5_ir_cnt_reg[3]/P0001  , \u5_lmr_ack_reg/NET0131  , \u5_lookup_ready1_reg/NET0131  , \u5_lookup_ready2_reg/NET0131  , \u5_mc_adv_r1_reg/NET0131  , \u5_mc_adv_r_reg/NET0131  , \u5_mc_c_oe_reg/NET0131  , \u5_mc_le_reg/NET0131  , \u5_mem_ack_r_reg/NET0131  , \u5_no_wb_cycle_reg/NET0131  , \u5_oe__reg/NET0131  , \u5_pack_le0_reg/P0001  , \u5_pack_le1_reg/P0001  , \u5_resume_req_r_reg/NET0131  , \u5_rfr_ack_r_reg/NET0131  , \u5_state_reg[0]/NET0131  , \u5_state_reg[10]/NET0131  , \u5_state_reg[11]/NET0131  , \u5_state_reg[12]/NET0131  , \u5_state_reg[13]/NET0131  , \u5_state_reg[14]/NET0131  , \u5_state_reg[15]/NET0131  , \u5_state_reg[16]/NET0131  , \u5_state_reg[17]/NET0131  , \u5_state_reg[18]/NET0131  , \u5_state_reg[19]/NET0131  , \u5_state_reg[1]/NET0131  , \u5_state_reg[20]/NET0131  , \u5_state_reg[21]/NET0131  , \u5_state_reg[22]/NET0131  , \u5_state_reg[23]/NET0131  , \u5_state_reg[24]/NET0131  , \u5_state_reg[25]/NET0131  , \u5_state_reg[26]/NET0131  , \u5_state_reg[27]/NET0131  , \u5_state_reg[28]/NET0131  , \u5_state_reg[29]/NET0131  , \u5_state_reg[2]/NET0131  , \u5_state_reg[30]/NET0131  , \u5_state_reg[31]/NET0131  , \u5_state_reg[32]/NET0131  , \u5_state_reg[33]/NET0131  , \u5_state_reg[34]/NET0131  , \u5_state_reg[35]/NET0131  , \u5_state_reg[36]/NET0131  , \u5_state_reg[37]/NET0131  , \u5_state_reg[38]/NET0131  , \u5_state_reg[39]/NET0131  , \u5_state_reg[3]/NET0131  , \u5_state_reg[40]/NET0131  , \u5_state_reg[41]/NET0131  , \u5_state_reg[42]/NET0131  , \u5_state_reg[43]/NET0131  , \u5_state_reg[44]/NET0131  , \u5_state_reg[45]/NET0131  , \u5_state_reg[46]/NET0131  , \u5_state_reg[47]/NET0131  , \u5_state_reg[48]/NET0131  , \u5_state_reg[49]/NET0131  , \u5_state_reg[4]/NET0131  , \u5_state_reg[50]/NET0131  , \u5_state_reg[51]/NET0131  , \u5_state_reg[52]/NET0131  , \u5_state_reg[53]/NET0131  , \u5_state_reg[54]/NET0131  , \u5_state_reg[55]/NET0131  , \u5_state_reg[56]/NET0131  , \u5_state_reg[57]/NET0131  , \u5_state_reg[58]/NET0131  , \u5_state_reg[59]/NET0131  , \u5_state_reg[5]/NET0131  , \u5_state_reg[60]/NET0131  , \u5_state_reg[61]/NET0131  , \u5_state_reg[62]/NET0131  , \u5_state_reg[63]/NET0131  , \u5_state_reg[64]/NET0131  , \u5_state_reg[65]/NET0131  , \u5_state_reg[6]/NET0131  , \u5_state_reg[7]/NET0131  , \u5_state_reg[8]/NET0131  , \u5_state_reg[9]/NET0131  , \u5_susp_req_r_reg/NET0131  , \u5_susp_sel_r_reg/NET0131  , \u5_timer2_reg[0]/P0001  , \u5_timer2_reg[1]/P0001  , \u5_timer2_reg[2]/P0001  , \u5_timer2_reg[3]/P0001  , \u5_timer2_reg[4]/P0001  , \u5_timer2_reg[5]/P0001  , \u5_timer2_reg[6]/P0001  , \u5_timer2_reg[7]/P0001  , \u5_timer2_reg[8]/P0001  , \u5_timer_reg[0]/NET0131  , \u5_timer_reg[1]/NET0131  , \u5_timer_reg[2]/NET0131  , \u5_timer_reg[3]/NET0131  , \u5_timer_reg[4]/NET0131  , \u5_timer_reg[5]/NET0131  , \u5_timer_reg[6]/NET0131  , \u5_timer_reg[7]/NET0131  , \u5_tmr2_done_reg/NET0131  , \u5_tmr_done_reg/NET0131  , \u5_wb_cycle_reg/NET0131  , \u5_wb_stb_first_reg/NET0131  , \u5_wb_wait_r_reg/P0001  , \u5_wb_write_go_r_reg/NET0131  , \u5_wr_cycle_reg/NET0131  , \u6_read_go_r1_reg/NET0131  , \u6_read_go_r_reg/NET0131  , \u6_rmw_en_reg/NET0131  , \u6_rmw_r_reg/NET0131  , \u6_wb_first_r_reg/NET0131  , \u6_wr_hold_reg/NET0131  , \u6_write_go_r1_reg/NET0131  , \u6_write_go_r_reg/NET0131  , \u7_mc_ack_r_reg/NET0131  , \u7_mc_br_r_reg/P0001  , \u7_mc_data_ir_reg[0]/P0001  , \u7_mc_data_ir_reg[10]/P0001  , \u7_mc_data_ir_reg[11]/P0001  , \u7_mc_data_ir_reg[12]/P0001  , \u7_mc_data_ir_reg[13]/P0001  , \u7_mc_data_ir_reg[14]/P0001  , \u7_mc_data_ir_reg[15]/P0001  , \u7_mc_data_ir_reg[16]/P0001  , \u7_mc_data_ir_reg[17]/P0001  , \u7_mc_data_ir_reg[18]/P0001  , \u7_mc_data_ir_reg[19]/P0001  , \u7_mc_data_ir_reg[1]/P0001  , \u7_mc_data_ir_reg[20]/P0001  , \u7_mc_data_ir_reg[21]/P0001  , \u7_mc_data_ir_reg[22]/P0001  , \u7_mc_data_ir_reg[23]/P0001  , \u7_mc_data_ir_reg[24]/P0001  , \u7_mc_data_ir_reg[25]/P0001  , \u7_mc_data_ir_reg[26]/P0001  , \u7_mc_data_ir_reg[27]/P0001  , \u7_mc_data_ir_reg[28]/P0001  , \u7_mc_data_ir_reg[29]/P0001  , \u7_mc_data_ir_reg[2]/P0001  , \u7_mc_data_ir_reg[30]/P0001  , \u7_mc_data_ir_reg[31]/P0001  , \u7_mc_data_ir_reg[3]/P0001  , \u7_mc_data_ir_reg[4]/P0001  , \u7_mc_data_ir_reg[5]/P0001  , \u7_mc_data_ir_reg[6]/P0001  , \u7_mc_data_ir_reg[7]/P0001  , \u7_mc_data_ir_reg[8]/P0001  , \u7_mc_data_ir_reg[9]/P0001  , \u7_mc_dqm_r2_reg[0]/P0001  , \u7_mc_dqm_r2_reg[1]/P0001  , \u7_mc_dqm_r2_reg[2]/P0001  , \u7_mc_dqm_r2_reg[3]/P0001  , \u7_mc_dqm_r_reg[0]/P0001  , \u7_mc_dqm_r_reg[1]/P0001  , \u7_mc_dqm_r_reg[2]/P0001  , \u7_mc_dqm_r_reg[3]/P0001  , wb_ack_o_pad , \wb_addr_i[0]_pad  , \wb_addr_i[10]_pad  , \wb_addr_i[11]_pad  , \wb_addr_i[12]_pad  , \wb_addr_i[13]_pad  , \wb_addr_i[14]_pad  , \wb_addr_i[15]_pad  , \wb_addr_i[16]_pad  , \wb_addr_i[17]_pad  , \wb_addr_i[18]_pad  , \wb_addr_i[19]_pad  , \wb_addr_i[1]_pad  , \wb_addr_i[20]_pad  , \wb_addr_i[21]_pad  , \wb_addr_i[22]_pad  , \wb_addr_i[23]_pad  , \wb_addr_i[24]_pad  , \wb_addr_i[25]_pad  , \wb_addr_i[26]_pad  , \wb_addr_i[27]_pad  , \wb_addr_i[28]_pad  , \wb_addr_i[29]_pad  , \wb_addr_i[2]_pad  , \wb_addr_i[30]_pad  , \wb_addr_i[31]_pad  , \wb_addr_i[3]_pad  , \wb_addr_i[4]_pad  , \wb_addr_i[5]_pad  , \wb_addr_i[6]_pad  , \wb_addr_i[7]_pad  , \wb_addr_i[8]_pad  , \wb_addr_i[9]_pad  , wb_cyc_i_pad , \wb_data_i[0]_pad  , \wb_data_i[10]_pad  , \wb_data_i[11]_pad  , \wb_data_i[12]_pad  , \wb_data_i[13]_pad  , \wb_data_i[14]_pad  , \wb_data_i[15]_pad  , \wb_data_i[16]_pad  , \wb_data_i[17]_pad  , \wb_data_i[18]_pad  , \wb_data_i[19]_pad  , \wb_data_i[1]_pad  , \wb_data_i[20]_pad  , \wb_data_i[21]_pad  , \wb_data_i[22]_pad  , \wb_data_i[23]_pad  , \wb_data_i[24]_pad  , \wb_data_i[25]_pad  , \wb_data_i[26]_pad  , \wb_data_i[27]_pad  , \wb_data_i[28]_pad  , \wb_data_i[29]_pad  , \wb_data_i[2]_pad  , \wb_data_i[30]_pad  , \wb_data_i[31]_pad  , \wb_data_i[3]_pad  , \wb_data_i[4]_pad  , \wb_data_i[5]_pad  , \wb_data_i[6]_pad  , \wb_data_i[7]_pad  , \wb_data_i[8]_pad  , \wb_data_i[9]_pad  , wb_err_o_pad , \wb_sel_i[0]_pad  , \wb_sel_i[1]_pad  , \wb_sel_i[2]_pad  , \wb_sel_i[3]_pad  , wb_stb_i_pad , wb_we_i_pad , \_al_n0  , \_al_n1  , \g22/_0_  , \g23/_0_  , \g25_dup61718/_2_  , \g43466/_0_  , \g43467/_0_  , \g43468/_0_  , \g43469/_0_  , \g43470/_0_  , \g43471/_0_  , \g43472/_0_  , \g43473/_0_  , \g43474/_0_  , \g43475/_0_  , \g43476/_0_  , \g43477/_0_  , \g43478/_0_  , \g43512/_0_  , \g43513/_0_  , \g43544/_3_  , \g43545/_0_  , \g43554/_0_  , \g43555/_0_  , \g43557/_0_  , \g43558/_0_  , \g43571/_2_  , \g43632/_0_  , \g43633/_0_  , \g43635/_0_  , \g43636/_0_  , \g43637/_0_  , \g43638/_0_  , \g43639/_0_  , \g43640/_0_  , \g43642/_0_  , \g43662/_0_  , \g43663/_0_  , \g43664/_0_  , \g43665/_0_  , \g43668/_0_  , \g43670/_0_  , \g43671/_0_  , \g43673/_0_  , \g43674/_0_  , \g43692/_0_  , \g43695/_0_  , \g43696/_0_  , \g43697/_0_  , \g43698/_0_  , \g43700/_0_  , \g43701/_0_  , \g43703/_0_  , \g43705/_0_  , \g43707/_0_  , \g43708/_0_  , \g43710/_0_  , \g43717/_0_  , \g43719/_0_  , \g43720/_0_  , \g43721/_0_  , \g43722/_1_  , \g43723/_0_  , \g43725/_0_  , \g43729/_0_  , \g43731/_0_  , \g43734/_0_  , \g43735/_0_  , \g43737/_0_  , \g43744/_0_  , \g43747/_0_  , \g43760/_2_  , \g43770/_1_  , \g43775/_2_  , \g43780/_2_  , \g43786/_0_  , \g43787/_1_  , \g43847/_0_  , \g43848/_1_  , \g43858/_1_  , \g43891/_3_  , \g43895/_0_  , \g43934/_0_  , \g43936/_3_  , \g43954/_3_  , \g43961/_0_  , \g44016/_1_  , \g44067/_0_  , \g44094/_0_  , \g44096/_0_  , \g44104/_0_  , \g44122/_0_  , \g44172/_0_  , \g44209/_0_  , \g44219/_0_  , \g44220/_0_  , \g44222/_0_  , \g44223/_0_  , \g44241/_2_  , \g44252/_0_  , \g44253/_0_  , \g44255/_2_  , \g44263/_2_  , \g44470/_0_  , \g44538/_0_  , \g44539/_0_  , \g44540/_0_  , \g44541/_0_  , \g44542/_0_  , \g44543/_0_  , \g44544/_0_  , \g44545/_0_  , \g44546/_0_  , \g44547/_0_  , \g44548/_0_  , \g44549/_0_  , \g44550/_0_  , \g44551/_0_  , \g44552/_0_  , \g44553/_0_  , \g44554/_0_  , \g44555/_0_  , \g44556/_0_  , \g44557/_0_  , \g44558/_0_  , \g44559/_0_  , \g44560/_0_  , \g44561/_0_  , \g44562/_0_  , \g44563/_0_  , \g44564/_0_  , \g44565/_0_  , \g44566/_0_  , \g44567/_0_  , \g44568/_0_  , \g44569/_0_  , \g44570/_0_  , \g44571/_0_  , \g44572/_0_  , \g44573/_0_  , \g44574/_0_  , \g44575/_0_  , \g44576/_0_  , \g44577/_0_  , \g44578/_0_  , \g44579/_0_  , \g44580/_0_  , \g44581/_0_  , \g44582/_0_  , \g44583/_0_  , \g44584/_0_  , \g44585/_0_  , \g44586/_0_  , \g44588/_0_  , \g44589/_0_  , \g44590/_0_  , \g44591/_0_  , \g44592/_0_  , \g44593/_0_  , \g44594/_0_  , \g44595/_0_  , \g44596/_0_  , \g44636/_2_  , \g44646/_0_  , \g44647/_0_  , \g44648/_0_  , \g44649/_0_  , \g44650/_0_  , \g44651/_0_  , \g44652/_0_  , \g44653/_0_  , \g44654/_0_  , \g44655/_0_  , \g44656/_0_  , \g44657/_0_  , \g44665/_0_  , \g44666/_0_  , \g44667/_0_  , \g44668/_0_  , \g44752/_0_  , \g44753/_0_  , \g44873/_0_  , \g44939/_0_  , \g44942/_0_  , \g44945/_0_  , \g45023/_2_  , \g45090/_0_  , \g45141/_0_  , \g45147/_3_  , \g45155/_0_  , \g45190/_0_  , \g45195/_2_  , \g45199/_2_  , \g45201/_2_  , \g45324/_0_  , \g45334/_2_  , \g45336/_0_  , \g45388/_0_  , \g45391/_0_  , \g45413/_2_  , \g45530/_0_  , \g45532/_0_  , \g45533/_0_  , \g45534/_0_  , \g45739/_2_  , \g45743/_2_  , \g45767/_0_  , \g45782/_0_  , \g45830/_3_  , \g45834/_3_  , \g45835/_3_  , \g45836/_3_  , \g45837/_3_  , \g45839/_3_  , \g45840/_3_  , \g45841/_3_  , \g45842/_3_  , \g45843/_3_  , \g45844/_3_  , \g45845/_3_  , \g46191/_0_  , \g46193/_3_  , \g46256/_3_  , \g46257/_3_  , \g46258/_3_  , \g46259/_3_  , \g46260/_3_  , \g46261/_3_  , \g46262/_3_  , \g46263/_3_  , \g46278/_0_  , \g46292/_0_  , \g46293/_0_  , \g46312/_0_  , \g46367/_2_  , \g46370/_2_  , \g46380/_2_  , \g46386/_2_  , \g46388/_2_  , \g46392/_2_  , \g46395/_2_  , \g46399/_2_  , \g46420/_0_  , \g46446/_0_  , \g46493/_0_  , \g46510/_0_  , \g46669/_2_  , \g46691/_0_  , \g46708/_0_  , \g46721/_00_  , \g46776/_0_  , \g46777/_0_  , \g46778/_0_  , \g46779/_0_  , \g46780/_0_  , \g46782/_0_  , \g46784/_0_  , \g46932/_0_  , \g47112/_0_  , \g47124/_0_  , \g47265/_0_  , \g47270/_0_  , \g47275/_0_  , \g47300/_1_  , \g47305/_1_  , \g47338/_0_  , \g47339/_0_  , \g47352/_0_  , \g47699/_3_  , \g47711/_0_  , \g47719/_3_  , \g47721/_3_  , \g47723/_3_  , \g47853/_0_  , \g48094/_0_  , \g48095/_0_  , \g48177/_2_  , \g48194/_0_  , \g48369/_2_  , \g48371/_2_  , \g48373/_2_  , \g48375/_2_  , \g48377/_2_  , \g48379/_2_  , \g48381/_2_  , \g48383/_2_  , \g48385/_2_  , \g48535/_0_  , \g48569/_0_  , \g48570/_0_  , \g48571/_0_  , \g48836/_0_  , \g48843/_0_  , \g49187/_3_  , \g49375/_2_  , \g49633/_0_  , \g49788/_1_  , \g49800/_1_  , \g49802/_1_  , \g49806/_1_  , \g49853/_1_  , \g49883/_0_  , \g49884/_0_  , \g49885/_0_  , \g49886/_0_  , \g49976/_1_  , \g50038/_0_  , \g50082/_0_  , \g50083/_0_  , \g50167/_3_  , \g50168/_3_  , \g50169/_3_  , \g50170/_3_  , \g50171/_3_  , \g50177/_0_  , \g50190/_0_  , \g50236/_0_  , \g50251/_3_  , \g50256/_0_  , \g50318/_3_  , \g50319/_3_  , \g50350/_3_  , \g50351/_3_  , \g50352/_3_  , \g50353/_3_  , \g50354/_3_  , \g50355/_3_  , \g50361/_2_  , \g50366/_0_  , \g50393/_0_  , \g50552/_1_  , \g51108/_0_  , \g51160/_0_  , \g51290/_1_  , \g51327/_3_  , \g51328/_3_  , \g51329/_3_  , \g51330/_3_  , \g51331/_3_  , \g51332/_3_  , \g51333/_3_  , \g51334/_3_  , \g51339/_3_  , \g51340/_3_  , \g51341/_3_  , \g51342/_3_  , \g51343/_3_  , \g51346/_0_  , \g51347/_0_  , \g51348/_0_  , \g51381/_3_  , \g51382/_3_  , \g51383/_3_  , \g51386/_3_  , \g51387/_3_  , \g51405/_3_  , \g51410/_3_  , \g51883/_0_  , \g51916/_0_  , \g51947/_0_  , \g51948/_0_  , \g51949/_0_  , \g51950/_0_  , \g51951/_0_  , \g51952/_0_  , \g51953/_0_  , \g51954/_0_  , \g51955/_0_  , \g51956/_0_  , \g51957/_0_  , \g51958/_0_  , \g51959/_0_  , \g51960/_0_  , \g51961/_0_  , \g51962/_0_  , \g51963/_0_  , \g51964/_0_  , \g51965/_0_  , \g51967/_0_  , \g51968/_0_  , \g51969/_0_  , \g51970/_0_  , \g51971/_0_  , \g51972/_0_  , \g51973/_0_  , \g51974/_0_  , \g51975/_0_  , \g51976/_0_  , \g51977/_0_  , \g51978/_0_  , \g51979/_0_  , \g51980/_0_  , \g51981/_0_  , \g51982/_0_  , \g51983/_0_  , \g51984/_0_  , \g51985/_0_  , \g51986/_0_  , \g51987/_0_  , \g51988/_0_  , \g51989/_0_  , \g51990/_0_  , \g51991/_0_  , \g51992/_0_  , \g51993/_0_  , \g51994/_0_  , \g51995/_0_  , \g51996/_0_  , \g51997/_0_  , \g51998/_0_  , \g51999/_0_  , \g52000/_0_  , \g52001/_0_  , \g52002/_0_  , \g52003/_0_  , \g52004/_0_  , \g52005/_0_  , \g52006/_0_  , \g52007/_0_  , \g52008/_0_  , \g52009/_0_  , \g52010/_0_  , \g52011/_0_  , \g52012/_0_  , \g52013/_0_  , \g52014/_0_  , \g52015/_0_  , \g52016/_0_  , \g52017/_0_  , \g52018/_0_  , \g52019/_0_  , \g52020/_0_  , \g52021/_0_  , \g52022/_0_  , \g52023/_0_  , \g52024/_0_  , \g52025/_0_  , \g52026/_0_  , \g52027/_0_  , \g52028/_0_  , \g52029/_0_  , \g52030/_0_  , \g52031/_0_  , \g52032/_0_  , \g52033/_0_  , \g52034/_0_  , \g52035/_0_  , \g52036/_0_  , \g52037/_0_  , \g52038/_0_  , \g52039/_0_  , \g52040/_0_  , \g52041/_0_  , \g52042/_0_  , \g52043/_0_  , \g52044/_0_  , \g52045/_0_  , \g52046/_0_  , \g52047/_0_  , \g52049/_0_  , \g52050/_0_  , \g52051/_0_  , \g52052/_0_  , \g52053/_0_  , \g52054/_0_  , \g52055/_0_  , \g52056/_0_  , \g52057/_0_  , \g52058/_0_  , \g52061/_0_  , \g52065/_0_  , \g52066/_0_  , \g52067/_0_  , \g52068/_0_  , \g52069/_0_  , \g52070/_0_  , \g52071/_0_  , \g52073/_0_  , \g52074/_0_  , \g52075/_0_  , \g52082/_0_  , \g52083/_0_  , \g52158/_0_  , \g52201/_0_  , \g52202/_0_  , \g52346/_0_  , \g52351/_0_  , \g52390/_0_  , \g52847/_0_  , \g52854/_0_  , \g52968/_0_  , \g52969/_0_  , \g52970/_0_  , \g52971/_0_  , \g52984/_0_  , \g52994/_0_  , \g53019/_0_  , \g53030/_0_  , \g53094/_1_  , \g53106/_0_  , \g53150/_0_  , \g53256/_0_  , \g53297/_0_  , \g53345/_0_  , \g53359/_0_  , \g53375/_0_  , \g53474/_1__syn_2  , \g53475/_2_  , \g53593/_0_  , \g53643/_1_  , \g53655/_0_  , \g53710/_0_  , \g53786/_0_  , \g53837/_0_  , \g53888/_1_  , \g53909/_0_  , \g54253/_2_  , \g54394/_3_  , \g54413/_0_  , \g55420/_0_  , \g55587/_0_  , \g55852/_0_  , \g57020/_0_  , \g59450/_0_  , \g59488/_2_  , \g59752/_0_  , \g59786/_0_  , \g59854/_0_  , \g59878/_0_  , \g59902/_0_  , \g59924/_0_  , \g59947/_0_  , \g59972/_0_  , \g59996/_0_  , \g60017/_0_  , \g60040/_0_  , \g60064/_0_  , \g60095/_0_  , \g60119/_0_  , \g60145/_1_  , \g60165/_0_  , \g60407/_2_  , \g60408/_0_  , \g60613/_2_  , \g60649/_0_  , \g60771/_0_  , \g60908/_1_  , \g60911/_0_  , \g60977/_0_  , \g61/_0_  , \g61002/_0_  , \g61308/_0_  , \g61312/_1_  , \g61314/_0_  , \g61319/_1_  , \g61342/_1_  , \g61360/_0_  , \g61377/_0_  , \g61423/_1_  , \g61426/_0_  , \g61479/_1_  , \g61523/_1_  , \g61558/_1_  , \g61652/_0_  , \g61866/_0_  , \g61868/_1_  , \g61887/_0_  , \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3  , \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3  , \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3  , \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3  , \u7_mc_we__reg/_05_  );
  input mc_cke_pad_o__pad ;
  input mc_vpen_pad_o_pad ;
  input \mem_ack_r_reg/P0001  ;
  input \poc_o[0]_pad  ;
  input \poc_o[10]_pad  ;
  input \poc_o[11]_pad  ;
  input \poc_o[12]_pad  ;
  input \poc_o[13]_pad  ;
  input \poc_o[14]_pad  ;
  input \poc_o[15]_pad  ;
  input \poc_o[16]_pad  ;
  input \poc_o[17]_pad  ;
  input \poc_o[18]_pad  ;
  input \poc_o[19]_pad  ;
  input \poc_o[1]_pad  ;
  input \poc_o[20]_pad  ;
  input \poc_o[21]_pad  ;
  input \poc_o[22]_pad  ;
  input \poc_o[23]_pad  ;
  input \poc_o[24]_pad  ;
  input \poc_o[25]_pad  ;
  input \poc_o[26]_pad  ;
  input \poc_o[27]_pad  ;
  input \poc_o[28]_pad  ;
  input \poc_o[29]_pad  ;
  input \poc_o[2]_pad  ;
  input \poc_o[30]_pad  ;
  input \poc_o[31]_pad  ;
  input \poc_o[3]_pad  ;
  input \poc_o[4]_pad  ;
  input \poc_o[5]_pad  ;
  input \poc_o[6]_pad  ;
  input \poc_o[7]_pad  ;
  input \poc_o[8]_pad  ;
  input \poc_o[9]_pad  ;
  input suspended_o_pad ;
  input \u0_cs_reg[0]/NET0131  ;
  input \u0_cs_reg[1]/NET0131  ;
  input \u0_csc_mask_r_reg[0]/NET0131  ;
  input \u0_csc_mask_r_reg[10]/NET0131  ;
  input \u0_csc_mask_r_reg[1]/NET0131  ;
  input \u0_csc_mask_r_reg[2]/NET0131  ;
  input \u0_csc_mask_r_reg[3]/NET0131  ;
  input \u0_csc_mask_r_reg[4]/NET0131  ;
  input \u0_csc_mask_r_reg[5]/NET0131  ;
  input \u0_csc_mask_r_reg[6]/NET0131  ;
  input \u0_csc_mask_r_reg[7]/NET0131  ;
  input \u0_csc_mask_r_reg[8]/NET0131  ;
  input \u0_csc_mask_r_reg[9]/NET0131  ;
  input \u0_csc_reg[10]/NET0131  ;
  input \u0_csc_reg[11]/NET0131  ;
  input \u0_csc_reg[1]/NET0131  ;
  input \u0_csc_reg[2]/NET0131  ;
  input \u0_csc_reg[3]/NET0131  ;
  input \u0_csc_reg[4]/NET0131  ;
  input \u0_csc_reg[5]/NET0131  ;
  input \u0_csc_reg[6]/NET0131  ;
  input \u0_csc_reg[7]/NET0131  ;
  input \u0_csc_reg[9]/NET0131  ;
  input \u0_csr_r2_reg[0]/NET0131  ;
  input \u0_csr_r2_reg[1]/NET0131  ;
  input \u0_csr_r2_reg[2]/NET0131  ;
  input \u0_csr_r2_reg[3]/NET0131  ;
  input \u0_csr_r2_reg[4]/NET0131  ;
  input \u0_csr_r2_reg[5]/NET0131  ;
  input \u0_csr_r2_reg[6]/NET0131  ;
  input \u0_csr_r2_reg[7]/NET0131  ;
  input \u0_csr_r_reg[0]/P0001  ;
  input \u0_csr_r_reg[10]/NET0131  ;
  input \u0_csr_r_reg[2]/NET0131  ;
  input \u0_csr_r_reg[3]/NET0131  ;
  input \u0_csr_r_reg[4]/NET0131  ;
  input \u0_csr_r_reg[5]/NET0131  ;
  input \u0_csr_r_reg[6]/NET0131  ;
  input \u0_csr_r_reg[7]/NET0131  ;
  input \u0_csr_r_reg[8]/NET0131  ;
  input \u0_csr_r_reg[9]/NET0131  ;
  input \u0_init_ack_r_reg/P0001  ;
  input \u0_init_req_reg/NET0131  ;
  input \u0_lmr_ack_r_reg/P0001  ;
  input \u0_lmr_req_reg/NET0131  ;
  input \u0_rf_we_reg/NET0131  ;
  input \u0_rst_r2_reg/NET0131  ;
  input \u0_sp_csc_reg[10]/NET0131  ;
  input \u0_sp_csc_reg[1]/NET0131  ;
  input \u0_sp_csc_reg[2]/NET0131  ;
  input \u0_sp_csc_reg[3]/NET0131  ;
  input \u0_sp_csc_reg[4]/NET0131  ;
  input \u0_sp_csc_reg[5]/NET0131  ;
  input \u0_sp_csc_reg[6]/NET0131  ;
  input \u0_sp_csc_reg[7]/NET0131  ;
  input \u0_sp_csc_reg[9]/NET0131  ;
  input \u0_sp_tms_reg[0]/NET0131  ;
  input \u0_sp_tms_reg[10]/NET0131  ;
  input \u0_sp_tms_reg[11]/NET0131  ;
  input \u0_sp_tms_reg[12]/NET0131  ;
  input \u0_sp_tms_reg[13]/NET0131  ;
  input \u0_sp_tms_reg[14]/NET0131  ;
  input \u0_sp_tms_reg[15]/NET0131  ;
  input \u0_sp_tms_reg[16]/NET0131  ;
  input \u0_sp_tms_reg[17]/NET0131  ;
  input \u0_sp_tms_reg[18]/NET0131  ;
  input \u0_sp_tms_reg[19]/NET0131  ;
  input \u0_sp_tms_reg[1]/NET0131  ;
  input \u0_sp_tms_reg[20]/NET0131  ;
  input \u0_sp_tms_reg[21]/NET0131  ;
  input \u0_sp_tms_reg[22]/NET0131  ;
  input \u0_sp_tms_reg[23]/NET0131  ;
  input \u0_sp_tms_reg[24]/NET0131  ;
  input \u0_sp_tms_reg[25]/NET0131  ;
  input \u0_sp_tms_reg[26]/NET0131  ;
  input \u0_sp_tms_reg[27]/NET0131  ;
  input \u0_sp_tms_reg[2]/NET0131  ;
  input \u0_sp_tms_reg[3]/NET0131  ;
  input \u0_sp_tms_reg[4]/NET0131  ;
  input \u0_sp_tms_reg[5]/NET0131  ;
  input \u0_sp_tms_reg[6]/NET0131  ;
  input \u0_sp_tms_reg[7]/NET0131  ;
  input \u0_sp_tms_reg[8]/NET0131  ;
  input \u0_sp_tms_reg[9]/NET0131  ;
  input \u0_spec_req_cs_reg[0]/NET0131  ;
  input \u0_spec_req_cs_reg[1]/NET0131  ;
  input \u0_sreq_cs_le_reg/NET0131  ;
  input \u0_tms_reg[0]/NET0131  ;
  input \u0_tms_reg[10]/NET0131  ;
  input \u0_tms_reg[11]/NET0131  ;
  input \u0_tms_reg[12]/NET0131  ;
  input \u0_tms_reg[13]/NET0131  ;
  input \u0_tms_reg[14]/NET0131  ;
  input \u0_tms_reg[15]/NET0131  ;
  input \u0_tms_reg[16]/NET0131  ;
  input \u0_tms_reg[17]/NET0131  ;
  input \u0_tms_reg[18]/NET0131  ;
  input \u0_tms_reg[19]/NET0131  ;
  input \u0_tms_reg[1]/NET0131  ;
  input \u0_tms_reg[20]/NET0131  ;
  input \u0_tms_reg[21]/NET0131  ;
  input \u0_tms_reg[22]/NET0131  ;
  input \u0_tms_reg[23]/NET0131  ;
  input \u0_tms_reg[24]/NET0131  ;
  input \u0_tms_reg[25]/NET0131  ;
  input \u0_tms_reg[26]/NET0131  ;
  input \u0_tms_reg[27]/NET0131  ;
  input \u0_tms_reg[2]/NET0131  ;
  input \u0_tms_reg[3]/NET0131  ;
  input \u0_tms_reg[4]/NET0131  ;
  input \u0_tms_reg[5]/NET0131  ;
  input \u0_tms_reg[6]/NET0131  ;
  input \u0_tms_reg[7]/NET0131  ;
  input \u0_tms_reg[8]/NET0131  ;
  input \u0_tms_reg[9]/NET0131  ;
  input \u0_u0_addr_r_reg[2]/P0001  ;
  input \u0_u0_addr_r_reg[3]/P0001  ;
  input \u0_u0_addr_r_reg[4]/P0001  ;
  input \u0_u0_addr_r_reg[5]/P0001  ;
  input \u0_u0_addr_r_reg[6]/P0001  ;
  input \u0_u0_csc_reg[0]/NET0131  ;
  input \u0_u0_csc_reg[10]/P0001  ;
  input \u0_u0_csc_reg[11]/P0001  ;
  input \u0_u0_csc_reg[12]/P0001  ;
  input \u0_u0_csc_reg[13]/P0001  ;
  input \u0_u0_csc_reg[14]/P0001  ;
  input \u0_u0_csc_reg[15]/P0001  ;
  input \u0_u0_csc_reg[16]/P0001  ;
  input \u0_u0_csc_reg[17]/P0001  ;
  input \u0_u0_csc_reg[18]/P0001  ;
  input \u0_u0_csc_reg[19]/P0001  ;
  input \u0_u0_csc_reg[1]/NET0131  ;
  input \u0_u0_csc_reg[20]/P0001  ;
  input \u0_u0_csc_reg[21]/P0001  ;
  input \u0_u0_csc_reg[22]/P0001  ;
  input \u0_u0_csc_reg[23]/P0001  ;
  input \u0_u0_csc_reg[24]/P0001  ;
  input \u0_u0_csc_reg[25]/P0001  ;
  input \u0_u0_csc_reg[26]/P0001  ;
  input \u0_u0_csc_reg[27]/P0001  ;
  input \u0_u0_csc_reg[28]/P0001  ;
  input \u0_u0_csc_reg[29]/P0001  ;
  input \u0_u0_csc_reg[2]/NET0131  ;
  input \u0_u0_csc_reg[30]/P0001  ;
  input \u0_u0_csc_reg[31]/P0001  ;
  input \u0_u0_csc_reg[3]/NET0131  ;
  input \u0_u0_csc_reg[4]/P0001  ;
  input \u0_u0_csc_reg[5]/P0001  ;
  input \u0_u0_csc_reg[6]/P0001  ;
  input \u0_u0_csc_reg[7]/P0001  ;
  input \u0_u0_csc_reg[8]/P0001  ;
  input \u0_u0_csc_reg[9]/P0001  ;
  input \u0_u0_init_req_reg/NET0131  ;
  input \u0_u0_init_req_we_reg/NET0131  ;
  input \u0_u0_inited_reg/NET0131  ;
  input \u0_u0_lmr_req_reg/NET0131  ;
  input \u0_u0_lmr_req_we_reg/NET0131  ;
  input \u0_u0_tms_reg[0]/P0001  ;
  input \u0_u0_tms_reg[10]/P0001  ;
  input \u0_u0_tms_reg[11]/P0001  ;
  input \u0_u0_tms_reg[12]/P0001  ;
  input \u0_u0_tms_reg[13]/P0001  ;
  input \u0_u0_tms_reg[14]/P0001  ;
  input \u0_u0_tms_reg[15]/P0001  ;
  input \u0_u0_tms_reg[16]/P0001  ;
  input \u0_u0_tms_reg[17]/P0001  ;
  input \u0_u0_tms_reg[18]/P0001  ;
  input \u0_u0_tms_reg[19]/P0001  ;
  input \u0_u0_tms_reg[1]/P0001  ;
  input \u0_u0_tms_reg[20]/P0001  ;
  input \u0_u0_tms_reg[21]/P0001  ;
  input \u0_u0_tms_reg[22]/P0001  ;
  input \u0_u0_tms_reg[23]/P0001  ;
  input \u0_u0_tms_reg[24]/P0001  ;
  input \u0_u0_tms_reg[25]/P0001  ;
  input \u0_u0_tms_reg[26]/P0001  ;
  input \u0_u0_tms_reg[27]/P0001  ;
  input \u0_u0_tms_reg[28]/P0001  ;
  input \u0_u0_tms_reg[29]/P0001  ;
  input \u0_u0_tms_reg[2]/P0001  ;
  input \u0_u0_tms_reg[30]/P0001  ;
  input \u0_u0_tms_reg[31]/P0001  ;
  input \u0_u0_tms_reg[3]/P0001  ;
  input \u0_u0_tms_reg[4]/P0001  ;
  input \u0_u0_tms_reg[5]/P0001  ;
  input \u0_u0_tms_reg[6]/P0001  ;
  input \u0_u0_tms_reg[7]/P0001  ;
  input \u0_u0_tms_reg[8]/P0001  ;
  input \u0_u0_tms_reg[9]/P0001  ;
  input \u0_u1_csc_reg[0]/NET0131  ;
  input \u0_u1_csc_reg[10]/P0001  ;
  input \u0_u1_csc_reg[11]/P0001  ;
  input \u0_u1_csc_reg[12]/P0001  ;
  input \u0_u1_csc_reg[13]/P0001  ;
  input \u0_u1_csc_reg[14]/P0001  ;
  input \u0_u1_csc_reg[15]/P0001  ;
  input \u0_u1_csc_reg[16]/P0001  ;
  input \u0_u1_csc_reg[17]/P0001  ;
  input \u0_u1_csc_reg[18]/P0001  ;
  input \u0_u1_csc_reg[19]/P0001  ;
  input \u0_u1_csc_reg[1]/NET0131  ;
  input \u0_u1_csc_reg[20]/P0001  ;
  input \u0_u1_csc_reg[21]/P0001  ;
  input \u0_u1_csc_reg[22]/P0001  ;
  input \u0_u1_csc_reg[23]/P0001  ;
  input \u0_u1_csc_reg[24]/P0001  ;
  input \u0_u1_csc_reg[25]/P0001  ;
  input \u0_u1_csc_reg[26]/P0001  ;
  input \u0_u1_csc_reg[27]/P0001  ;
  input \u0_u1_csc_reg[28]/P0001  ;
  input \u0_u1_csc_reg[29]/P0001  ;
  input \u0_u1_csc_reg[2]/NET0131  ;
  input \u0_u1_csc_reg[30]/P0001  ;
  input \u0_u1_csc_reg[31]/P0001  ;
  input \u0_u1_csc_reg[3]/NET0131  ;
  input \u0_u1_csc_reg[4]/P0001  ;
  input \u0_u1_csc_reg[5]/P0001  ;
  input \u0_u1_csc_reg[6]/P0001  ;
  input \u0_u1_csc_reg[7]/P0001  ;
  input \u0_u1_csc_reg[8]/P0001  ;
  input \u0_u1_csc_reg[9]/P0001  ;
  input \u0_u1_init_req_reg/NET0131  ;
  input \u0_u1_init_req_we_reg/NET0131  ;
  input \u0_u1_inited_reg/NET0131  ;
  input \u0_u1_lmr_req_reg/NET0131  ;
  input \u0_u1_lmr_req_we_reg/NET0131  ;
  input \u0_u1_tms_reg[0]/P0001  ;
  input \u0_u1_tms_reg[10]/P0001  ;
  input \u0_u1_tms_reg[11]/P0001  ;
  input \u0_u1_tms_reg[12]/P0001  ;
  input \u0_u1_tms_reg[13]/P0001  ;
  input \u0_u1_tms_reg[14]/P0001  ;
  input \u0_u1_tms_reg[15]/P0001  ;
  input \u0_u1_tms_reg[16]/P0001  ;
  input \u0_u1_tms_reg[17]/P0001  ;
  input \u0_u1_tms_reg[18]/P0001  ;
  input \u0_u1_tms_reg[19]/P0001  ;
  input \u0_u1_tms_reg[1]/P0001  ;
  input \u0_u1_tms_reg[20]/P0001  ;
  input \u0_u1_tms_reg[21]/P0001  ;
  input \u0_u1_tms_reg[22]/P0001  ;
  input \u0_u1_tms_reg[23]/P0001  ;
  input \u0_u1_tms_reg[24]/P0001  ;
  input \u0_u1_tms_reg[25]/P0001  ;
  input \u0_u1_tms_reg[26]/P0001  ;
  input \u0_u1_tms_reg[27]/P0001  ;
  input \u0_u1_tms_reg[28]/P0001  ;
  input \u0_u1_tms_reg[29]/P0001  ;
  input \u0_u1_tms_reg[2]/P0001  ;
  input \u0_u1_tms_reg[30]/P0001  ;
  input \u0_u1_tms_reg[31]/P0001  ;
  input \u0_u1_tms_reg[3]/P0001  ;
  input \u0_u1_tms_reg[4]/P0001  ;
  input \u0_u1_tms_reg[5]/P0001  ;
  input \u0_u1_tms_reg[6]/P0001  ;
  input \u0_u1_tms_reg[7]/P0001  ;
  input \u0_u1_tms_reg[8]/P0001  ;
  input \u0_u1_tms_reg[9]/P0001  ;
  input \u0_wp_err_reg/NET0131  ;
  input \u1_acs_addr_reg[0]/P0001  ;
  input \u1_acs_addr_reg[10]/P0001  ;
  input \u1_acs_addr_reg[11]/P0001  ;
  input \u1_acs_addr_reg[12]/P0001  ;
  input \u1_acs_addr_reg[13]/P0001  ;
  input \u1_acs_addr_reg[14]/P0001  ;
  input \u1_acs_addr_reg[15]/P0001  ;
  input \u1_acs_addr_reg[16]/P0001  ;
  input \u1_acs_addr_reg[17]/P0001  ;
  input \u1_acs_addr_reg[18]/P0001  ;
  input \u1_acs_addr_reg[19]/P0001  ;
  input \u1_acs_addr_reg[1]/P0001  ;
  input \u1_acs_addr_reg[20]/P0001  ;
  input \u1_acs_addr_reg[21]/P0001  ;
  input \u1_acs_addr_reg[22]/P0001  ;
  input \u1_acs_addr_reg[23]/P0001  ;
  input \u1_acs_addr_reg[2]/P0001  ;
  input \u1_acs_addr_reg[3]/P0001  ;
  input \u1_acs_addr_reg[4]/P0001  ;
  input \u1_acs_addr_reg[5]/P0001  ;
  input \u1_acs_addr_reg[6]/P0001  ;
  input \u1_acs_addr_reg[7]/P0001  ;
  input \u1_acs_addr_reg[8]/P0001  ;
  input \u1_acs_addr_reg[9]/P0001  ;
  input \u1_bank_adr_reg[0]/P0001  ;
  input \u1_bank_adr_reg[1]/P0001  ;
  input \u1_col_adr_reg[0]/P0001  ;
  input \u1_col_adr_reg[1]/P0001  ;
  input \u1_col_adr_reg[2]/P0001  ;
  input \u1_col_adr_reg[3]/P0001  ;
  input \u1_col_adr_reg[4]/P0001  ;
  input \u1_col_adr_reg[5]/P0001  ;
  input \u1_col_adr_reg[6]/P0001  ;
  input \u1_col_adr_reg[7]/P0001  ;
  input \u1_col_adr_reg[8]/P0001  ;
  input \u1_col_adr_reg[9]/P0001  ;
  input \u1_row_adr_reg[0]/P0001  ;
  input \u1_row_adr_reg[10]/P0001  ;
  input \u1_row_adr_reg[11]/P0001  ;
  input \u1_row_adr_reg[12]/P0001  ;
  input \u1_row_adr_reg[1]/P0001  ;
  input \u1_row_adr_reg[2]/P0001  ;
  input \u1_row_adr_reg[3]/P0001  ;
  input \u1_row_adr_reg[4]/P0001  ;
  input \u1_row_adr_reg[5]/P0001  ;
  input \u1_row_adr_reg[6]/P0001  ;
  input \u1_row_adr_reg[7]/P0001  ;
  input \u1_row_adr_reg[8]/P0001  ;
  input \u1_row_adr_reg[9]/P0001  ;
  input \u1_sram_addr_reg[0]/P0001  ;
  input \u1_sram_addr_reg[10]/P0001  ;
  input \u1_sram_addr_reg[11]/P0001  ;
  input \u1_sram_addr_reg[12]/P0001  ;
  input \u1_sram_addr_reg[13]/P0001  ;
  input \u1_sram_addr_reg[14]/P0001  ;
  input \u1_sram_addr_reg[15]/P0001  ;
  input \u1_sram_addr_reg[16]/P0001  ;
  input \u1_sram_addr_reg[17]/P0001  ;
  input \u1_sram_addr_reg[18]/P0001  ;
  input \u1_sram_addr_reg[19]/P0001  ;
  input \u1_sram_addr_reg[1]/P0001  ;
  input \u1_sram_addr_reg[20]/P0001  ;
  input \u1_sram_addr_reg[21]/P0001  ;
  input \u1_sram_addr_reg[22]/P0001  ;
  input \u1_sram_addr_reg[23]/P0001  ;
  input \u1_sram_addr_reg[2]/P0001  ;
  input \u1_sram_addr_reg[3]/P0001  ;
  input \u1_sram_addr_reg[4]/P0001  ;
  input \u1_sram_addr_reg[5]/P0001  ;
  input \u1_sram_addr_reg[6]/P0001  ;
  input \u1_sram_addr_reg[7]/P0001  ;
  input \u1_sram_addr_reg[8]/P0001  ;
  input \u1_sram_addr_reg[9]/P0001  ;
  input \u1_u0_out_r_reg[0]/P0001  ;
  input \u1_u0_out_r_reg[10]/P0001  ;
  input \u1_u0_out_r_reg[11]/P0001  ;
  input \u1_u0_out_r_reg[12]/P0001  ;
  input \u1_u0_out_r_reg[1]/P0001  ;
  input \u1_u0_out_r_reg[2]/P0001  ;
  input \u1_u0_out_r_reg[3]/P0001  ;
  input \u1_u0_out_r_reg[4]/P0001  ;
  input \u1_u0_out_r_reg[5]/P0001  ;
  input \u1_u0_out_r_reg[6]/P0001  ;
  input \u1_u0_out_r_reg[7]/P0001  ;
  input \u1_u0_out_r_reg[8]/P0001  ;
  input \u1_u0_out_r_reg[9]/P0001  ;
  input \u2_bank_open_reg/P0001  ;
  input \u2_row_same_reg/P0001  ;
  input \u2_u0_b0_last_row_reg[0]/P0001  ;
  input \u2_u0_b0_last_row_reg[10]/P0001  ;
  input \u2_u0_b0_last_row_reg[11]/P0001  ;
  input \u2_u0_b0_last_row_reg[12]/P0001  ;
  input \u2_u0_b0_last_row_reg[1]/P0001  ;
  input \u2_u0_b0_last_row_reg[2]/P0001  ;
  input \u2_u0_b0_last_row_reg[3]/P0001  ;
  input \u2_u0_b0_last_row_reg[4]/P0001  ;
  input \u2_u0_b0_last_row_reg[5]/P0001  ;
  input \u2_u0_b0_last_row_reg[6]/P0001  ;
  input \u2_u0_b0_last_row_reg[7]/P0001  ;
  input \u2_u0_b0_last_row_reg[8]/P0001  ;
  input \u2_u0_b0_last_row_reg[9]/P0001  ;
  input \u2_u0_b1_last_row_reg[0]/P0001  ;
  input \u2_u0_b1_last_row_reg[10]/P0001  ;
  input \u2_u0_b1_last_row_reg[11]/P0001  ;
  input \u2_u0_b1_last_row_reg[12]/P0001  ;
  input \u2_u0_b1_last_row_reg[1]/P0001  ;
  input \u2_u0_b1_last_row_reg[2]/P0001  ;
  input \u2_u0_b1_last_row_reg[3]/P0001  ;
  input \u2_u0_b1_last_row_reg[4]/P0001  ;
  input \u2_u0_b1_last_row_reg[5]/P0001  ;
  input \u2_u0_b1_last_row_reg[6]/P0001  ;
  input \u2_u0_b1_last_row_reg[7]/P0001  ;
  input \u2_u0_b1_last_row_reg[8]/P0001  ;
  input \u2_u0_b1_last_row_reg[9]/P0001  ;
  input \u2_u0_b2_last_row_reg[0]/P0001  ;
  input \u2_u0_b2_last_row_reg[10]/P0001  ;
  input \u2_u0_b2_last_row_reg[11]/P0001  ;
  input \u2_u0_b2_last_row_reg[12]/P0001  ;
  input \u2_u0_b2_last_row_reg[1]/P0001  ;
  input \u2_u0_b2_last_row_reg[2]/P0001  ;
  input \u2_u0_b2_last_row_reg[3]/P0001  ;
  input \u2_u0_b2_last_row_reg[4]/P0001  ;
  input \u2_u0_b2_last_row_reg[5]/P0001  ;
  input \u2_u0_b2_last_row_reg[6]/P0001  ;
  input \u2_u0_b2_last_row_reg[7]/P0001  ;
  input \u2_u0_b2_last_row_reg[8]/P0001  ;
  input \u2_u0_b2_last_row_reg[9]/P0001  ;
  input \u2_u0_b3_last_row_reg[0]/P0001  ;
  input \u2_u0_b3_last_row_reg[10]/P0001  ;
  input \u2_u0_b3_last_row_reg[11]/P0001  ;
  input \u2_u0_b3_last_row_reg[12]/P0001  ;
  input \u2_u0_b3_last_row_reg[1]/P0001  ;
  input \u2_u0_b3_last_row_reg[2]/P0001  ;
  input \u2_u0_b3_last_row_reg[3]/P0001  ;
  input \u2_u0_b3_last_row_reg[4]/P0001  ;
  input \u2_u0_b3_last_row_reg[5]/P0001  ;
  input \u2_u0_b3_last_row_reg[6]/P0001  ;
  input \u2_u0_b3_last_row_reg[7]/P0001  ;
  input \u2_u0_b3_last_row_reg[8]/P0001  ;
  input \u2_u0_b3_last_row_reg[9]/P0001  ;
  input \u2_u0_bank0_open_reg/NET0131  ;
  input \u2_u0_bank1_open_reg/NET0131  ;
  input \u2_u0_bank2_open_reg/NET0131  ;
  input \u2_u0_bank3_open_reg/NET0131  ;
  input \u2_u1_b0_last_row_reg[0]/P0001  ;
  input \u2_u1_b0_last_row_reg[10]/P0001  ;
  input \u2_u1_b0_last_row_reg[11]/P0001  ;
  input \u2_u1_b0_last_row_reg[12]/P0001  ;
  input \u2_u1_b0_last_row_reg[1]/P0001  ;
  input \u2_u1_b0_last_row_reg[2]/P0001  ;
  input \u2_u1_b0_last_row_reg[3]/P0001  ;
  input \u2_u1_b0_last_row_reg[4]/P0001  ;
  input \u2_u1_b0_last_row_reg[5]/P0001  ;
  input \u2_u1_b0_last_row_reg[6]/P0001  ;
  input \u2_u1_b0_last_row_reg[7]/P0001  ;
  input \u2_u1_b0_last_row_reg[8]/P0001  ;
  input \u2_u1_b0_last_row_reg[9]/P0001  ;
  input \u2_u1_b1_last_row_reg[0]/P0001  ;
  input \u2_u1_b1_last_row_reg[10]/P0001  ;
  input \u2_u1_b1_last_row_reg[11]/P0001  ;
  input \u2_u1_b1_last_row_reg[12]/P0001  ;
  input \u2_u1_b1_last_row_reg[1]/P0001  ;
  input \u2_u1_b1_last_row_reg[2]/P0001  ;
  input \u2_u1_b1_last_row_reg[3]/P0001  ;
  input \u2_u1_b1_last_row_reg[4]/P0001  ;
  input \u2_u1_b1_last_row_reg[5]/P0001  ;
  input \u2_u1_b1_last_row_reg[6]/P0001  ;
  input \u2_u1_b1_last_row_reg[7]/P0001  ;
  input \u2_u1_b1_last_row_reg[8]/P0001  ;
  input \u2_u1_b1_last_row_reg[9]/P0001  ;
  input \u2_u1_b2_last_row_reg[0]/P0001  ;
  input \u2_u1_b2_last_row_reg[10]/P0001  ;
  input \u2_u1_b2_last_row_reg[11]/P0001  ;
  input \u2_u1_b2_last_row_reg[12]/P0001  ;
  input \u2_u1_b2_last_row_reg[1]/P0001  ;
  input \u2_u1_b2_last_row_reg[2]/P0001  ;
  input \u2_u1_b2_last_row_reg[3]/P0001  ;
  input \u2_u1_b2_last_row_reg[4]/P0001  ;
  input \u2_u1_b2_last_row_reg[5]/P0001  ;
  input \u2_u1_b2_last_row_reg[6]/P0001  ;
  input \u2_u1_b2_last_row_reg[7]/P0001  ;
  input \u2_u1_b2_last_row_reg[8]/P0001  ;
  input \u2_u1_b2_last_row_reg[9]/P0001  ;
  input \u2_u1_b3_last_row_reg[0]/P0001  ;
  input \u2_u1_b3_last_row_reg[10]/P0001  ;
  input \u2_u1_b3_last_row_reg[11]/P0001  ;
  input \u2_u1_b3_last_row_reg[12]/P0001  ;
  input \u2_u1_b3_last_row_reg[1]/P0001  ;
  input \u2_u1_b3_last_row_reg[2]/P0001  ;
  input \u2_u1_b3_last_row_reg[3]/P0001  ;
  input \u2_u1_b3_last_row_reg[4]/P0001  ;
  input \u2_u1_b3_last_row_reg[5]/P0001  ;
  input \u2_u1_b3_last_row_reg[6]/P0001  ;
  input \u2_u1_b3_last_row_reg[7]/P0001  ;
  input \u2_u1_b3_last_row_reg[8]/P0001  ;
  input \u2_u1_b3_last_row_reg[9]/P0001  ;
  input \u2_u1_bank0_open_reg/NET0131  ;
  input \u2_u1_bank1_open_reg/NET0131  ;
  input \u2_u1_bank2_open_reg/NET0131  ;
  input \u2_u1_bank3_open_reg/NET0131  ;
  input \u3_byte0_reg[0]/P0001  ;
  input \u3_byte0_reg[1]/P0001  ;
  input \u3_byte0_reg[2]/P0001  ;
  input \u3_byte0_reg[3]/P0001  ;
  input \u3_byte0_reg[4]/P0001  ;
  input \u3_byte0_reg[5]/P0001  ;
  input \u3_byte0_reg[6]/P0001  ;
  input \u3_byte0_reg[7]/P0001  ;
  input \u3_byte1_reg[0]/P0001  ;
  input \u3_byte1_reg[1]/P0001  ;
  input \u3_byte1_reg[2]/P0001  ;
  input \u3_byte1_reg[3]/P0001  ;
  input \u3_byte1_reg[4]/P0001  ;
  input \u3_byte1_reg[5]/P0001  ;
  input \u3_byte1_reg[6]/P0001  ;
  input \u3_byte1_reg[7]/P0001  ;
  input \u3_byte2_reg[0]/P0001  ;
  input \u3_byte2_reg[1]/P0001  ;
  input \u3_byte2_reg[2]/P0001  ;
  input \u3_byte2_reg[3]/P0001  ;
  input \u3_byte2_reg[4]/P0001  ;
  input \u3_byte2_reg[5]/P0001  ;
  input \u3_byte2_reg[6]/P0001  ;
  input \u3_byte2_reg[7]/P0001  ;
  input \u3_u0_r0_reg[0]/P0001  ;
  input \u3_u0_r0_reg[10]/P0001  ;
  input \u3_u0_r0_reg[11]/P0001  ;
  input \u3_u0_r0_reg[12]/P0001  ;
  input \u3_u0_r0_reg[13]/P0001  ;
  input \u3_u0_r0_reg[14]/P0001  ;
  input \u3_u0_r0_reg[15]/P0001  ;
  input \u3_u0_r0_reg[16]/P0001  ;
  input \u3_u0_r0_reg[17]/P0001  ;
  input \u3_u0_r0_reg[18]/P0001  ;
  input \u3_u0_r0_reg[19]/P0001  ;
  input \u3_u0_r0_reg[1]/P0001  ;
  input \u3_u0_r0_reg[20]/P0001  ;
  input \u3_u0_r0_reg[21]/P0001  ;
  input \u3_u0_r0_reg[22]/P0001  ;
  input \u3_u0_r0_reg[23]/P0001  ;
  input \u3_u0_r0_reg[24]/P0001  ;
  input \u3_u0_r0_reg[25]/P0001  ;
  input \u3_u0_r0_reg[26]/P0001  ;
  input \u3_u0_r0_reg[27]/P0001  ;
  input \u3_u0_r0_reg[28]/P0001  ;
  input \u3_u0_r0_reg[29]/P0001  ;
  input \u3_u0_r0_reg[2]/P0001  ;
  input \u3_u0_r0_reg[30]/P0001  ;
  input \u3_u0_r0_reg[31]/P0001  ;
  input \u3_u0_r0_reg[32]/P0001  ;
  input \u3_u0_r0_reg[33]/P0001  ;
  input \u3_u0_r0_reg[34]/P0001  ;
  input \u3_u0_r0_reg[35]/P0001  ;
  input \u3_u0_r0_reg[3]/P0001  ;
  input \u3_u0_r0_reg[4]/P0001  ;
  input \u3_u0_r0_reg[5]/P0001  ;
  input \u3_u0_r0_reg[6]/P0001  ;
  input \u3_u0_r0_reg[7]/P0001  ;
  input \u3_u0_r0_reg[8]/P0001  ;
  input \u3_u0_r0_reg[9]/P0001  ;
  input \u3_u0_r1_reg[0]/P0001  ;
  input \u3_u0_r1_reg[10]/P0001  ;
  input \u3_u0_r1_reg[11]/P0001  ;
  input \u3_u0_r1_reg[12]/P0001  ;
  input \u3_u0_r1_reg[13]/P0001  ;
  input \u3_u0_r1_reg[14]/P0001  ;
  input \u3_u0_r1_reg[15]/P0001  ;
  input \u3_u0_r1_reg[16]/P0001  ;
  input \u3_u0_r1_reg[17]/P0001  ;
  input \u3_u0_r1_reg[18]/P0001  ;
  input \u3_u0_r1_reg[19]/P0001  ;
  input \u3_u0_r1_reg[1]/P0001  ;
  input \u3_u0_r1_reg[20]/P0001  ;
  input \u3_u0_r1_reg[21]/P0001  ;
  input \u3_u0_r1_reg[22]/P0001  ;
  input \u3_u0_r1_reg[23]/P0001  ;
  input \u3_u0_r1_reg[24]/P0001  ;
  input \u3_u0_r1_reg[25]/P0001  ;
  input \u3_u0_r1_reg[26]/P0001  ;
  input \u3_u0_r1_reg[27]/P0001  ;
  input \u3_u0_r1_reg[28]/P0001  ;
  input \u3_u0_r1_reg[29]/P0001  ;
  input \u3_u0_r1_reg[2]/P0001  ;
  input \u3_u0_r1_reg[30]/P0001  ;
  input \u3_u0_r1_reg[31]/P0001  ;
  input \u3_u0_r1_reg[32]/P0001  ;
  input \u3_u0_r1_reg[33]/P0001  ;
  input \u3_u0_r1_reg[34]/P0001  ;
  input \u3_u0_r1_reg[35]/P0001  ;
  input \u3_u0_r1_reg[3]/P0001  ;
  input \u3_u0_r1_reg[4]/P0001  ;
  input \u3_u0_r1_reg[5]/P0001  ;
  input \u3_u0_r1_reg[6]/P0001  ;
  input \u3_u0_r1_reg[7]/P0001  ;
  input \u3_u0_r1_reg[8]/P0001  ;
  input \u3_u0_r1_reg[9]/P0001  ;
  input \u3_u0_r2_reg[0]/P0001  ;
  input \u3_u0_r2_reg[10]/P0001  ;
  input \u3_u0_r2_reg[11]/P0001  ;
  input \u3_u0_r2_reg[12]/P0001  ;
  input \u3_u0_r2_reg[13]/P0001  ;
  input \u3_u0_r2_reg[14]/P0001  ;
  input \u3_u0_r2_reg[15]/P0001  ;
  input \u3_u0_r2_reg[16]/P0001  ;
  input \u3_u0_r2_reg[17]/P0001  ;
  input \u3_u0_r2_reg[18]/P0001  ;
  input \u3_u0_r2_reg[19]/P0001  ;
  input \u3_u0_r2_reg[1]/P0001  ;
  input \u3_u0_r2_reg[20]/P0001  ;
  input \u3_u0_r2_reg[21]/P0001  ;
  input \u3_u0_r2_reg[22]/P0001  ;
  input \u3_u0_r2_reg[23]/P0001  ;
  input \u3_u0_r2_reg[24]/P0001  ;
  input \u3_u0_r2_reg[25]/P0001  ;
  input \u3_u0_r2_reg[26]/P0001  ;
  input \u3_u0_r2_reg[27]/P0001  ;
  input \u3_u0_r2_reg[28]/P0001  ;
  input \u3_u0_r2_reg[29]/P0001  ;
  input \u3_u0_r2_reg[2]/P0001  ;
  input \u3_u0_r2_reg[30]/P0001  ;
  input \u3_u0_r2_reg[31]/P0001  ;
  input \u3_u0_r2_reg[32]/P0001  ;
  input \u3_u0_r2_reg[33]/P0001  ;
  input \u3_u0_r2_reg[34]/P0001  ;
  input \u3_u0_r2_reg[35]/P0001  ;
  input \u3_u0_r2_reg[3]/P0001  ;
  input \u3_u0_r2_reg[4]/P0001  ;
  input \u3_u0_r2_reg[5]/P0001  ;
  input \u3_u0_r2_reg[6]/P0001  ;
  input \u3_u0_r2_reg[7]/P0001  ;
  input \u3_u0_r2_reg[8]/P0001  ;
  input \u3_u0_r2_reg[9]/P0001  ;
  input \u3_u0_r3_reg[0]/P0001  ;
  input \u3_u0_r3_reg[10]/P0001  ;
  input \u3_u0_r3_reg[11]/P0001  ;
  input \u3_u0_r3_reg[12]/P0001  ;
  input \u3_u0_r3_reg[13]/P0001  ;
  input \u3_u0_r3_reg[14]/P0001  ;
  input \u3_u0_r3_reg[15]/P0001  ;
  input \u3_u0_r3_reg[16]/P0001  ;
  input \u3_u0_r3_reg[17]/P0001  ;
  input \u3_u0_r3_reg[18]/P0001  ;
  input \u3_u0_r3_reg[19]/P0001  ;
  input \u3_u0_r3_reg[1]/P0001  ;
  input \u3_u0_r3_reg[20]/P0001  ;
  input \u3_u0_r3_reg[21]/P0001  ;
  input \u3_u0_r3_reg[22]/P0001  ;
  input \u3_u0_r3_reg[23]/P0001  ;
  input \u3_u0_r3_reg[24]/P0001  ;
  input \u3_u0_r3_reg[25]/P0001  ;
  input \u3_u0_r3_reg[26]/P0001  ;
  input \u3_u0_r3_reg[27]/P0001  ;
  input \u3_u0_r3_reg[28]/P0001  ;
  input \u3_u0_r3_reg[29]/P0001  ;
  input \u3_u0_r3_reg[2]/P0001  ;
  input \u3_u0_r3_reg[30]/P0001  ;
  input \u3_u0_r3_reg[31]/P0001  ;
  input \u3_u0_r3_reg[32]/P0001  ;
  input \u3_u0_r3_reg[33]/P0001  ;
  input \u3_u0_r3_reg[34]/P0001  ;
  input \u3_u0_r3_reg[35]/P0001  ;
  input \u3_u0_r3_reg[3]/P0001  ;
  input \u3_u0_r3_reg[4]/P0001  ;
  input \u3_u0_r3_reg[5]/P0001  ;
  input \u3_u0_r3_reg[6]/P0001  ;
  input \u3_u0_r3_reg[7]/P0001  ;
  input \u3_u0_r3_reg[8]/P0001  ;
  input \u3_u0_r3_reg[9]/P0001  ;
  input \u3_u0_rd_adr_reg[0]/NET0131  ;
  input \u3_u0_rd_adr_reg[1]/NET0131  ;
  input \u3_u0_rd_adr_reg[2]/NET0131  ;
  input \u3_u0_rd_adr_reg[3]/NET0131  ;
  input \u3_u0_wr_adr_reg[0]/NET0131  ;
  input \u3_u0_wr_adr_reg[1]/NET0131  ;
  input \u3_u0_wr_adr_reg[2]/NET0131  ;
  input \u3_u0_wr_adr_reg[3]/NET0131  ;
  input \u4_ps_cnt_reg[0]/NET0131  ;
  input \u4_ps_cnt_reg[1]/NET0131  ;
  input \u4_ps_cnt_reg[2]/NET0131  ;
  input \u4_ps_cnt_reg[3]/NET0131  ;
  input \u4_ps_cnt_reg[4]/NET0131  ;
  input \u4_ps_cnt_reg[5]/NET0131  ;
  input \u4_ps_cnt_reg[6]/NET0131  ;
  input \u4_ps_cnt_reg[7]/NET0131  ;
  input \u4_rfr_ce_reg/NET0131  ;
  input \u4_rfr_clr_reg/P0001  ;
  input \u4_rfr_cnt_reg[0]/NET0131  ;
  input \u4_rfr_cnt_reg[1]/NET0131  ;
  input \u4_rfr_cnt_reg[2]/NET0131  ;
  input \u4_rfr_cnt_reg[3]/NET0131  ;
  input \u4_rfr_cnt_reg[4]/NET0131  ;
  input \u4_rfr_cnt_reg[5]/NET0131  ;
  input \u4_rfr_cnt_reg[6]/NET0131  ;
  input \u4_rfr_cnt_reg[7]/NET0131  ;
  input \u4_rfr_early_reg/NET0131  ;
  input \u4_rfr_en_reg/NET0131  ;
  input \u4_rfr_req_reg/NET0131  ;
  input \u5_ack_cnt_reg[0]/NET0131  ;
  input \u5_ack_cnt_reg[1]/NET0131  ;
  input \u5_ack_cnt_reg[2]/NET0131  ;
  input \u5_ack_cnt_reg[3]/NET0131  ;
  input \u5_ap_en_reg/NET0131  ;
  input \u5_burst_act_rd_reg/P0001  ;
  input \u5_burst_cnt_reg[0]/NET0131  ;
  input \u5_burst_cnt_reg[10]/NET0131  ;
  input \u5_burst_cnt_reg[1]/NET0131  ;
  input \u5_burst_cnt_reg[2]/NET0131  ;
  input \u5_burst_cnt_reg[3]/NET0131  ;
  input \u5_burst_cnt_reg[4]/NET0131  ;
  input \u5_burst_cnt_reg[5]/NET0131  ;
  input \u5_burst_cnt_reg[6]/NET0131  ;
  input \u5_burst_cnt_reg[7]/NET0131  ;
  input \u5_burst_cnt_reg[8]/NET0131  ;
  input \u5_burst_cnt_reg[9]/NET0131  ;
  input \u5_cke_o_del_reg/P0001  ;
  input \u5_cke_r_reg/NET0131  ;
  input \u5_cmd_a10_r_reg/P0001  ;
  input \u5_cmd_asserted2_reg/NET0131  ;
  input \u5_cmd_asserted_reg/NET0131  ;
  input \u5_cmd_del_reg[0]/NET0131  ;
  input \u5_cmd_del_reg[1]/NET0131  ;
  input \u5_cmd_del_reg[2]/NET0131  ;
  input \u5_cmd_del_reg[3]/NET0131  ;
  input \u5_cnt_reg/NET0131  ;
  input \u5_cs_le_r_reg/P0001  ;
  input \u5_cs_le_reg/P0001  ;
  input \u5_data_oe_r2_reg/NET0131  ;
  input \u5_data_oe_reg/NET0131  ;
  input \u5_dv_r_reg/NET0131  ;
  input \u5_ir_cnt_done_reg/P0001  ;
  input \u5_ir_cnt_reg[0]/P0001  ;
  input \u5_ir_cnt_reg[1]/P0001  ;
  input \u5_ir_cnt_reg[2]/P0001  ;
  input \u5_ir_cnt_reg[3]/P0001  ;
  input \u5_lmr_ack_reg/NET0131  ;
  input \u5_lookup_ready1_reg/NET0131  ;
  input \u5_lookup_ready2_reg/NET0131  ;
  input \u5_mc_adv_r1_reg/NET0131  ;
  input \u5_mc_adv_r_reg/NET0131  ;
  input \u5_mc_c_oe_reg/NET0131  ;
  input \u5_mc_le_reg/NET0131  ;
  input \u5_mem_ack_r_reg/NET0131  ;
  input \u5_no_wb_cycle_reg/NET0131  ;
  input \u5_oe__reg/NET0131  ;
  input \u5_pack_le0_reg/P0001  ;
  input \u5_pack_le1_reg/P0001  ;
  input \u5_resume_req_r_reg/NET0131  ;
  input \u5_rfr_ack_r_reg/NET0131  ;
  input \u5_state_reg[0]/NET0131  ;
  input \u5_state_reg[10]/NET0131  ;
  input \u5_state_reg[11]/NET0131  ;
  input \u5_state_reg[12]/NET0131  ;
  input \u5_state_reg[13]/NET0131  ;
  input \u5_state_reg[14]/NET0131  ;
  input \u5_state_reg[15]/NET0131  ;
  input \u5_state_reg[16]/NET0131  ;
  input \u5_state_reg[17]/NET0131  ;
  input \u5_state_reg[18]/NET0131  ;
  input \u5_state_reg[19]/NET0131  ;
  input \u5_state_reg[1]/NET0131  ;
  input \u5_state_reg[20]/NET0131  ;
  input \u5_state_reg[21]/NET0131  ;
  input \u5_state_reg[22]/NET0131  ;
  input \u5_state_reg[23]/NET0131  ;
  input \u5_state_reg[24]/NET0131  ;
  input \u5_state_reg[25]/NET0131  ;
  input \u5_state_reg[26]/NET0131  ;
  input \u5_state_reg[27]/NET0131  ;
  input \u5_state_reg[28]/NET0131  ;
  input \u5_state_reg[29]/NET0131  ;
  input \u5_state_reg[2]/NET0131  ;
  input \u5_state_reg[30]/NET0131  ;
  input \u5_state_reg[31]/NET0131  ;
  input \u5_state_reg[32]/NET0131  ;
  input \u5_state_reg[33]/NET0131  ;
  input \u5_state_reg[34]/NET0131  ;
  input \u5_state_reg[35]/NET0131  ;
  input \u5_state_reg[36]/NET0131  ;
  input \u5_state_reg[37]/NET0131  ;
  input \u5_state_reg[38]/NET0131  ;
  input \u5_state_reg[39]/NET0131  ;
  input \u5_state_reg[3]/NET0131  ;
  input \u5_state_reg[40]/NET0131  ;
  input \u5_state_reg[41]/NET0131  ;
  input \u5_state_reg[42]/NET0131  ;
  input \u5_state_reg[43]/NET0131  ;
  input \u5_state_reg[44]/NET0131  ;
  input \u5_state_reg[45]/NET0131  ;
  input \u5_state_reg[46]/NET0131  ;
  input \u5_state_reg[47]/NET0131  ;
  input \u5_state_reg[48]/NET0131  ;
  input \u5_state_reg[49]/NET0131  ;
  input \u5_state_reg[4]/NET0131  ;
  input \u5_state_reg[50]/NET0131  ;
  input \u5_state_reg[51]/NET0131  ;
  input \u5_state_reg[52]/NET0131  ;
  input \u5_state_reg[53]/NET0131  ;
  input \u5_state_reg[54]/NET0131  ;
  input \u5_state_reg[55]/NET0131  ;
  input \u5_state_reg[56]/NET0131  ;
  input \u5_state_reg[57]/NET0131  ;
  input \u5_state_reg[58]/NET0131  ;
  input \u5_state_reg[59]/NET0131  ;
  input \u5_state_reg[5]/NET0131  ;
  input \u5_state_reg[60]/NET0131  ;
  input \u5_state_reg[61]/NET0131  ;
  input \u5_state_reg[62]/NET0131  ;
  input \u5_state_reg[63]/NET0131  ;
  input \u5_state_reg[64]/NET0131  ;
  input \u5_state_reg[65]/NET0131  ;
  input \u5_state_reg[6]/NET0131  ;
  input \u5_state_reg[7]/NET0131  ;
  input \u5_state_reg[8]/NET0131  ;
  input \u5_state_reg[9]/NET0131  ;
  input \u5_susp_req_r_reg/NET0131  ;
  input \u5_susp_sel_r_reg/NET0131  ;
  input \u5_timer2_reg[0]/P0001  ;
  input \u5_timer2_reg[1]/P0001  ;
  input \u5_timer2_reg[2]/P0001  ;
  input \u5_timer2_reg[3]/P0001  ;
  input \u5_timer2_reg[4]/P0001  ;
  input \u5_timer2_reg[5]/P0001  ;
  input \u5_timer2_reg[6]/P0001  ;
  input \u5_timer2_reg[7]/P0001  ;
  input \u5_timer2_reg[8]/P0001  ;
  input \u5_timer_reg[0]/NET0131  ;
  input \u5_timer_reg[1]/NET0131  ;
  input \u5_timer_reg[2]/NET0131  ;
  input \u5_timer_reg[3]/NET0131  ;
  input \u5_timer_reg[4]/NET0131  ;
  input \u5_timer_reg[5]/NET0131  ;
  input \u5_timer_reg[6]/NET0131  ;
  input \u5_timer_reg[7]/NET0131  ;
  input \u5_tmr2_done_reg/NET0131  ;
  input \u5_tmr_done_reg/NET0131  ;
  input \u5_wb_cycle_reg/NET0131  ;
  input \u5_wb_stb_first_reg/NET0131  ;
  input \u5_wb_wait_r_reg/P0001  ;
  input \u5_wb_write_go_r_reg/NET0131  ;
  input \u5_wr_cycle_reg/NET0131  ;
  input \u6_read_go_r1_reg/NET0131  ;
  input \u6_read_go_r_reg/NET0131  ;
  input \u6_rmw_en_reg/NET0131  ;
  input \u6_rmw_r_reg/NET0131  ;
  input \u6_wb_first_r_reg/NET0131  ;
  input \u6_wr_hold_reg/NET0131  ;
  input \u6_write_go_r1_reg/NET0131  ;
  input \u6_write_go_r_reg/NET0131  ;
  input \u7_mc_ack_r_reg/NET0131  ;
  input \u7_mc_br_r_reg/P0001  ;
  input \u7_mc_data_ir_reg[0]/P0001  ;
  input \u7_mc_data_ir_reg[10]/P0001  ;
  input \u7_mc_data_ir_reg[11]/P0001  ;
  input \u7_mc_data_ir_reg[12]/P0001  ;
  input \u7_mc_data_ir_reg[13]/P0001  ;
  input \u7_mc_data_ir_reg[14]/P0001  ;
  input \u7_mc_data_ir_reg[15]/P0001  ;
  input \u7_mc_data_ir_reg[16]/P0001  ;
  input \u7_mc_data_ir_reg[17]/P0001  ;
  input \u7_mc_data_ir_reg[18]/P0001  ;
  input \u7_mc_data_ir_reg[19]/P0001  ;
  input \u7_mc_data_ir_reg[1]/P0001  ;
  input \u7_mc_data_ir_reg[20]/P0001  ;
  input \u7_mc_data_ir_reg[21]/P0001  ;
  input \u7_mc_data_ir_reg[22]/P0001  ;
  input \u7_mc_data_ir_reg[23]/P0001  ;
  input \u7_mc_data_ir_reg[24]/P0001  ;
  input \u7_mc_data_ir_reg[25]/P0001  ;
  input \u7_mc_data_ir_reg[26]/P0001  ;
  input \u7_mc_data_ir_reg[27]/P0001  ;
  input \u7_mc_data_ir_reg[28]/P0001  ;
  input \u7_mc_data_ir_reg[29]/P0001  ;
  input \u7_mc_data_ir_reg[2]/P0001  ;
  input \u7_mc_data_ir_reg[30]/P0001  ;
  input \u7_mc_data_ir_reg[31]/P0001  ;
  input \u7_mc_data_ir_reg[3]/P0001  ;
  input \u7_mc_data_ir_reg[4]/P0001  ;
  input \u7_mc_data_ir_reg[5]/P0001  ;
  input \u7_mc_data_ir_reg[6]/P0001  ;
  input \u7_mc_data_ir_reg[7]/P0001  ;
  input \u7_mc_data_ir_reg[8]/P0001  ;
  input \u7_mc_data_ir_reg[9]/P0001  ;
  input \u7_mc_dqm_r2_reg[0]/P0001  ;
  input \u7_mc_dqm_r2_reg[1]/P0001  ;
  input \u7_mc_dqm_r2_reg[2]/P0001  ;
  input \u7_mc_dqm_r2_reg[3]/P0001  ;
  input \u7_mc_dqm_r_reg[0]/P0001  ;
  input \u7_mc_dqm_r_reg[1]/P0001  ;
  input \u7_mc_dqm_r_reg[2]/P0001  ;
  input \u7_mc_dqm_r_reg[3]/P0001  ;
  input wb_ack_o_pad ;
  input \wb_addr_i[0]_pad  ;
  input \wb_addr_i[10]_pad  ;
  input \wb_addr_i[11]_pad  ;
  input \wb_addr_i[12]_pad  ;
  input \wb_addr_i[13]_pad  ;
  input \wb_addr_i[14]_pad  ;
  input \wb_addr_i[15]_pad  ;
  input \wb_addr_i[16]_pad  ;
  input \wb_addr_i[17]_pad  ;
  input \wb_addr_i[18]_pad  ;
  input \wb_addr_i[19]_pad  ;
  input \wb_addr_i[1]_pad  ;
  input \wb_addr_i[20]_pad  ;
  input \wb_addr_i[21]_pad  ;
  input \wb_addr_i[22]_pad  ;
  input \wb_addr_i[23]_pad  ;
  input \wb_addr_i[24]_pad  ;
  input \wb_addr_i[25]_pad  ;
  input \wb_addr_i[26]_pad  ;
  input \wb_addr_i[27]_pad  ;
  input \wb_addr_i[28]_pad  ;
  input \wb_addr_i[29]_pad  ;
  input \wb_addr_i[2]_pad  ;
  input \wb_addr_i[30]_pad  ;
  input \wb_addr_i[31]_pad  ;
  input \wb_addr_i[3]_pad  ;
  input \wb_addr_i[4]_pad  ;
  input \wb_addr_i[5]_pad  ;
  input \wb_addr_i[6]_pad  ;
  input \wb_addr_i[7]_pad  ;
  input \wb_addr_i[8]_pad  ;
  input \wb_addr_i[9]_pad  ;
  input wb_cyc_i_pad ;
  input \wb_data_i[0]_pad  ;
  input \wb_data_i[10]_pad  ;
  input \wb_data_i[11]_pad  ;
  input \wb_data_i[12]_pad  ;
  input \wb_data_i[13]_pad  ;
  input \wb_data_i[14]_pad  ;
  input \wb_data_i[15]_pad  ;
  input \wb_data_i[16]_pad  ;
  input \wb_data_i[17]_pad  ;
  input \wb_data_i[18]_pad  ;
  input \wb_data_i[19]_pad  ;
  input \wb_data_i[1]_pad  ;
  input \wb_data_i[20]_pad  ;
  input \wb_data_i[21]_pad  ;
  input \wb_data_i[22]_pad  ;
  input \wb_data_i[23]_pad  ;
  input \wb_data_i[24]_pad  ;
  input \wb_data_i[25]_pad  ;
  input \wb_data_i[26]_pad  ;
  input \wb_data_i[27]_pad  ;
  input \wb_data_i[28]_pad  ;
  input \wb_data_i[29]_pad  ;
  input \wb_data_i[2]_pad  ;
  input \wb_data_i[30]_pad  ;
  input \wb_data_i[31]_pad  ;
  input \wb_data_i[3]_pad  ;
  input \wb_data_i[4]_pad  ;
  input \wb_data_i[5]_pad  ;
  input \wb_data_i[6]_pad  ;
  input \wb_data_i[7]_pad  ;
  input \wb_data_i[8]_pad  ;
  input \wb_data_i[9]_pad  ;
  input wb_err_o_pad ;
  input \wb_sel_i[0]_pad  ;
  input \wb_sel_i[1]_pad  ;
  input \wb_sel_i[2]_pad  ;
  input \wb_sel_i[3]_pad  ;
  input wb_stb_i_pad ;
  input wb_we_i_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g22/_0_  ;
  output \g23/_0_  ;
  output \g25_dup61718/_2_  ;
  output \g43466/_0_  ;
  output \g43467/_0_  ;
  output \g43468/_0_  ;
  output \g43469/_0_  ;
  output \g43470/_0_  ;
  output \g43471/_0_  ;
  output \g43472/_0_  ;
  output \g43473/_0_  ;
  output \g43474/_0_  ;
  output \g43475/_0_  ;
  output \g43476/_0_  ;
  output \g43477/_0_  ;
  output \g43478/_0_  ;
  output \g43512/_0_  ;
  output \g43513/_0_  ;
  output \g43544/_3_  ;
  output \g43545/_0_  ;
  output \g43554/_0_  ;
  output \g43555/_0_  ;
  output \g43557/_0_  ;
  output \g43558/_0_  ;
  output \g43571/_2_  ;
  output \g43632/_0_  ;
  output \g43633/_0_  ;
  output \g43635/_0_  ;
  output \g43636/_0_  ;
  output \g43637/_0_  ;
  output \g43638/_0_  ;
  output \g43639/_0_  ;
  output \g43640/_0_  ;
  output \g43642/_0_  ;
  output \g43662/_0_  ;
  output \g43663/_0_  ;
  output \g43664/_0_  ;
  output \g43665/_0_  ;
  output \g43668/_0_  ;
  output \g43670/_0_  ;
  output \g43671/_0_  ;
  output \g43673/_0_  ;
  output \g43674/_0_  ;
  output \g43692/_0_  ;
  output \g43695/_0_  ;
  output \g43696/_0_  ;
  output \g43697/_0_  ;
  output \g43698/_0_  ;
  output \g43700/_0_  ;
  output \g43701/_0_  ;
  output \g43703/_0_  ;
  output \g43705/_0_  ;
  output \g43707/_0_  ;
  output \g43708/_0_  ;
  output \g43710/_0_  ;
  output \g43717/_0_  ;
  output \g43719/_0_  ;
  output \g43720/_0_  ;
  output \g43721/_0_  ;
  output \g43722/_1_  ;
  output \g43723/_0_  ;
  output \g43725/_0_  ;
  output \g43729/_0_  ;
  output \g43731/_0_  ;
  output \g43734/_0_  ;
  output \g43735/_0_  ;
  output \g43737/_0_  ;
  output \g43744/_0_  ;
  output \g43747/_0_  ;
  output \g43760/_2_  ;
  output \g43770/_1_  ;
  output \g43775/_2_  ;
  output \g43780/_2_  ;
  output \g43786/_0_  ;
  output \g43787/_1_  ;
  output \g43847/_0_  ;
  output \g43848/_1_  ;
  output \g43858/_1_  ;
  output \g43891/_3_  ;
  output \g43895/_0_  ;
  output \g43934/_0_  ;
  output \g43936/_3_  ;
  output \g43954/_3_  ;
  output \g43961/_0_  ;
  output \g44016/_1_  ;
  output \g44067/_0_  ;
  output \g44094/_0_  ;
  output \g44096/_0_  ;
  output \g44104/_0_  ;
  output \g44122/_0_  ;
  output \g44172/_0_  ;
  output \g44209/_0_  ;
  output \g44219/_0_  ;
  output \g44220/_0_  ;
  output \g44222/_0_  ;
  output \g44223/_0_  ;
  output \g44241/_2_  ;
  output \g44252/_0_  ;
  output \g44253/_0_  ;
  output \g44255/_2_  ;
  output \g44263/_2_  ;
  output \g44470/_0_  ;
  output \g44538/_0_  ;
  output \g44539/_0_  ;
  output \g44540/_0_  ;
  output \g44541/_0_  ;
  output \g44542/_0_  ;
  output \g44543/_0_  ;
  output \g44544/_0_  ;
  output \g44545/_0_  ;
  output \g44546/_0_  ;
  output \g44547/_0_  ;
  output \g44548/_0_  ;
  output \g44549/_0_  ;
  output \g44550/_0_  ;
  output \g44551/_0_  ;
  output \g44552/_0_  ;
  output \g44553/_0_  ;
  output \g44554/_0_  ;
  output \g44555/_0_  ;
  output \g44556/_0_  ;
  output \g44557/_0_  ;
  output \g44558/_0_  ;
  output \g44559/_0_  ;
  output \g44560/_0_  ;
  output \g44561/_0_  ;
  output \g44562/_0_  ;
  output \g44563/_0_  ;
  output \g44564/_0_  ;
  output \g44565/_0_  ;
  output \g44566/_0_  ;
  output \g44567/_0_  ;
  output \g44568/_0_  ;
  output \g44569/_0_  ;
  output \g44570/_0_  ;
  output \g44571/_0_  ;
  output \g44572/_0_  ;
  output \g44573/_0_  ;
  output \g44574/_0_  ;
  output \g44575/_0_  ;
  output \g44576/_0_  ;
  output \g44577/_0_  ;
  output \g44578/_0_  ;
  output \g44579/_0_  ;
  output \g44580/_0_  ;
  output \g44581/_0_  ;
  output \g44582/_0_  ;
  output \g44583/_0_  ;
  output \g44584/_0_  ;
  output \g44585/_0_  ;
  output \g44586/_0_  ;
  output \g44588/_0_  ;
  output \g44589/_0_  ;
  output \g44590/_0_  ;
  output \g44591/_0_  ;
  output \g44592/_0_  ;
  output \g44593/_0_  ;
  output \g44594/_0_  ;
  output \g44595/_0_  ;
  output \g44596/_0_  ;
  output \g44636/_2_  ;
  output \g44646/_0_  ;
  output \g44647/_0_  ;
  output \g44648/_0_  ;
  output \g44649/_0_  ;
  output \g44650/_0_  ;
  output \g44651/_0_  ;
  output \g44652/_0_  ;
  output \g44653/_0_  ;
  output \g44654/_0_  ;
  output \g44655/_0_  ;
  output \g44656/_0_  ;
  output \g44657/_0_  ;
  output \g44665/_0_  ;
  output \g44666/_0_  ;
  output \g44667/_0_  ;
  output \g44668/_0_  ;
  output \g44752/_0_  ;
  output \g44753/_0_  ;
  output \g44873/_0_  ;
  output \g44939/_0_  ;
  output \g44942/_0_  ;
  output \g44945/_0_  ;
  output \g45023/_2_  ;
  output \g45090/_0_  ;
  output \g45141/_0_  ;
  output \g45147/_3_  ;
  output \g45155/_0_  ;
  output \g45190/_0_  ;
  output \g45195/_2_  ;
  output \g45199/_2_  ;
  output \g45201/_2_  ;
  output \g45324/_0_  ;
  output \g45334/_2_  ;
  output \g45336/_0_  ;
  output \g45388/_0_  ;
  output \g45391/_0_  ;
  output \g45413/_2_  ;
  output \g45530/_0_  ;
  output \g45532/_0_  ;
  output \g45533/_0_  ;
  output \g45534/_0_  ;
  output \g45739/_2_  ;
  output \g45743/_2_  ;
  output \g45767/_0_  ;
  output \g45782/_0_  ;
  output \g45830/_3_  ;
  output \g45834/_3_  ;
  output \g45835/_3_  ;
  output \g45836/_3_  ;
  output \g45837/_3_  ;
  output \g45839/_3_  ;
  output \g45840/_3_  ;
  output \g45841/_3_  ;
  output \g45842/_3_  ;
  output \g45843/_3_  ;
  output \g45844/_3_  ;
  output \g45845/_3_  ;
  output \g46191/_0_  ;
  output \g46193/_3_  ;
  output \g46256/_3_  ;
  output \g46257/_3_  ;
  output \g46258/_3_  ;
  output \g46259/_3_  ;
  output \g46260/_3_  ;
  output \g46261/_3_  ;
  output \g46262/_3_  ;
  output \g46263/_3_  ;
  output \g46278/_0_  ;
  output \g46292/_0_  ;
  output \g46293/_0_  ;
  output \g46312/_0_  ;
  output \g46367/_2_  ;
  output \g46370/_2_  ;
  output \g46380/_2_  ;
  output \g46386/_2_  ;
  output \g46388/_2_  ;
  output \g46392/_2_  ;
  output \g46395/_2_  ;
  output \g46399/_2_  ;
  output \g46420/_0_  ;
  output \g46446/_0_  ;
  output \g46493/_0_  ;
  output \g46510/_0_  ;
  output \g46669/_2_  ;
  output \g46691/_0_  ;
  output \g46708/_0_  ;
  output \g46721/_00_  ;
  output \g46776/_0_  ;
  output \g46777/_0_  ;
  output \g46778/_0_  ;
  output \g46779/_0_  ;
  output \g46780/_0_  ;
  output \g46782/_0_  ;
  output \g46784/_0_  ;
  output \g46932/_0_  ;
  output \g47112/_0_  ;
  output \g47124/_0_  ;
  output \g47265/_0_  ;
  output \g47270/_0_  ;
  output \g47275/_0_  ;
  output \g47300/_1_  ;
  output \g47305/_1_  ;
  output \g47338/_0_  ;
  output \g47339/_0_  ;
  output \g47352/_0_  ;
  output \g47699/_3_  ;
  output \g47711/_0_  ;
  output \g47719/_3_  ;
  output \g47721/_3_  ;
  output \g47723/_3_  ;
  output \g47853/_0_  ;
  output \g48094/_0_  ;
  output \g48095/_0_  ;
  output \g48177/_2_  ;
  output \g48194/_0_  ;
  output \g48369/_2_  ;
  output \g48371/_2_  ;
  output \g48373/_2_  ;
  output \g48375/_2_  ;
  output \g48377/_2_  ;
  output \g48379/_2_  ;
  output \g48381/_2_  ;
  output \g48383/_2_  ;
  output \g48385/_2_  ;
  output \g48535/_0_  ;
  output \g48569/_0_  ;
  output \g48570/_0_  ;
  output \g48571/_0_  ;
  output \g48836/_0_  ;
  output \g48843/_0_  ;
  output \g49187/_3_  ;
  output \g49375/_2_  ;
  output \g49633/_0_  ;
  output \g49788/_1_  ;
  output \g49800/_1_  ;
  output \g49802/_1_  ;
  output \g49806/_1_  ;
  output \g49853/_1_  ;
  output \g49883/_0_  ;
  output \g49884/_0_  ;
  output \g49885/_0_  ;
  output \g49886/_0_  ;
  output \g49976/_1_  ;
  output \g50038/_0_  ;
  output \g50082/_0_  ;
  output \g50083/_0_  ;
  output \g50167/_3_  ;
  output \g50168/_3_  ;
  output \g50169/_3_  ;
  output \g50170/_3_  ;
  output \g50171/_3_  ;
  output \g50177/_0_  ;
  output \g50190/_0_  ;
  output \g50236/_0_  ;
  output \g50251/_3_  ;
  output \g50256/_0_  ;
  output \g50318/_3_  ;
  output \g50319/_3_  ;
  output \g50350/_3_  ;
  output \g50351/_3_  ;
  output \g50352/_3_  ;
  output \g50353/_3_  ;
  output \g50354/_3_  ;
  output \g50355/_3_  ;
  output \g50361/_2_  ;
  output \g50366/_0_  ;
  output \g50393/_0_  ;
  output \g50552/_1_  ;
  output \g51108/_0_  ;
  output \g51160/_0_  ;
  output \g51290/_1_  ;
  output \g51327/_3_  ;
  output \g51328/_3_  ;
  output \g51329/_3_  ;
  output \g51330/_3_  ;
  output \g51331/_3_  ;
  output \g51332/_3_  ;
  output \g51333/_3_  ;
  output \g51334/_3_  ;
  output \g51339/_3_  ;
  output \g51340/_3_  ;
  output \g51341/_3_  ;
  output \g51342/_3_  ;
  output \g51343/_3_  ;
  output \g51346/_0_  ;
  output \g51347/_0_  ;
  output \g51348/_0_  ;
  output \g51381/_3_  ;
  output \g51382/_3_  ;
  output \g51383/_3_  ;
  output \g51386/_3_  ;
  output \g51387/_3_  ;
  output \g51405/_3_  ;
  output \g51410/_3_  ;
  output \g51883/_0_  ;
  output \g51916/_0_  ;
  output \g51947/_0_  ;
  output \g51948/_0_  ;
  output \g51949/_0_  ;
  output \g51950/_0_  ;
  output \g51951/_0_  ;
  output \g51952/_0_  ;
  output \g51953/_0_  ;
  output \g51954/_0_  ;
  output \g51955/_0_  ;
  output \g51956/_0_  ;
  output \g51957/_0_  ;
  output \g51958/_0_  ;
  output \g51959/_0_  ;
  output \g51960/_0_  ;
  output \g51961/_0_  ;
  output \g51962/_0_  ;
  output \g51963/_0_  ;
  output \g51964/_0_  ;
  output \g51965/_0_  ;
  output \g51967/_0_  ;
  output \g51968/_0_  ;
  output \g51969/_0_  ;
  output \g51970/_0_  ;
  output \g51971/_0_  ;
  output \g51972/_0_  ;
  output \g51973/_0_  ;
  output \g51974/_0_  ;
  output \g51975/_0_  ;
  output \g51976/_0_  ;
  output \g51977/_0_  ;
  output \g51978/_0_  ;
  output \g51979/_0_  ;
  output \g51980/_0_  ;
  output \g51981/_0_  ;
  output \g51982/_0_  ;
  output \g51983/_0_  ;
  output \g51984/_0_  ;
  output \g51985/_0_  ;
  output \g51986/_0_  ;
  output \g51987/_0_  ;
  output \g51988/_0_  ;
  output \g51989/_0_  ;
  output \g51990/_0_  ;
  output \g51991/_0_  ;
  output \g51992/_0_  ;
  output \g51993/_0_  ;
  output \g51994/_0_  ;
  output \g51995/_0_  ;
  output \g51996/_0_  ;
  output \g51997/_0_  ;
  output \g51998/_0_  ;
  output \g51999/_0_  ;
  output \g52000/_0_  ;
  output \g52001/_0_  ;
  output \g52002/_0_  ;
  output \g52003/_0_  ;
  output \g52004/_0_  ;
  output \g52005/_0_  ;
  output \g52006/_0_  ;
  output \g52007/_0_  ;
  output \g52008/_0_  ;
  output \g52009/_0_  ;
  output \g52010/_0_  ;
  output \g52011/_0_  ;
  output \g52012/_0_  ;
  output \g52013/_0_  ;
  output \g52014/_0_  ;
  output \g52015/_0_  ;
  output \g52016/_0_  ;
  output \g52017/_0_  ;
  output \g52018/_0_  ;
  output \g52019/_0_  ;
  output \g52020/_0_  ;
  output \g52021/_0_  ;
  output \g52022/_0_  ;
  output \g52023/_0_  ;
  output \g52024/_0_  ;
  output \g52025/_0_  ;
  output \g52026/_0_  ;
  output \g52027/_0_  ;
  output \g52028/_0_  ;
  output \g52029/_0_  ;
  output \g52030/_0_  ;
  output \g52031/_0_  ;
  output \g52032/_0_  ;
  output \g52033/_0_  ;
  output \g52034/_0_  ;
  output \g52035/_0_  ;
  output \g52036/_0_  ;
  output \g52037/_0_  ;
  output \g52038/_0_  ;
  output \g52039/_0_  ;
  output \g52040/_0_  ;
  output \g52041/_0_  ;
  output \g52042/_0_  ;
  output \g52043/_0_  ;
  output \g52044/_0_  ;
  output \g52045/_0_  ;
  output \g52046/_0_  ;
  output \g52047/_0_  ;
  output \g52049/_0_  ;
  output \g52050/_0_  ;
  output \g52051/_0_  ;
  output \g52052/_0_  ;
  output \g52053/_0_  ;
  output \g52054/_0_  ;
  output \g52055/_0_  ;
  output \g52056/_0_  ;
  output \g52057/_0_  ;
  output \g52058/_0_  ;
  output \g52061/_0_  ;
  output \g52065/_0_  ;
  output \g52066/_0_  ;
  output \g52067/_0_  ;
  output \g52068/_0_  ;
  output \g52069/_0_  ;
  output \g52070/_0_  ;
  output \g52071/_0_  ;
  output \g52073/_0_  ;
  output \g52074/_0_  ;
  output \g52075/_0_  ;
  output \g52082/_0_  ;
  output \g52083/_0_  ;
  output \g52158/_0_  ;
  output \g52201/_0_  ;
  output \g52202/_0_  ;
  output \g52346/_0_  ;
  output \g52351/_0_  ;
  output \g52390/_0_  ;
  output \g52847/_0_  ;
  output \g52854/_0_  ;
  output \g52968/_0_  ;
  output \g52969/_0_  ;
  output \g52970/_0_  ;
  output \g52971/_0_  ;
  output \g52984/_0_  ;
  output \g52994/_0_  ;
  output \g53019/_0_  ;
  output \g53030/_0_  ;
  output \g53094/_1_  ;
  output \g53106/_0_  ;
  output \g53150/_0_  ;
  output \g53256/_0_  ;
  output \g53297/_0_  ;
  output \g53345/_0_  ;
  output \g53359/_0_  ;
  output \g53375/_0_  ;
  output \g53474/_1__syn_2  ;
  output \g53475/_2_  ;
  output \g53593/_0_  ;
  output \g53643/_1_  ;
  output \g53655/_0_  ;
  output \g53710/_0_  ;
  output \g53786/_0_  ;
  output \g53837/_0_  ;
  output \g53888/_1_  ;
  output \g53909/_0_  ;
  output \g54253/_2_  ;
  output \g54394/_3_  ;
  output \g54413/_0_  ;
  output \g55420/_0_  ;
  output \g55587/_0_  ;
  output \g55852/_0_  ;
  output \g57020/_0_  ;
  output \g59450/_0_  ;
  output \g59488/_2_  ;
  output \g59752/_0_  ;
  output \g59786/_0_  ;
  output \g59854/_0_  ;
  output \g59878/_0_  ;
  output \g59902/_0_  ;
  output \g59924/_0_  ;
  output \g59947/_0_  ;
  output \g59972/_0_  ;
  output \g59996/_0_  ;
  output \g60017/_0_  ;
  output \g60040/_0_  ;
  output \g60064/_0_  ;
  output \g60095/_0_  ;
  output \g60119/_0_  ;
  output \g60145/_1_  ;
  output \g60165/_0_  ;
  output \g60407/_2_  ;
  output \g60408/_0_  ;
  output \g60613/_2_  ;
  output \g60649/_0_  ;
  output \g60771/_0_  ;
  output \g60908/_1_  ;
  output \g60911/_0_  ;
  output \g60977/_0_  ;
  output \g61/_0_  ;
  output \g61002/_0_  ;
  output \g61308/_0_  ;
  output \g61312/_1_  ;
  output \g61314/_0_  ;
  output \g61319/_1_  ;
  output \g61342/_1_  ;
  output \g61360/_0_  ;
  output \g61377/_0_  ;
  output \g61423/_1_  ;
  output \g61426/_0_  ;
  output \g61479/_1_  ;
  output \g61523/_1_  ;
  output \g61558/_1_  ;
  output \g61652/_0_  ;
  output \g61866/_0_  ;
  output \g61868/_1_  ;
  output \g61887/_0_  ;
  output \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3  ;
  output \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3  ;
  output \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3  ;
  output \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3  ;
  output \u7_mc_we__reg/_05_  ;
  wire n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 ;
  assign n959 = ~\u5_state_reg[38]/NET0131  & ~\u5_state_reg[39]/NET0131  ;
  assign n960 = ~\u5_state_reg[40]/NET0131  & ~\u5_state_reg[41]/NET0131  ;
  assign n961 = n959 & n960 ;
  assign n962 = ~\u5_state_reg[43]/NET0131  & ~\u5_state_reg[45]/NET0131  ;
  assign n963 = ~\u5_state_reg[42]/NET0131  & ~\u5_state_reg[44]/NET0131  ;
  assign n964 = n962 & n963 ;
  assign n965 = n961 & n964 ;
  assign n966 = ~\u5_state_reg[34]/NET0131  & ~\u5_state_reg[35]/NET0131  ;
  assign n967 = ~\u5_state_reg[36]/NET0131  & ~\u5_state_reg[37]/NET0131  ;
  assign n968 = n966 & n967 ;
  assign n969 = ~\u5_state_reg[47]/NET0131  & ~\u5_state_reg[48]/NET0131  ;
  assign n970 = ~\u5_state_reg[46]/NET0131  & ~\u5_state_reg[49]/NET0131  ;
  assign n971 = n969 & n970 ;
  assign n972 = n968 & n971 ;
  assign n973 = n965 & n972 ;
  assign n974 = ~\u5_state_reg[28]/NET0131  & ~\u5_state_reg[29]/NET0131  ;
  assign n975 = ~\u5_state_reg[26]/NET0131  & ~\u5_state_reg[27]/NET0131  ;
  assign n976 = n974 & n975 ;
  assign n977 = ~\u5_state_reg[18]/NET0131  & ~\u5_state_reg[19]/NET0131  ;
  assign n978 = ~\u5_state_reg[20]/NET0131  & ~\u5_state_reg[21]/NET0131  ;
  assign n979 = n977 & n978 ;
  assign n980 = n976 & n979 ;
  assign n981 = ~\u5_state_reg[23]/NET0131  & ~\u5_state_reg[25]/NET0131  ;
  assign n982 = ~\u5_state_reg[22]/NET0131  & ~\u5_state_reg[24]/NET0131  ;
  assign n983 = n981 & n982 ;
  assign n984 = ~\u5_state_reg[32]/NET0131  & ~\u5_state_reg[33]/NET0131  ;
  assign n985 = ~\u5_state_reg[30]/NET0131  & ~\u5_state_reg[31]/NET0131  ;
  assign n986 = n984 & n985 ;
  assign n987 = n983 & n986 ;
  assign n988 = n980 & n987 ;
  assign n989 = n973 & n988 ;
  assign n990 = ~\u5_state_reg[15]/NET0131  & ~\u5_state_reg[16]/NET0131  ;
  assign n991 = ~\u5_state_reg[14]/NET0131  & ~\u5_state_reg[17]/NET0131  ;
  assign n992 = n990 & n991 ;
  assign n993 = ~\u5_state_reg[6]/NET0131  & ~\u5_state_reg[8]/NET0131  ;
  assign n994 = ~\u5_state_reg[7]/NET0131  & ~\u5_state_reg[9]/NET0131  ;
  assign n995 = n993 & n994 ;
  assign n996 = n992 & n995 ;
  assign n997 = ~\u5_state_reg[12]/NET0131  & ~\u5_state_reg[13]/NET0131  ;
  assign n998 = ~\u5_state_reg[10]/NET0131  & ~\u5_state_reg[11]/NET0131  ;
  assign n999 = n997 & n998 ;
  assign n1000 = ~\u5_state_reg[2]/NET0131  & ~\u5_state_reg[4]/NET0131  ;
  assign n1001 = ~\u5_state_reg[3]/NET0131  & ~\u5_state_reg[5]/NET0131  ;
  assign n1002 = n1000 & n1001 ;
  assign n1003 = n999 & n1002 ;
  assign n1004 = n996 & n1003 ;
  assign n1005 = ~\u5_state_reg[63]/NET0131  & ~\u5_state_reg[64]/NET0131  ;
  assign n1006 = ~\u5_state_reg[62]/NET0131  & ~\u5_state_reg[65]/NET0131  ;
  assign n1007 = n1005 & n1006 ;
  assign n1008 = ~\u5_state_reg[60]/NET0131  & ~\u5_state_reg[61]/NET0131  ;
  assign n1009 = ~\u5_state_reg[58]/NET0131  & ~\u5_state_reg[59]/NET0131  ;
  assign n1010 = n1008 & n1009 ;
  assign n1011 = n1007 & n1010 ;
  assign n1012 = ~\u5_state_reg[0]/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n1013 = n1011 & n1012 ;
  assign n1014 = n1004 & n1013 ;
  assign n1015 = n989 & n1014 ;
  assign n1016 = ~\u5_state_reg[52]/NET0131  & ~\u5_state_reg[53]/NET0131  ;
  assign n1017 = ~\u5_state_reg[50]/NET0131  & ~\u5_state_reg[51]/NET0131  ;
  assign n1018 = n1016 & n1017 ;
  assign n1019 = ~\u5_state_reg[56]/NET0131  & n1018 ;
  assign n1020 = \u5_state_reg[54]/NET0131  & ~\u5_state_reg[55]/NET0131  ;
  assign n1021 = ~\u5_state_reg[57]/NET0131  & n1020 ;
  assign n1022 = n1019 & n1021 ;
  assign n1023 = n1015 & n1022 ;
  assign n1024 = ~\u5_dv_r_reg/NET0131  & \u5_mc_adv_r_reg/NET0131  ;
  assign n1025 = n1023 & n1024 ;
  assign n1026 = ~\u5_state_reg[54]/NET0131  & ~\u5_state_reg[55]/NET0131  ;
  assign n1027 = ~\u5_state_reg[56]/NET0131  & ~\u5_state_reg[57]/NET0131  ;
  assign n1028 = n1026 & n1027 ;
  assign n1029 = n1018 & n1028 ;
  assign n1030 = n996 & n1029 ;
  assign n1031 = n1013 & n1030 ;
  assign n1032 = n989 & n1031 ;
  assign n1033 = ~\u5_state_reg[3]/NET0131  & n1000 ;
  assign n1034 = ~\u5_state_reg[5]/NET0131  & n997 ;
  assign n1035 = n1033 & n1034 ;
  assign n1036 = n1032 & n1035 ;
  assign n1037 = ~\u5_state_reg[10]/NET0131  & \u5_state_reg[11]/NET0131  ;
  assign n1038 = ~\u5_cnt_reg/NET0131  & \u5_wb_cycle_reg/NET0131  ;
  assign n1039 = \u5_burst_act_rd_reg/P0001  & \u5_cke_o_del_reg/P0001  ;
  assign n1040 = n1038 & n1039 ;
  assign n1041 = n1037 & n1040 ;
  assign n1042 = n1036 & n1041 ;
  assign n1043 = ~n1025 & ~n1042 ;
  assign n1044 = \u3_u0_wr_adr_reg[3]/NET0131  & ~n1043 ;
  assign n1045 = wb_cyc_i_pad & wb_stb_i_pad ;
  assign n1046 = wb_we_i_pad & n1045 ;
  assign n1047 = \u6_rmw_en_reg/NET0131  & ~\u6_wr_hold_reg/NET0131  ;
  assign n1048 = n1046 & n1047 ;
  assign n1049 = \u5_state_reg[6]/NET0131  & ~\u5_wb_wait_r_reg/P0001  ;
  assign n1050 = n971 & n1010 ;
  assign n1051 = n1029 & n1050 ;
  assign n1052 = n965 & n1051 ;
  assign n1053 = ~\u5_state_reg[8]/NET0131  & ~\u5_state_reg[9]/NET0131  ;
  assign n1054 = n998 & n1053 ;
  assign n1055 = n990 & n997 ;
  assign n1056 = n1054 & n1055 ;
  assign n1057 = ~\u5_state_reg[5]/NET0131  & ~\u5_state_reg[6]/NET0131  ;
  assign n1058 = \u5_state_reg[7]/NET0131  & n991 ;
  assign n1059 = n1057 & n1058 ;
  assign n1060 = n980 & n1059 ;
  assign n1061 = n1056 & n1060 ;
  assign n1062 = ~\u5_state_reg[32]/NET0131  & n985 ;
  assign n1063 = ~\u5_state_reg[1]/NET0131  & ~\u5_state_reg[3]/NET0131  ;
  assign n1064 = n1000 & n1063 ;
  assign n1065 = n1062 & n1064 ;
  assign n1066 = n983 & n1007 ;
  assign n1067 = ~\u5_state_reg[33]/NET0131  & n966 ;
  assign n1068 = ~\u5_state_reg[0]/NET0131  & ~\u5_state_reg[36]/NET0131  ;
  assign n1069 = ~\u5_state_reg[37]/NET0131  & n1068 ;
  assign n1070 = n1067 & n1069 ;
  assign n1071 = n1066 & n1070 ;
  assign n1072 = n1065 & n1071 ;
  assign n1073 = n1061 & n1072 ;
  assign n1074 = n1052 & n1073 ;
  assign n1075 = ~n1049 & ~n1074 ;
  assign n1076 = n1013 & n1029 ;
  assign n1077 = n973 & n976 ;
  assign n1078 = n1076 & n1077 ;
  assign n1079 = n979 & n983 ;
  assign n1080 = n1004 & n1079 ;
  assign n1081 = ~\u5_state_reg[32]/NET0131  & \u5_state_reg[33]/NET0131  ;
  assign n1082 = n985 & n1081 ;
  assign n1083 = n1080 & n1082 ;
  assign n1084 = n1078 & n1083 ;
  assign n1085 = n988 & n1004 ;
  assign n1086 = n965 & n1029 ;
  assign n1087 = n1013 & n1086 ;
  assign n1088 = n1085 & n1087 ;
  assign n1089 = \u5_state_reg[34]/NET0131  & ~\u5_state_reg[35]/NET0131  ;
  assign n1090 = n967 & n1089 ;
  assign n1091 = n971 & n1090 ;
  assign n1092 = n1088 & n1091 ;
  assign n1093 = ~n1084 & ~n1092 ;
  assign n1094 = n1036 & n1037 ;
  assign n1095 = n979 & n986 ;
  assign n1096 = n1004 & n1095 ;
  assign n1097 = \u5_state_reg[23]/NET0131  & ~\u5_state_reg[25]/NET0131  ;
  assign n1098 = n982 & n1097 ;
  assign n1099 = n1096 & n1098 ;
  assign n1100 = n1078 & n1099 ;
  assign n1101 = \u5_state_reg[30]/NET0131  & ~\u5_state_reg[31]/NET0131  ;
  assign n1102 = n984 & n1101 ;
  assign n1103 = n1080 & n1102 ;
  assign n1104 = n1078 & n1103 ;
  assign n1105 = ~n1100 & ~n1104 ;
  assign n1106 = ~n1094 & n1105 ;
  assign n1107 = n1093 & n1106 ;
  assign n1108 = ~\u5_state_reg[52]/NET0131  & \u5_state_reg[53]/NET0131  ;
  assign n1109 = n1017 & n1028 ;
  assign n1110 = n1108 & n1109 ;
  assign n1111 = n1015 & n1110 ;
  assign n1112 = ~n1023 & ~n1111 ;
  assign n1113 = n1012 & n1029 ;
  assign n1114 = n1004 & n1113 ;
  assign n1115 = n989 & n1114 ;
  assign n1116 = ~\u5_state_reg[62]/NET0131  & \u5_state_reg[65]/NET0131  ;
  assign n1117 = n1005 & n1116 ;
  assign n1118 = n1010 & n1117 ;
  assign n1119 = n1115 & n1118 ;
  assign n1120 = n972 & n1029 ;
  assign n1121 = n1013 & n1120 ;
  assign n1122 = n1085 & n1121 ;
  assign n1123 = \u5_state_reg[40]/NET0131  & ~\u5_state_reg[41]/NET0131  ;
  assign n1124 = n959 & n1123 ;
  assign n1125 = n964 & n1124 ;
  assign n1126 = n1122 & n1125 ;
  assign n1127 = ~n1119 & ~n1126 ;
  assign n1128 = n1112 & n1127 ;
  assign n1129 = n973 & n979 ;
  assign n1130 = n1076 & n1129 ;
  assign n1131 = n987 & n1004 ;
  assign n1132 = ~\u5_state_reg[28]/NET0131  & \u5_state_reg[29]/NET0131  ;
  assign n1133 = n975 & n1132 ;
  assign n1134 = n1131 & n1133 ;
  assign n1135 = n1130 & n1134 ;
  assign n1136 = n1128 & ~n1135 ;
  assign n1137 = n1107 & n1136 ;
  assign n1138 = \u5_state_reg[10]/NET0131  & ~\u5_state_reg[11]/NET0131  ;
  assign n1139 = n1036 & n1138 ;
  assign n1140 = \u5_state_reg[56]/NET0131  & ~\u5_state_reg[57]/NET0131  ;
  assign n1141 = n1026 & n1140 ;
  assign n1142 = n1018 & n1141 ;
  assign n1143 = n1015 & n1142 ;
  assign n1144 = \u5_state_reg[36]/NET0131  & ~\u5_state_reg[37]/NET0131  ;
  assign n1145 = n966 & n1144 ;
  assign n1146 = n971 & n1145 ;
  assign n1147 = n1088 & n1146 ;
  assign n1148 = ~n1143 & ~n1147 ;
  assign n1149 = ~n1139 & n1148 ;
  assign n1150 = \u5_state_reg[60]/NET0131  & ~\u5_state_reg[61]/NET0131  ;
  assign n1151 = n1007 & n1150 ;
  assign n1152 = n1009 & n1151 ;
  assign n1153 = n1115 & n1152 ;
  assign n1154 = ~\u5_state_reg[63]/NET0131  & \u5_state_reg[64]/NET0131  ;
  assign n1155 = n1006 & n1154 ;
  assign n1156 = n1010 & n1155 ;
  assign n1157 = n1115 & n1156 ;
  assign n1158 = ~n1153 & ~n1157 ;
  assign n1159 = n1149 & n1158 ;
  assign n1160 = ~\u5_state_reg[47]/NET0131  & \u5_state_reg[48]/NET0131  ;
  assign n1161 = n970 & n1160 ;
  assign n1162 = n968 & n1161 ;
  assign n1163 = n1088 & n1162 ;
  assign n1164 = ~\u5_state_reg[56]/NET0131  & \u5_state_reg[57]/NET0131  ;
  assign n1165 = n1026 & n1164 ;
  assign n1166 = n1018 & n1165 ;
  assign n1167 = n1015 & n1166 ;
  assign n1168 = ~\u5_state_reg[20]/NET0131  & \u5_state_reg[21]/NET0131  ;
  assign n1169 = n977 & n1168 ;
  assign n1170 = n1131 & n1169 ;
  assign n1171 = n1078 & n1170 ;
  assign n1172 = ~n1167 & ~n1171 ;
  assign n1173 = ~n1163 & n1172 ;
  assign n1174 = n1003 & n1029 ;
  assign n1175 = n1013 & n1174 ;
  assign n1176 = n989 & n1175 ;
  assign n1177 = ~\u5_state_reg[14]/NET0131  & \u5_state_reg[17]/NET0131  ;
  assign n1178 = n990 & n1177 ;
  assign n1179 = n995 & n1178 ;
  assign n1180 = n1176 & n1179 ;
  assign n1181 = ~\u5_state_reg[7]/NET0131  & \u5_state_reg[9]/NET0131  ;
  assign n1182 = n993 & n1181 ;
  assign n1183 = n992 & n1182 ;
  assign n1184 = n1176 & n1183 ;
  assign n1185 = ~n1180 & ~n1184 ;
  assign n1186 = ~\u5_state_reg[6]/NET0131  & \u5_state_reg[8]/NET0131  ;
  assign n1187 = n994 & n1186 ;
  assign n1188 = n992 & n1187 ;
  assign n1189 = n1176 & n1188 ;
  assign n1190 = \u5_state_reg[7]/NET0131  & ~\u5_state_reg[9]/NET0131  ;
  assign n1191 = n993 & n1190 ;
  assign n1192 = n992 & n1191 ;
  assign n1193 = n1176 & n1192 ;
  assign n1194 = ~n1189 & ~n1193 ;
  assign n1195 = n1185 & n1194 ;
  assign n1196 = n1173 & n1195 ;
  assign n1197 = n1159 & n1196 ;
  assign n1198 = n1137 & n1197 ;
  assign n1199 = ~\u5_lmr_ack_reg/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1200 = n983 & n1199 ;
  assign n1201 = \u0_sp_tms_reg[9]/NET0131  & ~n1200 ;
  assign n1202 = \u0_tms_reg[9]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1203 = ~\u5_lmr_ack_reg/NET0131  & n1202 ;
  assign n1204 = n983 & n1203 ;
  assign n1205 = ~n1201 & ~n1204 ;
  assign n1206 = \u0_sp_csc_reg[10]/NET0131  & ~n1200 ;
  assign n1207 = \u0_csc_reg[10]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1208 = ~\u5_lmr_ack_reg/NET0131  & n1207 ;
  assign n1209 = n983 & n1208 ;
  assign n1210 = ~n1206 & ~n1209 ;
  assign n1211 = ~n1205 & n1210 ;
  assign n1212 = \u0_sp_tms_reg[1]/NET0131  & ~n1200 ;
  assign n1213 = \u0_tms_reg[1]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1214 = ~\u5_lmr_ack_reg/NET0131  & n1213 ;
  assign n1215 = n983 & n1214 ;
  assign n1216 = ~n1212 & ~n1215 ;
  assign n1217 = \u0_sp_tms_reg[2]/NET0131  & ~n1200 ;
  assign n1218 = \u0_tms_reg[2]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1219 = ~\u5_lmr_ack_reg/NET0131  & n1218 ;
  assign n1220 = n983 & n1219 ;
  assign n1221 = ~n1217 & ~n1220 ;
  assign n1222 = n1216 & n1221 ;
  assign n1223 = \u0_sp_tms_reg[0]/NET0131  & ~n1200 ;
  assign n1224 = \u0_tms_reg[0]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1225 = ~\u5_lmr_ack_reg/NET0131  & n1224 ;
  assign n1226 = n983 & n1225 ;
  assign n1227 = ~n1223 & ~n1226 ;
  assign n1228 = n1210 & n1227 ;
  assign n1229 = n1222 & n1228 ;
  assign n1230 = ~n1211 & ~n1229 ;
  assign n1231 = wb_stb_i_pad & ~wb_we_i_pad ;
  assign n1232 = \u6_write_go_r1_reg/NET0131  & ~n1231 ;
  assign n1233 = wb_cyc_i_pad & ~wb_stb_i_pad ;
  assign n1234 = ~\u6_rmw_r_reg/NET0131  & wb_cyc_i_pad ;
  assign n1235 = ~n1233 & n1234 ;
  assign n1236 = n1232 & n1235 ;
  assign n1237 = ~n1048 & n1236 ;
  assign n1238 = n1189 & n1237 ;
  assign n1239 = ~n1230 & n1238 ;
  assign n1240 = ~n1198 & n1239 ;
  assign n1241 = ~\u5_ap_en_reg/NET0131  & ~n1240 ;
  assign n1242 = \u5_state_reg[14]/NET0131  & ~\u5_state_reg[17]/NET0131  ;
  assign n1243 = n990 & n1242 ;
  assign n1244 = n995 & n1243 ;
  assign n1245 = n1176 & n1244 ;
  assign n1246 = ~\u5_state_reg[5]/NET0131  & n998 ;
  assign n1247 = n1033 & n1246 ;
  assign n1248 = n1032 & n1247 ;
  assign n1249 = ~\u5_state_reg[12]/NET0131  & \u5_state_reg[13]/NET0131  ;
  assign n1250 = n1248 & n1249 ;
  assign n1251 = ~n1245 & ~n1250 ;
  assign n1252 = ~\u5_state_reg[18]/NET0131  & ~\u5_state_reg[21]/NET0131  ;
  assign n1253 = n1131 & n1252 ;
  assign n1254 = n1078 & n1253 ;
  assign n1255 = \u5_state_reg[19]/NET0131  & ~\u5_state_reg[20]/NET0131  ;
  assign n1256 = n1254 & n1255 ;
  assign n1257 = ~\u5_state_reg[46]/NET0131  & \u5_state_reg[49]/NET0131  ;
  assign n1258 = n969 & n1257 ;
  assign n1259 = n968 & n1258 ;
  assign n1260 = n1088 & n1259 ;
  assign n1261 = ~n1256 & ~n1260 ;
  assign n1262 = \u5_state_reg[26]/NET0131  & ~\u5_state_reg[27]/NET0131  ;
  assign n1263 = n974 & n1262 ;
  assign n1264 = n1131 & n1263 ;
  assign n1265 = n1130 & n1264 ;
  assign n1266 = \u5_state_reg[15]/NET0131  & ~\u5_state_reg[16]/NET0131  ;
  assign n1267 = n991 & n1266 ;
  assign n1268 = n995 & n1267 ;
  assign n1269 = n1176 & n1268 ;
  assign n1270 = \u5_state_reg[6]/NET0131  & ~\u5_state_reg[8]/NET0131  ;
  assign n1271 = n994 & n1270 ;
  assign n1272 = n992 & n1271 ;
  assign n1273 = n1176 & n1272 ;
  assign n1274 = ~n1269 & ~n1273 ;
  assign n1275 = ~n1265 & n1274 ;
  assign n1276 = n1261 & n1275 ;
  assign n1277 = n1251 & n1276 ;
  assign n1278 = \u5_state_reg[3]/NET0131  & n1000 ;
  assign n1279 = n999 & n1278 ;
  assign n1280 = ~\u5_state_reg[5]/NET0131  & n1279 ;
  assign n1281 = n1032 & n1280 ;
  assign n1282 = \u5_state_reg[32]/NET0131  & ~\u5_state_reg[33]/NET0131  ;
  assign n1283 = n985 & n1282 ;
  assign n1284 = n1080 & n1283 ;
  assign n1285 = n1078 & n1284 ;
  assign n1286 = ~n1281 & ~n1285 ;
  assign n1287 = \u5_state_reg[63]/NET0131  & ~\u5_state_reg[64]/NET0131  ;
  assign n1288 = n1006 & n1287 ;
  assign n1289 = n1010 & n1288 ;
  assign n1290 = n1115 & n1289 ;
  assign n1291 = n1004 & n1012 ;
  assign n1292 = n989 & n1291 ;
  assign n1293 = n1007 & n1008 ;
  assign n1294 = n1009 & n1016 ;
  assign n1295 = n1028 & n1294 ;
  assign n1296 = n1293 & n1295 ;
  assign n1297 = \u5_state_reg[50]/NET0131  & ~\u5_state_reg[51]/NET0131  ;
  assign n1298 = n1296 & n1297 ;
  assign n1299 = n1292 & n1298 ;
  assign n1300 = ~n1290 & ~n1299 ;
  assign n1301 = n1286 & n1300 ;
  assign n1302 = ~\u5_state_reg[3]/NET0131  & \u5_state_reg[5]/NET0131  ;
  assign n1303 = n1000 & n1302 ;
  assign n1304 = n999 & n1303 ;
  assign n1305 = n1032 & n1304 ;
  assign n1306 = n1011 & n1029 ;
  assign n1307 = n1004 & n1306 ;
  assign n1308 = n989 & n1307 ;
  assign n1309 = ~\u5_state_reg[0]/NET0131  & \u5_state_reg[1]/NET0131  ;
  assign n1310 = n1308 & n1309 ;
  assign n1311 = ~n1305 & ~n1310 ;
  assign n1312 = ~\u5_state_reg[58]/NET0131  & \u5_state_reg[59]/NET0131  ;
  assign n1313 = n1293 & n1312 ;
  assign n1314 = n1115 & n1313 ;
  assign n1315 = n1311 & ~n1314 ;
  assign n1316 = ~\u5_state_reg[19]/NET0131  & \u5_state_reg[20]/NET0131  ;
  assign n1317 = n1254 & n1316 ;
  assign n1318 = n1315 & ~n1317 ;
  assign n1319 = n1301 & n1318 ;
  assign n1320 = ~\u5_state_reg[36]/NET0131  & \u5_state_reg[37]/NET0131  ;
  assign n1321 = n966 & n1320 ;
  assign n1322 = n971 & n1321 ;
  assign n1323 = n1088 & n1322 ;
  assign n1324 = ~\u5_state_reg[30]/NET0131  & \u5_state_reg[31]/NET0131  ;
  assign n1325 = n984 & n1324 ;
  assign n1326 = n1080 & n1325 ;
  assign n1327 = n1078 & n1326 ;
  assign n1328 = \u5_state_reg[28]/NET0131  & ~\u5_state_reg[29]/NET0131  ;
  assign n1329 = n975 & n1328 ;
  assign n1330 = n1131 & n1329 ;
  assign n1331 = n1130 & n1330 ;
  assign n1332 = ~n1327 & ~n1331 ;
  assign n1333 = ~n1323 & n1332 ;
  assign n1334 = ~\u5_state_reg[38]/NET0131  & \u5_state_reg[39]/NET0131  ;
  assign n1335 = n960 & n1334 ;
  assign n1336 = n964 & n1335 ;
  assign n1337 = n1122 & n1336 ;
  assign n1338 = \u5_state_reg[0]/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n1339 = n1308 & n1338 ;
  assign n1340 = ~n1337 & ~n1339 ;
  assign n1341 = n1333 & n1340 ;
  assign n1342 = \u5_state_reg[58]/NET0131  & ~\u5_state_reg[59]/NET0131  ;
  assign n1343 = n1293 & n1342 ;
  assign n1344 = n1115 & n1343 ;
  assign n1345 = \u5_state_reg[52]/NET0131  & ~\u5_state_reg[53]/NET0131  ;
  assign n1346 = n1109 & n1345 ;
  assign n1347 = n1015 & n1346 ;
  assign n1348 = ~n1344 & ~n1347 ;
  assign n1349 = \u5_state_reg[47]/NET0131  & ~\u5_state_reg[48]/NET0131  ;
  assign n1350 = n970 & n1349 ;
  assign n1351 = n968 & n1350 ;
  assign n1352 = n1088 & n1351 ;
  assign n1353 = \u5_state_reg[38]/NET0131  & ~\u5_state_reg[39]/NET0131  ;
  assign n1354 = n960 & n1353 ;
  assign n1355 = ~\u5_state_reg[40]/NET0131  & \u5_state_reg[41]/NET0131  ;
  assign n1356 = n959 & n1355 ;
  assign n1357 = ~n1354 & ~n1356 ;
  assign n1358 = n964 & ~n1357 ;
  assign n1359 = n1122 & n1358 ;
  assign n1360 = ~\u5_state_reg[60]/NET0131  & \u5_state_reg[61]/NET0131  ;
  assign n1361 = n1007 & n1360 ;
  assign n1362 = n1009 & n1361 ;
  assign n1363 = n1115 & n1362 ;
  assign n1364 = ~n1359 & ~n1363 ;
  assign n1365 = ~n1352 & n1364 ;
  assign n1366 = n1348 & n1365 ;
  assign n1367 = n1341 & n1366 ;
  assign n1368 = n1319 & n1367 ;
  assign n1369 = n1277 & n1368 ;
  assign n1370 = ~\u5_state_reg[23]/NET0131  & \u5_state_reg[25]/NET0131  ;
  assign n1371 = n982 & n1370 ;
  assign n1372 = n1096 & n1371 ;
  assign n1373 = n1078 & n1372 ;
  assign n1374 = ~\u5_state_reg[50]/NET0131  & \u5_state_reg[51]/NET0131  ;
  assign n1375 = n1296 & n1374 ;
  assign n1376 = n1292 & n1375 ;
  assign n1377 = ~n1373 & ~n1376 ;
  assign n1378 = \u5_state_reg[44]/NET0131  & ~\u5_state_reg[45]/NET0131  ;
  assign n1379 = ~\u5_state_reg[42]/NET0131  & ~\u5_state_reg[43]/NET0131  ;
  assign n1380 = n961 & n1379 ;
  assign n1381 = n1378 & n1380 ;
  assign n1382 = n1122 & n1381 ;
  assign n1383 = ~\u5_state_reg[44]/NET0131  & ~\u5_state_reg[45]/NET0131  ;
  assign n1384 = n961 & n1383 ;
  assign n1385 = \u5_state_reg[42]/NET0131  & ~\u5_state_reg[43]/NET0131  ;
  assign n1386 = n1384 & n1385 ;
  assign n1387 = n1122 & n1386 ;
  assign n1388 = ~n1382 & ~n1387 ;
  assign n1389 = n1377 & n1388 ;
  assign n1390 = ~\u5_state_reg[44]/NET0131  & \u5_state_reg[45]/NET0131  ;
  assign n1391 = n1380 & n1390 ;
  assign n1392 = n1122 & n1391 ;
  assign n1393 = ~\u5_state_reg[42]/NET0131  & \u5_state_reg[43]/NET0131  ;
  assign n1394 = n1384 & n1393 ;
  assign n1395 = n1122 & n1394 ;
  assign n1396 = ~n1392 & ~n1395 ;
  assign n1397 = ~\u5_state_reg[54]/NET0131  & \u5_state_reg[55]/NET0131  ;
  assign n1398 = ~\u5_state_reg[57]/NET0131  & n1397 ;
  assign n1399 = n1019 & n1398 ;
  assign n1400 = n1015 & n1399 ;
  assign n1401 = \u5_state_reg[62]/NET0131  & ~\u5_state_reg[65]/NET0131  ;
  assign n1402 = n1005 & n1401 ;
  assign n1403 = n1010 & n1402 ;
  assign n1404 = n1115 & n1403 ;
  assign n1405 = ~n1400 & ~n1404 ;
  assign n1406 = n1396 & n1405 ;
  assign n1407 = n1389 & n1406 ;
  assign n1408 = ~\u5_state_reg[34]/NET0131  & \u5_state_reg[35]/NET0131  ;
  assign n1409 = n967 & n1408 ;
  assign n1410 = n971 & n1409 ;
  assign n1411 = n1088 & n1410 ;
  assign n1412 = \u5_state_reg[12]/NET0131  & ~\u5_state_reg[13]/NET0131  ;
  assign n1413 = n1248 & n1412 ;
  assign n1414 = \u5_state_reg[46]/NET0131  & ~\u5_state_reg[49]/NET0131  ;
  assign n1415 = n969 & n1414 ;
  assign n1416 = n968 & n1415 ;
  assign n1417 = n1088 & n1416 ;
  assign n1418 = ~\u5_state_reg[22]/NET0131  & \u5_state_reg[24]/NET0131  ;
  assign n1419 = n981 & n1418 ;
  assign n1420 = n1096 & n1419 ;
  assign n1421 = n1078 & n1420 ;
  assign n1422 = ~n1417 & ~n1421 ;
  assign n1423 = ~n1413 & n1422 ;
  assign n1424 = ~n1411 & n1423 ;
  assign n1425 = n1407 & n1424 ;
  assign n1426 = n1198 & n1425 ;
  assign n1427 = n1369 & n1426 ;
  assign n1428 = ~n1241 & ~n1427 ;
  assign n1429 = \u5_tmr_done_reg/NET0131  & n1234 ;
  assign n1430 = n1232 & n1429 ;
  assign n1431 = ~n1048 & n1430 ;
  assign n1432 = n1193 & n1431 ;
  assign n1433 = n1251 & ~n1432 ;
  assign n1434 = ~n1230 & ~n1433 ;
  assign n1435 = \u5_state_reg[2]/NET0131  & ~\u5_state_reg[4]/NET0131  ;
  assign n1436 = n1001 & n1435 ;
  assign n1437 = n999 & n1436 ;
  assign n1438 = n1032 & n1437 ;
  assign n1439 = \u5_cmd_a10_r_reg/P0001  & n1438 ;
  assign n1440 = ~\u5_state_reg[15]/NET0131  & \u5_state_reg[16]/NET0131  ;
  assign n1441 = n991 & n1440 ;
  assign n1442 = n995 & n1441 ;
  assign n1443 = n1176 & n1442 ;
  assign n1444 = \u5_tmr_done_reg/NET0131  & ~n1209 ;
  assign n1445 = ~n1206 & n1444 ;
  assign n1446 = \u5_cmd_a10_r_reg/P0001  & ~n1445 ;
  assign n1447 = n1443 & n1446 ;
  assign n1448 = ~n1439 & ~n1447 ;
  assign n1449 = \u5_state_reg[18]/NET0131  & ~\u5_state_reg[19]/NET0131  ;
  assign n1450 = ~\u5_state_reg[20]/NET0131  & n1449 ;
  assign n1451 = ~\u5_state_reg[21]/NET0131  & n1450 ;
  assign n1452 = n1131 & n1451 ;
  assign n1453 = n1078 & n1452 ;
  assign n1454 = \u5_state_reg[22]/NET0131  & ~\u5_state_reg[24]/NET0131  ;
  assign n1455 = n981 & n1454 ;
  assign n1456 = n1096 & n1455 ;
  assign n1457 = n1078 & n1456 ;
  assign n1458 = ~n1453 & ~n1457 ;
  assign n1459 = ~\u5_state_reg[26]/NET0131  & \u5_state_reg[27]/NET0131  ;
  assign n1460 = n974 & n1459 ;
  assign n1461 = n1131 & n1460 ;
  assign n1462 = n1130 & n1461 ;
  assign n1463 = ~\u5_state_reg[2]/NET0131  & \u5_state_reg[4]/NET0131  ;
  assign n1464 = n1001 & n1463 ;
  assign n1465 = n999 & n1464 ;
  assign n1466 = \u5_rfr_ack_r_reg/NET0131  & n1465 ;
  assign n1467 = n1032 & n1466 ;
  assign n1468 = ~n1462 & ~n1467 ;
  assign n1469 = n1458 & n1468 ;
  assign n1470 = n1448 & n1469 ;
  assign n1471 = ~n1434 & n1470 ;
  assign n1472 = ~n1428 & n1471 ;
  assign n1473 = n1075 & ~n1472 ;
  assign n1474 = n1315 & n1333 ;
  assign n1475 = ~n1273 & ~n1443 ;
  assign n1476 = n1474 & n1475 ;
  assign n1477 = \u5_wb_cycle_reg/NET0131  & ~n1205 ;
  assign n1478 = \u5_wb_cycle_reg/NET0131  & n1227 ;
  assign n1479 = n1222 & n1478 ;
  assign n1480 = ~n1477 & ~n1479 ;
  assign n1481 = n1245 & n1480 ;
  assign n1482 = n1032 & n1465 ;
  assign n1483 = ~n1462 & ~n1482 ;
  assign n1484 = ~n1285 & n1483 ;
  assign n1485 = ~n1481 & n1484 ;
  assign n1486 = n1107 & n1485 ;
  assign n1487 = ~n1413 & ~n1417 ;
  assign n1488 = ~n1269 & ~n1352 ;
  assign n1489 = n1487 & n1488 ;
  assign n1490 = n1340 & n1348 ;
  assign n1491 = n1489 & n1490 ;
  assign n1492 = n1486 & n1491 ;
  assign n1493 = n1476 & n1492 ;
  assign n1494 = ~n1189 & ~n1260 ;
  assign n1495 = ~n1256 & n1494 ;
  assign n1496 = ~n1163 & ~n1290 ;
  assign n1497 = ~n1167 & ~n1281 ;
  assign n1498 = n1496 & n1497 ;
  assign n1499 = n1495 & n1498 ;
  assign n1500 = n1128 & n1458 ;
  assign n1501 = n1499 & n1500 ;
  assign n1502 = n1407 & ~n1411 ;
  assign n1503 = ~n1193 & ~n1359 ;
  assign n1504 = ~n1363 & ~n1438 ;
  assign n1505 = ~n1171 & ~n1299 ;
  assign n1506 = n1504 & n1505 ;
  assign n1507 = n1503 & n1506 ;
  assign n1508 = n1159 & n1507 ;
  assign n1509 = n1502 & n1508 ;
  assign n1510 = n1501 & n1509 ;
  assign n1511 = n1493 & n1510 ;
  assign n1512 = ~\u5_wr_cycle_reg/NET0131  & ~n1511 ;
  assign n1513 = \u5_cmd_del_reg[1]/NET0131  & \u5_wr_cycle_reg/NET0131  ;
  assign n1514 = ~n1200 & ~n1513 ;
  assign n1515 = ~n1512 & n1514 ;
  assign n1516 = \u1_row_adr_reg[10]/P0001  & n1049 ;
  assign n1517 = \u1_row_adr_reg[10]/P0001  & n1052 ;
  assign n1518 = n1073 & n1517 ;
  assign n1519 = ~n1516 & ~n1518 ;
  assign n1520 = ~n1515 & n1519 ;
  assign n1521 = ~n1473 & n1520 ;
  assign n1522 = \u0_sp_csc_reg[1]/NET0131  & ~n1200 ;
  assign n1523 = \u0_csc_reg[1]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1524 = ~\u5_lmr_ack_reg/NET0131  & n1523 ;
  assign n1525 = n983 & n1524 ;
  assign n1526 = ~n1522 & ~n1525 ;
  assign n1527 = \u0_sp_csc_reg[3]/NET0131  & ~n1200 ;
  assign n1528 = \u0_csc_reg[3]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1529 = ~\u5_lmr_ack_reg/NET0131  & n1528 ;
  assign n1530 = n983 & n1529 ;
  assign n1531 = ~n1527 & ~n1530 ;
  assign n1532 = n1526 & n1531 ;
  assign n1533 = \u0_sp_csc_reg[2]/NET0131  & ~n1200 ;
  assign n1534 = \u0_csc_reg[2]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1535 = ~\u5_lmr_ack_reg/NET0131  & n1534 ;
  assign n1536 = n983 & n1535 ;
  assign n1537 = ~n1533 & ~n1536 ;
  assign n1538 = n1532 & n1537 ;
  assign n1539 = ~\u0_sp_tms_reg[10]/NET0131  & ~n1513 ;
  assign n1540 = ~n1200 & n1539 ;
  assign n1541 = ~n1512 & n1540 ;
  assign n1542 = n1538 & ~n1541 ;
  assign n1543 = ~n1521 & n1542 ;
  assign n1544 = ~n1526 & n1531 ;
  assign n1545 = \u6_wr_hold_reg/NET0131  & n1537 ;
  assign n1546 = n1544 & n1545 ;
  assign n1547 = ~\wb_addr_i[12]_pad  & ~n1546 ;
  assign n1548 = ~\u1_sram_addr_reg[10]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1549 = n1537 & n1548 ;
  assign n1550 = n1544 & n1549 ;
  assign n1551 = ~n1532 & ~n1550 ;
  assign n1552 = ~n1547 & n1551 ;
  assign n1553 = \u1_acs_addr_reg[10]/P0001  & ~n1537 ;
  assign n1554 = n1532 & n1553 ;
  assign n1555 = ~\u5_rfr_ack_r_reg/NET0131  & ~n1554 ;
  assign n1556 = ~n1552 & n1555 ;
  assign n1557 = ~n1543 & n1556 ;
  assign n1558 = ~\u1_col_adr_reg[0]/P0001  & ~n1049 ;
  assign n1559 = ~n1074 & n1558 ;
  assign n1560 = ~\u1_row_adr_reg[0]/P0001  & n1049 ;
  assign n1561 = ~\u1_row_adr_reg[0]/P0001  & n1052 ;
  assign n1562 = n1073 & n1561 ;
  assign n1563 = ~n1560 & ~n1562 ;
  assign n1564 = ~n1559 & n1563 ;
  assign n1565 = ~n1515 & ~n1564 ;
  assign n1566 = ~\u0_sp_tms_reg[0]/NET0131  & ~n1513 ;
  assign n1567 = ~n1200 & n1566 ;
  assign n1568 = ~n1512 & n1567 ;
  assign n1569 = n1538 & ~n1568 ;
  assign n1570 = ~n1565 & n1569 ;
  assign n1571 = \u1_acs_addr_reg[0]/P0001  & ~n1537 ;
  assign n1572 = n1532 & n1571 ;
  assign n1573 = ~\wb_addr_i[2]_pad  & ~n1546 ;
  assign n1574 = ~\u1_sram_addr_reg[0]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1575 = n1537 & n1574 ;
  assign n1576 = n1544 & n1575 ;
  assign n1577 = ~n1532 & ~n1576 ;
  assign n1578 = ~n1573 & n1577 ;
  assign n1579 = ~n1572 & ~n1578 ;
  assign n1580 = ~n1570 & n1579 ;
  assign n1581 = \u1_row_adr_reg[11]/P0001  & n1049 ;
  assign n1582 = \u1_row_adr_reg[11]/P0001  & n1052 ;
  assign n1583 = n1073 & n1582 ;
  assign n1584 = ~n1581 & ~n1583 ;
  assign n1585 = ~n1515 & n1584 ;
  assign n1586 = ~\u0_sp_tms_reg[11]/NET0131  & ~n1513 ;
  assign n1587 = ~n1200 & n1586 ;
  assign n1588 = ~n1512 & n1587 ;
  assign n1589 = n1538 & ~n1588 ;
  assign n1590 = ~n1585 & n1589 ;
  assign n1591 = \u1_acs_addr_reg[11]/P0001  & ~n1537 ;
  assign n1592 = n1532 & n1591 ;
  assign n1593 = ~\wb_addr_i[13]_pad  & ~n1546 ;
  assign n1594 = ~\u1_sram_addr_reg[11]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1595 = n1537 & n1594 ;
  assign n1596 = n1544 & n1595 ;
  assign n1597 = ~n1532 & ~n1596 ;
  assign n1598 = ~n1593 & n1597 ;
  assign n1599 = ~n1592 & ~n1598 ;
  assign n1600 = ~n1590 & n1599 ;
  assign n1601 = \u1_row_adr_reg[12]/P0001  & n1049 ;
  assign n1602 = \u1_row_adr_reg[12]/P0001  & n1052 ;
  assign n1603 = n1073 & n1602 ;
  assign n1604 = ~n1601 & ~n1603 ;
  assign n1605 = ~n1515 & n1604 ;
  assign n1606 = ~\u0_sp_tms_reg[12]/NET0131  & ~n1513 ;
  assign n1607 = ~n1200 & n1606 ;
  assign n1608 = ~n1512 & n1607 ;
  assign n1609 = n1538 & ~n1608 ;
  assign n1610 = ~n1605 & n1609 ;
  assign n1611 = \u1_acs_addr_reg[12]/P0001  & ~n1537 ;
  assign n1612 = n1532 & n1611 ;
  assign n1613 = ~\wb_addr_i[14]_pad  & ~n1546 ;
  assign n1614 = ~\u1_sram_addr_reg[12]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1615 = n1537 & n1614 ;
  assign n1616 = n1544 & n1615 ;
  assign n1617 = ~n1532 & ~n1616 ;
  assign n1618 = ~n1613 & n1617 ;
  assign n1619 = ~n1612 & ~n1618 ;
  assign n1620 = ~n1610 & n1619 ;
  assign n1621 = ~\u1_col_adr_reg[1]/P0001  & ~n1049 ;
  assign n1622 = ~n1074 & n1621 ;
  assign n1623 = ~\u1_row_adr_reg[1]/P0001  & n1049 ;
  assign n1624 = ~\u1_row_adr_reg[1]/P0001  & n1052 ;
  assign n1625 = n1073 & n1624 ;
  assign n1626 = ~n1623 & ~n1625 ;
  assign n1627 = ~n1622 & n1626 ;
  assign n1628 = ~n1515 & ~n1627 ;
  assign n1629 = ~\u0_sp_tms_reg[1]/NET0131  & ~n1513 ;
  assign n1630 = ~n1200 & n1629 ;
  assign n1631 = ~n1512 & n1630 ;
  assign n1632 = n1538 & ~n1631 ;
  assign n1633 = ~n1628 & n1632 ;
  assign n1634 = \u1_acs_addr_reg[1]/P0001  & ~n1537 ;
  assign n1635 = n1532 & n1634 ;
  assign n1636 = ~\wb_addr_i[3]_pad  & ~n1546 ;
  assign n1637 = ~\u1_sram_addr_reg[1]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1638 = n1537 & n1637 ;
  assign n1639 = n1544 & n1638 ;
  assign n1640 = ~n1532 & ~n1639 ;
  assign n1641 = ~n1636 & n1640 ;
  assign n1642 = ~n1635 & ~n1641 ;
  assign n1643 = ~n1633 & n1642 ;
  assign n1644 = ~\u1_col_adr_reg[2]/P0001  & ~n1049 ;
  assign n1645 = ~n1074 & n1644 ;
  assign n1646 = ~\u1_row_adr_reg[2]/P0001  & n1049 ;
  assign n1647 = ~\u1_row_adr_reg[2]/P0001  & n1052 ;
  assign n1648 = n1073 & n1647 ;
  assign n1649 = ~n1646 & ~n1648 ;
  assign n1650 = ~n1645 & n1649 ;
  assign n1651 = ~n1515 & ~n1650 ;
  assign n1652 = ~\u0_sp_tms_reg[2]/NET0131  & ~n1513 ;
  assign n1653 = ~n1200 & n1652 ;
  assign n1654 = ~n1512 & n1653 ;
  assign n1655 = n1538 & ~n1654 ;
  assign n1656 = ~n1651 & n1655 ;
  assign n1657 = \u1_acs_addr_reg[2]/P0001  & ~n1537 ;
  assign n1658 = n1532 & n1657 ;
  assign n1659 = ~\wb_addr_i[4]_pad  & ~n1546 ;
  assign n1660 = ~\u1_sram_addr_reg[2]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1661 = n1537 & n1660 ;
  assign n1662 = n1544 & n1661 ;
  assign n1663 = ~n1532 & ~n1662 ;
  assign n1664 = ~n1659 & n1663 ;
  assign n1665 = ~n1658 & ~n1664 ;
  assign n1666 = ~n1656 & n1665 ;
  assign n1667 = ~\u1_col_adr_reg[3]/P0001  & ~n1049 ;
  assign n1668 = ~n1074 & n1667 ;
  assign n1669 = ~\u1_row_adr_reg[3]/P0001  & n1049 ;
  assign n1670 = ~\u1_row_adr_reg[3]/P0001  & n1052 ;
  assign n1671 = n1073 & n1670 ;
  assign n1672 = ~n1669 & ~n1671 ;
  assign n1673 = ~n1668 & n1672 ;
  assign n1674 = ~n1515 & ~n1673 ;
  assign n1675 = ~\u0_sp_tms_reg[3]/NET0131  & ~n1513 ;
  assign n1676 = ~n1200 & n1675 ;
  assign n1677 = ~n1512 & n1676 ;
  assign n1678 = n1538 & ~n1677 ;
  assign n1679 = ~n1674 & n1678 ;
  assign n1680 = \u1_acs_addr_reg[3]/P0001  & ~n1537 ;
  assign n1681 = n1532 & n1680 ;
  assign n1682 = ~\wb_addr_i[5]_pad  & ~n1546 ;
  assign n1683 = ~\u1_sram_addr_reg[3]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1684 = n1537 & n1683 ;
  assign n1685 = n1544 & n1684 ;
  assign n1686 = ~n1532 & ~n1685 ;
  assign n1687 = ~n1682 & n1686 ;
  assign n1688 = ~n1681 & ~n1687 ;
  assign n1689 = ~n1679 & n1688 ;
  assign n1690 = ~\u1_col_adr_reg[4]/P0001  & ~n1049 ;
  assign n1691 = ~n1074 & n1690 ;
  assign n1692 = ~\u1_row_adr_reg[4]/P0001  & n1049 ;
  assign n1693 = ~\u1_row_adr_reg[4]/P0001  & n1052 ;
  assign n1694 = n1073 & n1693 ;
  assign n1695 = ~n1692 & ~n1694 ;
  assign n1696 = ~n1691 & n1695 ;
  assign n1697 = ~n1515 & ~n1696 ;
  assign n1698 = ~\u0_sp_tms_reg[4]/NET0131  & ~n1513 ;
  assign n1699 = ~n1200 & n1698 ;
  assign n1700 = ~n1512 & n1699 ;
  assign n1701 = n1538 & ~n1700 ;
  assign n1702 = ~n1697 & n1701 ;
  assign n1703 = \u1_acs_addr_reg[4]/P0001  & ~n1537 ;
  assign n1704 = n1532 & n1703 ;
  assign n1705 = ~\wb_addr_i[6]_pad  & ~n1546 ;
  assign n1706 = ~\u1_sram_addr_reg[4]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1707 = n1537 & n1706 ;
  assign n1708 = n1544 & n1707 ;
  assign n1709 = ~n1532 & ~n1708 ;
  assign n1710 = ~n1705 & n1709 ;
  assign n1711 = ~n1704 & ~n1710 ;
  assign n1712 = ~n1702 & n1711 ;
  assign n1713 = ~\u1_col_adr_reg[5]/P0001  & ~n1049 ;
  assign n1714 = ~n1074 & n1713 ;
  assign n1715 = ~\u1_row_adr_reg[5]/P0001  & n1049 ;
  assign n1716 = ~\u1_row_adr_reg[5]/P0001  & n1052 ;
  assign n1717 = n1073 & n1716 ;
  assign n1718 = ~n1715 & ~n1717 ;
  assign n1719 = ~n1714 & n1718 ;
  assign n1720 = ~n1515 & ~n1719 ;
  assign n1721 = ~\u0_sp_tms_reg[5]/NET0131  & ~n1513 ;
  assign n1722 = ~n1200 & n1721 ;
  assign n1723 = ~n1512 & n1722 ;
  assign n1724 = n1538 & ~n1723 ;
  assign n1725 = ~n1720 & n1724 ;
  assign n1726 = \u1_acs_addr_reg[5]/P0001  & ~n1537 ;
  assign n1727 = n1532 & n1726 ;
  assign n1728 = ~\wb_addr_i[7]_pad  & ~n1546 ;
  assign n1729 = ~\u1_sram_addr_reg[5]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1730 = n1537 & n1729 ;
  assign n1731 = n1544 & n1730 ;
  assign n1732 = ~n1532 & ~n1731 ;
  assign n1733 = ~n1728 & n1732 ;
  assign n1734 = ~n1727 & ~n1733 ;
  assign n1735 = ~n1725 & n1734 ;
  assign n1736 = ~\u1_col_adr_reg[6]/P0001  & ~n1049 ;
  assign n1737 = ~n1074 & n1736 ;
  assign n1738 = ~\u1_row_adr_reg[6]/P0001  & n1049 ;
  assign n1739 = ~\u1_row_adr_reg[6]/P0001  & n1052 ;
  assign n1740 = n1073 & n1739 ;
  assign n1741 = ~n1738 & ~n1740 ;
  assign n1742 = ~n1737 & n1741 ;
  assign n1743 = ~n1515 & ~n1742 ;
  assign n1744 = ~\u0_sp_tms_reg[6]/NET0131  & ~n1513 ;
  assign n1745 = ~n1200 & n1744 ;
  assign n1746 = ~n1512 & n1745 ;
  assign n1747 = n1538 & ~n1746 ;
  assign n1748 = ~n1743 & n1747 ;
  assign n1749 = \u1_acs_addr_reg[6]/P0001  & ~n1537 ;
  assign n1750 = n1532 & n1749 ;
  assign n1751 = ~\wb_addr_i[8]_pad  & ~n1546 ;
  assign n1752 = ~\u1_sram_addr_reg[6]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1753 = n1537 & n1752 ;
  assign n1754 = n1544 & n1753 ;
  assign n1755 = ~n1532 & ~n1754 ;
  assign n1756 = ~n1751 & n1755 ;
  assign n1757 = ~n1750 & ~n1756 ;
  assign n1758 = ~n1748 & n1757 ;
  assign n1759 = ~\u1_col_adr_reg[7]/P0001  & ~n1049 ;
  assign n1760 = ~n1074 & n1759 ;
  assign n1761 = ~\u1_row_adr_reg[7]/P0001  & n1049 ;
  assign n1762 = ~\u1_row_adr_reg[7]/P0001  & n1052 ;
  assign n1763 = n1073 & n1762 ;
  assign n1764 = ~n1761 & ~n1763 ;
  assign n1765 = ~n1760 & n1764 ;
  assign n1766 = ~n1515 & ~n1765 ;
  assign n1767 = ~\u0_sp_tms_reg[7]/NET0131  & ~n1513 ;
  assign n1768 = ~n1200 & n1767 ;
  assign n1769 = ~n1512 & n1768 ;
  assign n1770 = n1538 & ~n1769 ;
  assign n1771 = ~n1766 & n1770 ;
  assign n1772 = \u1_acs_addr_reg[7]/P0001  & ~n1537 ;
  assign n1773 = n1532 & n1772 ;
  assign n1774 = ~\wb_addr_i[9]_pad  & ~n1546 ;
  assign n1775 = ~\u1_sram_addr_reg[7]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1776 = n1537 & n1775 ;
  assign n1777 = n1544 & n1776 ;
  assign n1778 = ~n1532 & ~n1777 ;
  assign n1779 = ~n1774 & n1778 ;
  assign n1780 = ~n1773 & ~n1779 ;
  assign n1781 = ~n1771 & n1780 ;
  assign n1782 = ~\u1_col_adr_reg[8]/P0001  & ~n1049 ;
  assign n1783 = ~n1074 & n1782 ;
  assign n1784 = ~\u1_row_adr_reg[8]/P0001  & n1049 ;
  assign n1785 = ~\u1_row_adr_reg[8]/P0001  & n1052 ;
  assign n1786 = n1073 & n1785 ;
  assign n1787 = ~n1784 & ~n1786 ;
  assign n1788 = ~n1783 & n1787 ;
  assign n1789 = ~n1515 & ~n1788 ;
  assign n1790 = ~\u0_sp_tms_reg[8]/NET0131  & ~n1513 ;
  assign n1791 = ~n1200 & n1790 ;
  assign n1792 = ~n1512 & n1791 ;
  assign n1793 = n1538 & ~n1792 ;
  assign n1794 = ~n1789 & n1793 ;
  assign n1795 = \u1_acs_addr_reg[8]/P0001  & ~n1537 ;
  assign n1796 = n1532 & n1795 ;
  assign n1797 = ~\wb_addr_i[10]_pad  & ~n1546 ;
  assign n1798 = ~\u1_sram_addr_reg[8]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1799 = n1537 & n1798 ;
  assign n1800 = n1544 & n1799 ;
  assign n1801 = ~n1532 & ~n1800 ;
  assign n1802 = ~n1797 & n1801 ;
  assign n1803 = ~n1796 & ~n1802 ;
  assign n1804 = ~n1794 & n1803 ;
  assign n1805 = ~\u1_col_adr_reg[9]/P0001  & ~n1049 ;
  assign n1806 = ~n1074 & n1805 ;
  assign n1807 = ~\u1_row_adr_reg[9]/P0001  & n1049 ;
  assign n1808 = ~\u1_row_adr_reg[9]/P0001  & n1052 ;
  assign n1809 = n1073 & n1808 ;
  assign n1810 = ~n1807 & ~n1809 ;
  assign n1811 = ~n1806 & n1810 ;
  assign n1812 = ~n1515 & ~n1811 ;
  assign n1813 = ~\u0_sp_tms_reg[9]/NET0131  & ~n1513 ;
  assign n1814 = ~n1200 & n1813 ;
  assign n1815 = ~n1512 & n1814 ;
  assign n1816 = n1538 & ~n1815 ;
  assign n1817 = ~n1812 & n1816 ;
  assign n1818 = \u1_acs_addr_reg[9]/P0001  & ~n1537 ;
  assign n1819 = n1532 & n1818 ;
  assign n1820 = ~\wb_addr_i[11]_pad  & ~n1546 ;
  assign n1821 = ~\u1_sram_addr_reg[9]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n1822 = n1537 & n1821 ;
  assign n1823 = n1544 & n1822 ;
  assign n1824 = ~n1532 & ~n1823 ;
  assign n1825 = ~n1820 & n1824 ;
  assign n1826 = ~n1819 & ~n1825 ;
  assign n1827 = ~n1817 & n1826 ;
  assign n1828 = ~\u5_rfr_ack_r_reg/NET0131  & ~\u5_susp_sel_r_reg/NET0131  ;
  assign n1829 = ~\u0_cs_reg[0]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1830 = ~\u5_lmr_ack_reg/NET0131  & n1829 ;
  assign n1831 = n983 & n1830 ;
  assign n1832 = n1828 & n1831 ;
  assign n1833 = ~\u0_spec_req_cs_reg[0]/NET0131  & n1828 ;
  assign n1834 = ~n1200 & n1833 ;
  assign n1835 = ~n1832 & ~n1834 ;
  assign n1836 = ~\u0_u0_csc_reg[1]/NET0131  & ~\u0_u0_csc_reg[2]/NET0131  ;
  assign n1837 = \u0_u0_csc_reg[0]/NET0131  & ~\u0_u0_csc_reg[3]/NET0131  ;
  assign n1838 = n1836 & n1837 ;
  assign n1839 = ~n1828 & ~n1838 ;
  assign n1840 = n1835 & ~n1839 ;
  assign n1841 = \u5_cmd_del_reg[3]/NET0131  & \u5_wr_cycle_reg/NET0131  ;
  assign n1842 = \u5_wr_cycle_reg/NET0131  & ~n1841 ;
  assign n1843 = ~n1304 & ~n1465 ;
  assign n1844 = n1032 & ~n1843 ;
  assign n1845 = ~\u4_rfr_req_reg/NET0131  & ~n1844 ;
  assign n1846 = ~\u5_rfr_ack_r_reg/NET0131  & n1844 ;
  assign n1847 = ~n1311 & ~n1846 ;
  assign n1848 = ~n1845 & n1847 ;
  assign n1849 = ~n1135 & ~n1180 ;
  assign n1850 = \u5_mc_c_oe_reg/NET0131  & n1828 ;
  assign n1851 = n1849 & n1850 ;
  assign n1852 = \u0_tms_reg[19]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1853 = ~\u5_lmr_ack_reg/NET0131  & n1852 ;
  assign n1854 = n983 & n1853 ;
  assign n1855 = \u0_sp_tms_reg[19]/NET0131  & ~n1200 ;
  assign n1856 = ~n1854 & ~n1855 ;
  assign n1857 = \u0_tms_reg[18]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1858 = ~\u5_lmr_ack_reg/NET0131  & n1857 ;
  assign n1859 = n983 & n1858 ;
  assign n1860 = \u0_sp_tms_reg[18]/NET0131  & ~n1200 ;
  assign n1861 = ~n1859 & ~n1860 ;
  assign n1862 = n1856 & n1861 ;
  assign n1863 = n1851 & n1862 ;
  assign n1864 = ~n1848 & n1863 ;
  assign n1865 = \u0_tms_reg[17]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1866 = ~\u5_lmr_ack_reg/NET0131  & n1865 ;
  assign n1867 = n983 & n1866 ;
  assign n1868 = \u0_sp_tms_reg[17]/NET0131  & ~n1200 ;
  assign n1869 = ~n1867 & ~n1868 ;
  assign n1870 = ~\u0_tms_reg[16]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1871 = ~\u5_lmr_ack_reg/NET0131  & n1870 ;
  assign n1872 = n983 & n1871 ;
  assign n1873 = ~\u0_sp_tms_reg[16]/NET0131  & ~n1200 ;
  assign n1874 = ~n1872 & ~n1873 ;
  assign n1875 = n1869 & ~n1874 ;
  assign n1876 = n1851 & n1875 ;
  assign n1877 = ~n1848 & n1876 ;
  assign n1878 = n1864 & n1877 ;
  assign n1879 = n1260 & ~n1878 ;
  assign n1880 = n1496 & ~n1879 ;
  assign n1881 = ~n1337 & n1396 ;
  assign n1882 = ~n1382 & ~n1417 ;
  assign n1883 = ~n1250 & n1882 ;
  assign n1884 = n1881 & n1883 ;
  assign n1885 = ~n1153 & n1185 ;
  assign n1886 = ~n1387 & ~n1421 ;
  assign n1887 = ~\u5_tmr2_done_reg/NET0131  & n1297 ;
  assign n1888 = n1296 & n1887 ;
  assign n1889 = n1292 & n1888 ;
  assign n1890 = ~n1135 & ~n1889 ;
  assign n1891 = n1886 & n1890 ;
  assign n1892 = n1885 & n1891 ;
  assign n1893 = n1884 & n1892 ;
  assign n1894 = n1232 & n1234 ;
  assign n1895 = ~n1048 & n1894 ;
  assign n1896 = \u6_read_go_r1_reg/NET0131  & n1234 ;
  assign n1897 = ~n1048 & n1896 ;
  assign n1898 = ~n1895 & ~n1897 ;
  assign n1899 = n1233 & ~n1898 ;
  assign n1900 = ~n1526 & ~n1537 ;
  assign n1901 = n1531 & n1900 ;
  assign n1902 = ~n1899 & n1901 ;
  assign n1903 = ~n1233 & ~n1895 ;
  assign n1904 = ~n1898 & ~n1903 ;
  assign n1905 = n1544 & ~n1904 ;
  assign n1906 = n1537 & n1905 ;
  assign n1907 = ~n1902 & ~n1906 ;
  assign n1908 = \u0_cs_reg[1]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n1909 = ~\u5_lmr_ack_reg/NET0131  & n1908 ;
  assign n1910 = n983 & n1909 ;
  assign n1911 = n1828 & n1910 ;
  assign n1912 = \u0_spec_req_cs_reg[1]/NET0131  & n1828 ;
  assign n1913 = ~n1200 & n1912 ;
  assign n1914 = ~n1911 & ~n1913 ;
  assign n1915 = ~\u0_u1_csc_reg[1]/NET0131  & ~\u0_u1_csc_reg[2]/NET0131  ;
  assign n1916 = \u0_u1_csc_reg[0]/NET0131  & ~\u0_u1_csc_reg[3]/NET0131  ;
  assign n1917 = n1915 & n1916 ;
  assign n1918 = ~n1828 & n1917 ;
  assign n1919 = n1914 & ~n1918 ;
  assign n1920 = ~n1840 & n1919 ;
  assign n1921 = \u5_lookup_ready2_reg/NET0131  & ~n1898 ;
  assign n1922 = ~n1920 & n1921 ;
  assign n1923 = \u0_lmr_req_reg/NET0131  & \u5_lookup_ready2_reg/NET0131  ;
  assign n1924 = ~\u0_init_req_reg/NET0131  & ~n1923 ;
  assign n1925 = \u5_susp_req_r_reg/NET0131  & ~\u5_wb_cycle_reg/NET0131  ;
  assign n1926 = ~\u4_rfr_req_reg/NET0131  & ~n1925 ;
  assign n1927 = n1924 & n1926 ;
  assign n1928 = n1309 & n1927 ;
  assign n1929 = n1308 & n1928 ;
  assign n1930 = n1922 & n1929 ;
  assign n1931 = ~n1907 & n1930 ;
  assign n1932 = n1366 & ~n1931 ;
  assign n1933 = n1893 & n1932 ;
  assign n1934 = ~\u5_wb_wait_r_reg/P0001  & n1273 ;
  assign n1935 = ~n1269 & n1458 ;
  assign n1936 = n1443 & n1445 ;
  assign n1937 = n1483 & ~n1936 ;
  assign n1938 = n1935 & n1937 ;
  assign n1939 = ~n1934 & n1938 ;
  assign n1940 = ~n1265 & ~n1317 ;
  assign n1941 = ~n1147 & ~n1323 ;
  assign n1942 = ~\u5_tmr_done_reg/NET0131  & n1157 ;
  assign n1943 = n1941 & ~n1942 ;
  assign n1944 = n1940 & n1943 ;
  assign n1945 = n1939 & n1944 ;
  assign n1946 = n1933 & n1945 ;
  assign n1947 = n1880 & n1946 ;
  assign n1948 = n1245 & ~n1480 ;
  assign n1949 = n1311 & n1467 ;
  assign n1950 = n1227 & n1850 ;
  assign n1951 = n1222 & n1950 ;
  assign n1952 = n1849 & n1951 ;
  assign n1953 = ~n1949 & n1952 ;
  assign n1954 = ~n1848 & n1953 ;
  assign n1955 = n1222 & n1227 ;
  assign n1956 = n1205 & ~n1955 ;
  assign n1957 = ~\u5_burst_cnt_reg[0]/NET0131  & ~\u5_burst_cnt_reg[1]/NET0131  ;
  assign n1958 = ~\u5_burst_cnt_reg[2]/NET0131  & n1957 ;
  assign n1959 = ~\u5_burst_cnt_reg[3]/NET0131  & ~\u5_burst_cnt_reg[4]/NET0131  ;
  assign n1960 = ~\u5_burst_cnt_reg[5]/NET0131  & ~\u5_burst_cnt_reg[6]/NET0131  ;
  assign n1961 = n1959 & n1960 ;
  assign n1962 = n1958 & n1961 ;
  assign n1963 = ~\u5_burst_cnt_reg[7]/NET0131  & ~\u5_burst_cnt_reg[8]/NET0131  ;
  assign n1964 = ~\u5_burst_cnt_reg[10]/NET0131  & ~\u5_burst_cnt_reg[9]/NET0131  ;
  assign n1965 = n1963 & n1964 ;
  assign n1966 = n1962 & n1965 ;
  assign n1967 = ~\u5_wb_write_go_r_reg/NET0131  & ~n1966 ;
  assign n1968 = n1956 & n1967 ;
  assign n1969 = ~n1954 & n1968 ;
  assign n1970 = ~\u5_cnt_reg/NET0131  & n1205 ;
  assign n1971 = ~n1955 & n1970 ;
  assign n1972 = \u5_cke_r_reg/NET0131  & ~n1971 ;
  assign n1973 = ~n1899 & n1970 ;
  assign n1974 = ~n1955 & n1973 ;
  assign n1975 = ~n1972 & ~n1974 ;
  assign n1976 = n1245 & ~n1975 ;
  assign n1977 = n1969 & n1976 ;
  assign n1978 = ~n1948 & ~n1977 ;
  assign n1979 = ~n1841 & n1978 ;
  assign n1980 = n1947 & n1979 ;
  assign n1981 = ~n1842 & ~n1980 ;
  assign n1982 = n1840 & n1981 ;
  assign n1983 = ~n1919 & n1981 ;
  assign n1984 = n1481 & ~n1975 ;
  assign n1985 = ~n1969 & n1984 ;
  assign n1986 = n1497 & n1503 ;
  assign n1987 = n1443 & ~n1445 ;
  assign n1988 = ~n1305 & ~n1314 ;
  assign n1989 = ~n1987 & n1988 ;
  assign n1990 = n1986 & n1989 ;
  assign n1991 = n1495 & n1990 ;
  assign n1992 = n1149 & n1341 ;
  assign n1993 = n1991 & n1992 ;
  assign n1994 = n1137 & n1993 ;
  assign n1995 = n1924 & ~n1925 ;
  assign n1996 = \u5_lookup_ready2_reg/NET0131  & n1995 ;
  assign n1997 = ~n1898 & n1996 ;
  assign n1998 = ~n1920 & n1997 ;
  assign n1999 = n1237 & n1900 ;
  assign n2000 = n1531 & ~n1999 ;
  assign n2001 = n1998 & ~n2000 ;
  assign n2002 = n1310 & ~n2001 ;
  assign n2003 = \u4_rfr_req_reg/NET0131  & n1309 ;
  assign n2004 = n1308 & n2003 ;
  assign n2005 = ~n1285 & ~n2004 ;
  assign n2006 = ~n1273 & ~n1347 ;
  assign n2007 = n2005 & n2006 ;
  assign n2008 = n1506 & n2007 ;
  assign n2009 = \u5_tmr_done_reg/NET0131  & n1157 ;
  assign n2010 = n1885 & ~n2009 ;
  assign n2011 = n2008 & n2010 ;
  assign n2012 = ~n2002 & n2011 ;
  assign n2013 = n1245 & ~n1974 ;
  assign n2014 = ~n1972 & n2013 ;
  assign n2015 = n1480 & n2014 ;
  assign n2016 = n1425 & ~n2015 ;
  assign n2017 = n2012 & n2016 ;
  assign n2018 = n1994 & n2017 ;
  assign n2019 = ~n1985 & n2018 ;
  assign n2020 = \u5_cmd_asserted_reg/NET0131  & \u5_mc_le_reg/NET0131  ;
  assign n2021 = \u5_mc_le_reg/NET0131  & ~n2020 ;
  assign n2022 = n1978 & ~n2020 ;
  assign n2023 = n1947 & n2022 ;
  assign n2024 = ~n2021 & ~n2023 ;
  assign n2025 = ~n1848 & n1851 ;
  assign n2026 = n1237 & n1531 ;
  assign n2027 = n1900 & n2026 ;
  assign n2028 = n1929 & n2027 ;
  assign n2029 = n1922 & n2028 ;
  assign n2030 = ~n1290 & ~n2029 ;
  assign n2031 = ~n2025 & ~n2030 ;
  assign n2032 = \u0_sp_tms_reg[14]/NET0131  & ~n1200 ;
  assign n2033 = \u0_tms_reg[14]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2034 = ~\u5_lmr_ack_reg/NET0131  & n2033 ;
  assign n2035 = n983 & n2034 ;
  assign n2036 = ~n2032 & ~n2035 ;
  assign n2037 = ~n2030 & n2036 ;
  assign n2038 = ~n2031 & n2037 ;
  assign n2039 = ~n1363 & n1404 ;
  assign n2040 = \u5_tmr_done_reg/NET0131  & n1009 ;
  assign n2041 = n1361 & n2040 ;
  assign n2042 = n1115 & n2041 ;
  assign n2043 = ~n2039 & ~n2042 ;
  assign n2044 = \u0_sp_tms_reg[10]/NET0131  & ~n1200 ;
  assign n2045 = \u0_tms_reg[10]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2046 = ~\u5_lmr_ack_reg/NET0131  & n2045 ;
  assign n2047 = n983 & n2046 ;
  assign n2048 = ~n2044 & ~n2047 ;
  assign n2049 = ~n2043 & n2048 ;
  assign n2050 = ~n1537 & n1905 ;
  assign n2051 = n1930 & n2050 ;
  assign n2052 = ~n1153 & ~n2051 ;
  assign n2053 = n1221 & n1851 ;
  assign n2054 = ~n1848 & n2053 ;
  assign n2055 = ~n2052 & ~n2054 ;
  assign n2056 = n2043 & ~n2055 ;
  assign n2057 = ~n2049 & ~n2056 ;
  assign n2058 = ~\u5_state_reg[9]/NET0131  & ~n1934 ;
  assign n2059 = n1938 & n2058 ;
  assign n2060 = ~\u5_state_reg[17]/NET0131  & ~\u5_state_reg[20]/NET0131  ;
  assign n2061 = ~\u5_state_reg[24]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2062 = n2060 & n2061 ;
  assign n2063 = ~\u5_timer_reg[2]/NET0131  & ~\u5_timer_reg[3]/NET0131  ;
  assign n2064 = ~\u5_timer_reg[4]/NET0131  & ~\u5_timer_reg[5]/NET0131  ;
  assign n2065 = n2063 & n2064 ;
  assign n2066 = ~\u5_timer_reg[0]/NET0131  & ~\u5_timer_reg[1]/NET0131  ;
  assign n2067 = ~\u5_timer_reg[6]/NET0131  & ~\u5_timer_reg[7]/NET0131  ;
  assign n2068 = n2066 & n2067 ;
  assign n2069 = n2065 & n2068 ;
  assign n2070 = ~\u5_mc_le_reg/NET0131  & ~\u5_timer_reg[1]/NET0131  ;
  assign n2071 = ~\u5_timer_reg[0]/NET0131  & n2070 ;
  assign n2072 = ~n2069 & n2071 ;
  assign n2073 = ~\u5_timer_reg[2]/NET0131  & n985 ;
  assign n2074 = ~n2072 & n2073 ;
  assign n2075 = \u5_timer_reg[2]/NET0131  & n985 ;
  assign n2076 = n2072 & n2075 ;
  assign n2077 = ~n2074 & ~n2076 ;
  assign n2078 = ~\u5_state_reg[35]/NET0131  & n2077 ;
  assign n2079 = n2062 & ~n2078 ;
  assign n2080 = \u0_sp_tms_reg[26]/NET0131  & ~n1200 ;
  assign n2081 = \u0_tms_reg[26]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2082 = ~\u5_lmr_ack_reg/NET0131  & n2081 ;
  assign n2083 = n983 & n2082 ;
  assign n2084 = ~n2062 & ~n2083 ;
  assign n2085 = ~n2080 & n2084 ;
  assign n2086 = n1851 & n2085 ;
  assign n2087 = ~n1848 & n2086 ;
  assign n2088 = ~n2079 & ~n2087 ;
  assign n2089 = n2059 & n2088 ;
  assign n2090 = \u0_tms_reg[22]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2091 = ~\u5_lmr_ack_reg/NET0131  & n2090 ;
  assign n2092 = n983 & n2091 ;
  assign n2093 = \u0_sp_tms_reg[22]/NET0131  & ~n1200 ;
  assign n2094 = ~n2092 & ~n2093 ;
  assign n2095 = n1851 & n2094 ;
  assign n2096 = ~n1848 & n2095 ;
  assign n2097 = ~n1938 & ~n2096 ;
  assign n2098 = ~\u5_state_reg[13]/NET0131  & ~\u5_state_reg[14]/NET0131  ;
  assign n2099 = n1851 & n1856 ;
  assign n2100 = ~n1848 & n2099 ;
  assign n2101 = n1934 & n1938 ;
  assign n2102 = ~n2100 & n2101 ;
  assign n2103 = n2098 & ~n2102 ;
  assign n2104 = ~n2097 & n2103 ;
  assign n2105 = ~n2089 & n2104 ;
  assign n2106 = n2052 & ~n2105 ;
  assign n2107 = ~\u0_tms_reg[21]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2108 = ~\u5_lmr_ack_reg/NET0131  & n2107 ;
  assign n2109 = n983 & n2108 ;
  assign n2110 = ~\u0_sp_tms_reg[21]/NET0131  & ~n1200 ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = n1874 & n2111 ;
  assign n2113 = n1851 & ~n2112 ;
  assign n2114 = ~n1848 & n2113 ;
  assign n2115 = ~n1874 & ~n2111 ;
  assign n2116 = n1851 & n2115 ;
  assign n2117 = ~n1848 & n2116 ;
  assign n2118 = \u0_sp_tms_reg[15]/NET0131  & ~n1200 ;
  assign n2119 = \u0_tms_reg[15]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2120 = ~\u5_lmr_ack_reg/NET0131  & n2119 ;
  assign n2121 = n983 & n2120 ;
  assign n2122 = ~n2118 & ~n2121 ;
  assign n2123 = \u0_sp_tms_reg[20]/NET0131  & ~n1200 ;
  assign n2124 = \u0_tms_reg[20]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2125 = ~\u5_lmr_ack_reg/NET0131  & n2124 ;
  assign n2126 = n983 & n2125 ;
  assign n2127 = ~n2123 & ~n2126 ;
  assign n2128 = ~n2122 & ~n2127 ;
  assign n2129 = n1851 & ~n2128 ;
  assign n2130 = ~n1848 & n2129 ;
  assign n2131 = ~n2117 & ~n2130 ;
  assign n2132 = n2114 & ~n2131 ;
  assign n2133 = ~n2096 & ~n2098 ;
  assign n2134 = ~n2132 & n2133 ;
  assign n2135 = n2096 & ~n2098 ;
  assign n2136 = n2132 & n2135 ;
  assign n2137 = ~n2134 & ~n2136 ;
  assign n2138 = ~n2049 & n2137 ;
  assign n2139 = n2106 & n2138 ;
  assign n2140 = ~n2057 & ~n2139 ;
  assign n2141 = ~n2025 & ~n2043 ;
  assign n2142 = n2030 & ~n2141 ;
  assign n2143 = ~n2031 & n2142 ;
  assign n2144 = n2140 & n2143 ;
  assign n2145 = ~n2038 & ~n2144 ;
  assign n2146 = \u5_cmd_asserted_reg/NET0131  & n1249 ;
  assign n2147 = ~\u5_mem_ack_r_reg/NET0131  & \u5_wb_cycle_reg/NET0131  ;
  assign n2148 = n1237 & n2147 ;
  assign n2149 = n2146 & n2148 ;
  assign n2150 = n1248 & n2149 ;
  assign n2151 = ~n1966 & n2150 ;
  assign n2152 = ~n1954 & n2151 ;
  assign n2153 = ~\u5_mem_ack_r_reg/NET0131  & \u5_wr_cycle_reg/NET0131  ;
  assign n2154 = n1237 & n2153 ;
  assign n2155 = n1245 & n2154 ;
  assign n2156 = ~n1966 & n2155 ;
  assign n2157 = ~n1954 & n2156 ;
  assign n2158 = n1127 & ~n1376 ;
  assign n2159 = ~n1157 & ~n1363 ;
  assign n2160 = \u5_tmr_done_reg/NET0131  & ~n2159 ;
  assign n2161 = ~\u5_mem_ack_r_reg/NET0131  & n1237 ;
  assign n2162 = n1189 & n2161 ;
  assign n2163 = ~n2160 & ~n2162 ;
  assign n2164 = n2158 & n2163 ;
  assign n2165 = wb_stb_i_pad & wb_we_i_pad ;
  assign n2166 = ~\u5_ack_cnt_reg[0]/NET0131  & ~\u5_ack_cnt_reg[1]/NET0131  ;
  assign n2167 = ~\u5_ack_cnt_reg[2]/NET0131  & ~\u5_ack_cnt_reg[3]/NET0131  ;
  assign n2168 = n2166 & n2167 ;
  assign n2169 = n1896 & ~n2168 ;
  assign n2170 = ~n1048 & n2169 ;
  assign n2171 = ~n2165 & n2170 ;
  assign n2172 = ~\u5_mem_ack_r_reg/NET0131  & n2171 ;
  assign n2173 = ~n1899 & n2172 ;
  assign n2174 = n1237 & n1537 ;
  assign n2175 = n1544 & n2174 ;
  assign n2176 = n1929 & n2175 ;
  assign n2177 = n1922 & n2176 ;
  assign n2178 = \u5_cmd_asserted_reg/NET0131  & n1342 ;
  assign n2179 = n1293 & n2178 ;
  assign n2180 = n1115 & n2179 ;
  assign n2181 = n2161 & n2180 ;
  assign n2182 = ~\u5_mem_ack_r_reg/NET0131  & n1431 ;
  assign n2183 = n1193 & n2182 ;
  assign n2184 = ~n2181 & ~n2183 ;
  assign n2185 = ~n2177 & n2184 ;
  assign n2186 = ~n2173 & n2185 ;
  assign n2187 = n2164 & n2186 ;
  assign n2188 = ~n2157 & n2187 ;
  assign n2189 = ~n2152 & n2188 ;
  assign n2190 = ~\wb_addr_i[29]_pad  & ~\wb_addr_i[30]_pad  ;
  assign n2191 = ~\wb_addr_i[31]_pad  & n2190 ;
  assign n2192 = ~n1898 & n2191 ;
  assign n2193 = ~n2189 & n2192 ;
  assign n2194 = ~n1045 & n2193 ;
  assign n2195 = ~\u3_u0_rd_adr_reg[2]/NET0131  & ~\u3_u0_rd_adr_reg[3]/NET0131  ;
  assign n2196 = \u3_u0_rd_adr_reg[0]/NET0131  & ~\u3_u0_rd_adr_reg[1]/NET0131  ;
  assign n2197 = n2195 & n2196 ;
  assign n2198 = \u3_u0_r0_reg[13]/P0001  & n2197 ;
  assign n2199 = ~\u3_u0_rd_adr_reg[0]/NET0131  & \u3_u0_rd_adr_reg[1]/NET0131  ;
  assign n2200 = n2195 & n2199 ;
  assign n2201 = \u3_u0_r1_reg[13]/P0001  & n2200 ;
  assign n2202 = ~n2198 & ~n2201 ;
  assign n2203 = ~\u3_u0_rd_adr_reg[0]/NET0131  & ~\u3_u0_rd_adr_reg[1]/NET0131  ;
  assign n2204 = ~\u3_u0_rd_adr_reg[2]/NET0131  & \u3_u0_rd_adr_reg[3]/NET0131  ;
  assign n2205 = n2203 & n2204 ;
  assign n2206 = \u3_u0_r3_reg[13]/P0001  & n2205 ;
  assign n2207 = \u3_u0_rd_adr_reg[2]/NET0131  & ~\u3_u0_rd_adr_reg[3]/NET0131  ;
  assign n2208 = n2203 & n2207 ;
  assign n2209 = \u3_u0_r2_reg[13]/P0001  & n2208 ;
  assign n2210 = ~n2206 & ~n2209 ;
  assign n2211 = n2202 & n2210 ;
  assign n2212 = \u3_u0_r0_reg[9]/P0001  & n2197 ;
  assign n2213 = \u3_u0_r1_reg[9]/P0001  & n2200 ;
  assign n2214 = ~n2212 & ~n2213 ;
  assign n2215 = \u3_u0_r3_reg[9]/P0001  & n2205 ;
  assign n2216 = \u3_u0_r2_reg[9]/P0001  & n2208 ;
  assign n2217 = ~n2215 & ~n2216 ;
  assign n2218 = n2214 & n2217 ;
  assign n2219 = n2211 & ~n2218 ;
  assign n2220 = ~n2211 & n2218 ;
  assign n2221 = ~n2219 & ~n2220 ;
  assign n2222 = \u3_u0_r0_reg[14]/P0001  & n2197 ;
  assign n2223 = \u3_u0_r1_reg[14]/P0001  & n2200 ;
  assign n2224 = ~n2222 & ~n2223 ;
  assign n2225 = \u3_u0_r3_reg[14]/P0001  & n2205 ;
  assign n2226 = \u3_u0_r2_reg[14]/P0001  & n2208 ;
  assign n2227 = ~n2225 & ~n2226 ;
  assign n2228 = n2224 & n2227 ;
  assign n2229 = \u3_u0_r0_reg[11]/P0001  & n2197 ;
  assign n2230 = \u3_u0_r1_reg[11]/P0001  & n2200 ;
  assign n2231 = ~n2229 & ~n2230 ;
  assign n2232 = \u3_u0_r3_reg[11]/P0001  & n2205 ;
  assign n2233 = \u3_u0_r2_reg[11]/P0001  & n2208 ;
  assign n2234 = ~n2232 & ~n2233 ;
  assign n2235 = n2231 & n2234 ;
  assign n2236 = \u3_u0_r0_reg[12]/P0001  & n2197 ;
  assign n2237 = \u3_u0_r1_reg[12]/P0001  & n2200 ;
  assign n2238 = ~n2236 & ~n2237 ;
  assign n2239 = \u3_u0_r3_reg[12]/P0001  & n2205 ;
  assign n2240 = \u3_u0_r2_reg[12]/P0001  & n2208 ;
  assign n2241 = ~n2239 & ~n2240 ;
  assign n2242 = n2238 & n2241 ;
  assign n2243 = ~n2235 & ~n2242 ;
  assign n2244 = n2235 & n2242 ;
  assign n2245 = ~n2243 & ~n2244 ;
  assign n2246 = n2228 & ~n2245 ;
  assign n2247 = ~n2228 & n2245 ;
  assign n2248 = ~n2246 & ~n2247 ;
  assign n2249 = n2221 & n2248 ;
  assign n2250 = ~n2221 & ~n2248 ;
  assign n2251 = ~n2249 & ~n2250 ;
  assign n2252 = \u3_u0_r0_reg[8]/P0001  & n2197 ;
  assign n2253 = \u3_u0_r1_reg[8]/P0001  & n2200 ;
  assign n2254 = ~n2252 & ~n2253 ;
  assign n2255 = \u3_u0_r3_reg[8]/P0001  & n2205 ;
  assign n2256 = \u3_u0_r2_reg[8]/P0001  & n2208 ;
  assign n2257 = ~n2255 & ~n2256 ;
  assign n2258 = n2254 & n2257 ;
  assign n2259 = \u3_u0_r0_reg[15]/P0001  & n2197 ;
  assign n2260 = \u3_u0_r1_reg[15]/P0001  & n2200 ;
  assign n2261 = ~n2259 & ~n2260 ;
  assign n2262 = \u3_u0_r3_reg[15]/P0001  & n2205 ;
  assign n2263 = \u3_u0_r2_reg[15]/P0001  & n2208 ;
  assign n2264 = ~n2262 & ~n2263 ;
  assign n2265 = n2261 & n2264 ;
  assign n2266 = n2258 & ~n2265 ;
  assign n2267 = ~n2258 & n2265 ;
  assign n2268 = ~n2266 & ~n2267 ;
  assign n2269 = \u3_u0_r0_reg[33]/P0001  & n2197 ;
  assign n2270 = \u3_u0_r1_reg[33]/P0001  & n2200 ;
  assign n2271 = ~n2269 & ~n2270 ;
  assign n2272 = \u3_u0_r3_reg[33]/P0001  & n2205 ;
  assign n2273 = \u3_u0_r2_reg[33]/P0001  & n2208 ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = n2271 & n2274 ;
  assign n2276 = \u3_u0_r0_reg[10]/P0001  & n2197 ;
  assign n2277 = \u3_u0_r1_reg[10]/P0001  & n2200 ;
  assign n2278 = ~n2276 & ~n2277 ;
  assign n2279 = \u3_u0_r3_reg[10]/P0001  & n2205 ;
  assign n2280 = \u3_u0_r2_reg[10]/P0001  & n2208 ;
  assign n2281 = ~n2279 & ~n2280 ;
  assign n2282 = n2278 & n2281 ;
  assign n2283 = n2275 & ~n2282 ;
  assign n2284 = ~n2275 & n2282 ;
  assign n2285 = ~n2283 & ~n2284 ;
  assign n2286 = n2268 & n2285 ;
  assign n2287 = ~n2268 & ~n2285 ;
  assign n2288 = ~n2286 & ~n2287 ;
  assign n2289 = n2251 & ~n2288 ;
  assign n2290 = \wb_sel_i[1]_pad  & ~n2221 ;
  assign n2291 = n2248 & n2290 ;
  assign n2292 = \wb_sel_i[1]_pad  & ~n2288 ;
  assign n2293 = \wb_sel_i[1]_pad  & n2221 ;
  assign n2294 = ~n2248 & n2293 ;
  assign n2295 = ~n2292 & ~n2294 ;
  assign n2296 = ~n2291 & n2295 ;
  assign n2297 = ~n2289 & ~n2296 ;
  assign n2298 = \u3_u0_r0_reg[30]/P0001  & n2197 ;
  assign n2299 = \u3_u0_r1_reg[30]/P0001  & n2200 ;
  assign n2300 = ~n2298 & ~n2299 ;
  assign n2301 = \u3_u0_r3_reg[30]/P0001  & n2205 ;
  assign n2302 = \u3_u0_r2_reg[30]/P0001  & n2208 ;
  assign n2303 = ~n2301 & ~n2302 ;
  assign n2304 = n2300 & n2303 ;
  assign n2305 = \u3_u0_r3_reg[29]/P0001  & n2205 ;
  assign n2306 = \u3_u0_r2_reg[29]/P0001  & n2208 ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2308 = \u3_u0_r1_reg[29]/P0001  & n2200 ;
  assign n2309 = \u3_u0_r0_reg[29]/P0001  & n2197 ;
  assign n2310 = ~n2308 & ~n2309 ;
  assign n2311 = n2307 & n2310 ;
  assign n2312 = n2304 & ~n2311 ;
  assign n2313 = ~n2304 & n2311 ;
  assign n2314 = ~n2312 & ~n2313 ;
  assign n2315 = \u3_u0_r0_reg[27]/P0001  & n2197 ;
  assign n2316 = \u3_u0_r3_reg[27]/P0001  & n2205 ;
  assign n2317 = ~n2315 & ~n2316 ;
  assign n2318 = \u3_u0_r1_reg[27]/P0001  & n2200 ;
  assign n2319 = \u3_u0_r2_reg[27]/P0001  & n2208 ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2321 = n2317 & n2320 ;
  assign n2322 = \u3_u0_r0_reg[25]/P0001  & n2197 ;
  assign n2323 = \u3_u0_r1_reg[25]/P0001  & n2200 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = \u3_u0_r3_reg[25]/P0001  & n2205 ;
  assign n2326 = \u3_u0_r2_reg[25]/P0001  & n2208 ;
  assign n2327 = ~n2325 & ~n2326 ;
  assign n2328 = n2324 & n2327 ;
  assign n2329 = \u3_u0_r0_reg[28]/P0001  & n2197 ;
  assign n2330 = \u3_u0_r1_reg[28]/P0001  & n2200 ;
  assign n2331 = ~n2329 & ~n2330 ;
  assign n2332 = \u3_u0_r3_reg[28]/P0001  & n2205 ;
  assign n2333 = \u3_u0_r2_reg[28]/P0001  & n2208 ;
  assign n2334 = ~n2332 & ~n2333 ;
  assign n2335 = n2331 & n2334 ;
  assign n2336 = ~n2328 & ~n2335 ;
  assign n2337 = n2328 & n2335 ;
  assign n2338 = ~n2336 & ~n2337 ;
  assign n2339 = n2321 & ~n2338 ;
  assign n2340 = ~n2321 & n2338 ;
  assign n2341 = ~n2339 & ~n2340 ;
  assign n2342 = n2314 & n2341 ;
  assign n2343 = ~n2314 & ~n2341 ;
  assign n2344 = ~n2342 & ~n2343 ;
  assign n2345 = \u3_u0_r0_reg[24]/P0001  & n2197 ;
  assign n2346 = \u3_u0_r2_reg[24]/P0001  & n2208 ;
  assign n2347 = ~n2345 & ~n2346 ;
  assign n2348 = \u3_u0_r1_reg[24]/P0001  & n2200 ;
  assign n2349 = \u3_u0_r3_reg[24]/P0001  & n2205 ;
  assign n2350 = ~n2348 & ~n2349 ;
  assign n2351 = n2347 & n2350 ;
  assign n2352 = \u3_u0_r0_reg[31]/P0001  & n2197 ;
  assign n2353 = \u3_u0_r1_reg[31]/P0001  & n2200 ;
  assign n2354 = ~n2352 & ~n2353 ;
  assign n2355 = \u3_u0_r3_reg[31]/P0001  & n2205 ;
  assign n2356 = \u3_u0_r2_reg[31]/P0001  & n2208 ;
  assign n2357 = ~n2355 & ~n2356 ;
  assign n2358 = n2354 & n2357 ;
  assign n2359 = n2351 & ~n2358 ;
  assign n2360 = ~n2351 & n2358 ;
  assign n2361 = ~n2359 & ~n2360 ;
  assign n2362 = \u3_u0_r1_reg[35]/P0001  & n2200 ;
  assign n2363 = \u3_u0_r3_reg[35]/P0001  & n2205 ;
  assign n2364 = ~n2362 & ~n2363 ;
  assign n2365 = \u3_u0_r0_reg[35]/P0001  & n2197 ;
  assign n2366 = \u3_u0_r2_reg[35]/P0001  & n2208 ;
  assign n2367 = ~n2365 & ~n2366 ;
  assign n2368 = n2364 & n2367 ;
  assign n2369 = \u3_u0_r0_reg[26]/P0001  & n2197 ;
  assign n2370 = \u3_u0_r1_reg[26]/P0001  & n2200 ;
  assign n2371 = ~n2369 & ~n2370 ;
  assign n2372 = \u3_u0_r3_reg[26]/P0001  & n2205 ;
  assign n2373 = \u3_u0_r2_reg[26]/P0001  & n2208 ;
  assign n2374 = ~n2372 & ~n2373 ;
  assign n2375 = n2371 & n2374 ;
  assign n2376 = n2368 & ~n2375 ;
  assign n2377 = ~n2368 & n2375 ;
  assign n2378 = ~n2376 & ~n2377 ;
  assign n2379 = n2361 & n2378 ;
  assign n2380 = ~n2361 & ~n2378 ;
  assign n2381 = ~n2379 & ~n2380 ;
  assign n2382 = n2344 & ~n2381 ;
  assign n2383 = \wb_sel_i[3]_pad  & ~n2314 ;
  assign n2384 = n2341 & n2383 ;
  assign n2385 = \wb_sel_i[3]_pad  & ~n2381 ;
  assign n2386 = \wb_sel_i[3]_pad  & n2314 ;
  assign n2387 = ~n2341 & n2386 ;
  assign n2388 = ~n2385 & ~n2387 ;
  assign n2389 = ~n2384 & n2388 ;
  assign n2390 = ~n2382 & ~n2389 ;
  assign n2391 = ~n2297 & ~n2390 ;
  assign n2392 = \u3_u0_r1_reg[21]/P0001  & n2200 ;
  assign n2393 = \u3_u0_r0_reg[21]/P0001  & n2197 ;
  assign n2394 = ~n2392 & ~n2393 ;
  assign n2395 = \u3_u0_r2_reg[21]/P0001  & n2208 ;
  assign n2396 = \u3_u0_r3_reg[21]/P0001  & n2205 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = n2394 & n2397 ;
  assign n2399 = \u3_u0_r0_reg[17]/P0001  & n2197 ;
  assign n2400 = \u3_u0_r1_reg[17]/P0001  & n2200 ;
  assign n2401 = ~n2399 & ~n2400 ;
  assign n2402 = \u3_u0_r3_reg[17]/P0001  & n2205 ;
  assign n2403 = \u3_u0_r2_reg[17]/P0001  & n2208 ;
  assign n2404 = ~n2402 & ~n2403 ;
  assign n2405 = n2401 & n2404 ;
  assign n2406 = n2398 & ~n2405 ;
  assign n2407 = ~n2398 & n2405 ;
  assign n2408 = ~n2406 & ~n2407 ;
  assign n2409 = \u3_u0_r0_reg[22]/P0001  & n2197 ;
  assign n2410 = \u3_u0_r1_reg[22]/P0001  & n2200 ;
  assign n2411 = ~n2409 & ~n2410 ;
  assign n2412 = \u3_u0_r3_reg[22]/P0001  & n2205 ;
  assign n2413 = \u3_u0_r2_reg[22]/P0001  & n2208 ;
  assign n2414 = ~n2412 & ~n2413 ;
  assign n2415 = n2411 & n2414 ;
  assign n2416 = \u3_u0_r0_reg[19]/P0001  & n2197 ;
  assign n2417 = \u3_u0_r2_reg[19]/P0001  & n2208 ;
  assign n2418 = ~n2416 & ~n2417 ;
  assign n2419 = \u3_u0_r1_reg[19]/P0001  & n2200 ;
  assign n2420 = \u3_u0_r3_reg[19]/P0001  & n2205 ;
  assign n2421 = ~n2419 & ~n2420 ;
  assign n2422 = n2418 & n2421 ;
  assign n2423 = \u3_u0_r0_reg[20]/P0001  & n2197 ;
  assign n2424 = \u3_u0_r3_reg[20]/P0001  & n2205 ;
  assign n2425 = ~n2423 & ~n2424 ;
  assign n2426 = \u3_u0_r1_reg[20]/P0001  & n2200 ;
  assign n2427 = \u3_u0_r2_reg[20]/P0001  & n2208 ;
  assign n2428 = ~n2426 & ~n2427 ;
  assign n2429 = n2425 & n2428 ;
  assign n2430 = ~n2422 & ~n2429 ;
  assign n2431 = n2422 & n2429 ;
  assign n2432 = ~n2430 & ~n2431 ;
  assign n2433 = n2415 & ~n2432 ;
  assign n2434 = ~n2415 & n2432 ;
  assign n2435 = ~n2433 & ~n2434 ;
  assign n2436 = n2408 & n2435 ;
  assign n2437 = ~n2408 & ~n2435 ;
  assign n2438 = ~n2436 & ~n2437 ;
  assign n2439 = \u3_u0_r0_reg[16]/P0001  & n2197 ;
  assign n2440 = \u3_u0_r1_reg[16]/P0001  & n2200 ;
  assign n2441 = ~n2439 & ~n2440 ;
  assign n2442 = \u3_u0_r3_reg[16]/P0001  & n2205 ;
  assign n2443 = \u3_u0_r2_reg[16]/P0001  & n2208 ;
  assign n2444 = ~n2442 & ~n2443 ;
  assign n2445 = n2441 & n2444 ;
  assign n2446 = \u3_u0_r0_reg[23]/P0001  & n2197 ;
  assign n2447 = \u3_u0_r1_reg[23]/P0001  & n2200 ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2449 = \u3_u0_r3_reg[23]/P0001  & n2205 ;
  assign n2450 = \u3_u0_r2_reg[23]/P0001  & n2208 ;
  assign n2451 = ~n2449 & ~n2450 ;
  assign n2452 = n2448 & n2451 ;
  assign n2453 = n2445 & ~n2452 ;
  assign n2454 = ~n2445 & n2452 ;
  assign n2455 = ~n2453 & ~n2454 ;
  assign n2456 = \u3_u0_r0_reg[34]/P0001  & n2197 ;
  assign n2457 = \u3_u0_r1_reg[34]/P0001  & n2200 ;
  assign n2458 = ~n2456 & ~n2457 ;
  assign n2459 = \u3_u0_r3_reg[34]/P0001  & n2205 ;
  assign n2460 = \u3_u0_r2_reg[34]/P0001  & n2208 ;
  assign n2461 = ~n2459 & ~n2460 ;
  assign n2462 = n2458 & n2461 ;
  assign n2463 = \u3_u0_r0_reg[18]/P0001  & n2197 ;
  assign n2464 = \u3_u0_r1_reg[18]/P0001  & n2200 ;
  assign n2465 = ~n2463 & ~n2464 ;
  assign n2466 = \u3_u0_r3_reg[18]/P0001  & n2205 ;
  assign n2467 = \u3_u0_r2_reg[18]/P0001  & n2208 ;
  assign n2468 = ~n2466 & ~n2467 ;
  assign n2469 = n2465 & n2468 ;
  assign n2470 = n2462 & ~n2469 ;
  assign n2471 = ~n2462 & n2469 ;
  assign n2472 = ~n2470 & ~n2471 ;
  assign n2473 = n2455 & n2472 ;
  assign n2474 = ~n2455 & ~n2472 ;
  assign n2475 = ~n2473 & ~n2474 ;
  assign n2476 = n2438 & ~n2475 ;
  assign n2477 = \wb_sel_i[2]_pad  & ~n2408 ;
  assign n2478 = n2435 & n2477 ;
  assign n2479 = \wb_sel_i[2]_pad  & ~n2475 ;
  assign n2480 = \wb_sel_i[2]_pad  & n2408 ;
  assign n2481 = ~n2435 & n2480 ;
  assign n2482 = ~n2479 & ~n2481 ;
  assign n2483 = ~n2478 & n2482 ;
  assign n2484 = ~n2476 & ~n2483 ;
  assign n2485 = \u3_u0_r0_reg[0]/P0001  & n2197 ;
  assign n2486 = \u3_u0_r2_reg[0]/P0001  & n2208 ;
  assign n2487 = ~n2485 & ~n2486 ;
  assign n2488 = \u3_u0_r1_reg[0]/P0001  & n2200 ;
  assign n2489 = \u3_u0_r3_reg[0]/P0001  & n2205 ;
  assign n2490 = ~n2488 & ~n2489 ;
  assign n2491 = n2487 & n2490 ;
  assign n2492 = \u3_u0_r0_reg[2]/P0001  & n2197 ;
  assign n2493 = \u3_u0_r1_reg[2]/P0001  & n2200 ;
  assign n2494 = ~n2492 & ~n2493 ;
  assign n2495 = \u3_u0_r3_reg[2]/P0001  & n2205 ;
  assign n2496 = \u3_u0_r2_reg[2]/P0001  & n2208 ;
  assign n2497 = ~n2495 & ~n2496 ;
  assign n2498 = n2494 & n2497 ;
  assign n2499 = n2491 & ~n2498 ;
  assign n2500 = ~n2491 & n2498 ;
  assign n2501 = ~n2499 & ~n2500 ;
  assign n2502 = \u3_u0_r0_reg[4]/P0001  & n2197 ;
  assign n2503 = \u3_u0_r1_reg[4]/P0001  & n2200 ;
  assign n2504 = ~n2502 & ~n2503 ;
  assign n2505 = \u3_u0_r3_reg[4]/P0001  & n2205 ;
  assign n2506 = \u3_u0_r2_reg[4]/P0001  & n2208 ;
  assign n2507 = ~n2505 & ~n2506 ;
  assign n2508 = n2504 & n2507 ;
  assign n2509 = \u3_u0_r3_reg[7]/P0001  & n2205 ;
  assign n2510 = \u3_u0_r2_reg[7]/P0001  & n2208 ;
  assign n2511 = ~n2509 & ~n2510 ;
  assign n2512 = \u3_u0_r0_reg[7]/P0001  & n2197 ;
  assign n2513 = \u3_u0_r1_reg[7]/P0001  & n2200 ;
  assign n2514 = ~n2512 & ~n2513 ;
  assign n2515 = n2511 & n2514 ;
  assign n2516 = \u3_u0_r1_reg[6]/P0001  & n2200 ;
  assign n2517 = \u3_u0_r2_reg[6]/P0001  & n2208 ;
  assign n2518 = ~n2516 & ~n2517 ;
  assign n2519 = \u3_u0_r0_reg[6]/P0001  & n2197 ;
  assign n2520 = \u3_u0_r3_reg[6]/P0001  & n2205 ;
  assign n2521 = ~n2519 & ~n2520 ;
  assign n2522 = n2518 & n2521 ;
  assign n2523 = ~n2515 & ~n2522 ;
  assign n2524 = n2515 & n2522 ;
  assign n2525 = ~n2523 & ~n2524 ;
  assign n2526 = n2508 & ~n2525 ;
  assign n2527 = ~n2508 & n2525 ;
  assign n2528 = ~n2526 & ~n2527 ;
  assign n2529 = n2501 & n2528 ;
  assign n2530 = ~n2501 & ~n2528 ;
  assign n2531 = ~n2529 & ~n2530 ;
  assign n2532 = \u3_u0_r3_reg[5]/P0001  & n2205 ;
  assign n2533 = \u3_u0_r2_reg[5]/P0001  & n2208 ;
  assign n2534 = ~n2532 & ~n2533 ;
  assign n2535 = \u3_u0_r0_reg[5]/P0001  & n2197 ;
  assign n2536 = \u3_u0_r1_reg[5]/P0001  & n2200 ;
  assign n2537 = ~n2535 & ~n2536 ;
  assign n2538 = n2534 & n2537 ;
  assign n2539 = \u3_u0_r0_reg[3]/P0001  & n2197 ;
  assign n2540 = \u3_u0_r2_reg[3]/P0001  & n2208 ;
  assign n2541 = ~n2539 & ~n2540 ;
  assign n2542 = \u3_u0_r1_reg[3]/P0001  & n2200 ;
  assign n2543 = \u3_u0_r3_reg[3]/P0001  & n2205 ;
  assign n2544 = ~n2542 & ~n2543 ;
  assign n2545 = n2541 & n2544 ;
  assign n2546 = n2538 & ~n2545 ;
  assign n2547 = ~n2538 & n2545 ;
  assign n2548 = ~n2546 & ~n2547 ;
  assign n2549 = \u3_u0_r3_reg[32]/P0001  & n2205 ;
  assign n2550 = \u3_u0_r2_reg[32]/P0001  & n2208 ;
  assign n2551 = ~n2549 & ~n2550 ;
  assign n2552 = \u3_u0_r0_reg[32]/P0001  & n2197 ;
  assign n2553 = \u3_u0_r1_reg[32]/P0001  & n2200 ;
  assign n2554 = ~n2552 & ~n2553 ;
  assign n2555 = n2551 & n2554 ;
  assign n2556 = \u3_u0_r0_reg[1]/P0001  & n2197 ;
  assign n2557 = \u3_u0_r1_reg[1]/P0001  & n2200 ;
  assign n2558 = ~n2556 & ~n2557 ;
  assign n2559 = \u3_u0_r3_reg[1]/P0001  & n2205 ;
  assign n2560 = \u3_u0_r2_reg[1]/P0001  & n2208 ;
  assign n2561 = ~n2559 & ~n2560 ;
  assign n2562 = n2558 & n2561 ;
  assign n2563 = n2555 & ~n2562 ;
  assign n2564 = ~n2555 & n2562 ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = n2548 & n2565 ;
  assign n2567 = ~n2548 & ~n2565 ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = n2531 & ~n2568 ;
  assign n2570 = \wb_sel_i[0]_pad  & ~n2501 ;
  assign n2571 = n2528 & n2570 ;
  assign n2572 = \wb_sel_i[0]_pad  & ~n2568 ;
  assign n2573 = \wb_sel_i[0]_pad  & n2501 ;
  assign n2574 = ~n2528 & n2573 ;
  assign n2575 = ~n2572 & ~n2574 ;
  assign n2576 = ~n2571 & n2575 ;
  assign n2577 = ~n2569 & ~n2576 ;
  assign n2578 = ~n2484 & ~n2577 ;
  assign n2579 = n2391 & n2578 ;
  assign n2580 = \u0_csc_reg[11]/NET0131  & ~wb_we_i_pad ;
  assign n2581 = ~n1898 & n2580 ;
  assign n2582 = ~n2189 & n2581 ;
  assign n2583 = ~n2579 & n2582 ;
  assign n2584 = ~\u0_wp_err_reg/NET0131  & ~\u5_state_reg[65]/NET0131  ;
  assign n2585 = n2193 & n2584 ;
  assign n2586 = ~n2583 & n2585 ;
  assign n2587 = ~n2194 & ~n2586 ;
  assign n2588 = \wb_addr_i[29]_pad  & \wb_addr_i[30]_pad  ;
  assign n2589 = ~\wb_addr_i[31]_pad  & n2588 ;
  assign n2590 = ~wb_ack_o_pad & n1045 ;
  assign n2591 = n2589 & n2590 ;
  assign n2592 = n2587 & ~n2591 ;
  assign n2593 = n1947 & n1978 ;
  assign n2594 = n1851 & n2122 ;
  assign n2595 = ~n1848 & n2594 ;
  assign n2596 = ~n2030 & ~n2595 ;
  assign n2597 = \u0_tms_reg[11]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2598 = ~\u5_lmr_ack_reg/NET0131  & n2597 ;
  assign n2599 = n983 & n2598 ;
  assign n2600 = \u0_sp_tms_reg[11]/NET0131  & ~n1200 ;
  assign n2601 = ~n2599 & ~n2600 ;
  assign n2602 = n1851 & n2601 ;
  assign n2603 = ~n1848 & n2602 ;
  assign n2604 = ~n2043 & n2603 ;
  assign n2605 = n2030 & ~n2604 ;
  assign n2606 = ~n2596 & ~n2605 ;
  assign n2607 = \u0_tms_reg[23]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2608 = ~\u5_lmr_ack_reg/NET0131  & n2607 ;
  assign n2609 = n983 & n2608 ;
  assign n2610 = \u0_sp_tms_reg[23]/NET0131  & ~n1200 ;
  assign n2611 = ~n2609 & ~n2610 ;
  assign n2612 = n1851 & n2611 ;
  assign n2613 = ~n1848 & n2612 ;
  assign n2614 = ~n1938 & ~n2613 ;
  assign n2615 = n2063 & n2072 ;
  assign n2616 = ~\u5_state_reg[35]/NET0131  & n985 ;
  assign n2617 = n2062 & n2616 ;
  assign n2618 = n2615 & n2617 ;
  assign n2619 = ~\u5_timer_reg[2]/NET0131  & n2072 ;
  assign n2620 = \u5_timer_reg[3]/NET0131  & n2617 ;
  assign n2621 = ~n2619 & n2620 ;
  assign n2622 = ~n2618 & ~n2621 ;
  assign n2623 = \u0_sp_tms_reg[27]/NET0131  & ~n1200 ;
  assign n2624 = \u0_tms_reg[27]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2625 = ~\u5_lmr_ack_reg/NET0131  & n2624 ;
  assign n2626 = n983 & n2625 ;
  assign n2627 = ~n2623 & ~n2626 ;
  assign n2628 = n1851 & n2627 ;
  assign n2629 = ~n1848 & n2628 ;
  assign n2630 = ~n2062 & ~n2629 ;
  assign n2631 = n2622 & ~n2630 ;
  assign n2632 = ~\u5_state_reg[9]/NET0131  & n2098 ;
  assign n2633 = ~n1934 & n2632 ;
  assign n2634 = n1938 & n2633 ;
  assign n2635 = ~n2631 & n2634 ;
  assign n2636 = ~n2614 & ~n2635 ;
  assign n2637 = n2052 & ~n2636 ;
  assign n2638 = ~n2096 & ~n2613 ;
  assign n2639 = ~n2132 & n2638 ;
  assign n2640 = ~n2098 & ~n2639 ;
  assign n2641 = n2096 & n2613 ;
  assign n2642 = n2114 & n2613 ;
  assign n2643 = ~n2131 & n2642 ;
  assign n2644 = ~n2641 & ~n2643 ;
  assign n2645 = n2052 & n2644 ;
  assign n2646 = n2640 & n2645 ;
  assign n2647 = ~n2637 & ~n2646 ;
  assign n2648 = \u0_tms_reg[3]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2649 = ~\u5_lmr_ack_reg/NET0131  & n2648 ;
  assign n2650 = n983 & n2649 ;
  assign n2651 = \u0_sp_tms_reg[3]/NET0131  & ~n1200 ;
  assign n2652 = ~n2650 & ~n2651 ;
  assign n2653 = n1851 & n2652 ;
  assign n2654 = ~n1848 & n2653 ;
  assign n2655 = ~n2052 & ~n2654 ;
  assign n2656 = n2043 & ~n2655 ;
  assign n2657 = ~n2596 & n2656 ;
  assign n2658 = n2647 & n2657 ;
  assign n2659 = ~n2606 & ~n2658 ;
  assign n2660 = \u5_state_reg[16]/NET0131  & ~n1974 ;
  assign n2661 = ~n1972 & n2660 ;
  assign n2662 = n1245 & n2661 ;
  assign n2663 = ~\u5_wb_cycle_reg/NET0131  & ~n1205 ;
  assign n2664 = ~\u5_wb_cycle_reg/NET0131  & n1227 ;
  assign n2665 = n1222 & n2664 ;
  assign n2666 = ~n2663 & ~n2665 ;
  assign n2667 = ~\u5_wb_write_go_r_reg/NET0131  & \u6_read_go_r1_reg/NET0131  ;
  assign n2668 = n1234 & n2667 ;
  assign n2669 = ~n1048 & n2668 ;
  assign n2670 = \u5_state_reg[16]/NET0131  & ~n2669 ;
  assign n2671 = ~n1966 & n2670 ;
  assign n2672 = ~n1954 & n2671 ;
  assign n2673 = n2666 & n2672 ;
  assign n2674 = ~n1954 & ~n1966 ;
  assign n2675 = ~\u5_ap_en_reg/NET0131  & n2666 ;
  assign n2676 = ~n2674 & n2675 ;
  assign n2677 = ~n2673 & ~n2676 ;
  assign n2678 = ~n1969 & ~n1975 ;
  assign n2679 = n1245 & n2678 ;
  assign n2680 = ~n2677 & n2679 ;
  assign n2681 = ~n2662 & ~n2680 ;
  assign n2682 = n1956 & ~n1966 ;
  assign n2683 = ~n1954 & n2682 ;
  assign n2684 = ~n1895 & ~n2683 ;
  assign n2685 = ~\u5_ap_en_reg/NET0131  & \u5_cmd_asserted_reg/NET0131  ;
  assign n2686 = n1249 & n2685 ;
  assign n2687 = n1248 & n2686 ;
  assign n2688 = ~\u5_wb_cycle_reg/NET0131  & n2687 ;
  assign n2689 = ~n1966 & n2687 ;
  assign n2690 = ~n1954 & n2689 ;
  assign n2691 = ~n2688 & ~n2690 ;
  assign n2692 = n2684 & ~n2691 ;
  assign n2693 = \u5_mem_ack_r_reg/NET0131  & \u5_state_reg[16]/NET0131  ;
  assign n2694 = \u5_state_reg[16]/NET0131  & n1233 ;
  assign n2695 = ~n1898 & n2694 ;
  assign n2696 = ~n2693 & ~n2695 ;
  assign n2697 = ~\u5_ap_en_reg/NET0131  & ~n1209 ;
  assign n2698 = ~n1206 & n2697 ;
  assign n2699 = n2696 & ~n2698 ;
  assign n2700 = ~n1895 & ~n2168 ;
  assign n2701 = n1412 & ~n2700 ;
  assign n2702 = n1248 & n2701 ;
  assign n2703 = ~n2699 & n2702 ;
  assign n2704 = \u5_cmd_asserted_reg/NET0131  & n1269 ;
  assign n2705 = \u5_tmr_done_reg/NET0131  & n1209 ;
  assign n2706 = \u0_sp_csc_reg[10]/NET0131  & \u5_tmr_done_reg/NET0131  ;
  assign n2707 = ~n1200 & n2706 ;
  assign n2708 = ~n2705 & ~n2707 ;
  assign n2709 = \u5_cmd_asserted_reg/NET0131  & \u5_tmr_done_reg/NET0131  ;
  assign n2710 = ~n1209 & n2709 ;
  assign n2711 = ~n1206 & n2710 ;
  assign n2712 = \u5_state_reg[16]/NET0131  & ~n2711 ;
  assign n2713 = n2708 & n2712 ;
  assign n2714 = n1443 & n2713 ;
  assign n2715 = ~n2704 & ~n2714 ;
  assign n2716 = ~n2703 & n2715 ;
  assign n2717 = ~n2692 & n2716 ;
  assign n2718 = n2681 & n2717 ;
  assign n2719 = \u0_sp_csc_reg[7]/NET0131  & ~n1200 ;
  assign n2720 = \u0_csc_reg[7]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2721 = ~\u5_lmr_ack_reg/NET0131  & n2720 ;
  assign n2722 = n983 & n2721 ;
  assign n2723 = ~n2719 & ~n2722 ;
  assign n2724 = \u0_sp_csc_reg[6]/NET0131  & ~n1200 ;
  assign n2725 = \u0_csc_reg[6]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2726 = ~\u5_lmr_ack_reg/NET0131  & n2725 ;
  assign n2727 = n983 & n2726 ;
  assign n2728 = ~n2724 & ~n2727 ;
  assign n2729 = n2723 & n2728 ;
  assign n2730 = \u0_sp_csc_reg[4]/NET0131  & ~n1200 ;
  assign n2731 = \u0_csc_reg[4]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2732 = ~\u5_lmr_ack_reg/NET0131  & n2731 ;
  assign n2733 = n983 & n2732 ;
  assign n2734 = ~n2730 & ~n2733 ;
  assign n2735 = n2729 & ~n2734 ;
  assign n2736 = \u0_sp_csc_reg[5]/NET0131  & ~n1200 ;
  assign n2737 = \u0_csc_reg[5]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2738 = ~\u5_lmr_ack_reg/NET0131  & n2737 ;
  assign n2739 = n983 & n2738 ;
  assign n2740 = ~n2736 & ~n2739 ;
  assign n2741 = ~n2735 & n2740 ;
  assign n2742 = \u5_state_reg[1]/NET0131  & ~n2741 ;
  assign n2743 = ~n2054 & n2742 ;
  assign n2744 = \u5_wr_cycle_reg/NET0131  & n2185 ;
  assign n2745 = n2164 & n2744 ;
  assign n2746 = ~n2157 & n2745 ;
  assign n2747 = ~n2152 & n2746 ;
  assign n2748 = n1962 & n1963 ;
  assign n2749 = ~\u5_wr_cycle_reg/NET0131  & n1043 ;
  assign n2750 = n2748 & ~n2749 ;
  assign n2751 = ~n2747 & n2750 ;
  assign n2752 = ~\u5_state_reg[1]/NET0131  & n2751 ;
  assign n2753 = ~\u5_burst_cnt_reg[7]/NET0131  & n1962 ;
  assign n2754 = ~n2749 & n2753 ;
  assign n2755 = ~n2747 & n2754 ;
  assign n2756 = \u5_burst_cnt_reg[8]/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n2757 = ~n2755 & n2756 ;
  assign n2758 = ~n2752 & ~n2757 ;
  assign n2759 = ~n2743 & n2758 ;
  assign n2760 = ~\u5_state_reg[52]/NET0131  & ~n2759 ;
  assign n2761 = n1966 & ~n2749 ;
  assign n2762 = ~n2747 & n2761 ;
  assign n2763 = ~\u5_state_reg[1]/NET0131  & n2762 ;
  assign n2764 = ~\u5_burst_cnt_reg[9]/NET0131  & n2748 ;
  assign n2765 = ~n2749 & n2764 ;
  assign n2766 = ~n2747 & n2765 ;
  assign n2767 = \u5_burst_cnt_reg[10]/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n2768 = ~n2766 & n2767 ;
  assign n2769 = ~n2763 & ~n2768 ;
  assign n2770 = n2734 & n2740 ;
  assign n2771 = ~n2729 & n2770 ;
  assign n2772 = \u5_state_reg[1]/NET0131  & n2771 ;
  assign n2773 = ~n2054 & n2772 ;
  assign n2774 = n2769 & ~n2773 ;
  assign n2775 = ~\u5_state_reg[52]/NET0131  & ~n2774 ;
  assign n2776 = \u5_state_reg[1]/NET0131  & n1227 ;
  assign n2777 = n1851 & n2776 ;
  assign n2778 = ~n1848 & n2777 ;
  assign n2779 = n1222 & n2778 ;
  assign n2780 = ~\u5_state_reg[52]/NET0131  & n2779 ;
  assign n2781 = ~\u5_burst_cnt_reg[0]/NET0131  & ~n2749 ;
  assign n2782 = ~n2747 & n2781 ;
  assign n2783 = \u5_burst_cnt_reg[0]/NET0131  & n2749 ;
  assign n2784 = \u5_burst_cnt_reg[0]/NET0131  & ~n2152 ;
  assign n2785 = n2746 & n2784 ;
  assign n2786 = ~n2783 & ~n2785 ;
  assign n2787 = ~n2782 & n2786 ;
  assign n2788 = ~\u5_state_reg[1]/NET0131  & ~\u5_state_reg[52]/NET0131  ;
  assign n2789 = ~n2787 & n2788 ;
  assign n2790 = ~n2780 & ~n2789 ;
  assign n2791 = ~\u5_state_reg[17]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n2792 = ~\u5_rfr_ack_r_reg/NET0131  & \u5_tmr_done_reg/NET0131  ;
  assign n2793 = n1304 & ~n2792 ;
  assign n2794 = n1032 & n2793 ;
  assign n2795 = ~n1285 & ~n2794 ;
  assign n2796 = ~n2791 & ~n2795 ;
  assign n2797 = ~\u5_cmd_asserted_reg/NET0131  & n1180 ;
  assign n2798 = ~n2796 & ~n2797 ;
  assign n2799 = ~n2583 & n2584 ;
  assign n2800 = ~\wb_addr_i[31]_pad  & ~wb_err_o_pad ;
  assign n2801 = n2190 & n2800 ;
  assign n2802 = n1045 & n2801 ;
  assign n2803 = ~n2799 & n2802 ;
  assign n2804 = \u5_lookup_ready2_reg/NET0131  & ~n1899 ;
  assign n2805 = n1538 & ~n2804 ;
  assign n2806 = n1526 & n1537 ;
  assign n2807 = n1531 & ~n2806 ;
  assign n2808 = n1899 & n2807 ;
  assign n2809 = ~n2805 & ~n2808 ;
  assign n2810 = n1922 & n2809 ;
  assign n2811 = ~\u5_cmd_asserted2_reg/NET0131  & \u7_mc_br_r_reg/P0001  ;
  assign n2812 = ~n1922 & n2811 ;
  assign n2813 = n1929 & ~n2812 ;
  assign n2814 = ~n2810 & n2813 ;
  assign n2815 = n1443 & ~n2708 ;
  assign n2816 = ~\u5_state_reg[1]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n2817 = ~n1339 & ~n1438 ;
  assign n2818 = ~n2816 & ~n2817 ;
  assign n2819 = \u5_wb_cycle_reg/NET0131  & n1233 ;
  assign n2820 = ~n1898 & n2819 ;
  assign n2821 = ~\u5_cs_le_r_reg/P0001  & \u5_wb_cycle_reg/NET0131  ;
  assign n2822 = ~\u5_state_reg[1]/NET0131  & n2821 ;
  assign n2823 = \u5_tmr2_done_reg/NET0131  & ~n2822 ;
  assign n2824 = ~n2820 & n2823 ;
  assign n2825 = n1281 & n2824 ;
  assign n2826 = ~n1167 & ~n2825 ;
  assign n2827 = ~n2818 & n2826 ;
  assign n2828 = ~n2815 & n2827 ;
  assign n2829 = ~n2814 & n2828 ;
  assign n2830 = n1958 & ~n2749 ;
  assign n2831 = ~n2747 & n2830 ;
  assign n2832 = ~\u5_state_reg[1]/NET0131  & n2831 ;
  assign n2833 = n1957 & ~n2749 ;
  assign n2834 = ~n2747 & n2833 ;
  assign n2835 = \u5_burst_cnt_reg[2]/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n2836 = ~n2834 & n2835 ;
  assign n2837 = ~n2832 & ~n2836 ;
  assign n2838 = ~n1216 & n1221 ;
  assign n2839 = n1851 & n2838 ;
  assign n2840 = ~n1848 & n2839 ;
  assign n2841 = n2778 & n2840 ;
  assign n2842 = ~\u5_state_reg[52]/NET0131  & ~n2841 ;
  assign n2843 = n2837 & n2842 ;
  assign n2844 = \u5_burst_cnt_reg[9]/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n2845 = ~n2751 & n2844 ;
  assign n2846 = ~\u5_burst_cnt_reg[9]/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n2847 = n2751 & n2846 ;
  assign n2848 = ~n2845 & ~n2847 ;
  assign n2849 = n2729 & ~n2770 ;
  assign n2850 = ~n2729 & n2734 ;
  assign n2851 = ~n2849 & ~n2850 ;
  assign n2852 = \u5_state_reg[1]/NET0131  & n2851 ;
  assign n2853 = ~n2054 & n2852 ;
  assign n2854 = n2848 & ~n2853 ;
  assign n2855 = ~\u5_state_reg[52]/NET0131  & ~n2854 ;
  assign n2856 = \u5_wb_cycle_reg/NET0131  & ~\u5_wr_cycle_reg/NET0131  ;
  assign n2857 = ~\u5_data_oe_reg/NET0131  & ~n2856 ;
  assign n2858 = \u5_data_oe_reg/NET0131  & ~\u7_mc_dqm_r2_reg[0]/P0001  ;
  assign n2859 = ~\u5_susp_sel_r_reg/NET0131  & ~n2858 ;
  assign n2860 = ~n2857 & n2859 ;
  assign n2861 = \u5_data_oe_reg/NET0131  & ~\u7_mc_dqm_r2_reg[1]/P0001  ;
  assign n2862 = ~\u5_susp_sel_r_reg/NET0131  & ~n2861 ;
  assign n2863 = ~n2857 & n2862 ;
  assign n2864 = \u5_data_oe_reg/NET0131  & ~\u7_mc_dqm_r2_reg[2]/P0001  ;
  assign n2865 = ~\u5_susp_sel_r_reg/NET0131  & ~n2864 ;
  assign n2866 = ~n2857 & n2865 ;
  assign n2867 = \u5_data_oe_reg/NET0131  & ~\u7_mc_dqm_r2_reg[3]/P0001  ;
  assign n2868 = ~\u5_susp_sel_r_reg/NET0131  & ~n2867 ;
  assign n2869 = ~n2857 & n2868 ;
  assign n2870 = \u5_state_reg[2]/NET0131  & ~n1974 ;
  assign n2871 = ~n1972 & n2870 ;
  assign n2872 = ~n1975 & ~n2666 ;
  assign n2873 = ~n2871 & ~n2872 ;
  assign n2874 = n1245 & ~n2873 ;
  assign n2875 = ~\u5_ap_en_reg/NET0131  & ~n2674 ;
  assign n2876 = ~\u5_state_reg[2]/NET0131  & ~n2669 ;
  assign n2877 = ~n1966 & n2876 ;
  assign n2878 = ~n1954 & n2877 ;
  assign n2879 = ~n2875 & ~n2878 ;
  assign n2880 = n2679 & n2879 ;
  assign n2881 = ~n2874 & ~n2880 ;
  assign n2882 = n1248 & n2146 ;
  assign n2883 = \u5_wb_cycle_reg/NET0131  & ~n2674 ;
  assign n2884 = \u5_ap_en_reg/NET0131  & ~n1895 ;
  assign n2885 = ~n2683 & n2884 ;
  assign n2886 = ~n2883 & ~n2885 ;
  assign n2887 = n2882 & ~n2886 ;
  assign n2888 = \u5_mem_ack_r_reg/NET0131  & ~\u5_state_reg[2]/NET0131  ;
  assign n2889 = ~\u5_state_reg[2]/NET0131  & n1233 ;
  assign n2890 = ~n1898 & n2889 ;
  assign n2891 = ~n2888 & ~n2890 ;
  assign n2892 = ~n2698 & n2891 ;
  assign n2893 = n2702 & n2892 ;
  assign n2894 = ~n1404 & ~n2009 ;
  assign n2895 = ~\u5_state_reg[2]/NET0131  & \u7_mc_br_r_reg/P0001  ;
  assign n2896 = n1411 & ~n2895 ;
  assign n2897 = ~\u5_state_reg[2]/NET0131  & ~n2711 ;
  assign n2898 = n2708 & ~n2897 ;
  assign n2899 = n1443 & n2898 ;
  assign n2900 = ~n2896 & ~n2899 ;
  assign n2901 = n2894 & n2900 ;
  assign n2902 = ~n2893 & n2901 ;
  assign n2903 = ~\u5_tmr_done_reg/NET0131  & ~n1504 ;
  assign n2904 = n1940 & ~n2903 ;
  assign n2905 = \u5_state_reg[2]/NET0131  & ~n2904 ;
  assign n2906 = ~n1180 & ~n1265 ;
  assign n2907 = ~n1317 & n2906 ;
  assign n2908 = \u5_cmd_asserted_reg/NET0131  & ~n2907 ;
  assign n2909 = ~n2905 & ~n2908 ;
  assign n2910 = n2902 & n2909 ;
  assign n2911 = ~n2887 & n2910 ;
  assign n2912 = n2881 & n2911 ;
  assign n2913 = n1314 & ~n1904 ;
  assign n2914 = \u5_state_reg[57]/NET0131  & n1233 ;
  assign n2915 = n1896 & ~n2914 ;
  assign n2916 = ~n1048 & n2915 ;
  assign n2917 = n1142 & ~n2916 ;
  assign n2918 = n1015 & n2917 ;
  assign n2919 = ~n2913 & ~n2918 ;
  assign n2920 = ~\u5_state_reg[57]/NET0131  & n1234 ;
  assign n2921 = n1232 & n2920 ;
  assign n2922 = ~n1048 & n2921 ;
  assign n2923 = ~n1899 & ~n2922 ;
  assign n2924 = n2180 & n2923 ;
  assign n2925 = \u5_state_reg[57]/NET0131  & ~n2168 ;
  assign n2926 = n1897 & ~n2925 ;
  assign n2927 = n1400 & ~n2926 ;
  assign n2928 = ~n2924 & ~n2927 ;
  assign n2929 = n2919 & n2928 ;
  assign n2930 = ~n1314 & ~n2180 ;
  assign n2931 = n1899 & ~n2930 ;
  assign n2932 = \u5_state_reg[59]/NET0131  & n1234 ;
  assign n2933 = n1232 & n2932 ;
  assign n2934 = ~n1048 & n2933 ;
  assign n2935 = n2180 & n2934 ;
  assign n2936 = ~n2931 & ~n2935 ;
  assign n2937 = n1227 & n1851 ;
  assign n2938 = ~n1848 & n2937 ;
  assign n2939 = ~n2052 & ~n2938 ;
  assign n2940 = n2043 & n2939 ;
  assign n2941 = ~\u0_tms_reg[24]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2942 = ~\u5_lmr_ack_reg/NET0131  & n2941 ;
  assign n2943 = n983 & n2942 ;
  assign n2944 = ~\u0_sp_tms_reg[24]/NET0131  & ~n1200 ;
  assign n2945 = ~n2943 & ~n2944 ;
  assign n2946 = ~n2062 & ~n2945 ;
  assign n2947 = n1851 & n2946 ;
  assign n2948 = ~n1848 & n2947 ;
  assign n2949 = ~\u5_mc_le_reg/NET0131  & ~n2069 ;
  assign n2950 = \u5_timer_reg[0]/NET0131  & ~n2949 ;
  assign n2951 = ~\u5_mc_le_reg/NET0131  & ~\u5_timer_reg[0]/NET0131  ;
  assign n2952 = ~n2069 & n2951 ;
  assign n2953 = n2617 & ~n2952 ;
  assign n2954 = ~n2950 & n2953 ;
  assign n2955 = ~n2948 & ~n2954 ;
  assign n2956 = ~\u5_state_reg[9]/NET0131  & ~n2955 ;
  assign n2957 = \u0_tms_reg[4]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2958 = ~\u5_lmr_ack_reg/NET0131  & n2957 ;
  assign n2959 = n983 & n2958 ;
  assign n2960 = \u0_sp_tms_reg[4]/NET0131  & ~n1200 ;
  assign n2961 = ~n2959 & ~n2960 ;
  assign n2962 = \u5_state_reg[9]/NET0131  & n2961 ;
  assign n2963 = n1851 & n2962 ;
  assign n2964 = ~n1848 & n2963 ;
  assign n2965 = n1939 & ~n2964 ;
  assign n2966 = ~n2956 & n2965 ;
  assign n2967 = n1851 & n2127 ;
  assign n2968 = ~n1848 & n2967 ;
  assign n2969 = ~n1938 & ~n2968 ;
  assign n2970 = n1851 & n1869 ;
  assign n2971 = ~n1848 & n2970 ;
  assign n2972 = n2101 & ~n2971 ;
  assign n2973 = n2098 & ~n2972 ;
  assign n2974 = ~n2969 & n2973 ;
  assign n2975 = ~n2966 & n2974 ;
  assign n2976 = n2122 & n2127 ;
  assign n2977 = n1851 & n2976 ;
  assign n2978 = ~n1848 & n2977 ;
  assign n2979 = n2130 & ~n2978 ;
  assign n2980 = ~n2098 & ~n2979 ;
  assign n2981 = n2052 & ~n2980 ;
  assign n2982 = n2043 & n2981 ;
  assign n2983 = ~n2975 & n2982 ;
  assign n2984 = ~n2940 & ~n2983 ;
  assign n2985 = \u0_tms_reg[8]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2986 = ~\u5_lmr_ack_reg/NET0131  & n2985 ;
  assign n2987 = n983 & n2986 ;
  assign n2988 = \u0_sp_tms_reg[8]/NET0131  & ~n1200 ;
  assign n2989 = ~n2987 & ~n2988 ;
  assign n2990 = n1851 & n2989 ;
  assign n2991 = ~n1848 & n2990 ;
  assign n2992 = ~n2043 & ~n2991 ;
  assign n2993 = n2984 & ~n2992 ;
  assign n2994 = n2030 & ~n2993 ;
  assign n2995 = \u0_tms_reg[12]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n2996 = ~\u5_lmr_ack_reg/NET0131  & n2995 ;
  assign n2997 = n983 & n2996 ;
  assign n2998 = \u0_sp_tms_reg[12]/NET0131  & ~n1200 ;
  assign n2999 = ~n2997 & ~n2998 ;
  assign n3000 = n1851 & n2999 ;
  assign n3001 = ~n1848 & n3000 ;
  assign n3002 = ~n2030 & ~n3001 ;
  assign n3003 = ~n2994 & ~n3002 ;
  assign n3004 = \u0_sp_tms_reg[13]/NET0131  & ~n1200 ;
  assign n3005 = \u0_tms_reg[13]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n3006 = ~\u5_lmr_ack_reg/NET0131  & n3005 ;
  assign n3007 = n983 & n3006 ;
  assign n3008 = ~n3004 & ~n3007 ;
  assign n3009 = ~n2030 & n3008 ;
  assign n3010 = ~n2031 & n3009 ;
  assign n3011 = n1216 & n1851 ;
  assign n3012 = ~n1848 & n3011 ;
  assign n3013 = ~n2052 & n3012 ;
  assign n3014 = n2043 & ~n3013 ;
  assign n3015 = ~n2052 & n3014 ;
  assign n3016 = ~\u0_tms_reg[25]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n3017 = ~\u5_lmr_ack_reg/NET0131  & n3016 ;
  assign n3018 = n983 & n3017 ;
  assign n3019 = ~\u0_sp_tms_reg[25]/NET0131  & ~n1200 ;
  assign n3020 = ~n3018 & ~n3019 ;
  assign n3021 = ~n2062 & ~n3020 ;
  assign n3022 = n1851 & n3021 ;
  assign n3023 = ~n1848 & n3022 ;
  assign n3024 = \u5_timer_reg[1]/NET0131  & ~n2952 ;
  assign n3025 = ~n2072 & n2617 ;
  assign n3026 = ~n3024 & n3025 ;
  assign n3027 = ~n3023 & ~n3026 ;
  assign n3028 = ~\u5_state_reg[9]/NET0131  & ~n3027 ;
  assign n3029 = \u0_tms_reg[5]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n3030 = ~\u5_lmr_ack_reg/NET0131  & n3029 ;
  assign n3031 = n983 & n3030 ;
  assign n3032 = \u0_sp_tms_reg[5]/NET0131  & ~n1200 ;
  assign n3033 = ~n3031 & ~n3032 ;
  assign n3034 = \u5_state_reg[9]/NET0131  & n3033 ;
  assign n3035 = n1851 & n3034 ;
  assign n3036 = ~n1848 & n3035 ;
  assign n3037 = n1939 & ~n3036 ;
  assign n3038 = ~n3028 & n3037 ;
  assign n3039 = n1851 & n1861 ;
  assign n3040 = ~n1848 & n3039 ;
  assign n3041 = n2101 & ~n3040 ;
  assign n3042 = n1851 & ~n2111 ;
  assign n3043 = ~n1848 & n3042 ;
  assign n3044 = ~n1938 & ~n3043 ;
  assign n3045 = n2098 & ~n3044 ;
  assign n3046 = ~n3041 & n3045 ;
  assign n3047 = ~n3038 & n3046 ;
  assign n3048 = n2114 & ~n2117 ;
  assign n3049 = ~n2098 & n2130 ;
  assign n3050 = ~n3048 & n3049 ;
  assign n3051 = ~n2098 & ~n2130 ;
  assign n3052 = n3048 & n3051 ;
  assign n3053 = ~n3050 & ~n3052 ;
  assign n3054 = n3014 & n3053 ;
  assign n3055 = ~n3047 & n3054 ;
  assign n3056 = ~n3015 & ~n3055 ;
  assign n3057 = n1205 & n1851 ;
  assign n3058 = ~n1848 & n3057 ;
  assign n3059 = ~n2043 & ~n3058 ;
  assign n3060 = n2030 & ~n3059 ;
  assign n3061 = ~n2031 & n3060 ;
  assign n3062 = n3056 & n3061 ;
  assign n3063 = ~n3010 & ~n3062 ;
  assign n3064 = ~\u5_state_reg[41]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3065 = \u5_tmr2_done_reg/NET0131  & ~n2770 ;
  assign n3066 = ~n3064 & ~n3065 ;
  assign n3067 = n1323 & n3066 ;
  assign n3068 = ~\u5_state_reg[45]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3069 = ~n2734 & n2740 ;
  assign n3070 = \u5_tmr2_done_reg/NET0131  & ~n3069 ;
  assign n3071 = n1323 & ~n3070 ;
  assign n3072 = ~n1382 & ~n3071 ;
  assign n3073 = ~n3068 & ~n3072 ;
  assign n3074 = \u5_state_reg[46]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3075 = ~n1882 & n3074 ;
  assign n3076 = ~n1392 & ~n3075 ;
  assign n3077 = n1237 & ~n1537 ;
  assign n3078 = n1532 & n3077 ;
  assign n3079 = n1922 & n3078 ;
  assign n3080 = \u5_state_reg[47]/NET0131  & n1922 ;
  assign n3081 = ~n2809 & n3080 ;
  assign n3082 = ~n3079 & ~n3081 ;
  assign n3083 = \u5_state_reg[47]/NET0131  & ~n2811 ;
  assign n3084 = ~n1922 & n3083 ;
  assign n3085 = n3082 & ~n3084 ;
  assign n3086 = n1929 & ~n3085 ;
  assign n3087 = ~\u5_cmd_asserted_reg/NET0131  & n1345 ;
  assign n3088 = n1109 & n3087 ;
  assign n3089 = n1015 & n3088 ;
  assign n3090 = \u6_read_go_r1_reg/NET0131  & ~n1233 ;
  assign n3091 = n1234 & n3090 ;
  assign n3092 = ~n1048 & n3091 ;
  assign n3093 = n1142 & n3092 ;
  assign n3094 = n1015 & n3093 ;
  assign n3095 = ~n3089 & ~n3094 ;
  assign n3096 = ~n1929 & n3095 ;
  assign n3097 = \u5_state_reg[52]/NET0131  & ~n2812 ;
  assign n3098 = ~n2810 & n3097 ;
  assign n3099 = n1906 & n1922 ;
  assign n3100 = n3095 & ~n3099 ;
  assign n3101 = ~n3098 & n3100 ;
  assign n3102 = ~n3096 & ~n3101 ;
  assign n3103 = ~\u5_cmd_asserted_reg/NET0131  & n1342 ;
  assign n3104 = n1293 & n3103 ;
  assign n3105 = n1115 & n3104 ;
  assign n3106 = ~n1312 & ~n1342 ;
  assign n3107 = n1293 & ~n3106 ;
  assign n3108 = n1115 & n3107 ;
  assign n3109 = n1237 & n3108 ;
  assign n3110 = ~n3105 & ~n3109 ;
  assign n3111 = ~n1929 & n3110 ;
  assign n3112 = n1922 & n2175 ;
  assign n3113 = \u5_state_reg[58]/NET0131  & n1922 ;
  assign n3114 = ~n2809 & n3113 ;
  assign n3115 = ~n3112 & ~n3114 ;
  assign n3116 = \u5_state_reg[58]/NET0131  & ~n2811 ;
  assign n3117 = ~n1922 & n3116 ;
  assign n3118 = n3110 & ~n3117 ;
  assign n3119 = n3115 & n3118 ;
  assign n3120 = ~n3111 & ~n3119 ;
  assign n3121 = ~\u5_cmd_asserted_reg/NET0131  & ~\u5_state_reg[5]/NET0131  ;
  assign n3122 = n1465 & ~n3121 ;
  assign n3123 = n1032 & n3122 ;
  assign n3124 = ~n1305 & ~n1331 ;
  assign n3125 = \u5_state_reg[5]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n3126 = ~n3124 & n3125 ;
  assign n3127 = ~n3123 & ~n3126 ;
  assign n3128 = \u5_state_reg[60]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3129 = ~\u7_mc_ack_r_reg/NET0131  & n3128 ;
  assign n3130 = n1009 & n3129 ;
  assign n3131 = n1151 & n3130 ;
  assign n3132 = n1115 & n3131 ;
  assign n3133 = ~n1929 & ~n3132 ;
  assign n3134 = n1922 & n2050 ;
  assign n3135 = \u5_state_reg[60]/NET0131  & n1922 ;
  assign n3136 = ~n2809 & n3135 ;
  assign n3137 = ~n3134 & ~n3136 ;
  assign n3138 = \u5_state_reg[60]/NET0131  & ~n2811 ;
  assign n3139 = ~n1922 & n3138 ;
  assign n3140 = ~n3132 & ~n3139 ;
  assign n3141 = n3137 & n3140 ;
  assign n3142 = ~n3133 & ~n3141 ;
  assign n3143 = \u5_state_reg[63]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3144 = ~\u7_mc_ack_r_reg/NET0131  & n3143 ;
  assign n3145 = n1290 & n3144 ;
  assign n3146 = ~n1929 & ~n3145 ;
  assign n3147 = n1922 & n2027 ;
  assign n3148 = \u5_state_reg[63]/NET0131  & n1922 ;
  assign n3149 = ~n2809 & n3148 ;
  assign n3150 = ~n3147 & ~n3149 ;
  assign n3151 = \u5_state_reg[63]/NET0131  & ~n2811 ;
  assign n3152 = ~n1922 & n3151 ;
  assign n3153 = ~n3145 & ~n3152 ;
  assign n3154 = n3150 & n3153 ;
  assign n3155 = ~n3146 & ~n3154 ;
  assign n3156 = ~\u5_cmd_asserted_reg/NET0131  & ~\u5_state_reg[7]/NET0131  ;
  assign n3157 = n1273 & ~n3156 ;
  assign n3158 = \u5_tmr_done_reg/NET0131  & ~\u5_wb_wait_r_reg/P0001  ;
  assign n3159 = ~\u5_state_reg[7]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n3160 = ~n3158 & ~n3159 ;
  assign n3161 = ~n1431 & n3160 ;
  assign n3162 = n1193 & n3161 ;
  assign n3163 = ~n3157 & ~n3162 ;
  assign n3164 = \u5_wb_wait_r_reg/P0001  & n1209 ;
  assign n3165 = \u0_sp_csc_reg[10]/NET0131  & \u5_wb_wait_r_reg/P0001  ;
  assign n3166 = ~n1200 & n3165 ;
  assign n3167 = ~n3164 & ~n3166 ;
  assign n3168 = ~n1899 & n3167 ;
  assign n3169 = n1189 & ~n1237 ;
  assign n3170 = ~n3168 & n3169 ;
  assign n3171 = ~n1929 & ~n3170 ;
  assign n3172 = n1538 & n2804 ;
  assign n3173 = \u2_bank_open_reg/P0001  & n1209 ;
  assign n3174 = \u0_sp_csc_reg[10]/NET0131  & \u2_bank_open_reg/P0001  ;
  assign n3175 = ~n1200 & n3174 ;
  assign n3176 = ~n3173 & ~n3175 ;
  assign n3177 = \u2_row_same_reg/P0001  & ~n3176 ;
  assign n3178 = n3172 & n3177 ;
  assign n3179 = n1922 & n3178 ;
  assign n3180 = \u5_state_reg[8]/NET0131  & n1922 ;
  assign n3181 = ~n2809 & n3180 ;
  assign n3182 = ~n3179 & ~n3181 ;
  assign n3183 = \u5_state_reg[8]/NET0131  & ~n2811 ;
  assign n3184 = ~n1922 & n3183 ;
  assign n3185 = ~n3170 & ~n3184 ;
  assign n3186 = n3182 & n3185 ;
  assign n3187 = ~n3171 & ~n3186 ;
  assign n3188 = \u5_state_reg[9]/NET0131  & n3169 ;
  assign n3189 = ~\u5_cmd_asserted_reg/NET0131  & \u5_state_reg[9]/NET0131  ;
  assign n3190 = ~n1185 & n3189 ;
  assign n3191 = ~n3188 & ~n3190 ;
  assign n3192 = n1193 & n3158 ;
  assign n3193 = n1189 & n3168 ;
  assign n3194 = ~n3192 & ~n3193 ;
  assign n3195 = ~n1895 & ~n3194 ;
  assign n3196 = n3191 & ~n3195 ;
  assign n3197 = n964 & n1356 ;
  assign n3198 = n1122 & n3197 ;
  assign n3199 = ~\u5_tmr2_done_reg/NET0131  & n1385 ;
  assign n3200 = n1384 & n3199 ;
  assign n3201 = n1122 & n3200 ;
  assign n3202 = ~n3198 & ~n3201 ;
  assign n3203 = \u7_mc_ack_r_reg/NET0131  & n1290 ;
  assign n3204 = ~n1942 & ~n3203 ;
  assign n3205 = ~n1153 & ~n1290 ;
  assign n3206 = ~\u5_state_reg[65]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3207 = ~\u7_mc_ack_r_reg/NET0131  & ~n3206 ;
  assign n3208 = ~n3205 & n3207 ;
  assign n3209 = ~\u5_cmd_asserted_reg/NET0131  & n1273 ;
  assign n3210 = \u5_state_reg[6]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n3211 = ~n2792 & ~n3210 ;
  assign n3212 = n1304 & ~n3211 ;
  assign n3213 = n1032 & n3212 ;
  assign n3214 = ~n3209 & ~n3213 ;
  assign n3215 = ~n1929 & n3214 ;
  assign n3216 = n1537 & n3176 ;
  assign n3217 = n1532 & n3216 ;
  assign n3218 = n2804 & n3217 ;
  assign n3219 = n1922 & n3218 ;
  assign n3220 = \u5_state_reg[6]/NET0131  & n1922 ;
  assign n3221 = ~n2809 & n3220 ;
  assign n3222 = ~n3219 & ~n3221 ;
  assign n3223 = \u5_state_reg[6]/NET0131  & ~n2811 ;
  assign n3224 = ~n1922 & n3223 ;
  assign n3225 = n3214 & ~n3224 ;
  assign n3226 = n3222 & n3225 ;
  assign n3227 = ~n3215 & ~n3226 ;
  assign n3228 = \u5_wb_cycle_reg/NET0131  & ~n1895 ;
  assign n3229 = n1094 & n3228 ;
  assign n3230 = n2674 & n3229 ;
  assign n3231 = \u5_tmr_done_reg/NET0131  & n1138 ;
  assign n3232 = n1036 & n3231 ;
  assign n3233 = ~n3230 & ~n3232 ;
  assign n3234 = \u5_burst_cnt_reg[1]/NET0131  & n2788 ;
  assign n3235 = ~n2782 & n3234 ;
  assign n3236 = ~\u5_burst_cnt_reg[1]/NET0131  & n2788 ;
  assign n3237 = n2782 & n3236 ;
  assign n3238 = ~n3235 & ~n3237 ;
  assign n3239 = \u5_state_reg[1]/NET0131  & ~\u5_state_reg[52]/NET0131  ;
  assign n3240 = ~n2938 & n3239 ;
  assign n3241 = n1222 & n1851 ;
  assign n3242 = ~n1848 & n3241 ;
  assign n3243 = n3240 & n3242 ;
  assign n3244 = n3238 & ~n3243 ;
  assign n3245 = n2840 & n3240 ;
  assign n3246 = \u5_burst_cnt_reg[3]/NET0131  & n2788 ;
  assign n3247 = ~n2831 & n3246 ;
  assign n3248 = ~\u5_burst_cnt_reg[3]/NET0131  & n2788 ;
  assign n3249 = n2831 & n3248 ;
  assign n3250 = ~n3247 & ~n3249 ;
  assign n3251 = ~n3245 & n3250 ;
  assign n3252 = \u5_resume_req_r_reg/NET0131  & n1104 ;
  assign n3253 = \u5_cmd_asserted_reg/NET0131  & n1345 ;
  assign n3254 = n1109 & n3253 ;
  assign n3255 = n1015 & n3254 ;
  assign n3256 = ~\u5_tmr2_done_reg/NET0131  & n1108 ;
  assign n3257 = n1109 & n3256 ;
  assign n3258 = n1015 & n3257 ;
  assign n3259 = ~n3255 & ~n3258 ;
  assign n3260 = ~\u5_burst_cnt_reg[3]/NET0131  & n1958 ;
  assign n3261 = ~n2749 & n3260 ;
  assign n3262 = ~n2747 & n3261 ;
  assign n3263 = ~\u5_burst_cnt_reg[4]/NET0131  & n3262 ;
  assign n3264 = \u5_burst_cnt_reg[5]/NET0131  & n2788 ;
  assign n3265 = ~n3263 & n3264 ;
  assign n3266 = ~\u5_burst_cnt_reg[5]/NET0131  & n2788 ;
  assign n3267 = n3263 & n3266 ;
  assign n3268 = ~n3265 & ~n3267 ;
  assign n3269 = n1962 & ~n2749 ;
  assign n3270 = ~n2747 & n3269 ;
  assign n3271 = n2788 & n3270 ;
  assign n3272 = ~\u5_burst_cnt_reg[4]/NET0131  & ~\u5_burst_cnt_reg[5]/NET0131  ;
  assign n3273 = n3262 & n3272 ;
  assign n3274 = \u5_burst_cnt_reg[6]/NET0131  & n2788 ;
  assign n3275 = ~n3273 & n3274 ;
  assign n3276 = ~n3271 & ~n3275 ;
  assign n3277 = ~\u5_oe__reg/NET0131  & ~\u5_susp_sel_r_reg/NET0131  ;
  assign n3278 = \u5_burst_cnt_reg[7]/NET0131  & n2788 ;
  assign n3279 = ~n3270 & n3278 ;
  assign n3280 = ~\u5_burst_cnt_reg[7]/NET0131  & n2788 ;
  assign n3281 = n3270 & n3280 ;
  assign n3282 = ~n3279 & ~n3281 ;
  assign n3283 = \u5_burst_cnt_reg[4]/NET0131  & n2788 ;
  assign n3284 = ~n3262 & n3283 ;
  assign n3285 = ~\u5_burst_cnt_reg[4]/NET0131  & n2788 ;
  assign n3286 = n3262 & n3285 ;
  assign n3287 = ~n3284 & ~n3286 ;
  assign n3288 = ~n1111 & ~n1163 ;
  assign n3289 = \u5_state_reg[48]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3290 = ~n3288 & n3289 ;
  assign n3291 = ~n1352 & ~n3290 ;
  assign n3292 = \u5_wb_cycle_reg/NET0131  & ~n3228 ;
  assign n3293 = ~n1966 & ~n3228 ;
  assign n3294 = ~n1954 & n3293 ;
  assign n3295 = ~n3292 & ~n3294 ;
  assign n3296 = \u5_state_reg[15]/NET0131  & ~n1966 ;
  assign n3297 = ~n1954 & n3296 ;
  assign n3298 = n3295 & ~n3297 ;
  assign n3299 = n1094 & ~n3298 ;
  assign n3300 = ~\u5_cmd_asserted_reg/NET0131  & n1269 ;
  assign n3301 = ~n1895 & n2146 ;
  assign n3302 = n1248 & n3301 ;
  assign n3303 = n2682 & n3302 ;
  assign n3304 = ~n1954 & n3303 ;
  assign n3305 = ~n3300 & ~n3304 ;
  assign n3306 = ~n1977 & n3305 ;
  assign n3307 = ~n3299 & n3306 ;
  assign n3308 = n1400 & n2170 ;
  assign n3309 = n1897 & ~n1966 ;
  assign n3310 = ~n1954 & n3309 ;
  assign n3311 = n1023 & ~n3310 ;
  assign n3312 = ~n3308 & ~n3311 ;
  assign n3313 = n1245 & ~n2669 ;
  assign n3314 = n2666 & n3313 ;
  assign n3315 = ~n1966 & n3314 ;
  assign n3316 = ~n1954 & n3315 ;
  assign n3317 = n2678 & n3316 ;
  assign n3318 = ~n1250 & ~n2014 ;
  assign n3319 = \u5_cmd_asserted_reg/NET0131  & n1234 ;
  assign n3320 = n1232 & n3319 ;
  assign n3321 = ~n1048 & n3320 ;
  assign n3322 = ~\u5_wb_cycle_reg/NET0131  & n3321 ;
  assign n3323 = ~n1966 & n3321 ;
  assign n3324 = ~n1954 & n3323 ;
  assign n3325 = ~n3322 & ~n3324 ;
  assign n3326 = ~\u5_cmd_asserted_reg/NET0131  & \u5_state_reg[14]/NET0131  ;
  assign n3327 = ~n2014 & ~n3326 ;
  assign n3328 = n3325 & n3327 ;
  assign n3329 = ~n3318 & ~n3328 ;
  assign n3330 = ~n3317 & ~n3329 ;
  assign n3331 = \u5_data_oe_reg/NET0131  & \u5_mc_c_oe_reg/NET0131  ;
  assign n3332 = ~\u5_susp_sel_r_reg/NET0131  & n3331 ;
  assign n3333 = ~\u5_state_reg[24]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n3334 = n982 & n1096 ;
  assign n3335 = n1078 & n3334 ;
  assign n3336 = \u5_ir_cnt_done_reg/P0001  & \u5_tmr_done_reg/NET0131  ;
  assign n3337 = ~\u5_state_reg[23]/NET0131  & n3336 ;
  assign n3338 = \u5_state_reg[23]/NET0131  & \u5_state_reg[25]/NET0131  ;
  assign n3339 = ~n981 & ~n3338 ;
  assign n3340 = ~n3337 & n3339 ;
  assign n3341 = n3335 & n3340 ;
  assign n3342 = ~n3333 & n3341 ;
  assign n3343 = ~\u5_cmd_asserted_reg/NET0131  & n1419 ;
  assign n3344 = n1096 & n3343 ;
  assign n3345 = n1078 & n3344 ;
  assign n3346 = ~n3342 & ~n3345 ;
  assign n3347 = ~\u5_wb_stb_first_reg/NET0131  & ~wb_stb_i_pad ;
  assign n3348 = ~\u6_read_go_r_reg/NET0131  & ~\u6_write_go_r_reg/NET0131  ;
  assign n3349 = n1045 & n3348 ;
  assign n3350 = n2191 & n3349 ;
  assign n3351 = \u6_wb_first_r_reg/NET0131  & ~wb_ack_o_pad ;
  assign n3352 = ~wb_err_o_pad & n3351 ;
  assign n3353 = ~\u5_wb_stb_first_reg/NET0131  & ~n3352 ;
  assign n3354 = ~n3350 & n3353 ;
  assign n3355 = ~n3347 & ~n3354 ;
  assign n3356 = n1898 & n3355 ;
  assign n3357 = ~n2152 & n3355 ;
  assign n3358 = n2188 & n3357 ;
  assign n3359 = ~n3356 & ~n3358 ;
  assign n3360 = ~\u5_cmd_asserted_reg/NET0131  & ~\u5_state_reg[19]/NET0131  ;
  assign n3361 = n1453 & ~n3360 ;
  assign n3362 = ~\u5_tmr_done_reg/NET0131  & n1255 ;
  assign n3363 = n1254 & n3362 ;
  assign n3364 = ~n3361 & ~n3363 ;
  assign n3365 = n1023 & n3309 ;
  assign n3366 = ~n1954 & n3365 ;
  assign n3367 = ~\u5_state_reg[54]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n3368 = n1108 & ~n3367 ;
  assign n3369 = n1109 & n3368 ;
  assign n3370 = n1015 & n3369 ;
  assign n3371 = ~n3366 & ~n3370 ;
  assign n3372 = n1310 & n1901 ;
  assign n3373 = n1861 & n3372 ;
  assign n3374 = n1851 & n3373 ;
  assign n3375 = ~n1848 & n3374 ;
  assign n3376 = n968 & n970 ;
  assign n3377 = n1088 & n3376 ;
  assign n3378 = ~n1160 & ~n1349 ;
  assign n3379 = \u5_cmd_asserted_reg/NET0131  & ~n1349 ;
  assign n3380 = ~n3378 & ~n3379 ;
  assign n3381 = n3377 & n3380 ;
  assign n3382 = n2036 & n3381 ;
  assign n3383 = n1851 & n3382 ;
  assign n3384 = ~n1848 & n3383 ;
  assign n3385 = \u5_state_reg[51]/NET0131  & ~n2096 ;
  assign n3386 = ~n3381 & ~n3385 ;
  assign n3387 = ~n3384 & ~n3386 ;
  assign n3388 = \u5_state_reg[40]/NET0131  & ~\u5_state_reg[51]/NET0131  ;
  assign n3389 = ~n3058 & n3388 ;
  assign n3390 = ~\u5_state_reg[40]/NET0131  & ~\u5_state_reg[51]/NET0131  ;
  assign n3391 = ~\u5_timer2_reg[0]/P0001  & ~\u5_timer2_reg[1]/P0001  ;
  assign n3392 = ~\u5_timer2_reg[2]/P0001  & ~\u5_timer2_reg[3]/P0001  ;
  assign n3393 = n3391 & n3392 ;
  assign n3394 = ~\u5_timer2_reg[4]/P0001  & ~\u5_timer2_reg[6]/P0001  ;
  assign n3395 = ~\u5_timer2_reg[5]/P0001  & n3394 ;
  assign n3396 = n3393 & n3395 ;
  assign n3397 = ~\u5_timer2_reg[7]/P0001  & ~\u5_timer2_reg[8]/P0001  ;
  assign n3398 = n3396 & n3397 ;
  assign n3399 = ~\u5_state_reg[36]/NET0131  & ~\u5_state_reg[41]/NET0131  ;
  assign n3400 = n962 & n3399 ;
  assign n3401 = ~\u5_timer2_reg[2]/P0001  & n3391 ;
  assign n3402 = \u5_timer2_reg[2]/P0001  & ~n3391 ;
  assign n3403 = ~n3401 & ~n3402 ;
  assign n3404 = n3400 & ~n3403 ;
  assign n3405 = ~n3398 & n3404 ;
  assign n3406 = n3390 & n3405 ;
  assign n3407 = n3390 & ~n3400 ;
  assign n3408 = ~n3012 & n3407 ;
  assign n3409 = ~n3406 & ~n3408 ;
  assign n3410 = ~n3389 & n3409 ;
  assign n3411 = \u5_tmr2_done_reg/NET0131  & n1163 ;
  assign n3412 = ~n3384 & ~n3411 ;
  assign n3413 = ~n3410 & n3412 ;
  assign n3414 = ~n3387 & ~n3413 ;
  assign n3415 = ~n3381 & n3411 ;
  assign n3416 = ~n2971 & n3415 ;
  assign n3417 = n1310 & n1544 ;
  assign n3418 = ~n1347 & ~n3417 ;
  assign n3419 = ~n3416 & n3418 ;
  assign n3420 = n3414 & n3419 ;
  assign n3421 = ~n3375 & ~n3420 ;
  assign n3422 = \u5_state_reg[37]/NET0131  & ~n2739 ;
  assign n3423 = ~n2736 & n3422 ;
  assign n3424 = n963 & ~n3423 ;
  assign n3425 = \u1_acs_addr_reg[12]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n3426 = \u1_u0_out_r_reg[12]/P0001  & n3425 ;
  assign n3427 = ~n3424 & n3426 ;
  assign n3428 = \u1_acs_addr_reg[13]/P0001  & \u1_acs_addr_reg[15]/P0001  ;
  assign n3429 = \u1_acs_addr_reg[14]/P0001  & n3428 ;
  assign n3430 = n3427 & n3429 ;
  assign n3431 = \u1_acs_addr_reg[16]/P0001  & \u1_acs_addr_reg[18]/P0001  ;
  assign n3432 = \u1_acs_addr_reg[17]/P0001  & n3431 ;
  assign n3433 = n3430 & n3432 ;
  assign n3434 = \u1_acs_addr_reg[19]/P0001  & \u1_acs_addr_reg[21]/P0001  ;
  assign n3435 = \u1_acs_addr_reg[20]/P0001  & n3434 ;
  assign n3436 = n3433 & n3435 ;
  assign n3437 = \u1_acs_addr_reg[22]/P0001  & ~\u1_acs_addr_reg[23]/P0001  ;
  assign n3438 = n3436 & n3437 ;
  assign n3439 = ~\u5_cs_le_reg/P0001  & ~wb_we_i_pad ;
  assign n3440 = ~\u1_acs_addr_reg[23]/P0001  & n3439 ;
  assign n3441 = \u1_acs_addr_reg[22]/P0001  & n3439 ;
  assign n3442 = n3436 & n3441 ;
  assign n3443 = ~n3440 & ~n3442 ;
  assign n3444 = ~n3438 & ~n3443 ;
  assign n3445 = \wb_addr_i[25]_pad  & ~n2733 ;
  assign n3446 = ~n2730 & n3445 ;
  assign n3447 = ~n2740 & n3446 ;
  assign n3448 = ~n3439 & ~n3447 ;
  assign n3449 = \wb_addr_i[24]_pad  & ~n2739 ;
  assign n3450 = ~n2736 & n3449 ;
  assign n3451 = ~n2734 & n3450 ;
  assign n3452 = \wb_addr_i[23]_pad  & ~n2733 ;
  assign n3453 = ~n2730 & n3452 ;
  assign n3454 = n2740 & n3453 ;
  assign n3455 = ~n3451 & ~n3454 ;
  assign n3456 = n3448 & n3455 ;
  assign n3457 = ~n3444 & ~n3456 ;
  assign n3458 = ~n2971 & n3372 ;
  assign n3459 = ~n3418 & ~n3458 ;
  assign n3460 = n3008 & n3381 ;
  assign n3461 = n1851 & n3460 ;
  assign n3462 = ~n1848 & n3461 ;
  assign n3463 = \u5_state_reg[51]/NET0131  & ~n3043 ;
  assign n3464 = ~n3381 & ~n3463 ;
  assign n3465 = ~n3462 & ~n3464 ;
  assign n3466 = \u5_timer2_reg[0]/P0001  & \u5_timer2_reg[1]/P0001  ;
  assign n3467 = ~n3391 & ~n3466 ;
  assign n3468 = n3400 & ~n3467 ;
  assign n3469 = ~n3398 & n3468 ;
  assign n3470 = n3390 & n3469 ;
  assign n3471 = ~n2938 & n3407 ;
  assign n3472 = ~n3470 & ~n3471 ;
  assign n3473 = ~n2991 & n3388 ;
  assign n3474 = n3472 & ~n3473 ;
  assign n3475 = ~n3411 & ~n3462 ;
  assign n3476 = ~n3474 & n3475 ;
  assign n3477 = ~n3465 & ~n3476 ;
  assign n3478 = n1851 & ~n1874 ;
  assign n3479 = ~n1848 & n3478 ;
  assign n3480 = n3415 & ~n3479 ;
  assign n3481 = ~n3458 & ~n3480 ;
  assign n3482 = n3477 & n3481 ;
  assign n3483 = ~n3459 & ~n3482 ;
  assign n3484 = ~n2100 & n3372 ;
  assign n3485 = n1851 & n2048 ;
  assign n3486 = ~n1848 & n3485 ;
  assign n3487 = n3388 & ~n3486 ;
  assign n3488 = n1221 & ~n3400 ;
  assign n3489 = n1851 & n3488 ;
  assign n3490 = ~n1848 & n3489 ;
  assign n3491 = ~n3398 & n3401 ;
  assign n3492 = \u5_timer2_reg[3]/P0001  & ~n3491 ;
  assign n3493 = n3393 & ~n3398 ;
  assign n3494 = n3400 & ~n3493 ;
  assign n3495 = ~n3492 & n3494 ;
  assign n3496 = n3390 & ~n3495 ;
  assign n3497 = ~n3490 & n3496 ;
  assign n3498 = ~n3487 & ~n3497 ;
  assign n3499 = ~n3411 & ~n3498 ;
  assign n3500 = \u5_state_reg[51]/NET0131  & ~n2613 ;
  assign n3501 = ~n3040 & n3411 ;
  assign n3502 = ~n3381 & ~n3501 ;
  assign n3503 = ~n3500 & n3502 ;
  assign n3504 = ~n3499 & n3503 ;
  assign n3505 = n2122 & n3381 ;
  assign n3506 = n1851 & n3505 ;
  assign n3507 = ~n1848 & n3506 ;
  assign n3508 = n3418 & ~n3507 ;
  assign n3509 = ~n3504 & n3508 ;
  assign n3510 = ~n3484 & ~n3509 ;
  assign n3511 = n1929 & n2807 ;
  assign n3512 = n1922 & n3511 ;
  assign n3513 = ~n1189 & ~n1314 ;
  assign n3514 = ~n3512 & n3513 ;
  assign n3515 = n1237 & ~n3514 ;
  assign n3516 = ~n1344 & ~n1352 ;
  assign n3517 = ~n1157 & n3516 ;
  assign n3518 = n1251 & n3517 ;
  assign n3519 = ~n3515 & n3518 ;
  assign n3520 = n1496 & n3519 ;
  assign n3521 = ~n1879 & n3520 ;
  assign n3522 = ~\u5_wr_cycle_reg/NET0131  & ~n3521 ;
  assign n3523 = \u5_data_oe_r2_reg/NET0131  & \u5_wr_cycle_reg/NET0131  ;
  assign n3524 = ~n3522 & ~n3523 ;
  assign n3525 = \u5_cnt_reg/NET0131  & \u5_wb_cycle_reg/NET0131  ;
  assign n3526 = ~n1966 & n3525 ;
  assign n3527 = ~n1954 & n3526 ;
  assign n3528 = ~mc_cke_pad_o__pad & ~n3527 ;
  assign n3529 = n1899 & n3526 ;
  assign n3530 = ~n1954 & n3529 ;
  assign n3531 = n1094 & ~n3530 ;
  assign n3532 = ~n3528 & n3531 ;
  assign n3533 = \u5_cke_r_reg/NET0131  & n3532 ;
  assign n3534 = ~n1482 & n2907 ;
  assign n3535 = n1501 & n3534 ;
  assign n3536 = ~n1421 & ~n1462 ;
  assign n3537 = n1158 & ~n1184 ;
  assign n3538 = n1149 & n3537 ;
  assign n3539 = n1507 & n3538 ;
  assign n3540 = n3536 & n3539 ;
  assign n3541 = n3535 & n3540 ;
  assign n3542 = ~n1250 & n1488 ;
  assign n3543 = n1487 & n3542 ;
  assign n3544 = n1407 & n3543 ;
  assign n3545 = ~n1100 & ~n1285 ;
  assign n3546 = ~n1094 & ~n1245 ;
  assign n3547 = n3545 & n3546 ;
  assign n3548 = n1093 & ~n1411 ;
  assign n3549 = n1490 & n3548 ;
  assign n3550 = n3547 & n3549 ;
  assign n3551 = n3544 & n3550 ;
  assign n3552 = ~n1135 & n1475 ;
  assign n3553 = n1474 & n3552 ;
  assign n3554 = n3551 & n3553 ;
  assign n3555 = n3541 & n3554 ;
  assign n3556 = \u5_cke_r_reg/NET0131  & ~n1094 ;
  assign n3557 = ~n3555 & n3556 ;
  assign n3558 = ~n3533 & ~n3557 ;
  assign n3559 = ~n1339 & n3545 ;
  assign n3560 = \u5_state_reg[0]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n3561 = ~n3559 & n3560 ;
  assign n3562 = \wb_addr_i[21]_pad  & ~n2733 ;
  assign n3563 = ~n2730 & n3562 ;
  assign n3564 = ~n2740 & n3563 ;
  assign n3565 = \wb_addr_i[20]_pad  & ~n2739 ;
  assign n3566 = ~n2736 & n3565 ;
  assign n3567 = ~n2734 & n3566 ;
  assign n3568 = \wb_addr_i[19]_pad  & ~n2733 ;
  assign n3569 = ~n2730 & n3568 ;
  assign n3570 = n2740 & n3569 ;
  assign n3571 = ~n3567 & ~n3570 ;
  assign n3572 = ~n3564 & n3571 ;
  assign n3573 = ~n3439 & ~n3572 ;
  assign n3574 = \u1_acs_addr_reg[19]/P0001  & n3439 ;
  assign n3575 = ~n3433 & n3574 ;
  assign n3576 = ~\u1_acs_addr_reg[19]/P0001  & n3439 ;
  assign n3577 = n3433 & n3576 ;
  assign n3578 = ~n3575 & ~n3577 ;
  assign n3579 = ~n3573 & n3578 ;
  assign n3580 = \wb_addr_i[23]_pad  & ~n2739 ;
  assign n3581 = ~n2736 & n3580 ;
  assign n3582 = ~n2734 & n3581 ;
  assign n3583 = \wb_addr_i[22]_pad  & ~n2733 ;
  assign n3584 = ~n2730 & n3583 ;
  assign n3585 = n2740 & n3584 ;
  assign n3586 = \wb_addr_i[24]_pad  & ~n2733 ;
  assign n3587 = ~n2730 & n3586 ;
  assign n3588 = ~n2740 & n3587 ;
  assign n3589 = ~n3585 & ~n3588 ;
  assign n3590 = ~n3582 & n3589 ;
  assign n3591 = ~n3439 & ~n3590 ;
  assign n3592 = ~n3436 & n3441 ;
  assign n3593 = ~\u1_acs_addr_reg[22]/P0001  & n3439 ;
  assign n3594 = n3436 & n3593 ;
  assign n3595 = ~n3592 & ~n3594 ;
  assign n3596 = ~n3591 & n3595 ;
  assign n3597 = n1038 & ~n1966 ;
  assign n3598 = ~n1954 & n3597 ;
  assign n3599 = ~\u5_cke_r_reg/NET0131  & ~n3598 ;
  assign n3600 = n1899 & n3597 ;
  assign n3601 = ~n1954 & n3600 ;
  assign n3602 = ~n1245 & ~n3601 ;
  assign n3603 = ~n3599 & n3602 ;
  assign n3604 = \u5_cke_r_reg/NET0131  & \u5_cnt_reg/NET0131  ;
  assign n3605 = \u5_cnt_reg/NET0131  & ~n3604 ;
  assign n3606 = n1233 & ~n3604 ;
  assign n3607 = ~n1898 & n3606 ;
  assign n3608 = ~n3605 & ~n3607 ;
  assign n3609 = n1245 & ~n3608 ;
  assign n3610 = ~n1250 & ~n3609 ;
  assign n3611 = ~n3603 & ~n3610 ;
  assign n3612 = n1251 & n1475 ;
  assign n3613 = n1474 & n3612 ;
  assign n3614 = ~n1104 & n3613 ;
  assign n3615 = n3551 & n3614 ;
  assign n3616 = n3541 & n3615 ;
  assign n3617 = ~n3611 & ~n3616 ;
  assign n3618 = ~n3043 & n3372 ;
  assign n3619 = n1851 & n2961 ;
  assign n3620 = ~n1848 & n3619 ;
  assign n3621 = ~\u5_state_reg[40]/NET0131  & ~n3400 ;
  assign n3622 = ~n3620 & n3621 ;
  assign n3623 = ~n3398 & n3400 ;
  assign n3624 = ~\u5_timer2_reg[4]/P0001  & n3393 ;
  assign n3625 = ~\u5_state_reg[40]/NET0131  & \u5_timer2_reg[5]/P0001  ;
  assign n3626 = ~n3624 & n3625 ;
  assign n3627 = ~\u5_state_reg[40]/NET0131  & ~\u5_timer2_reg[5]/P0001  ;
  assign n3628 = n3624 & n3627 ;
  assign n3629 = ~n3626 & ~n3628 ;
  assign n3630 = n3623 & ~n3629 ;
  assign n3631 = ~\u5_state_reg[51]/NET0131  & ~n3630 ;
  assign n3632 = ~n3622 & n3631 ;
  assign n3633 = ~n3381 & ~n3411 ;
  assign n3634 = n3418 & n3633 ;
  assign n3635 = \u5_state_reg[51]/NET0131  & ~n3020 ;
  assign n3636 = n1851 & n3635 ;
  assign n3637 = ~n1848 & n3636 ;
  assign n3638 = n3634 & ~n3637 ;
  assign n3639 = ~n3632 & n3638 ;
  assign n3640 = ~n3618 & ~n3639 ;
  assign n3641 = \u1_acs_addr_reg[19]/P0001  & n3433 ;
  assign n3642 = ~\u1_acs_addr_reg[20]/P0001  & n3439 ;
  assign n3643 = ~n3641 & n3642 ;
  assign n3644 = \u1_acs_addr_reg[20]/P0001  & n3439 ;
  assign n3645 = n3641 & n3644 ;
  assign n3646 = ~n3643 & ~n3645 ;
  assign n3647 = ~n2740 & n3584 ;
  assign n3648 = ~n3439 & ~n3647 ;
  assign n3649 = \wb_addr_i[21]_pad  & ~n2739 ;
  assign n3650 = ~n2736 & n3649 ;
  assign n3651 = ~n2734 & n3650 ;
  assign n3652 = \wb_addr_i[20]_pad  & ~n2733 ;
  assign n3653 = ~n2730 & n3652 ;
  assign n3654 = n2740 & n3653 ;
  assign n3655 = ~n3651 & ~n3654 ;
  assign n3656 = n3648 & n3655 ;
  assign n3657 = n3646 & ~n3656 ;
  assign n3658 = ~n3381 & n3418 ;
  assign n3659 = ~n2100 & n3411 ;
  assign n3660 = n1851 & ~n2945 ;
  assign n3661 = ~n1848 & n3660 ;
  assign n3662 = \u5_state_reg[51]/NET0131  & ~n3661 ;
  assign n3663 = ~n3659 & ~n3662 ;
  assign n3664 = n3658 & ~n3663 ;
  assign n3665 = \u5_state_reg[40]/NET0131  & ~n2603 ;
  assign n3666 = ~n2654 & n3621 ;
  assign n3667 = \u5_timer2_reg[4]/P0001  & n3393 ;
  assign n3668 = ~n3398 & n3667 ;
  assign n3669 = ~\u5_state_reg[36]/NET0131  & n962 ;
  assign n3670 = n960 & n3669 ;
  assign n3671 = \u5_timer2_reg[4]/P0001  & n3670 ;
  assign n3672 = n3393 & n3670 ;
  assign n3673 = ~n3398 & n3672 ;
  assign n3674 = ~n3671 & ~n3673 ;
  assign n3675 = ~n3668 & ~n3674 ;
  assign n3676 = ~n3666 & ~n3675 ;
  assign n3677 = ~n3665 & n3676 ;
  assign n3678 = ~\u5_state_reg[51]/NET0131  & ~n3411 ;
  assign n3679 = n3658 & n3678 ;
  assign n3680 = ~n3677 & n3679 ;
  assign n3681 = ~n3664 & ~n3680 ;
  assign n3682 = ~n2968 & n3372 ;
  assign n3683 = n3681 & ~n3682 ;
  assign n3684 = \u1_bank_adr_reg[0]/P0001  & ~\u1_bank_adr_reg[1]/P0001  ;
  assign n3685 = \u5_state_reg[7]/NET0131  & n1209 ;
  assign n3686 = \u0_sp_csc_reg[10]/NET0131  & \u5_state_reg[7]/NET0131  ;
  assign n3687 = ~n1200 & n3686 ;
  assign n3688 = ~n3685 & ~n3687 ;
  assign n3689 = n3684 & ~n3688 ;
  assign n3690 = n1840 & n3689 ;
  assign n3691 = \u5_state_reg[22]/NET0131  & ~n975 ;
  assign n3692 = ~\u5_state_reg[24]/NET0131  & n981 ;
  assign n3693 = n986 & n3692 ;
  assign n3694 = ~n3691 & n3693 ;
  assign n3695 = ~\u5_state_reg[22]/NET0131  & ~n1459 ;
  assign n3696 = ~n1262 & n3695 ;
  assign n3697 = ~\u5_state_reg[21]/NET0131  & n966 ;
  assign n3698 = n974 & n3697 ;
  assign n3699 = ~n3696 & n3698 ;
  assign n3700 = n3694 & n3699 ;
  assign n3701 = n971 & n1017 ;
  assign n3702 = n967 & n1383 ;
  assign n3703 = n961 & n3702 ;
  assign n3704 = n3701 & n3703 ;
  assign n3705 = n1008 & n1379 ;
  assign n3706 = n1007 & n3705 ;
  assign n3707 = n1295 & n3706 ;
  assign n3708 = n3704 & n3707 ;
  assign n3709 = n3700 & n3708 ;
  assign n3710 = ~\u5_state_reg[20]/NET0131  & n977 ;
  assign n3711 = n3709 & n3710 ;
  assign n3712 = ~\u5_state_reg[7]/NET0131  & n997 ;
  assign n3713 = n1012 & n1057 ;
  assign n3714 = n3712 & n3713 ;
  assign n3715 = n992 & n1033 ;
  assign n3716 = n1054 & n3715 ;
  assign n3717 = n3714 & n3716 ;
  assign n3718 = n3711 & n3717 ;
  assign n3719 = ~n977 & ~n1450 ;
  assign n3720 = ~\u5_state_reg[20]/NET0131  & ~n1450 ;
  assign n3721 = ~n3709 & n3720 ;
  assign n3722 = ~n3719 & ~n3721 ;
  assign n3723 = ~\u5_state_reg[27]/NET0131  & n974 ;
  assign n3724 = n3707 & n3723 ;
  assign n3725 = ~\u5_state_reg[21]/NET0131  & ~\u5_state_reg[23]/NET0131  ;
  assign n3726 = n982 & n3725 ;
  assign n3727 = n1067 & n3726 ;
  assign n3728 = ~\u5_state_reg[25]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n3729 = n1062 & n3728 ;
  assign n3730 = n3727 & n3729 ;
  assign n3731 = n3704 & n3730 ;
  assign n3732 = n3724 & n3731 ;
  assign n3733 = n3717 & n3732 ;
  assign n3734 = n3722 & n3733 ;
  assign n3735 = ~n3718 & ~n3734 ;
  assign n3736 = n1840 & ~n3735 ;
  assign n3737 = ~\u5_rfr_ack_r_reg/NET0131  & ~\u5_state_reg[16]/NET0131  ;
  assign n3738 = \u5_state_reg[4]/NET0131  & n3737 ;
  assign n3739 = \u5_state_reg[16]/NET0131  & ~\u5_state_reg[4]/NET0131  ;
  assign n3740 = \u5_tmr_done_reg/NET0131  & n3739 ;
  assign n3741 = ~n1209 & n3740 ;
  assign n3742 = ~n1206 & n3741 ;
  assign n3743 = ~n3738 & ~n3742 ;
  assign n3744 = ~n1839 & n3684 ;
  assign n3745 = n1835 & n3744 ;
  assign n3746 = ~n3743 & n3745 ;
  assign n3747 = \u2_u0_bank1_open_reg/NET0131  & ~n3746 ;
  assign n3748 = ~\u5_rfr_ack_r_reg/NET0131  & n3747 ;
  assign n3749 = ~n3736 & n3748 ;
  assign n3750 = ~n3690 & ~n3749 ;
  assign n3751 = ~\u1_bank_adr_reg[0]/P0001  & \u1_bank_adr_reg[1]/P0001  ;
  assign n3752 = ~n3688 & n3751 ;
  assign n3753 = n1840 & n3752 ;
  assign n3754 = ~n1839 & n3751 ;
  assign n3755 = n1835 & n3754 ;
  assign n3756 = ~n3743 & n3755 ;
  assign n3757 = \u2_u0_bank2_open_reg/NET0131  & ~n3756 ;
  assign n3758 = ~\u5_rfr_ack_r_reg/NET0131  & n3757 ;
  assign n3759 = ~n3736 & n3758 ;
  assign n3760 = ~n3753 & ~n3759 ;
  assign n3761 = ~n1919 & n3752 ;
  assign n3762 = ~n1919 & ~n3735 ;
  assign n3763 = ~n1919 & ~n3743 ;
  assign n3764 = n3751 & n3763 ;
  assign n3765 = \u2_u1_bank2_open_reg/NET0131  & ~n3764 ;
  assign n3766 = ~\u5_rfr_ack_r_reg/NET0131  & n3765 ;
  assign n3767 = ~n3762 & n3766 ;
  assign n3768 = ~n3761 & ~n3767 ;
  assign n3769 = ~n1919 & n3689 ;
  assign n3770 = n3684 & n3763 ;
  assign n3771 = \u2_u1_bank1_open_reg/NET0131  & ~n3770 ;
  assign n3772 = ~\u5_rfr_ack_r_reg/NET0131  & n3771 ;
  assign n3773 = ~n3762 & n3772 ;
  assign n3774 = ~n3769 & ~n3773 ;
  assign n3775 = ~\u1_acs_addr_reg[16]/P0001  & n3439 ;
  assign n3776 = ~n3430 & n3775 ;
  assign n3777 = \u1_acs_addr_reg[16]/P0001  & n3439 ;
  assign n3778 = n3430 & n3777 ;
  assign n3779 = ~n3776 & ~n3778 ;
  assign n3780 = \wb_addr_i[16]_pad  & ~n2733 ;
  assign n3781 = ~n2730 & n3780 ;
  assign n3782 = n2740 & n3781 ;
  assign n3783 = ~n3439 & ~n3782 ;
  assign n3784 = \wb_addr_i[18]_pad  & ~n2733 ;
  assign n3785 = ~n2730 & n3784 ;
  assign n3786 = ~n2740 & n3785 ;
  assign n3787 = \wb_addr_i[17]_pad  & ~n2739 ;
  assign n3788 = ~n2736 & n3787 ;
  assign n3789 = ~n2734 & n3788 ;
  assign n3790 = ~n3786 & ~n3789 ;
  assign n3791 = n3783 & n3790 ;
  assign n3792 = n3779 & ~n3791 ;
  assign n3793 = \u1_bank_adr_reg[0]/P0001  & \u1_bank_adr_reg[1]/P0001  ;
  assign n3794 = ~n3688 & n3793 ;
  assign n3795 = n1840 & n3794 ;
  assign n3796 = ~n1839 & n3793 ;
  assign n3797 = n1835 & n3796 ;
  assign n3798 = ~n3743 & n3797 ;
  assign n3799 = \u2_u0_bank3_open_reg/NET0131  & ~n3798 ;
  assign n3800 = ~\u5_rfr_ack_r_reg/NET0131  & n3799 ;
  assign n3801 = ~n3736 & n3800 ;
  assign n3802 = ~n3795 & ~n3801 ;
  assign n3803 = ~n1919 & n3794 ;
  assign n3804 = n3763 & n3793 ;
  assign n3805 = \u2_u1_bank3_open_reg/NET0131  & ~n3804 ;
  assign n3806 = ~\u5_rfr_ack_r_reg/NET0131  & n3805 ;
  assign n3807 = ~n3762 & n3806 ;
  assign n3808 = ~n3803 & ~n3807 ;
  assign n3809 = \wb_addr_i[19]_pad  & ~n2739 ;
  assign n3810 = ~n2736 & n3809 ;
  assign n3811 = ~n2734 & n3810 ;
  assign n3812 = n2740 & n3785 ;
  assign n3813 = ~n2740 & n3653 ;
  assign n3814 = ~n3812 & ~n3813 ;
  assign n3815 = ~n3811 & n3814 ;
  assign n3816 = ~n3439 & ~n3815 ;
  assign n3817 = \u1_acs_addr_reg[16]/P0001  & \u1_acs_addr_reg[17]/P0001  ;
  assign n3818 = n3430 & n3817 ;
  assign n3819 = ~\u1_acs_addr_reg[18]/P0001  & ~n3818 ;
  assign n3820 = ~n3433 & n3439 ;
  assign n3821 = ~n3819 & n3820 ;
  assign n3822 = ~n3816 & ~n3821 ;
  assign n3823 = n3372 & ~n3479 ;
  assign n3824 = \u5_state_reg[51]/NET0131  & n2127 ;
  assign n3825 = n1851 & n3824 ;
  assign n3826 = ~n1848 & n3825 ;
  assign n3827 = ~\u5_timer2_reg[0]/P0001  & ~n3398 ;
  assign n3828 = \u5_timer2_reg[0]/P0001  & ~\u5_timer2_reg[8]/P0001  ;
  assign n3829 = ~\u5_timer2_reg[7]/P0001  & n3828 ;
  assign n3830 = n3396 & n3829 ;
  assign n3831 = n3390 & n3400 ;
  assign n3832 = ~n3830 & n3831 ;
  assign n3833 = ~n3827 & n3832 ;
  assign n3834 = ~n3411 & ~n3833 ;
  assign n3835 = ~n3826 & n3834 ;
  assign n3836 = ~n3381 & ~n3835 ;
  assign n3837 = n2999 & n3381 ;
  assign n3838 = n1851 & n3837 ;
  assign n3839 = ~n1848 & n3838 ;
  assign n3840 = n3418 & ~n3839 ;
  assign n3841 = ~n3836 & n3840 ;
  assign n3842 = ~n3823 & ~n3841 ;
  assign n3843 = ~n2096 & n3372 ;
  assign n3844 = n3033 & ~n3400 ;
  assign n3845 = n1851 & n3844 ;
  assign n3846 = ~n1848 & n3845 ;
  assign n3847 = n3396 & ~n3398 ;
  assign n3848 = ~\u5_timer2_reg[4]/P0001  & ~\u5_timer2_reg[5]/P0001  ;
  assign n3849 = n3393 & n3848 ;
  assign n3850 = \u5_timer2_reg[6]/P0001  & ~n3849 ;
  assign n3851 = n3400 & ~n3850 ;
  assign n3852 = ~n3847 & n3851 ;
  assign n3853 = n3390 & ~n3852 ;
  assign n3854 = n3634 & n3853 ;
  assign n3855 = ~n3846 & n3854 ;
  assign n3856 = ~n3843 & ~n3855 ;
  assign n3857 = \u0_sp_tms_reg[0]/NET0131  & ~n1045 ;
  assign n3858 = ~\u4_rfr_req_reg/NET0131  & n1309 ;
  assign n3859 = n1308 & n3858 ;
  assign n3860 = ~n1531 & n1921 ;
  assign n3861 = ~n1920 & n3860 ;
  assign n3862 = \u5_wb_stb_first_reg/NET0131  & ~n3861 ;
  assign n3863 = \u5_lookup_ready2_reg/NET0131  & ~n1920 ;
  assign n3864 = ~n1233 & ~n1898 ;
  assign n3865 = n2807 & n3864 ;
  assign n3866 = n3863 & n3865 ;
  assign n3867 = n1995 & ~n3866 ;
  assign n3868 = ~n3862 & n3867 ;
  assign n3869 = n3859 & ~n3868 ;
  assign n3870 = \u5_tmr2_done_reg/NET0131  & ~n2820 ;
  assign n3871 = n1281 & n3870 ;
  assign n3872 = \u5_tmr_done_reg/NET0131  & ~n1899 ;
  assign n3873 = n1438 & n3872 ;
  assign n3874 = ~n1167 & ~n3873 ;
  assign n3875 = ~n3871 & n3874 ;
  assign n3876 = \u5_wb_cycle_reg/NET0131  & ~n3875 ;
  assign n3877 = ~n1092 & ~n1411 ;
  assign n3878 = ~n3094 & n3877 ;
  assign n3879 = ~n2708 & n3864 ;
  assign n3880 = n1443 & n3879 ;
  assign n3881 = \u4_rfr_req_reg/NET0131  & \u5_wb_stb_first_reg/NET0131  ;
  assign n3882 = n1309 & n3881 ;
  assign n3883 = n1308 & n3882 ;
  assign n3884 = ~n1171 & ~n1180 ;
  assign n3885 = ~n3883 & n3884 ;
  assign n3886 = ~n3880 & n3885 ;
  assign n3887 = n3878 & n3886 ;
  assign n3888 = ~n3876 & n3887 ;
  assign n3889 = ~n3869 & n3888 ;
  assign n3890 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[0]/NET0131  ;
  assign n3891 = n3889 & n3890 ;
  assign n3892 = ~n3857 & ~n3891 ;
  assign n3893 = ~\u0_rf_we_reg/NET0131  & n3889 ;
  assign n3894 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[0]/P0001  ;
  assign n3895 = ~\u0_spec_req_cs_reg[0]/NET0131  & \u0_spec_req_cs_reg[1]/NET0131  ;
  assign n3896 = \u0_u1_tms_reg[0]/P0001  & n3895 ;
  assign n3897 = ~n3894 & ~n3896 ;
  assign n3898 = n1045 & ~n3897 ;
  assign n3899 = ~n3893 & n3898 ;
  assign n3900 = n3892 & ~n3899 ;
  assign n3901 = \u0_sp_tms_reg[10]/NET0131  & ~n1045 ;
  assign n3902 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[10]/NET0131  ;
  assign n3903 = n3889 & n3902 ;
  assign n3904 = ~n3901 & ~n3903 ;
  assign n3905 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[10]/P0001  ;
  assign n3906 = \u0_u1_tms_reg[10]/P0001  & n3895 ;
  assign n3907 = ~n3905 & ~n3906 ;
  assign n3908 = n1045 & ~n3907 ;
  assign n3909 = ~n3893 & n3908 ;
  assign n3910 = n3904 & ~n3909 ;
  assign n3911 = \u0_sp_tms_reg[11]/NET0131  & ~n1045 ;
  assign n3912 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[11]/NET0131  ;
  assign n3913 = n3889 & n3912 ;
  assign n3914 = ~n3911 & ~n3913 ;
  assign n3915 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[11]/P0001  ;
  assign n3916 = \u0_u1_tms_reg[11]/P0001  & n3895 ;
  assign n3917 = ~n3915 & ~n3916 ;
  assign n3918 = n1045 & ~n3917 ;
  assign n3919 = ~n3893 & n3918 ;
  assign n3920 = n3914 & ~n3919 ;
  assign n3921 = \u0_sp_tms_reg[12]/NET0131  & ~n1045 ;
  assign n3922 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[12]/NET0131  ;
  assign n3923 = n3889 & n3922 ;
  assign n3924 = ~n3921 & ~n3923 ;
  assign n3925 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[12]/P0001  ;
  assign n3926 = \u0_u1_tms_reg[12]/P0001  & n3895 ;
  assign n3927 = ~n3925 & ~n3926 ;
  assign n3928 = n1045 & ~n3927 ;
  assign n3929 = ~n3893 & n3928 ;
  assign n3930 = n3924 & ~n3929 ;
  assign n3931 = \u0_sp_tms_reg[14]/NET0131  & ~n1045 ;
  assign n3932 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[14]/NET0131  ;
  assign n3933 = n3889 & n3932 ;
  assign n3934 = ~n3931 & ~n3933 ;
  assign n3935 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[14]/P0001  ;
  assign n3936 = \u0_u1_tms_reg[14]/P0001  & n3895 ;
  assign n3937 = ~n3935 & ~n3936 ;
  assign n3938 = n1045 & ~n3937 ;
  assign n3939 = ~n3893 & n3938 ;
  assign n3940 = n3934 & ~n3939 ;
  assign n3941 = \u0_sp_tms_reg[13]/NET0131  & ~n1045 ;
  assign n3942 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[13]/NET0131  ;
  assign n3943 = n3889 & n3942 ;
  assign n3944 = ~n3941 & ~n3943 ;
  assign n3945 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[13]/P0001  ;
  assign n3946 = \u0_u1_tms_reg[13]/P0001  & n3895 ;
  assign n3947 = ~n3945 & ~n3946 ;
  assign n3948 = n1045 & ~n3947 ;
  assign n3949 = ~n3893 & n3948 ;
  assign n3950 = n3944 & ~n3949 ;
  assign n3951 = \u0_sp_tms_reg[16]/NET0131  & ~n1045 ;
  assign n3952 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[16]/NET0131  ;
  assign n3953 = n3889 & n3952 ;
  assign n3954 = ~n3951 & ~n3953 ;
  assign n3955 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[16]/P0001  ;
  assign n3956 = \u0_u1_tms_reg[16]/P0001  & n3895 ;
  assign n3957 = ~n3955 & ~n3956 ;
  assign n3958 = n1045 & ~n3957 ;
  assign n3959 = ~n3893 & n3958 ;
  assign n3960 = n3954 & ~n3959 ;
  assign n3961 = \u0_sp_tms_reg[17]/NET0131  & ~n1045 ;
  assign n3962 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[17]/NET0131  ;
  assign n3963 = n3889 & n3962 ;
  assign n3964 = ~n3961 & ~n3963 ;
  assign n3965 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[17]/P0001  ;
  assign n3966 = \u0_u1_tms_reg[17]/P0001  & n3895 ;
  assign n3967 = ~n3965 & ~n3966 ;
  assign n3968 = n1045 & ~n3967 ;
  assign n3969 = ~n3893 & n3968 ;
  assign n3970 = n3964 & ~n3969 ;
  assign n3971 = \u0_sp_tms_reg[18]/NET0131  & ~n1045 ;
  assign n3972 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[18]/NET0131  ;
  assign n3973 = n3889 & n3972 ;
  assign n3974 = ~n3971 & ~n3973 ;
  assign n3975 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[18]/P0001  ;
  assign n3976 = \u0_u1_tms_reg[18]/P0001  & n3895 ;
  assign n3977 = ~n3975 & ~n3976 ;
  assign n3978 = n1045 & ~n3977 ;
  assign n3979 = ~n3893 & n3978 ;
  assign n3980 = n3974 & ~n3979 ;
  assign n3981 = \u0_sp_tms_reg[19]/NET0131  & ~n1045 ;
  assign n3982 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[19]/NET0131  ;
  assign n3983 = n3889 & n3982 ;
  assign n3984 = ~n3981 & ~n3983 ;
  assign n3985 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[19]/P0001  ;
  assign n3986 = \u0_u1_tms_reg[19]/P0001  & n3895 ;
  assign n3987 = ~n3985 & ~n3986 ;
  assign n3988 = n1045 & ~n3987 ;
  assign n3989 = ~n3893 & n3988 ;
  assign n3990 = n3984 & ~n3989 ;
  assign n3991 = \u0_sp_tms_reg[15]/NET0131  & ~n1045 ;
  assign n3992 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[15]/NET0131  ;
  assign n3993 = n3889 & n3992 ;
  assign n3994 = ~n3991 & ~n3993 ;
  assign n3995 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[15]/P0001  ;
  assign n3996 = \u0_u1_tms_reg[15]/P0001  & n3895 ;
  assign n3997 = ~n3995 & ~n3996 ;
  assign n3998 = n1045 & ~n3997 ;
  assign n3999 = ~n3893 & n3998 ;
  assign n4000 = n3994 & ~n3999 ;
  assign n4001 = \u0_sp_tms_reg[1]/NET0131  & ~n1045 ;
  assign n4002 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[1]/NET0131  ;
  assign n4003 = n3889 & n4002 ;
  assign n4004 = ~n4001 & ~n4003 ;
  assign n4005 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[1]/P0001  ;
  assign n4006 = \u0_u1_tms_reg[1]/P0001  & n3895 ;
  assign n4007 = ~n4005 & ~n4006 ;
  assign n4008 = n1045 & ~n4007 ;
  assign n4009 = ~n3893 & n4008 ;
  assign n4010 = n4004 & ~n4009 ;
  assign n4011 = \u0_sp_tms_reg[21]/NET0131  & ~n1045 ;
  assign n4012 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[21]/NET0131  ;
  assign n4013 = n3889 & n4012 ;
  assign n4014 = ~n4011 & ~n4013 ;
  assign n4015 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[21]/P0001  ;
  assign n4016 = \u0_u1_tms_reg[21]/P0001  & n3895 ;
  assign n4017 = ~n4015 & ~n4016 ;
  assign n4018 = n1045 & ~n4017 ;
  assign n4019 = ~n3893 & n4018 ;
  assign n4020 = n4014 & ~n4019 ;
  assign n4021 = \u0_sp_tms_reg[20]/NET0131  & ~n1045 ;
  assign n4022 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[20]/NET0131  ;
  assign n4023 = n3889 & n4022 ;
  assign n4024 = ~n4021 & ~n4023 ;
  assign n4025 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[20]/P0001  ;
  assign n4026 = \u0_u1_tms_reg[20]/P0001  & n3895 ;
  assign n4027 = ~n4025 & ~n4026 ;
  assign n4028 = n1045 & ~n4027 ;
  assign n4029 = ~n3893 & n4028 ;
  assign n4030 = n4024 & ~n4029 ;
  assign n4031 = \u0_sp_tms_reg[22]/NET0131  & ~n1045 ;
  assign n4032 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[22]/NET0131  ;
  assign n4033 = n3889 & n4032 ;
  assign n4034 = ~n4031 & ~n4033 ;
  assign n4035 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[22]/P0001  ;
  assign n4036 = \u0_u1_tms_reg[22]/P0001  & n3895 ;
  assign n4037 = ~n4035 & ~n4036 ;
  assign n4038 = n1045 & ~n4037 ;
  assign n4039 = ~n3893 & n4038 ;
  assign n4040 = n4034 & ~n4039 ;
  assign n4041 = \u0_sp_tms_reg[23]/NET0131  & ~n1045 ;
  assign n4042 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[23]/NET0131  ;
  assign n4043 = n3889 & n4042 ;
  assign n4044 = ~n4041 & ~n4043 ;
  assign n4045 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[23]/P0001  ;
  assign n4046 = \u0_u1_tms_reg[23]/P0001  & n3895 ;
  assign n4047 = ~n4045 & ~n4046 ;
  assign n4048 = n1045 & ~n4047 ;
  assign n4049 = ~n3893 & n4048 ;
  assign n4050 = n4044 & ~n4049 ;
  assign n4051 = \u0_sp_tms_reg[24]/NET0131  & ~n1045 ;
  assign n4052 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[24]/NET0131  ;
  assign n4053 = n3889 & n4052 ;
  assign n4054 = ~n4051 & ~n4053 ;
  assign n4055 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[24]/P0001  ;
  assign n4056 = \u0_u1_tms_reg[24]/P0001  & n3895 ;
  assign n4057 = ~n4055 & ~n4056 ;
  assign n4058 = n1045 & ~n4057 ;
  assign n4059 = ~n3893 & n4058 ;
  assign n4060 = n4054 & ~n4059 ;
  assign n4061 = \u0_sp_tms_reg[25]/NET0131  & ~n1045 ;
  assign n4062 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[25]/NET0131  ;
  assign n4063 = n3889 & n4062 ;
  assign n4064 = ~n4061 & ~n4063 ;
  assign n4065 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[25]/P0001  ;
  assign n4066 = \u0_u1_tms_reg[25]/P0001  & n3895 ;
  assign n4067 = ~n4065 & ~n4066 ;
  assign n4068 = n1045 & ~n4067 ;
  assign n4069 = ~n3893 & n4068 ;
  assign n4070 = n4064 & ~n4069 ;
  assign n4071 = \u0_sp_tms_reg[26]/NET0131  & ~n1045 ;
  assign n4072 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[26]/NET0131  ;
  assign n4073 = n3889 & n4072 ;
  assign n4074 = ~n4071 & ~n4073 ;
  assign n4075 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[26]/P0001  ;
  assign n4076 = \u0_u1_tms_reg[26]/P0001  & n3895 ;
  assign n4077 = ~n4075 & ~n4076 ;
  assign n4078 = n1045 & ~n4077 ;
  assign n4079 = ~n3893 & n4078 ;
  assign n4080 = n4074 & ~n4079 ;
  assign n4081 = \u0_sp_tms_reg[27]/NET0131  & ~n1045 ;
  assign n4082 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[27]/NET0131  ;
  assign n4083 = n3889 & n4082 ;
  assign n4084 = ~n4081 & ~n4083 ;
  assign n4085 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[27]/P0001  ;
  assign n4086 = \u0_u1_tms_reg[27]/P0001  & n3895 ;
  assign n4087 = ~n4085 & ~n4086 ;
  assign n4088 = n1045 & ~n4087 ;
  assign n4089 = ~n3893 & n4088 ;
  assign n4090 = n4084 & ~n4089 ;
  assign n4091 = \u0_sp_tms_reg[2]/NET0131  & ~n1045 ;
  assign n4092 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[2]/NET0131  ;
  assign n4093 = n3889 & n4092 ;
  assign n4094 = ~n4091 & ~n4093 ;
  assign n4095 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[2]/P0001  ;
  assign n4096 = \u0_u1_tms_reg[2]/P0001  & n3895 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4098 = n1045 & ~n4097 ;
  assign n4099 = ~n3893 & n4098 ;
  assign n4100 = n4094 & ~n4099 ;
  assign n4101 = \u0_sp_tms_reg[3]/NET0131  & ~n1045 ;
  assign n4102 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[3]/NET0131  ;
  assign n4103 = n3889 & n4102 ;
  assign n4104 = ~n4101 & ~n4103 ;
  assign n4105 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[3]/P0001  ;
  assign n4106 = \u0_u1_tms_reg[3]/P0001  & n3895 ;
  assign n4107 = ~n4105 & ~n4106 ;
  assign n4108 = n1045 & ~n4107 ;
  assign n4109 = ~n3893 & n4108 ;
  assign n4110 = n4104 & ~n4109 ;
  assign n4111 = \u0_sp_tms_reg[4]/NET0131  & ~n1045 ;
  assign n4112 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[4]/NET0131  ;
  assign n4113 = n3889 & n4112 ;
  assign n4114 = ~n4111 & ~n4113 ;
  assign n4115 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[4]/P0001  ;
  assign n4116 = \u0_u1_tms_reg[4]/P0001  & n3895 ;
  assign n4117 = ~n4115 & ~n4116 ;
  assign n4118 = n1045 & ~n4117 ;
  assign n4119 = ~n3893 & n4118 ;
  assign n4120 = n4114 & ~n4119 ;
  assign n4121 = \u0_sp_tms_reg[5]/NET0131  & ~n1045 ;
  assign n4122 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[5]/NET0131  ;
  assign n4123 = n3889 & n4122 ;
  assign n4124 = ~n4121 & ~n4123 ;
  assign n4125 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[5]/P0001  ;
  assign n4126 = \u0_u1_tms_reg[5]/P0001  & n3895 ;
  assign n4127 = ~n4125 & ~n4126 ;
  assign n4128 = n1045 & ~n4127 ;
  assign n4129 = ~n3893 & n4128 ;
  assign n4130 = n4124 & ~n4129 ;
  assign n4131 = \u0_sp_tms_reg[7]/NET0131  & ~n1045 ;
  assign n4132 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[7]/NET0131  ;
  assign n4133 = n3889 & n4132 ;
  assign n4134 = ~n4131 & ~n4133 ;
  assign n4135 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[7]/P0001  ;
  assign n4136 = \u0_u1_tms_reg[7]/P0001  & n3895 ;
  assign n4137 = ~n4135 & ~n4136 ;
  assign n4138 = n1045 & ~n4137 ;
  assign n4139 = ~n3893 & n4138 ;
  assign n4140 = n4134 & ~n4139 ;
  assign n4141 = \u0_sp_tms_reg[6]/NET0131  & ~n1045 ;
  assign n4142 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[6]/NET0131  ;
  assign n4143 = n3889 & n4142 ;
  assign n4144 = ~n4141 & ~n4143 ;
  assign n4145 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[6]/P0001  ;
  assign n4146 = \u0_u1_tms_reg[6]/P0001  & n3895 ;
  assign n4147 = ~n4145 & ~n4146 ;
  assign n4148 = n1045 & ~n4147 ;
  assign n4149 = ~n3893 & n4148 ;
  assign n4150 = n4144 & ~n4149 ;
  assign n4151 = \u0_sp_tms_reg[8]/NET0131  & ~n1045 ;
  assign n4152 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[8]/NET0131  ;
  assign n4153 = n3889 & n4152 ;
  assign n4154 = ~n4151 & ~n4153 ;
  assign n4155 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[8]/P0001  ;
  assign n4156 = \u0_u1_tms_reg[8]/P0001  & n3895 ;
  assign n4157 = ~n4155 & ~n4156 ;
  assign n4158 = n1045 & ~n4157 ;
  assign n4159 = ~n3893 & n4158 ;
  assign n4160 = n4154 & ~n4159 ;
  assign n4161 = \u0_sp_tms_reg[9]/NET0131  & ~n1045 ;
  assign n4162 = ~\u0_rf_we_reg/NET0131  & \u0_sp_tms_reg[9]/NET0131  ;
  assign n4163 = n3889 & n4162 ;
  assign n4164 = ~n4161 & ~n4163 ;
  assign n4165 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_tms_reg[9]/P0001  ;
  assign n4166 = \u0_u1_tms_reg[9]/P0001  & n3895 ;
  assign n4167 = ~n4165 & ~n4166 ;
  assign n4168 = n1045 & ~n4167 ;
  assign n4169 = ~n3893 & n4168 ;
  assign n4170 = n4164 & ~n4169 ;
  assign n4171 = \u0_tms_reg[10]/NET0131  & ~n1045 ;
  assign n4172 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[10]/NET0131  ;
  assign n4173 = n3889 & n4172 ;
  assign n4174 = ~n4171 & ~n4173 ;
  assign n4175 = \u0_u0_csc_reg[18]/P0001  & \wb_addr_i[23]_pad  ;
  assign n4176 = ~\u0_u0_csc_reg[18]/P0001  & ~\wb_addr_i[23]_pad  ;
  assign n4177 = \u0_csc_mask_r_reg[2]/NET0131  & ~n4176 ;
  assign n4178 = ~n4175 & n4177 ;
  assign n4179 = \u0_u0_csc_reg[0]/NET0131  & ~n4178 ;
  assign n4180 = \u0_u0_csc_reg[20]/P0001  & ~\wb_addr_i[25]_pad  ;
  assign n4181 = ~\u0_u0_csc_reg[20]/P0001  & \wb_addr_i[25]_pad  ;
  assign n4182 = ~n4180 & ~n4181 ;
  assign n4183 = \u0_csc_mask_r_reg[4]/NET0131  & ~n4182 ;
  assign n4184 = \u0_u0_csc_reg[22]/P0001  & \wb_addr_i[27]_pad  ;
  assign n4185 = ~\u0_u0_csc_reg[22]/P0001  & ~\wb_addr_i[27]_pad  ;
  assign n4186 = \u0_csc_mask_r_reg[6]/NET0131  & ~n4185 ;
  assign n4187 = ~n4184 & n4186 ;
  assign n4188 = ~n4183 & ~n4187 ;
  assign n4189 = \u0_u0_csc_reg[23]/P0001  & \wb_addr_i[28]_pad  ;
  assign n4190 = ~\u0_u0_csc_reg[23]/P0001  & ~\wb_addr_i[28]_pad  ;
  assign n4191 = \u0_csc_mask_r_reg[7]/NET0131  & ~n4190 ;
  assign n4192 = ~n4189 & n4191 ;
  assign n4193 = \u0_u0_csc_reg[17]/P0001  & \wb_addr_i[22]_pad  ;
  assign n4194 = ~\u0_u0_csc_reg[17]/P0001  & ~\wb_addr_i[22]_pad  ;
  assign n4195 = \u0_csc_mask_r_reg[1]/NET0131  & ~n4194 ;
  assign n4196 = ~n4193 & n4195 ;
  assign n4197 = ~n4192 & ~n4196 ;
  assign n4198 = n4188 & n4197 ;
  assign n4199 = n4179 & n4198 ;
  assign n4200 = \u0_u0_csc_reg[8]/P0001  & wb_we_i_pad ;
  assign n4201 = \u0_u0_csc_reg[21]/P0001  & \wb_addr_i[26]_pad  ;
  assign n4202 = ~\u0_u0_csc_reg[21]/P0001  & ~\wb_addr_i[26]_pad  ;
  assign n4203 = \u0_csc_mask_r_reg[5]/NET0131  & ~n4202 ;
  assign n4204 = ~n4201 & n4203 ;
  assign n4205 = \u0_u0_csc_reg[16]/P0001  & \wb_addr_i[21]_pad  ;
  assign n4206 = ~\u0_u0_csc_reg[16]/P0001  & ~\wb_addr_i[21]_pad  ;
  assign n4207 = \u0_csc_mask_r_reg[0]/NET0131  & ~n4206 ;
  assign n4208 = ~n4205 & n4207 ;
  assign n4209 = \u0_u0_csc_reg[19]/P0001  & \wb_addr_i[24]_pad  ;
  assign n4210 = ~\u0_u0_csc_reg[19]/P0001  & ~\wb_addr_i[24]_pad  ;
  assign n4211 = \u0_csc_mask_r_reg[3]/NET0131  & ~n4210 ;
  assign n4212 = ~n4209 & n4211 ;
  assign n4213 = ~n4208 & ~n4212 ;
  assign n4214 = ~n4204 & n4213 ;
  assign n4215 = ~n4200 & n4214 ;
  assign n4216 = n4199 & n4215 ;
  assign n4217 = \u0_u1_csc_reg[17]/P0001  & \wb_addr_i[22]_pad  ;
  assign n4218 = ~\u0_u1_csc_reg[17]/P0001  & ~\wb_addr_i[22]_pad  ;
  assign n4219 = \u0_csc_mask_r_reg[1]/NET0131  & ~n4218 ;
  assign n4220 = ~n4217 & n4219 ;
  assign n4221 = \u0_u1_csc_reg[0]/NET0131  & ~n4220 ;
  assign n4222 = \u0_u1_csc_reg[21]/P0001  & ~\wb_addr_i[26]_pad  ;
  assign n4223 = ~\u0_u1_csc_reg[21]/P0001  & \wb_addr_i[26]_pad  ;
  assign n4224 = ~n4222 & ~n4223 ;
  assign n4225 = \u0_csc_mask_r_reg[5]/NET0131  & ~n4224 ;
  assign n4226 = \u0_u1_csc_reg[22]/P0001  & \wb_addr_i[27]_pad  ;
  assign n4227 = ~\u0_u1_csc_reg[22]/P0001  & ~\wb_addr_i[27]_pad  ;
  assign n4228 = \u0_csc_mask_r_reg[6]/NET0131  & ~n4227 ;
  assign n4229 = ~n4226 & n4228 ;
  assign n4230 = ~n4225 & ~n4229 ;
  assign n4231 = \u0_u1_csc_reg[19]/P0001  & \wb_addr_i[24]_pad  ;
  assign n4232 = ~\u0_u1_csc_reg[19]/P0001  & ~\wb_addr_i[24]_pad  ;
  assign n4233 = \u0_csc_mask_r_reg[3]/NET0131  & ~n4232 ;
  assign n4234 = ~n4231 & n4233 ;
  assign n4235 = \u0_u1_csc_reg[16]/P0001  & \wb_addr_i[21]_pad  ;
  assign n4236 = ~\u0_u1_csc_reg[16]/P0001  & ~\wb_addr_i[21]_pad  ;
  assign n4237 = \u0_csc_mask_r_reg[0]/NET0131  & ~n4236 ;
  assign n4238 = ~n4235 & n4237 ;
  assign n4239 = ~n4234 & ~n4238 ;
  assign n4240 = n4230 & n4239 ;
  assign n4241 = n4221 & n4240 ;
  assign n4242 = \u0_u1_csc_reg[8]/P0001  & wb_we_i_pad ;
  assign n4243 = \u0_u1_csc_reg[20]/P0001  & \wb_addr_i[25]_pad  ;
  assign n4244 = ~\u0_u1_csc_reg[20]/P0001  & ~\wb_addr_i[25]_pad  ;
  assign n4245 = \u0_csc_mask_r_reg[4]/NET0131  & ~n4244 ;
  assign n4246 = ~n4243 & n4245 ;
  assign n4247 = \u0_u1_csc_reg[18]/P0001  & \wb_addr_i[23]_pad  ;
  assign n4248 = ~\u0_u1_csc_reg[18]/P0001  & ~\wb_addr_i[23]_pad  ;
  assign n4249 = \u0_csc_mask_r_reg[2]/NET0131  & ~n4248 ;
  assign n4250 = ~n4247 & n4249 ;
  assign n4251 = \u0_u1_csc_reg[23]/P0001  & \wb_addr_i[28]_pad  ;
  assign n4252 = ~\u0_u1_csc_reg[23]/P0001  & ~\wb_addr_i[28]_pad  ;
  assign n4253 = \u0_csc_mask_r_reg[7]/NET0131  & ~n4252 ;
  assign n4254 = ~n4251 & n4253 ;
  assign n4255 = ~n4250 & ~n4254 ;
  assign n4256 = ~n4246 & n4255 ;
  assign n4257 = ~n4242 & n4256 ;
  assign n4258 = n4241 & n4257 ;
  assign n4259 = ~n4216 & n4258 ;
  assign n4260 = \u0_u1_tms_reg[10]/P0001  & n4259 ;
  assign n4261 = \u0_u0_tms_reg[10]/P0001  & ~n4200 ;
  assign n4262 = n4214 & n4261 ;
  assign n4263 = n4199 & n4262 ;
  assign n4264 = ~n4260 & ~n4263 ;
  assign n4265 = n1045 & ~n4264 ;
  assign n4266 = ~n3893 & n4265 ;
  assign n4267 = n4174 & ~n4266 ;
  assign n4268 = \u0_tms_reg[11]/NET0131  & ~n1045 ;
  assign n4269 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[11]/NET0131  ;
  assign n4270 = n3889 & n4269 ;
  assign n4271 = ~n4268 & ~n4270 ;
  assign n4272 = \u0_u1_tms_reg[11]/P0001  & n4259 ;
  assign n4273 = \u0_u0_tms_reg[11]/P0001  & ~n4200 ;
  assign n4274 = n4214 & n4273 ;
  assign n4275 = n4199 & n4274 ;
  assign n4276 = ~n4272 & ~n4275 ;
  assign n4277 = n1045 & ~n4276 ;
  assign n4278 = ~n3893 & n4277 ;
  assign n4279 = n4271 & ~n4278 ;
  assign n4280 = \u0_tms_reg[12]/NET0131  & ~n1045 ;
  assign n4281 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[12]/NET0131  ;
  assign n4282 = n3889 & n4281 ;
  assign n4283 = ~n4280 & ~n4282 ;
  assign n4284 = \u0_u1_tms_reg[12]/P0001  & n4259 ;
  assign n4285 = \u0_u0_tms_reg[12]/P0001  & ~n4200 ;
  assign n4286 = n4214 & n4285 ;
  assign n4287 = n4199 & n4286 ;
  assign n4288 = ~n4284 & ~n4287 ;
  assign n4289 = n1045 & ~n4288 ;
  assign n4290 = ~n3893 & n4289 ;
  assign n4291 = n4283 & ~n4290 ;
  assign n4292 = \u0_tms_reg[13]/NET0131  & ~n1045 ;
  assign n4293 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[13]/NET0131  ;
  assign n4294 = n3889 & n4293 ;
  assign n4295 = ~n4292 & ~n4294 ;
  assign n4296 = \u0_u1_tms_reg[13]/P0001  & n4259 ;
  assign n4297 = \u0_u0_tms_reg[13]/P0001  & ~n4200 ;
  assign n4298 = n4214 & n4297 ;
  assign n4299 = n4199 & n4298 ;
  assign n4300 = ~n4296 & ~n4299 ;
  assign n4301 = n1045 & ~n4300 ;
  assign n4302 = ~n3893 & n4301 ;
  assign n4303 = n4295 & ~n4302 ;
  assign n4304 = \u0_tms_reg[0]/NET0131  & ~n1045 ;
  assign n4305 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[0]/NET0131  ;
  assign n4306 = n3889 & n4305 ;
  assign n4307 = ~n4304 & ~n4306 ;
  assign n4308 = \u0_u1_tms_reg[0]/P0001  & n4259 ;
  assign n4309 = \u0_u0_tms_reg[0]/P0001  & ~n4200 ;
  assign n4310 = n4214 & n4309 ;
  assign n4311 = n4199 & n4310 ;
  assign n4312 = ~n4308 & ~n4311 ;
  assign n4313 = n1045 & ~n4312 ;
  assign n4314 = ~n3893 & n4313 ;
  assign n4315 = n4307 & ~n4314 ;
  assign n4316 = \u0_tms_reg[14]/NET0131  & ~n1045 ;
  assign n4317 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[14]/NET0131  ;
  assign n4318 = n3889 & n4317 ;
  assign n4319 = ~n4316 & ~n4318 ;
  assign n4320 = \u0_u1_tms_reg[14]/P0001  & n4259 ;
  assign n4321 = \u0_u0_tms_reg[14]/P0001  & ~n4200 ;
  assign n4322 = n4214 & n4321 ;
  assign n4323 = n4199 & n4322 ;
  assign n4324 = ~n4320 & ~n4323 ;
  assign n4325 = n1045 & ~n4324 ;
  assign n4326 = ~n3893 & n4325 ;
  assign n4327 = n4319 & ~n4326 ;
  assign n4328 = \u0_tms_reg[15]/NET0131  & ~n1045 ;
  assign n4329 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[15]/NET0131  ;
  assign n4330 = n3889 & n4329 ;
  assign n4331 = ~n4328 & ~n4330 ;
  assign n4332 = \u0_u1_tms_reg[15]/P0001  & n4259 ;
  assign n4333 = \u0_u0_tms_reg[15]/P0001  & ~n4200 ;
  assign n4334 = n4214 & n4333 ;
  assign n4335 = n4199 & n4334 ;
  assign n4336 = ~n4332 & ~n4335 ;
  assign n4337 = n1045 & ~n4336 ;
  assign n4338 = ~n3893 & n4337 ;
  assign n4339 = n4331 & ~n4338 ;
  assign n4340 = \u0_tms_reg[16]/NET0131  & ~n1045 ;
  assign n4341 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[16]/NET0131  ;
  assign n4342 = n3889 & n4341 ;
  assign n4343 = ~n4340 & ~n4342 ;
  assign n4344 = \u0_u1_tms_reg[16]/P0001  & n4259 ;
  assign n4345 = \u0_u0_tms_reg[16]/P0001  & ~n4200 ;
  assign n4346 = n4214 & n4345 ;
  assign n4347 = n4199 & n4346 ;
  assign n4348 = ~n4344 & ~n4347 ;
  assign n4349 = n1045 & ~n4348 ;
  assign n4350 = ~n3893 & n4349 ;
  assign n4351 = n4343 & ~n4350 ;
  assign n4352 = \u0_tms_reg[17]/NET0131  & ~n1045 ;
  assign n4353 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[17]/NET0131  ;
  assign n4354 = n3889 & n4353 ;
  assign n4355 = ~n4352 & ~n4354 ;
  assign n4356 = \u0_u1_tms_reg[17]/P0001  & n4259 ;
  assign n4357 = \u0_u0_tms_reg[17]/P0001  & ~n4200 ;
  assign n4358 = n4214 & n4357 ;
  assign n4359 = n4199 & n4358 ;
  assign n4360 = ~n4356 & ~n4359 ;
  assign n4361 = n1045 & ~n4360 ;
  assign n4362 = ~n3893 & n4361 ;
  assign n4363 = n4355 & ~n4362 ;
  assign n4364 = \u0_tms_reg[18]/NET0131  & ~n1045 ;
  assign n4365 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[18]/NET0131  ;
  assign n4366 = n3889 & n4365 ;
  assign n4367 = ~n4364 & ~n4366 ;
  assign n4368 = \u0_u1_tms_reg[18]/P0001  & n4259 ;
  assign n4369 = \u0_u0_tms_reg[18]/P0001  & ~n4200 ;
  assign n4370 = n4214 & n4369 ;
  assign n4371 = n4199 & n4370 ;
  assign n4372 = ~n4368 & ~n4371 ;
  assign n4373 = n1045 & ~n4372 ;
  assign n4374 = ~n3893 & n4373 ;
  assign n4375 = n4367 & ~n4374 ;
  assign n4376 = \u0_tms_reg[19]/NET0131  & ~n1045 ;
  assign n4377 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[19]/NET0131  ;
  assign n4378 = n3889 & n4377 ;
  assign n4379 = ~n4376 & ~n4378 ;
  assign n4380 = \u0_u1_tms_reg[19]/P0001  & n4259 ;
  assign n4381 = \u0_u0_tms_reg[19]/P0001  & ~n4200 ;
  assign n4382 = n4214 & n4381 ;
  assign n4383 = n4199 & n4382 ;
  assign n4384 = ~n4380 & ~n4383 ;
  assign n4385 = n1045 & ~n4384 ;
  assign n4386 = ~n3893 & n4385 ;
  assign n4387 = n4379 & ~n4386 ;
  assign n4388 = \u0_tms_reg[1]/NET0131  & ~n1045 ;
  assign n4389 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[1]/NET0131  ;
  assign n4390 = n3889 & n4389 ;
  assign n4391 = ~n4388 & ~n4390 ;
  assign n4392 = \u0_u1_tms_reg[1]/P0001  & n4259 ;
  assign n4393 = \u0_u0_tms_reg[1]/P0001  & ~n4200 ;
  assign n4394 = n4214 & n4393 ;
  assign n4395 = n4199 & n4394 ;
  assign n4396 = ~n4392 & ~n4395 ;
  assign n4397 = n1045 & ~n4396 ;
  assign n4398 = ~n3893 & n4397 ;
  assign n4399 = n4391 & ~n4398 ;
  assign n4400 = \u0_tms_reg[20]/NET0131  & ~n1045 ;
  assign n4401 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[20]/NET0131  ;
  assign n4402 = n3889 & n4401 ;
  assign n4403 = ~n4400 & ~n4402 ;
  assign n4404 = \u0_u1_tms_reg[20]/P0001  & n4259 ;
  assign n4405 = \u0_u0_tms_reg[20]/P0001  & ~n4200 ;
  assign n4406 = n4214 & n4405 ;
  assign n4407 = n4199 & n4406 ;
  assign n4408 = ~n4404 & ~n4407 ;
  assign n4409 = n1045 & ~n4408 ;
  assign n4410 = ~n3893 & n4409 ;
  assign n4411 = n4403 & ~n4410 ;
  assign n4412 = \u0_tms_reg[21]/NET0131  & ~n1045 ;
  assign n4413 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[21]/NET0131  ;
  assign n4414 = n3889 & n4413 ;
  assign n4415 = ~n4412 & ~n4414 ;
  assign n4416 = \u0_u1_tms_reg[21]/P0001  & n4259 ;
  assign n4417 = \u0_u0_tms_reg[21]/P0001  & ~n4200 ;
  assign n4418 = n4214 & n4417 ;
  assign n4419 = n4199 & n4418 ;
  assign n4420 = ~n4416 & ~n4419 ;
  assign n4421 = n1045 & ~n4420 ;
  assign n4422 = ~n3893 & n4421 ;
  assign n4423 = n4415 & ~n4422 ;
  assign n4424 = \u0_tms_reg[23]/NET0131  & ~n1045 ;
  assign n4425 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[23]/NET0131  ;
  assign n4426 = n3889 & n4425 ;
  assign n4427 = ~n4424 & ~n4426 ;
  assign n4428 = \u0_u1_tms_reg[23]/P0001  & n4259 ;
  assign n4429 = \u0_u0_tms_reg[23]/P0001  & ~n4200 ;
  assign n4430 = n4214 & n4429 ;
  assign n4431 = n4199 & n4430 ;
  assign n4432 = ~n4428 & ~n4431 ;
  assign n4433 = n1045 & ~n4432 ;
  assign n4434 = ~n3893 & n4433 ;
  assign n4435 = n4427 & ~n4434 ;
  assign n4436 = \u0_tms_reg[24]/NET0131  & ~n1045 ;
  assign n4437 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[24]/NET0131  ;
  assign n4438 = n3889 & n4437 ;
  assign n4439 = ~n4436 & ~n4438 ;
  assign n4440 = \u0_u1_tms_reg[24]/P0001  & n4259 ;
  assign n4441 = \u0_u0_tms_reg[24]/P0001  & ~n4200 ;
  assign n4442 = n4214 & n4441 ;
  assign n4443 = n4199 & n4442 ;
  assign n4444 = ~n4440 & ~n4443 ;
  assign n4445 = n1045 & ~n4444 ;
  assign n4446 = ~n3893 & n4445 ;
  assign n4447 = n4439 & ~n4446 ;
  assign n4448 = \u0_tms_reg[22]/NET0131  & ~n1045 ;
  assign n4449 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[22]/NET0131  ;
  assign n4450 = n3889 & n4449 ;
  assign n4451 = ~n4448 & ~n4450 ;
  assign n4452 = \u0_u1_tms_reg[22]/P0001  & n4259 ;
  assign n4453 = \u0_u0_tms_reg[22]/P0001  & ~n4200 ;
  assign n4454 = n4214 & n4453 ;
  assign n4455 = n4199 & n4454 ;
  assign n4456 = ~n4452 & ~n4455 ;
  assign n4457 = n1045 & ~n4456 ;
  assign n4458 = ~n3893 & n4457 ;
  assign n4459 = n4451 & ~n4458 ;
  assign n4460 = \u0_tms_reg[25]/NET0131  & ~n1045 ;
  assign n4461 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[25]/NET0131  ;
  assign n4462 = n3889 & n4461 ;
  assign n4463 = ~n4460 & ~n4462 ;
  assign n4464 = \u0_u1_tms_reg[25]/P0001  & n4259 ;
  assign n4465 = \u0_u0_tms_reg[25]/P0001  & ~n4200 ;
  assign n4466 = n4214 & n4465 ;
  assign n4467 = n4199 & n4466 ;
  assign n4468 = ~n4464 & ~n4467 ;
  assign n4469 = n1045 & ~n4468 ;
  assign n4470 = ~n3893 & n4469 ;
  assign n4471 = n4463 & ~n4470 ;
  assign n4472 = \u0_tms_reg[26]/NET0131  & ~n1045 ;
  assign n4473 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[26]/NET0131  ;
  assign n4474 = n3889 & n4473 ;
  assign n4475 = ~n4472 & ~n4474 ;
  assign n4476 = \u0_u1_tms_reg[26]/P0001  & n4259 ;
  assign n4477 = \u0_u0_tms_reg[26]/P0001  & ~n4200 ;
  assign n4478 = n4214 & n4477 ;
  assign n4479 = n4199 & n4478 ;
  assign n4480 = ~n4476 & ~n4479 ;
  assign n4481 = n1045 & ~n4480 ;
  assign n4482 = ~n3893 & n4481 ;
  assign n4483 = n4475 & ~n4482 ;
  assign n4484 = \u0_tms_reg[27]/NET0131  & ~n1045 ;
  assign n4485 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[27]/NET0131  ;
  assign n4486 = n3889 & n4485 ;
  assign n4487 = ~n4484 & ~n4486 ;
  assign n4488 = \u0_u1_tms_reg[27]/P0001  & n4259 ;
  assign n4489 = \u0_u0_tms_reg[27]/P0001  & ~n4200 ;
  assign n4490 = n4214 & n4489 ;
  assign n4491 = n4199 & n4490 ;
  assign n4492 = ~n4488 & ~n4491 ;
  assign n4493 = n1045 & ~n4492 ;
  assign n4494 = ~n3893 & n4493 ;
  assign n4495 = n4487 & ~n4494 ;
  assign n4496 = \u0_tms_reg[2]/NET0131  & ~n1045 ;
  assign n4497 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[2]/NET0131  ;
  assign n4498 = n3889 & n4497 ;
  assign n4499 = ~n4496 & ~n4498 ;
  assign n4500 = \u0_u1_tms_reg[2]/P0001  & n4259 ;
  assign n4501 = \u0_u0_tms_reg[2]/P0001  & ~n4200 ;
  assign n4502 = n4214 & n4501 ;
  assign n4503 = n4199 & n4502 ;
  assign n4504 = ~n4500 & ~n4503 ;
  assign n4505 = n1045 & ~n4504 ;
  assign n4506 = ~n3893 & n4505 ;
  assign n4507 = n4499 & ~n4506 ;
  assign n4508 = \u0_tms_reg[3]/NET0131  & ~n1045 ;
  assign n4509 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[3]/NET0131  ;
  assign n4510 = n3889 & n4509 ;
  assign n4511 = ~n4508 & ~n4510 ;
  assign n4512 = \u0_u1_tms_reg[3]/P0001  & n4259 ;
  assign n4513 = \u0_u0_tms_reg[3]/P0001  & ~n4200 ;
  assign n4514 = n4214 & n4513 ;
  assign n4515 = n4199 & n4514 ;
  assign n4516 = ~n4512 & ~n4515 ;
  assign n4517 = n1045 & ~n4516 ;
  assign n4518 = ~n3893 & n4517 ;
  assign n4519 = n4511 & ~n4518 ;
  assign n4520 = \u0_tms_reg[4]/NET0131  & ~n1045 ;
  assign n4521 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[4]/NET0131  ;
  assign n4522 = n3889 & n4521 ;
  assign n4523 = ~n4520 & ~n4522 ;
  assign n4524 = \u0_u1_tms_reg[4]/P0001  & n4259 ;
  assign n4525 = \u0_u0_tms_reg[4]/P0001  & ~n4200 ;
  assign n4526 = n4214 & n4525 ;
  assign n4527 = n4199 & n4526 ;
  assign n4528 = ~n4524 & ~n4527 ;
  assign n4529 = n1045 & ~n4528 ;
  assign n4530 = ~n3893 & n4529 ;
  assign n4531 = n4523 & ~n4530 ;
  assign n4532 = \u0_tms_reg[5]/NET0131  & ~n1045 ;
  assign n4533 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[5]/NET0131  ;
  assign n4534 = n3889 & n4533 ;
  assign n4535 = ~n4532 & ~n4534 ;
  assign n4536 = \u0_u1_tms_reg[5]/P0001  & n4259 ;
  assign n4537 = \u0_u0_tms_reg[5]/P0001  & ~n4200 ;
  assign n4538 = n4214 & n4537 ;
  assign n4539 = n4199 & n4538 ;
  assign n4540 = ~n4536 & ~n4539 ;
  assign n4541 = n1045 & ~n4540 ;
  assign n4542 = ~n3893 & n4541 ;
  assign n4543 = n4535 & ~n4542 ;
  assign n4544 = \u0_tms_reg[6]/NET0131  & ~n1045 ;
  assign n4545 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[6]/NET0131  ;
  assign n4546 = n3889 & n4545 ;
  assign n4547 = ~n4544 & ~n4546 ;
  assign n4548 = \u0_u1_tms_reg[6]/P0001  & n4259 ;
  assign n4549 = \u0_u0_tms_reg[6]/P0001  & ~n4200 ;
  assign n4550 = n4214 & n4549 ;
  assign n4551 = n4199 & n4550 ;
  assign n4552 = ~n4548 & ~n4551 ;
  assign n4553 = n1045 & ~n4552 ;
  assign n4554 = ~n3893 & n4553 ;
  assign n4555 = n4547 & ~n4554 ;
  assign n4556 = \u0_tms_reg[7]/NET0131  & ~n1045 ;
  assign n4557 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[7]/NET0131  ;
  assign n4558 = n3889 & n4557 ;
  assign n4559 = ~n4556 & ~n4558 ;
  assign n4560 = \u0_u1_tms_reg[7]/P0001  & n4259 ;
  assign n4561 = \u0_u0_tms_reg[7]/P0001  & ~n4200 ;
  assign n4562 = n4214 & n4561 ;
  assign n4563 = n4199 & n4562 ;
  assign n4564 = ~n4560 & ~n4563 ;
  assign n4565 = n1045 & ~n4564 ;
  assign n4566 = ~n3893 & n4565 ;
  assign n4567 = n4559 & ~n4566 ;
  assign n4568 = \u0_tms_reg[8]/NET0131  & ~n1045 ;
  assign n4569 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[8]/NET0131  ;
  assign n4570 = n3889 & n4569 ;
  assign n4571 = ~n4568 & ~n4570 ;
  assign n4572 = \u0_u1_tms_reg[8]/P0001  & n4259 ;
  assign n4573 = \u0_u0_tms_reg[8]/P0001  & ~n4200 ;
  assign n4574 = n4214 & n4573 ;
  assign n4575 = n4199 & n4574 ;
  assign n4576 = ~n4572 & ~n4575 ;
  assign n4577 = n1045 & ~n4576 ;
  assign n4578 = ~n3893 & n4577 ;
  assign n4579 = n4571 & ~n4578 ;
  assign n4580 = \u0_tms_reg[9]/NET0131  & ~n1045 ;
  assign n4581 = ~\u0_rf_we_reg/NET0131  & \u0_tms_reg[9]/NET0131  ;
  assign n4582 = n3889 & n4581 ;
  assign n4583 = ~n4580 & ~n4582 ;
  assign n4584 = \u0_u1_tms_reg[9]/P0001  & n4259 ;
  assign n4585 = \u0_u0_tms_reg[9]/P0001  & ~n4200 ;
  assign n4586 = n4214 & n4585 ;
  assign n4587 = n4199 & n4586 ;
  assign n4588 = ~n4584 & ~n4587 ;
  assign n4589 = n1045 & ~n4588 ;
  assign n4590 = ~n3893 & n4589 ;
  assign n4591 = n4583 & ~n4590 ;
  assign n4592 = ~n2613 & n3372 ;
  assign n4593 = \u0_tms_reg[6]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n4594 = ~\u5_lmr_ack_reg/NET0131  & n4593 ;
  assign n4595 = n983 & n4594 ;
  assign n4596 = \u0_sp_tms_reg[6]/NET0131  & ~n1200 ;
  assign n4597 = ~n4595 & ~n4596 ;
  assign n4598 = ~n3400 & n4597 ;
  assign n4599 = n1851 & n4598 ;
  assign n4600 = ~n1848 & n4599 ;
  assign n4601 = \u5_timer2_reg[7]/P0001  & ~n3396 ;
  assign n4602 = ~\u5_timer2_reg[7]/P0001  & \u5_timer2_reg[8]/P0001  ;
  assign n4603 = n3396 & n4602 ;
  assign n4604 = ~n4601 & ~n4603 ;
  assign n4605 = n3400 & n4604 ;
  assign n4606 = n3390 & ~n4605 ;
  assign n4607 = n3634 & n4606 ;
  assign n4608 = ~n4600 & n4607 ;
  assign n4609 = ~n4592 & ~n4608 ;
  assign n4610 = n3372 & ~n3661 ;
  assign n4611 = \u0_tms_reg[7]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n4612 = ~\u5_lmr_ack_reg/NET0131  & n4611 ;
  assign n4613 = n983 & n4612 ;
  assign n4614 = \u0_sp_tms_reg[7]/NET0131  & ~n1200 ;
  assign n4615 = ~n4613 & ~n4614 ;
  assign n4616 = ~n3400 & n4615 ;
  assign n4617 = n1851 & n4616 ;
  assign n4618 = ~n1848 & n4617 ;
  assign n4619 = ~\u5_timer2_reg[8]/P0001  & n3400 ;
  assign n4620 = ~\u5_timer2_reg[7]/P0001  & n3400 ;
  assign n4621 = n3396 & n4620 ;
  assign n4622 = ~n4619 & ~n4621 ;
  assign n4623 = n3390 & n4622 ;
  assign n4624 = n3634 & n4623 ;
  assign n4625 = ~n4618 & n4624 ;
  assign n4626 = ~n4610 & ~n4625 ;
  assign n4627 = \wb_addr_i[16]_pad  & ~n2739 ;
  assign n4628 = ~n2736 & n4627 ;
  assign n4629 = ~n2734 & n4628 ;
  assign n4630 = \wb_addr_i[15]_pad  & ~n2733 ;
  assign n4631 = ~n2730 & n4630 ;
  assign n4632 = n2740 & n4631 ;
  assign n4633 = \wb_addr_i[17]_pad  & ~n2733 ;
  assign n4634 = ~n2730 & n4633 ;
  assign n4635 = ~n2740 & n4634 ;
  assign n4636 = ~n4632 & ~n4635 ;
  assign n4637 = ~n4629 & n4636 ;
  assign n4638 = ~n3439 & ~n4637 ;
  assign n4639 = \u1_acs_addr_reg[13]/P0001  & \u1_acs_addr_reg[14]/P0001  ;
  assign n4640 = n3427 & n4639 ;
  assign n4641 = ~\u1_acs_addr_reg[15]/P0001  & ~n4640 ;
  assign n4642 = ~n3430 & n3439 ;
  assign n4643 = ~n4641 & n4642 ;
  assign n4644 = ~n4638 & ~n4643 ;
  assign n4645 = n1045 & ~n3889 ;
  assign n4646 = \u0_csc_reg[4]/NET0131  & ~n4645 ;
  assign n4647 = \u0_u1_csc_reg[4]/P0001  & n1045 ;
  assign n4648 = n4259 & n4647 ;
  assign n4649 = ~n3889 & n4648 ;
  assign n4650 = \u0_u0_csc_reg[4]/P0001  & n1045 ;
  assign n4651 = n4216 & n4650 ;
  assign n4652 = ~n3889 & n4651 ;
  assign n4653 = ~n4649 & ~n4652 ;
  assign n4654 = ~n4646 & n4653 ;
  assign n4655 = \u0_csc_reg[5]/NET0131  & ~n4645 ;
  assign n4656 = \u0_u1_csc_reg[5]/P0001  & n1045 ;
  assign n4657 = n4259 & n4656 ;
  assign n4658 = ~n3889 & n4657 ;
  assign n4659 = \u0_u0_csc_reg[5]/P0001  & n1045 ;
  assign n4660 = n4216 & n4659 ;
  assign n4661 = ~n3889 & n4660 ;
  assign n4662 = ~n4658 & ~n4661 ;
  assign n4663 = ~n4655 & n4662 ;
  assign n4664 = \u0_csc_reg[6]/NET0131  & ~n4645 ;
  assign n4665 = \u0_u0_csc_reg[6]/P0001  & n1045 ;
  assign n4666 = n4216 & n4665 ;
  assign n4667 = ~n3889 & n4666 ;
  assign n4668 = \u0_u1_csc_reg[6]/P0001  & n1045 ;
  assign n4669 = n4259 & n4668 ;
  assign n4670 = ~n3889 & n4669 ;
  assign n4671 = ~n4667 & ~n4670 ;
  assign n4672 = ~n4664 & n4671 ;
  assign n4673 = \u0_csc_reg[9]/NET0131  & ~n4645 ;
  assign n4674 = \u0_u0_csc_reg[9]/P0001  & n1045 ;
  assign n4675 = n4216 & n4674 ;
  assign n4676 = ~n3889 & n4675 ;
  assign n4677 = \u0_u1_csc_reg[9]/P0001  & n1045 ;
  assign n4678 = n4259 & n4677 ;
  assign n4679 = ~n3889 & n4678 ;
  assign n4680 = ~n4676 & ~n4679 ;
  assign n4681 = ~n4673 & n4680 ;
  assign n4682 = \u0_csc_reg[7]/NET0131  & ~n4645 ;
  assign n4683 = \u0_u0_csc_reg[7]/P0001  & n1045 ;
  assign n4684 = n4216 & n4683 ;
  assign n4685 = ~n3889 & n4684 ;
  assign n4686 = \u0_u1_csc_reg[7]/P0001  & n1045 ;
  assign n4687 = n4259 & n4686 ;
  assign n4688 = ~n3889 & n4687 ;
  assign n4689 = ~n4685 & ~n4688 ;
  assign n4690 = ~n4682 & n4689 ;
  assign n4691 = \u0_sp_csc_reg[10]/NET0131  & ~n4645 ;
  assign n4692 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[10]/P0001  ;
  assign n4693 = n1045 & n4692 ;
  assign n4694 = ~n3889 & n4693 ;
  assign n4695 = \u0_u1_csc_reg[10]/P0001  & n1045 ;
  assign n4696 = n3895 & n4695 ;
  assign n4697 = ~n3889 & n4696 ;
  assign n4698 = ~n4694 & ~n4697 ;
  assign n4699 = ~n4691 & n4698 ;
  assign n4700 = \u0_sp_csc_reg[4]/NET0131  & ~n4645 ;
  assign n4701 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[4]/P0001  ;
  assign n4702 = n1045 & n4701 ;
  assign n4703 = ~n3889 & n4702 ;
  assign n4704 = n3895 & n4647 ;
  assign n4705 = ~n3889 & n4704 ;
  assign n4706 = ~n4703 & ~n4705 ;
  assign n4707 = ~n4700 & n4706 ;
  assign n4708 = \u0_sp_csc_reg[5]/NET0131  & ~n4645 ;
  assign n4709 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[5]/P0001  ;
  assign n4710 = n1045 & n4709 ;
  assign n4711 = ~n3889 & n4710 ;
  assign n4712 = n3895 & n4656 ;
  assign n4713 = ~n3889 & n4712 ;
  assign n4714 = ~n4711 & ~n4713 ;
  assign n4715 = ~n4708 & n4714 ;
  assign n4716 = \u0_sp_csc_reg[6]/NET0131  & ~n4645 ;
  assign n4717 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[6]/P0001  ;
  assign n4718 = n1045 & n4717 ;
  assign n4719 = ~n3889 & n4718 ;
  assign n4720 = n3895 & n4668 ;
  assign n4721 = ~n3889 & n4720 ;
  assign n4722 = ~n4719 & ~n4721 ;
  assign n4723 = ~n4716 & n4722 ;
  assign n4724 = \u0_sp_csc_reg[7]/NET0131  & ~n4645 ;
  assign n4725 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[7]/P0001  ;
  assign n4726 = n1045 & n4725 ;
  assign n4727 = ~n3889 & n4726 ;
  assign n4728 = n3895 & n4686 ;
  assign n4729 = ~n3889 & n4728 ;
  assign n4730 = ~n4727 & ~n4729 ;
  assign n4731 = ~n4724 & n4730 ;
  assign n4732 = \u0_sp_csc_reg[9]/NET0131  & ~n4645 ;
  assign n4733 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[9]/P0001  ;
  assign n4734 = n1045 & n4733 ;
  assign n4735 = ~n3889 & n4734 ;
  assign n4736 = n3895 & n4677 ;
  assign n4737 = ~n3889 & n4736 ;
  assign n4738 = ~n4735 & ~n4737 ;
  assign n4739 = ~n4732 & n4738 ;
  assign n4740 = \u0_csc_reg[10]/NET0131  & ~n4645 ;
  assign n4741 = n4259 & n4695 ;
  assign n4742 = ~n3889 & n4741 ;
  assign n4743 = \u0_u0_csc_reg[10]/P0001  & n1045 ;
  assign n4744 = n4216 & n4743 ;
  assign n4745 = ~n3889 & n4744 ;
  assign n4746 = ~n4742 & ~n4745 ;
  assign n4747 = ~n4740 & n4746 ;
  assign n4748 = \u5_ap_en_reg/NET0131  & ~\u5_state_reg[1]/NET0131  ;
  assign n4749 = n1210 & n1222 ;
  assign n4750 = n2778 & n4749 ;
  assign n4751 = ~n4748 & ~n4750 ;
  assign n4752 = \u0_sp_csc_reg[2]/NET0131  & ~n4645 ;
  assign n4753 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[2]/NET0131  ;
  assign n4754 = n1045 & n4753 ;
  assign n4755 = ~n3889 & n4754 ;
  assign n4756 = \u0_u1_csc_reg[2]/NET0131  & n3895 ;
  assign n4757 = n1045 & n4756 ;
  assign n4758 = ~n3889 & n4757 ;
  assign n4759 = ~n4755 & ~n4758 ;
  assign n4760 = ~n4752 & n4759 ;
  assign n4761 = \u0_sp_csc_reg[1]/NET0131  & ~n4645 ;
  assign n4762 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[1]/NET0131  ;
  assign n4763 = n1045 & n4762 ;
  assign n4764 = ~n3889 & n4763 ;
  assign n4765 = \u0_u1_csc_reg[1]/NET0131  & n3895 ;
  assign n4766 = n1045 & n4765 ;
  assign n4767 = ~n3889 & n4766 ;
  assign n4768 = ~n4764 & ~n4767 ;
  assign n4769 = ~n4761 & n4768 ;
  assign n4770 = \u0_sp_csc_reg[3]/NET0131  & ~n4645 ;
  assign n4771 = \u0_spec_req_cs_reg[0]/NET0131  & \u0_u0_csc_reg[3]/NET0131  ;
  assign n4772 = n1045 & n4771 ;
  assign n4773 = ~n3889 & n4772 ;
  assign n4774 = \u0_u1_csc_reg[3]/NET0131  & n3895 ;
  assign n4775 = n1045 & n4774 ;
  assign n4776 = ~n3889 & n4775 ;
  assign n4777 = ~n4773 & ~n4776 ;
  assign n4778 = ~n4770 & n4777 ;
  assign n4779 = ~n1290 & ~n2042 ;
  assign n4780 = ~n2039 & n4779 ;
  assign n4781 = ~n2029 & n4780 ;
  assign n4782 = ~n2052 & ~n3620 ;
  assign n4783 = n4781 & n4782 ;
  assign n4784 = ~n1153 & n2617 ;
  assign n4785 = ~n2051 & n4784 ;
  assign n4786 = n2634 & n4785 ;
  assign n4787 = \u5_timer_reg[4]/NET0131  & ~n2615 ;
  assign n4788 = ~\u5_timer_reg[4]/NET0131  & n2063 ;
  assign n4789 = n2072 & n4788 ;
  assign n4790 = ~n4787 & ~n4789 ;
  assign n4791 = n4781 & ~n4790 ;
  assign n4792 = n4786 & n4791 ;
  assign n4793 = ~n4783 & ~n4792 ;
  assign n4794 = n1851 & n3033 ;
  assign n4795 = ~n1848 & n4794 ;
  assign n4796 = ~n2052 & ~n4795 ;
  assign n4797 = n4781 & n4796 ;
  assign n4798 = \u5_timer_reg[5]/NET0131  & ~n4789 ;
  assign n4799 = n2065 & n2072 ;
  assign n4800 = ~n4798 & ~n4799 ;
  assign n4801 = n4781 & ~n4800 ;
  assign n4802 = n4786 & n4801 ;
  assign n4803 = ~n4797 & ~n4802 ;
  assign n4804 = n1851 & n4597 ;
  assign n4805 = ~n1848 & n4804 ;
  assign n4806 = ~n2052 & ~n4805 ;
  assign n4807 = n4781 & n4806 ;
  assign n4808 = \u5_timer_reg[6]/NET0131  & ~n4799 ;
  assign n4809 = ~\u5_mc_le_reg/NET0131  & ~\u5_timer_reg[6]/NET0131  ;
  assign n4810 = n2066 & n4809 ;
  assign n4811 = n2065 & n4810 ;
  assign n4812 = ~n2069 & n4811 ;
  assign n4813 = ~n4808 & ~n4812 ;
  assign n4814 = n4781 & ~n4813 ;
  assign n4815 = n4786 & n4814 ;
  assign n4816 = ~n4807 & ~n4815 ;
  assign n4817 = n1851 & n4615 ;
  assign n4818 = ~n1848 & n4817 ;
  assign n4819 = ~n2052 & ~n4818 ;
  assign n4820 = n4781 & n4819 ;
  assign n4821 = \u5_timer_reg[7]/NET0131  & ~n4811 ;
  assign n4822 = n4781 & n4821 ;
  assign n4823 = n4786 & n4822 ;
  assign n4824 = ~n4820 & ~n4823 ;
  assign n4825 = \u0_csc_reg[11]/NET0131  & ~n4645 ;
  assign n4826 = \u0_u1_csc_reg[11]/P0001  & n4259 ;
  assign n4827 = \u0_u0_csc_reg[11]/P0001  & ~n4200 ;
  assign n4828 = n4214 & n4827 ;
  assign n4829 = n4199 & n4828 ;
  assign n4830 = ~n4826 & ~n4829 ;
  assign n4831 = n1045 & ~n4830 ;
  assign n4832 = ~n3889 & n4831 ;
  assign n4833 = ~n4825 & ~n4832 ;
  assign n4834 = \wb_addr_i[15]_pad  & ~n2739 ;
  assign n4835 = ~n2736 & n4834 ;
  assign n4836 = ~n2734 & n4835 ;
  assign n4837 = \wb_addr_i[14]_pad  & ~n2733 ;
  assign n4838 = ~n2730 & n4837 ;
  assign n4839 = n2740 & n4838 ;
  assign n4840 = ~n2740 & n3781 ;
  assign n4841 = ~n4839 & ~n4840 ;
  assign n4842 = ~n4836 & n4841 ;
  assign n4843 = ~n3439 & ~n4842 ;
  assign n4844 = \u1_acs_addr_reg[13]/P0001  & n3427 ;
  assign n4845 = ~\u1_acs_addr_reg[14]/P0001  & ~n4844 ;
  assign n4846 = n3439 & ~n4640 ;
  assign n4847 = ~n4845 & n4846 ;
  assign n4848 = ~n4843 & ~n4847 ;
  assign n4849 = n1906 & n1930 ;
  assign n4850 = ~n1167 & n1348 ;
  assign n4851 = ~n4849 & n4850 ;
  assign n4852 = ~n1143 & ~n1400 ;
  assign n4853 = ~n1897 & ~n4852 ;
  assign n4854 = ~n1400 & n1904 ;
  assign n4855 = n1314 & ~n4854 ;
  assign n4856 = ~n4853 & ~n4855 ;
  assign n4857 = n4851 & n4856 ;
  assign n4858 = \u5_cmd_del_reg[2]/NET0131  & \u5_wr_cycle_reg/NET0131  ;
  assign n4859 = ~n1104 & n3551 ;
  assign n4860 = n1128 & n1499 ;
  assign n4861 = \u5_wb_wait_r_reg/P0001  & n1273 ;
  assign n4862 = ~n1987 & ~n4861 ;
  assign n4863 = n1474 & n4862 ;
  assign n4864 = n4860 & n4863 ;
  assign n4865 = n3539 & n4864 ;
  assign n4866 = n4859 & n4865 ;
  assign n4867 = ~\u5_wr_cycle_reg/NET0131  & ~n4866 ;
  assign n4868 = ~n4858 & ~n4867 ;
  assign n4869 = \wb_addr_i[22]_pad  & ~n2739 ;
  assign n4870 = ~n2736 & n4869 ;
  assign n4871 = ~n2734 & n4870 ;
  assign n4872 = n2740 & n3563 ;
  assign n4873 = ~n2740 & n3453 ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = ~n4871 & n4874 ;
  assign n4876 = ~n3439 & ~n4875 ;
  assign n4877 = \u1_acs_addr_reg[19]/P0001  & \u1_acs_addr_reg[20]/P0001  ;
  assign n4878 = n3433 & n4877 ;
  assign n4879 = ~\u1_acs_addr_reg[21]/P0001  & ~n4878 ;
  assign n4880 = ~n3436 & n3439 ;
  assign n4881 = ~n4879 & n4880 ;
  assign n4882 = ~n4876 & ~n4881 ;
  assign n4883 = ~\u4_rfr_clr_reg/P0001  & ~\u4_rfr_req_reg/NET0131  ;
  assign n4884 = ~\u5_rfr_ack_r_reg/NET0131  & ~n4883 ;
  assign n4885 = \wb_addr_i[14]_pad  & ~n2739 ;
  assign n4886 = ~n2736 & n4885 ;
  assign n4887 = ~n2734 & n4886 ;
  assign n4888 = \wb_addr_i[13]_pad  & ~n2733 ;
  assign n4889 = ~n2730 & n4888 ;
  assign n4890 = n2740 & n4889 ;
  assign n4891 = ~n2740 & n4631 ;
  assign n4892 = ~n4890 & ~n4891 ;
  assign n4893 = ~n4887 & n4892 ;
  assign n4894 = ~n3439 & ~n4893 ;
  assign n4895 = \u1_acs_addr_reg[13]/P0001  & n3439 ;
  assign n4896 = ~n3427 & n4895 ;
  assign n4897 = ~\u1_acs_addr_reg[13]/P0001  & n3439 ;
  assign n4898 = n3427 & n4897 ;
  assign n4899 = ~n4896 & ~n4898 ;
  assign n4900 = ~n4894 & n4899 ;
  assign n4901 = ~\u1_u0_out_r_reg[11]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n4902 = ~n3424 & n4901 ;
  assign n4903 = ~\u1_acs_addr_reg[11]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n4904 = ~\u1_acs_addr_reg[11]/P0001  & n963 ;
  assign n4905 = ~n3423 & n4904 ;
  assign n4906 = ~n4903 & ~n4905 ;
  assign n4907 = n3439 & n4906 ;
  assign n4908 = ~n4902 & n4907 ;
  assign n4909 = ~n2740 & n4889 ;
  assign n4910 = \wb_addr_i[11]_pad  & ~n2733 ;
  assign n4911 = ~n2730 & n4910 ;
  assign n4912 = n2740 & n4911 ;
  assign n4913 = \wb_addr_i[12]_pad  & ~n2739 ;
  assign n4914 = ~n2736 & n4913 ;
  assign n4915 = ~n2734 & n4914 ;
  assign n4916 = ~n4912 & ~n4915 ;
  assign n4917 = ~n4909 & n4916 ;
  assign n4918 = ~n3439 & ~n4917 ;
  assign n4919 = ~n4908 & ~n4918 ;
  assign n4920 = \wb_addr_i[18]_pad  & ~n2739 ;
  assign n4921 = ~n2736 & n4920 ;
  assign n4922 = ~n2734 & n4921 ;
  assign n4923 = n2740 & n4634 ;
  assign n4924 = ~n2740 & n3569 ;
  assign n4925 = ~n4923 & ~n4924 ;
  assign n4926 = ~n4922 & n4925 ;
  assign n4927 = ~n3439 & ~n4926 ;
  assign n4928 = \u1_acs_addr_reg[16]/P0001  & n3430 ;
  assign n4929 = ~\u1_acs_addr_reg[17]/P0001  & ~n4928 ;
  assign n4930 = n3439 & ~n3818 ;
  assign n4931 = ~n4929 & n4930 ;
  assign n4932 = ~n4927 & ~n4931 ;
  assign n4933 = n3535 & n3539 ;
  assign n4934 = n1490 & n3547 ;
  assign n4935 = n1927 & n2811 ;
  assign n4936 = ~n1922 & n4935 ;
  assign n4937 = n1310 & ~n4936 ;
  assign n4938 = n4934 & ~n4937 ;
  assign n4939 = n1333 & n3552 ;
  assign n4940 = ~n1104 & n1988 ;
  assign n4941 = \u7_mc_br_r_reg/P0001  & n1411 ;
  assign n4942 = n3536 & ~n4941 ;
  assign n4943 = n4940 & n4942 ;
  assign n4944 = n4939 & n4943 ;
  assign n4945 = n3544 & n4944 ;
  assign n4946 = n4938 & n4945 ;
  assign n4947 = n4933 & n4946 ;
  assign n4948 = \wb_addr_i[7]_pad  & ~n2733 ;
  assign n4949 = ~n2730 & n4948 ;
  assign n4950 = n2740 & n4949 ;
  assign n4951 = \wb_addr_i[8]_pad  & ~n2739 ;
  assign n4952 = ~n2736 & n4951 ;
  assign n4953 = ~n2734 & n4952 ;
  assign n4954 = \wb_addr_i[9]_pad  & ~n2733 ;
  assign n4955 = ~n2730 & n4954 ;
  assign n4956 = ~n2740 & n4955 ;
  assign n4957 = ~n4953 & ~n4956 ;
  assign n4958 = ~n4950 & n4957 ;
  assign n4959 = ~n3439 & ~n4958 ;
  assign n4960 = ~\u1_u0_out_r_reg[7]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n4961 = ~n3424 & n4960 ;
  assign n4962 = ~\u1_acs_addr_reg[7]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n4963 = ~\u1_acs_addr_reg[7]/P0001  & n963 ;
  assign n4964 = ~n3423 & n4963 ;
  assign n4965 = ~n4962 & ~n4964 ;
  assign n4966 = n3439 & n4965 ;
  assign n4967 = ~n4961 & n4966 ;
  assign n4968 = ~n4959 & ~n4967 ;
  assign n4969 = ~\u5_state_reg[1]/NET0131  & \u5_wr_cycle_reg/NET0131  ;
  assign n4970 = ~n1895 & ~n2165 ;
  assign n4971 = ~n1194 & ~n4970 ;
  assign n4972 = n3172 & ~n4970 ;
  assign n4973 = n1930 & n4972 ;
  assign n4974 = ~n4971 & ~n4973 ;
  assign n4975 = ~n4969 & n4974 ;
  assign n4976 = \u0_csr_r_reg[8]/NET0131  & ~\u4_rfr_cnt_reg[1]/NET0131  ;
  assign n4977 = ~\u0_csr_r_reg[10]/NET0131  & ~\u0_csr_r_reg[9]/NET0131  ;
  assign n4978 = ~n4976 & n4977 ;
  assign n4979 = \u0_csr_r_reg[8]/NET0131  & ~\u4_rfr_cnt_reg[3]/NET0131  ;
  assign n4980 = ~\u0_csr_r_reg[10]/NET0131  & ~n4979 ;
  assign n4981 = \u4_rfr_cnt_reg[1]/NET0131  & \u4_rfr_cnt_reg[2]/NET0131  ;
  assign n4982 = n4980 & n4981 ;
  assign n4983 = \u0_csr_r_reg[8]/NET0131  & ~\u4_rfr_cnt_reg[5]/NET0131  ;
  assign n4984 = ~\u0_csr_r_reg[9]/NET0131  & ~n4983 ;
  assign n4985 = \u0_csr_r_reg[8]/NET0131  & ~\u4_rfr_cnt_reg[7]/NET0131  ;
  assign n4986 = \u4_rfr_cnt_reg[5]/NET0131  & \u4_rfr_cnt_reg[6]/NET0131  ;
  assign n4987 = ~n4985 & n4986 ;
  assign n4988 = ~n4984 & ~n4987 ;
  assign n4989 = \u4_rfr_cnt_reg[3]/NET0131  & \u4_rfr_cnt_reg[4]/NET0131  ;
  assign n4990 = n4981 & n4989 ;
  assign n4991 = ~n4988 & n4990 ;
  assign n4992 = ~n4982 & ~n4991 ;
  assign n4993 = ~n4978 & n4992 ;
  assign n4994 = \u4_rfr_cnt_reg[0]/NET0131  & \u4_rfr_early_reg/NET0131  ;
  assign n4995 = ~n4993 & n4994 ;
  assign n4996 = \wb_addr_i[13]_pad  & ~n2739 ;
  assign n4997 = ~n2736 & n4996 ;
  assign n4998 = ~n2734 & n4997 ;
  assign n4999 = \wb_addr_i[12]_pad  & ~n2733 ;
  assign n5000 = ~n2730 & n4999 ;
  assign n5001 = n2740 & n5000 ;
  assign n5002 = ~n2740 & n4838 ;
  assign n5003 = ~n5001 & ~n5002 ;
  assign n5004 = ~n4998 & n5003 ;
  assign n5005 = ~n3439 & ~n5004 ;
  assign n5006 = \u1_u0_out_r_reg[12]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5007 = ~n3424 & n5006 ;
  assign n5008 = ~\u1_acs_addr_reg[12]/P0001  & ~n5007 ;
  assign n5009 = ~n3427 & n3439 ;
  assign n5010 = ~n5008 & n5009 ;
  assign n5011 = ~n5005 & ~n5010 ;
  assign n5012 = ~\u5_ack_cnt_reg[0]/NET0131  & ~\u5_no_wb_cycle_reg/NET0131  ;
  assign n5013 = ~n2173 & n5012 ;
  assign n5014 = ~n1043 & n5013 ;
  assign n5015 = \u5_ack_cnt_reg[0]/NET0131  & ~\u5_no_wb_cycle_reg/NET0131  ;
  assign n5016 = n2173 & n5015 ;
  assign n5017 = ~n1043 & n5016 ;
  assign n5018 = ~n5014 & ~n5017 ;
  assign n5019 = ~n2173 & n5015 ;
  assign n5020 = n1043 & n5019 ;
  assign n5021 = n2173 & n5012 ;
  assign n5022 = n1043 & n5021 ;
  assign n5023 = ~n5020 & ~n5022 ;
  assign n5024 = n5018 & n5023 ;
  assign n5025 = n1043 & n2173 ;
  assign n5026 = ~\u5_ack_cnt_reg[0]/NET0131  & ~n5025 ;
  assign n5027 = ~n1043 & ~n2173 ;
  assign n5028 = \u5_ack_cnt_reg[0]/NET0131  & \u5_ack_cnt_reg[1]/NET0131  ;
  assign n5029 = ~n2166 & ~n5028 ;
  assign n5030 = ~n5027 & n5029 ;
  assign n5031 = ~n5026 & n5030 ;
  assign n5032 = n5027 & ~n5029 ;
  assign n5033 = ~\u5_ack_cnt_reg[0]/NET0131  & ~n5029 ;
  assign n5034 = ~n5025 & n5033 ;
  assign n5035 = ~n5032 & ~n5034 ;
  assign n5036 = ~\u5_no_wb_cycle_reg/NET0131  & n5035 ;
  assign n5037 = ~n5031 & n5036 ;
  assign n5038 = n2166 & n2173 ;
  assign n5039 = n1043 & n5038 ;
  assign n5040 = \u5_ack_cnt_reg[2]/NET0131  & ~n5039 ;
  assign n5041 = ~\u5_ack_cnt_reg[2]/NET0131  & n2166 ;
  assign n5042 = n2173 & n5041 ;
  assign n5043 = n1043 & n5042 ;
  assign n5044 = ~n5027 & ~n5043 ;
  assign n5045 = ~n5040 & n5044 ;
  assign n5046 = ~\u5_ack_cnt_reg[2]/NET0131  & ~n5028 ;
  assign n5047 = \u5_ack_cnt_reg[2]/NET0131  & n5028 ;
  assign n5048 = ~n5046 & ~n5047 ;
  assign n5049 = ~n2173 & ~n5048 ;
  assign n5050 = ~n1043 & n5049 ;
  assign n5051 = ~\u5_no_wb_cycle_reg/NET0131  & ~n5050 ;
  assign n5052 = ~n5045 & n5051 ;
  assign n5053 = \u5_ack_cnt_reg[3]/NET0131  & ~n5043 ;
  assign n5054 = n2168 & n2173 ;
  assign n5055 = n1043 & n5054 ;
  assign n5056 = ~n5027 & ~n5055 ;
  assign n5057 = ~n5053 & n5056 ;
  assign n5058 = \u5_ack_cnt_reg[3]/NET0131  & ~n5047 ;
  assign n5059 = \u5_ack_cnt_reg[2]/NET0131  & ~\u5_ack_cnt_reg[3]/NET0131  ;
  assign n5060 = n5028 & n5059 ;
  assign n5061 = ~n5058 & ~n5060 ;
  assign n5062 = ~n2173 & n5061 ;
  assign n5063 = ~n1043 & n5062 ;
  assign n5064 = ~\u5_no_wb_cycle_reg/NET0131  & ~n5063 ;
  assign n5065 = ~n5057 & n5064 ;
  assign n5066 = \wb_addr_i[4]_pad  & ~n2733 ;
  assign n5067 = ~n2730 & n5066 ;
  assign n5068 = n2740 & n5067 ;
  assign n5069 = \wb_addr_i[5]_pad  & ~n2739 ;
  assign n5070 = ~n2736 & n5069 ;
  assign n5071 = ~n2734 & n5070 ;
  assign n5072 = \wb_addr_i[6]_pad  & ~n2733 ;
  assign n5073 = ~n2730 & n5072 ;
  assign n5074 = ~n2740 & n5073 ;
  assign n5075 = ~n5071 & ~n5074 ;
  assign n5076 = ~n5068 & n5075 ;
  assign n5077 = ~n3439 & ~n5076 ;
  assign n5078 = ~\u1_u0_out_r_reg[4]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5079 = ~n3424 & n5078 ;
  assign n5080 = ~\u1_acs_addr_reg[4]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5081 = ~\u1_acs_addr_reg[4]/P0001  & n963 ;
  assign n5082 = ~n3423 & n5081 ;
  assign n5083 = ~n5080 & ~n5082 ;
  assign n5084 = n3439 & n5083 ;
  assign n5085 = ~n5079 & n5084 ;
  assign n5086 = ~n5077 & ~n5085 ;
  assign n5087 = ~\u1_u0_out_r_reg[8]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5088 = ~n3424 & n5087 ;
  assign n5089 = ~\u1_acs_addr_reg[8]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5090 = ~\u1_acs_addr_reg[8]/P0001  & n963 ;
  assign n5091 = ~n3423 & n5090 ;
  assign n5092 = ~n5089 & ~n5091 ;
  assign n5093 = n3439 & n5092 ;
  assign n5094 = ~n5088 & n5093 ;
  assign n5095 = \wb_addr_i[8]_pad  & ~n2733 ;
  assign n5096 = ~n2730 & n5095 ;
  assign n5097 = n2740 & n5096 ;
  assign n5098 = \wb_addr_i[9]_pad  & ~n2739 ;
  assign n5099 = ~n2736 & n5098 ;
  assign n5100 = ~n2734 & n5099 ;
  assign n5101 = \wb_addr_i[10]_pad  & ~n2733 ;
  assign n5102 = ~n2730 & n5101 ;
  assign n5103 = ~n2740 & n5102 ;
  assign n5104 = ~n5100 & ~n5103 ;
  assign n5105 = ~n5097 & n5104 ;
  assign n5106 = ~n3439 & ~n5105 ;
  assign n5107 = ~n5094 & ~n5106 ;
  assign n5108 = ~n3654 & ~n3811 ;
  assign n5109 = n2729 & ~n5108 ;
  assign n5110 = ~n2723 & ~n2728 ;
  assign n5111 = n4924 & ~n5110 ;
  assign n5112 = ~n5109 & ~n5111 ;
  assign n5113 = n2723 & ~n2728 ;
  assign n5114 = ~n2723 & n2728 ;
  assign n5115 = ~n5113 & ~n5114 ;
  assign n5116 = ~n3567 & ~n4872 ;
  assign n5117 = ~n5115 & ~n5116 ;
  assign n5118 = \u0_sp_csc_reg[9]/NET0131  & ~n1200 ;
  assign n5119 = \u0_csc_reg[9]/NET0131  & ~\u5_state_reg[26]/NET0131  ;
  assign n5120 = ~\u5_lmr_ack_reg/NET0131  & n5119 ;
  assign n5121 = n983 & n5120 ;
  assign n5122 = ~n5118 & ~n5121 ;
  assign n5123 = ~n5117 & ~n5122 ;
  assign n5124 = n5112 & n5123 ;
  assign n5125 = \wb_addr_i[22]_pad  & ~n2722 ;
  assign n5126 = ~n2719 & n5125 ;
  assign n5127 = n2728 & n5126 ;
  assign n5128 = n2770 & n5127 ;
  assign n5129 = \wb_addr_i[23]_pad  & n2770 ;
  assign n5130 = ~n5115 & n5129 ;
  assign n5131 = ~n5128 & ~n5130 ;
  assign n5132 = n2729 & n3651 ;
  assign n5133 = ~n3564 & ~n4871 ;
  assign n5134 = ~n5115 & ~n5133 ;
  assign n5135 = ~n5132 & ~n5134 ;
  assign n5136 = n5131 & n5135 ;
  assign n5137 = n2729 & n3564 ;
  assign n5138 = n5122 & ~n5137 ;
  assign n5139 = n5136 & n5138 ;
  assign n5140 = ~n5124 & ~n5139 ;
  assign n5141 = \u1_acs_addr_reg[0]/P0001  & \u1_acs_addr_reg[1]/P0001  ;
  assign n5142 = \u1_acs_addr_reg[2]/P0001  & \u1_acs_addr_reg[3]/P0001  ;
  assign n5143 = n5141 & n5142 ;
  assign n5144 = \u1_acs_addr_reg[4]/P0001  & \u1_acs_addr_reg[6]/P0001  ;
  assign n5145 = \u1_acs_addr_reg[5]/P0001  & n5144 ;
  assign n5146 = n5143 & n5145 ;
  assign n5147 = \u1_acs_addr_reg[7]/P0001  & \u1_acs_addr_reg[9]/P0001  ;
  assign n5148 = \u1_acs_addr_reg[8]/P0001  & n5147 ;
  assign n5149 = n5146 & n5148 ;
  assign n5150 = \u1_acs_addr_reg[10]/P0001  & \u1_acs_addr_reg[11]/P0001  ;
  assign n5151 = n5149 & n5150 ;
  assign n5152 = \u1_acs_addr_reg[10]/P0001  & n5149 ;
  assign n5153 = ~\u1_acs_addr_reg[11]/P0001  & ~n5152 ;
  assign n5154 = ~n5151 & ~n5153 ;
  assign n5155 = \wb_addr_i[10]_pad  & ~n2739 ;
  assign n5156 = ~n2736 & n5155 ;
  assign n5157 = ~n2734 & n5156 ;
  assign n5158 = ~n4912 & ~n5157 ;
  assign n5159 = n2729 & ~n5158 ;
  assign n5160 = n5103 & ~n5110 ;
  assign n5161 = \wb_addr_i[11]_pad  & ~n2739 ;
  assign n5162 = ~n2736 & n5161 ;
  assign n5163 = ~n2734 & n5162 ;
  assign n5164 = ~n5001 & ~n5163 ;
  assign n5165 = ~n5115 & ~n5164 ;
  assign n5166 = ~n5160 & ~n5165 ;
  assign n5167 = ~n5159 & n5166 ;
  assign n5168 = n5122 & ~n5167 ;
  assign n5169 = n2740 & n3446 ;
  assign n5170 = ~n3451 & ~n4873 ;
  assign n5171 = ~n5169 & n5170 ;
  assign n5172 = n5114 & ~n5171 ;
  assign n5173 = ~n3454 & ~n4871 ;
  assign n5174 = n2729 & ~n5173 ;
  assign n5175 = n2740 & n3587 ;
  assign n5176 = ~n3582 & ~n5175 ;
  assign n5177 = n5113 & ~n5176 ;
  assign n5178 = ~n5174 & ~n5177 ;
  assign n5179 = n3647 & n5113 ;
  assign n5180 = ~n5137 & ~n5179 ;
  assign n5181 = n5178 & n5180 ;
  assign n5182 = ~n5172 & n5181 ;
  assign n5183 = ~n5122 & ~n5182 ;
  assign n5184 = ~n5168 & ~n5183 ;
  assign n5185 = ~n4890 & ~n4915 ;
  assign n5186 = ~n5115 & ~n5185 ;
  assign n5187 = n2729 & ~n5164 ;
  assign n5188 = ~n2740 & n4911 ;
  assign n5189 = ~n5110 & n5188 ;
  assign n5190 = ~n5187 & ~n5189 ;
  assign n5191 = ~n5186 & n5190 ;
  assign n5192 = n5122 & ~n5191 ;
  assign n5193 = n2729 & n3582 ;
  assign n5194 = n5113 & ~n5171 ;
  assign n5195 = ~n5193 & ~n5194 ;
  assign n5196 = ~n3647 & ~n5175 ;
  assign n5197 = n2729 & ~n5196 ;
  assign n5198 = \wb_addr_i[25]_pad  & ~n2739 ;
  assign n5199 = ~n2736 & n5198 ;
  assign n5200 = ~n2734 & n5199 ;
  assign n5201 = \wb_addr_i[26]_pad  & ~n2733 ;
  assign n5202 = ~n2730 & n5201 ;
  assign n5203 = n2740 & n5202 ;
  assign n5204 = ~n3588 & ~n5203 ;
  assign n5205 = ~n5200 & n5204 ;
  assign n5206 = n5114 & ~n5205 ;
  assign n5207 = ~n5197 & ~n5206 ;
  assign n5208 = n5195 & n5207 ;
  assign n5209 = ~n5122 & ~n5208 ;
  assign n5210 = ~n5192 & ~n5209 ;
  assign n5211 = ~n4839 & ~n4998 ;
  assign n5212 = ~n5115 & ~n5211 ;
  assign n5213 = n2729 & ~n5185 ;
  assign n5214 = ~n2740 & n5000 ;
  assign n5215 = ~n5110 & n5214 ;
  assign n5216 = ~n5213 & ~n5215 ;
  assign n5217 = ~n5212 & n5216 ;
  assign n5218 = n5122 & ~n5217 ;
  assign n5219 = ~n5122 & ~n5167 ;
  assign n5220 = ~n5218 & ~n5219 ;
  assign n5221 = ~n3585 & ~n3651 ;
  assign n5222 = ~n5115 & ~n5221 ;
  assign n5223 = n3813 & ~n5110 ;
  assign n5224 = n2729 & ~n5116 ;
  assign n5225 = ~n5223 & ~n5224 ;
  assign n5226 = ~n5222 & n5225 ;
  assign n5227 = ~n5122 & ~n5226 ;
  assign n5228 = ~n3647 & n5176 ;
  assign n5229 = n5114 & ~n5228 ;
  assign n5230 = n2723 & n3647 ;
  assign n5231 = n5178 & ~n5230 ;
  assign n5232 = ~n5229 & n5231 ;
  assign n5233 = n5122 & ~n5232 ;
  assign n5234 = ~n5227 & ~n5233 ;
  assign n5235 = ~n4632 & ~n4887 ;
  assign n5236 = ~n5115 & ~n5235 ;
  assign n5237 = n2729 & ~n5211 ;
  assign n5238 = n4909 & ~n5110 ;
  assign n5239 = ~n5237 & ~n5238 ;
  assign n5240 = ~n5236 & n5239 ;
  assign n5241 = n5122 & ~n5240 ;
  assign n5242 = ~n5122 & ~n5191 ;
  assign n5243 = ~n5241 & ~n5242 ;
  assign n5244 = ~n3782 & ~n4836 ;
  assign n5245 = ~n5115 & ~n5244 ;
  assign n5246 = n2729 & ~n5235 ;
  assign n5247 = n5002 & ~n5110 ;
  assign n5248 = ~n5246 & ~n5247 ;
  assign n5249 = ~n5245 & n5248 ;
  assign n5250 = n5122 & ~n5249 ;
  assign n5251 = ~n5122 & ~n5217 ;
  assign n5252 = ~n5250 & ~n5251 ;
  assign n5253 = ~n4629 & ~n4923 ;
  assign n5254 = ~n5115 & ~n5253 ;
  assign n5255 = n2729 & ~n5244 ;
  assign n5256 = n4891 & ~n5110 ;
  assign n5257 = ~n5255 & ~n5256 ;
  assign n5258 = ~n5254 & n5257 ;
  assign n5259 = n5122 & ~n5258 ;
  assign n5260 = ~n5122 & ~n5240 ;
  assign n5261 = ~n5259 & ~n5260 ;
  assign n5262 = ~n3789 & ~n3812 ;
  assign n5263 = ~n5115 & ~n5262 ;
  assign n5264 = n2729 & ~n5253 ;
  assign n5265 = n4840 & ~n5110 ;
  assign n5266 = ~n5264 & ~n5265 ;
  assign n5267 = ~n5263 & n5266 ;
  assign n5268 = n5122 & ~n5267 ;
  assign n5269 = ~n5122 & ~n5249 ;
  assign n5270 = ~n5268 & ~n5269 ;
  assign n5271 = ~n3570 & ~n4922 ;
  assign n5272 = ~n5115 & ~n5271 ;
  assign n5273 = n2729 & ~n5262 ;
  assign n5274 = n4635 & ~n5110 ;
  assign n5275 = ~n5273 & ~n5274 ;
  assign n5276 = ~n5272 & n5275 ;
  assign n5277 = n5122 & ~n5276 ;
  assign n5278 = ~n5122 & ~n5258 ;
  assign n5279 = ~n5277 & ~n5278 ;
  assign n5280 = ~n5108 & ~n5115 ;
  assign n5281 = n2729 & ~n5271 ;
  assign n5282 = n3786 & ~n5110 ;
  assign n5283 = ~n5281 & ~n5282 ;
  assign n5284 = ~n5280 & n5283 ;
  assign n5285 = n5122 & ~n5284 ;
  assign n5286 = ~n5122 & ~n5267 ;
  assign n5287 = ~n5285 & ~n5286 ;
  assign n5288 = ~n5122 & ~n5272 ;
  assign n5289 = n5275 & n5288 ;
  assign n5290 = ~n5117 & n5122 ;
  assign n5291 = n5112 & n5290 ;
  assign n5292 = ~n5289 & ~n5291 ;
  assign n5293 = ~n5122 & ~n5284 ;
  assign n5294 = n5122 & ~n5226 ;
  assign n5295 = ~n5293 & ~n5294 ;
  assign n5296 = n1849 & ~n1949 ;
  assign n5297 = ~n1848 & n5296 ;
  assign n5298 = ~n5122 & ~n5136 ;
  assign n5299 = n2729 & n5175 ;
  assign n5300 = ~n5172 & ~n5299 ;
  assign n5301 = n5195 & n5300 ;
  assign n5302 = n5122 & ~n5301 ;
  assign n5303 = ~n5298 & ~n5302 ;
  assign n5304 = ~\u0_csc_reg[4]/NET0131  & ~\u0_csc_reg[5]/NET0131  ;
  assign n5305 = \u5_pack_le1_reg/P0001  & n5304 ;
  assign n5306 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[0]/P0001  ;
  assign n5307 = n5304 & n5306 ;
  assign n5308 = n5305 & ~n5307 ;
  assign n5309 = \u0_csc_reg[4]/NET0131  & ~\u0_csc_reg[5]/NET0131  ;
  assign n5310 = \u5_pack_le0_reg/P0001  & n5309 ;
  assign n5311 = \u3_byte1_reg[0]/P0001  & ~n5310 ;
  assign n5312 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[8]/P0001  ;
  assign n5313 = n5309 & n5312 ;
  assign n5314 = ~n5307 & ~n5313 ;
  assign n5315 = ~n5311 & n5314 ;
  assign n5316 = ~n5308 & ~n5315 ;
  assign n5317 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[2]/P0001  ;
  assign n5318 = n5304 & n5317 ;
  assign n5319 = n5305 & ~n5318 ;
  assign n5320 = \u3_byte1_reg[2]/P0001  & ~n5310 ;
  assign n5321 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[10]/P0001  ;
  assign n5322 = n5309 & n5321 ;
  assign n5323 = ~n5318 & ~n5322 ;
  assign n5324 = ~n5320 & n5323 ;
  assign n5325 = ~n5319 & ~n5324 ;
  assign n5326 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[1]/P0001  ;
  assign n5327 = n5304 & n5326 ;
  assign n5328 = n5305 & ~n5327 ;
  assign n5329 = \u3_byte1_reg[1]/P0001  & ~n5310 ;
  assign n5330 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[9]/P0001  ;
  assign n5331 = n5309 & n5330 ;
  assign n5332 = ~n5327 & ~n5331 ;
  assign n5333 = ~n5329 & n5332 ;
  assign n5334 = ~n5328 & ~n5333 ;
  assign n5335 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[3]/P0001  ;
  assign n5336 = n5304 & n5335 ;
  assign n5337 = n5305 & ~n5336 ;
  assign n5338 = \u3_byte1_reg[3]/P0001  & ~n5310 ;
  assign n5339 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[11]/P0001  ;
  assign n5340 = n5309 & n5339 ;
  assign n5341 = ~n5336 & ~n5340 ;
  assign n5342 = ~n5338 & n5341 ;
  assign n5343 = ~n5337 & ~n5342 ;
  assign n5344 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[4]/P0001  ;
  assign n5345 = n5304 & n5344 ;
  assign n5346 = n5305 & ~n5345 ;
  assign n5347 = \u3_byte1_reg[4]/P0001  & ~n5310 ;
  assign n5348 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[12]/P0001  ;
  assign n5349 = n5309 & n5348 ;
  assign n5350 = ~n5345 & ~n5349 ;
  assign n5351 = ~n5347 & n5350 ;
  assign n5352 = ~n5346 & ~n5351 ;
  assign n5353 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[5]/P0001  ;
  assign n5354 = n5304 & n5353 ;
  assign n5355 = n5305 & ~n5354 ;
  assign n5356 = \u3_byte1_reg[5]/P0001  & ~n5310 ;
  assign n5357 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[13]/P0001  ;
  assign n5358 = n5309 & n5357 ;
  assign n5359 = ~n5354 & ~n5358 ;
  assign n5360 = ~n5356 & n5359 ;
  assign n5361 = ~n5355 & ~n5360 ;
  assign n5362 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[6]/P0001  ;
  assign n5363 = n5304 & n5362 ;
  assign n5364 = n5305 & ~n5363 ;
  assign n5365 = \u3_byte1_reg[6]/P0001  & ~n5310 ;
  assign n5366 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[14]/P0001  ;
  assign n5367 = n5309 & n5366 ;
  assign n5368 = ~n5363 & ~n5367 ;
  assign n5369 = ~n5365 & n5368 ;
  assign n5370 = ~n5364 & ~n5369 ;
  assign n5371 = \u5_pack_le1_reg/P0001  & \u7_mc_data_ir_reg[7]/P0001  ;
  assign n5372 = n5304 & n5371 ;
  assign n5373 = n5305 & ~n5372 ;
  assign n5374 = \u3_byte1_reg[7]/P0001  & ~n5310 ;
  assign n5375 = \u5_pack_le0_reg/P0001  & \u7_mc_data_ir_reg[15]/P0001  ;
  assign n5376 = n5309 & n5375 ;
  assign n5377 = ~n5372 & ~n5376 ;
  assign n5378 = ~n5374 & n5377 ;
  assign n5379 = ~n5373 & ~n5378 ;
  assign n5380 = wb_cyc_i_pad & ~n2165 ;
  assign n5381 = ~\u3_u0_wr_adr_reg[3]/NET0131  & n5380 ;
  assign n5382 = ~n1043 & n5381 ;
  assign n5383 = ~\u3_u0_wr_adr_reg[0]/NET0131  & n5380 ;
  assign n5384 = n1043 & n5383 ;
  assign n5385 = ~n5382 & ~n5384 ;
  assign n5386 = \u3_u0_wr_adr_reg[1]/NET0131  & n5380 ;
  assign n5387 = ~n1043 & n5386 ;
  assign n5388 = \u3_u0_wr_adr_reg[2]/NET0131  & n5380 ;
  assign n5389 = n1043 & n5388 ;
  assign n5390 = ~n5387 & ~n5389 ;
  assign n5391 = ~n1043 & n5388 ;
  assign n5392 = \u3_u0_wr_adr_reg[3]/NET0131  & n5380 ;
  assign n5393 = n1043 & n5392 ;
  assign n5394 = ~n5391 & ~n5393 ;
  assign n5395 = ~\u0_init_req_reg/NET0131  & n1923 ;
  assign n5396 = ~\u4_rfr_req_reg/NET0131  & \u5_state_reg[1]/NET0131  ;
  assign n5397 = n5395 & n5396 ;
  assign n5398 = ~n1255 & ~n1316 ;
  assign n5399 = ~\u5_state_reg[18]/NET0131  & ~n5398 ;
  assign n5400 = ~n1450 & ~n5399 ;
  assign n5401 = n3717 & ~n5400 ;
  assign n5402 = n3732 & n5401 ;
  assign n5403 = ~n5397 & ~n5402 ;
  assign n5404 = \wb_addr_i[0]_pad  & ~n2733 ;
  assign n5405 = ~n2730 & n5404 ;
  assign n5406 = n2740 & n5405 ;
  assign n5407 = \wb_addr_i[2]_pad  & ~n2733 ;
  assign n5408 = ~n2730 & n5407 ;
  assign n5409 = ~n2740 & n5408 ;
  assign n5410 = \wb_addr_i[1]_pad  & ~n2739 ;
  assign n5411 = ~n2736 & n5410 ;
  assign n5412 = ~n2734 & n5411 ;
  assign n5413 = ~n5409 & ~n5412 ;
  assign n5414 = ~n5406 & n5413 ;
  assign n5415 = ~n3439 & ~n5414 ;
  assign n5416 = ~\u1_u0_out_r_reg[0]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5417 = ~n3424 & n5416 ;
  assign n5418 = ~\u1_acs_addr_reg[0]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5419 = ~\u1_acs_addr_reg[0]/P0001  & n963 ;
  assign n5420 = ~n3423 & n5419 ;
  assign n5421 = ~n5418 & ~n5420 ;
  assign n5422 = n3439 & n5421 ;
  assign n5423 = ~n5417 & n5422 ;
  assign n5424 = ~n5415 & ~n5423 ;
  assign n5425 = ~\u1_u0_out_r_reg[10]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5426 = ~n3424 & n5425 ;
  assign n5427 = ~\u1_acs_addr_reg[10]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5428 = ~\u1_acs_addr_reg[10]/P0001  & n963 ;
  assign n5429 = ~n3423 & n5428 ;
  assign n5430 = ~n5427 & ~n5429 ;
  assign n5431 = n3439 & n5430 ;
  assign n5432 = ~n5426 & n5431 ;
  assign n5433 = n2740 & n5102 ;
  assign n5434 = ~n5163 & ~n5214 ;
  assign n5435 = ~n5433 & n5434 ;
  assign n5436 = ~n3439 & ~n5435 ;
  assign n5437 = ~n5432 & ~n5436 ;
  assign n5438 = \wb_addr_i[2]_pad  & ~n2739 ;
  assign n5439 = ~n2736 & n5438 ;
  assign n5440 = ~n2734 & n5439 ;
  assign n5441 = \wb_addr_i[3]_pad  & ~n2733 ;
  assign n5442 = ~n2730 & n5441 ;
  assign n5443 = ~n2740 & n5442 ;
  assign n5444 = \wb_addr_i[1]_pad  & ~n2733 ;
  assign n5445 = ~n2730 & n5444 ;
  assign n5446 = n2740 & n5445 ;
  assign n5447 = ~n5443 & ~n5446 ;
  assign n5448 = ~n5440 & n5447 ;
  assign n5449 = ~n3439 & ~n5448 ;
  assign n5450 = ~\u1_u0_out_r_reg[1]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5451 = ~n3424 & n5450 ;
  assign n5452 = ~\u1_acs_addr_reg[1]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5453 = ~\u1_acs_addr_reg[1]/P0001  & n963 ;
  assign n5454 = ~n3423 & n5453 ;
  assign n5455 = ~n5452 & ~n5454 ;
  assign n5456 = n3439 & n5455 ;
  assign n5457 = ~n5451 & n5456 ;
  assign n5458 = ~n5449 & ~n5457 ;
  assign n5459 = n2740 & n5408 ;
  assign n5460 = \wb_addr_i[3]_pad  & ~n2739 ;
  assign n5461 = ~n2736 & n5460 ;
  assign n5462 = ~n2734 & n5461 ;
  assign n5463 = ~n2740 & n5067 ;
  assign n5464 = ~n5462 & ~n5463 ;
  assign n5465 = ~n5459 & n5464 ;
  assign n5466 = ~n3439 & ~n5465 ;
  assign n5467 = ~\u1_u0_out_r_reg[2]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5468 = ~n3424 & n5467 ;
  assign n5469 = ~\u1_acs_addr_reg[2]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5470 = ~\u1_acs_addr_reg[2]/P0001  & n963 ;
  assign n5471 = ~n3423 & n5470 ;
  assign n5472 = ~n5469 & ~n5471 ;
  assign n5473 = n3439 & n5472 ;
  assign n5474 = ~n5468 & n5473 ;
  assign n5475 = ~n5466 & ~n5474 ;
  assign n5476 = n2740 & n5442 ;
  assign n5477 = \wb_addr_i[4]_pad  & ~n2739 ;
  assign n5478 = ~n2736 & n5477 ;
  assign n5479 = ~n2734 & n5478 ;
  assign n5480 = \wb_addr_i[5]_pad  & ~n2733 ;
  assign n5481 = ~n2730 & n5480 ;
  assign n5482 = ~n2740 & n5481 ;
  assign n5483 = ~n5479 & ~n5482 ;
  assign n5484 = ~n5476 & n5483 ;
  assign n5485 = ~n3439 & ~n5484 ;
  assign n5486 = ~\u1_u0_out_r_reg[3]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5487 = ~n3424 & n5486 ;
  assign n5488 = ~\u1_acs_addr_reg[3]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5489 = ~\u1_acs_addr_reg[3]/P0001  & n963 ;
  assign n5490 = ~n3423 & n5489 ;
  assign n5491 = ~n5488 & ~n5490 ;
  assign n5492 = n3439 & n5491 ;
  assign n5493 = ~n5487 & n5492 ;
  assign n5494 = ~n5485 & ~n5493 ;
  assign n5495 = n2740 & n5481 ;
  assign n5496 = \wb_addr_i[6]_pad  & ~n2739 ;
  assign n5497 = ~n2736 & n5496 ;
  assign n5498 = ~n2734 & n5497 ;
  assign n5499 = ~n2740 & n4949 ;
  assign n5500 = ~n5498 & ~n5499 ;
  assign n5501 = ~n5495 & n5500 ;
  assign n5502 = ~n3439 & ~n5501 ;
  assign n5503 = ~\u1_u0_out_r_reg[5]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5504 = ~n3424 & n5503 ;
  assign n5505 = ~\u1_acs_addr_reg[5]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5506 = ~\u1_acs_addr_reg[5]/P0001  & n963 ;
  assign n5507 = ~n3423 & n5506 ;
  assign n5508 = ~n5505 & ~n5507 ;
  assign n5509 = n3439 & n5508 ;
  assign n5510 = ~n5504 & n5509 ;
  assign n5511 = ~n5502 & ~n5510 ;
  assign n5512 = n2740 & n5073 ;
  assign n5513 = \wb_addr_i[7]_pad  & ~n2739 ;
  assign n5514 = ~n2736 & n5513 ;
  assign n5515 = ~n2734 & n5514 ;
  assign n5516 = ~n2740 & n5096 ;
  assign n5517 = ~n5515 & ~n5516 ;
  assign n5518 = ~n5512 & n5517 ;
  assign n5519 = ~n3439 & ~n5518 ;
  assign n5520 = ~\u1_u0_out_r_reg[6]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5521 = ~n3424 & n5520 ;
  assign n5522 = ~\u1_acs_addr_reg[6]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5523 = ~\u1_acs_addr_reg[6]/P0001  & n963 ;
  assign n5524 = ~n3423 & n5523 ;
  assign n5525 = ~n5522 & ~n5524 ;
  assign n5526 = n3439 & n5525 ;
  assign n5527 = ~n5521 & n5526 ;
  assign n5528 = ~n5519 & ~n5527 ;
  assign n5529 = ~\u1_u0_out_r_reg[9]/P0001  & \u5_tmr2_done_reg/NET0131  ;
  assign n5530 = ~n3424 & n5529 ;
  assign n5531 = ~\u1_acs_addr_reg[9]/P0001  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5532 = ~\u1_acs_addr_reg[9]/P0001  & n963 ;
  assign n5533 = ~n3423 & n5532 ;
  assign n5534 = ~n5531 & ~n5533 ;
  assign n5535 = n3439 & n5534 ;
  assign n5536 = ~n5530 & n5535 ;
  assign n5537 = n2740 & n4955 ;
  assign n5538 = ~n5157 & ~n5188 ;
  assign n5539 = ~n5537 & n5538 ;
  assign n5540 = ~n3439 & ~n5539 ;
  assign n5541 = ~n5536 & ~n5540 ;
  assign n5542 = ~n1094 & n1251 ;
  assign n5543 = ~\u5_cnt_reg/NET0131  & ~n5542 ;
  assign n5544 = wb_stb_i_pad & ~n2191 ;
  assign n5545 = \u5_wb_cycle_reg/NET0131  & wb_cyc_i_pad ;
  assign n5546 = ~n5544 & n5545 ;
  assign n5547 = ~n1930 & ~n5546 ;
  assign n5548 = \mem_ack_r_reg/P0001  & \u5_wr_cycle_reg/NET0131  ;
  assign n5549 = ~\u5_wr_cycle_reg/NET0131  & wb_stb_i_pad ;
  assign n5550 = ~n5548 & ~n5549 ;
  assign n5551 = \u1_col_adr_reg[8]/P0001  & n5550 ;
  assign n5552 = \wb_addr_i[10]_pad  & ~n5550 ;
  assign n5553 = n2740 & n5552 ;
  assign n5554 = ~n5110 & n5553 ;
  assign n5555 = ~n2735 & n5554 ;
  assign n5556 = ~n5551 & ~n5555 ;
  assign n5557 = \u1_acs_addr_reg[7]/P0001  & n5146 ;
  assign n5558 = ~\u1_acs_addr_reg[7]/P0001  & ~n5146 ;
  assign n5559 = ~n5557 & ~n5558 ;
  assign n5560 = \u5_state_reg[61]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n5561 = ~\u7_mc_ack_r_reg/NET0131  & ~n5560 ;
  assign n5562 = n1009 & ~n5561 ;
  assign n5563 = n1151 & n5562 ;
  assign n5564 = n1115 & n5563 ;
  assign n5565 = \u5_state_reg[61]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n5566 = ~n5564 & ~n5565 ;
  assign n5567 = ~n1157 & ~n5564 ;
  assign n5568 = n1504 & n5567 ;
  assign n5569 = ~n5566 & ~n5568 ;
  assign n5570 = ~\u0_csr_r2_reg[1]/NET0131  & \u4_ps_cnt_reg[1]/NET0131  ;
  assign n5571 = \u0_csr_r2_reg[4]/NET0131  & ~\u4_ps_cnt_reg[4]/NET0131  ;
  assign n5572 = ~n5570 & ~n5571 ;
  assign n5573 = ~\u0_csr_r2_reg[4]/NET0131  & \u4_ps_cnt_reg[4]/NET0131  ;
  assign n5574 = ~\u0_csr_r2_reg[2]/NET0131  & \u4_ps_cnt_reg[2]/NET0131  ;
  assign n5575 = ~n5573 & ~n5574 ;
  assign n5576 = n5572 & n5575 ;
  assign n5577 = ~\u0_csr_r2_reg[5]/NET0131  & ~\u4_ps_cnt_reg[5]/NET0131  ;
  assign n5578 = \u0_csr_r2_reg[5]/NET0131  & \u4_ps_cnt_reg[5]/NET0131  ;
  assign n5579 = ~n5577 & ~n5578 ;
  assign n5580 = ~\u0_csr_r2_reg[7]/NET0131  & ~\u4_ps_cnt_reg[7]/NET0131  ;
  assign n5581 = \u0_csr_r2_reg[7]/NET0131  & \u4_ps_cnt_reg[7]/NET0131  ;
  assign n5582 = ~n5580 & ~n5581 ;
  assign n5583 = ~n5579 & ~n5582 ;
  assign n5584 = n5576 & n5583 ;
  assign n5585 = \u0_csr_r2_reg[0]/NET0131  & ~\u4_ps_cnt_reg[0]/NET0131  ;
  assign n5586 = \u0_csr_r2_reg[3]/NET0131  & ~\u4_ps_cnt_reg[3]/NET0131  ;
  assign n5587 = ~n5585 & ~n5586 ;
  assign n5588 = ~\u0_csr_r2_reg[0]/NET0131  & \u4_ps_cnt_reg[0]/NET0131  ;
  assign n5589 = \u0_csr_r2_reg[1]/NET0131  & ~\u4_ps_cnt_reg[1]/NET0131  ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5591 = n5587 & n5590 ;
  assign n5592 = \u0_csr_r2_reg[2]/NET0131  & ~\u4_ps_cnt_reg[2]/NET0131  ;
  assign n5593 = \u0_csr_r2_reg[6]/NET0131  & ~\u4_ps_cnt_reg[6]/NET0131  ;
  assign n5594 = ~n5592 & ~n5593 ;
  assign n5595 = ~\u0_csr_r2_reg[6]/NET0131  & \u4_ps_cnt_reg[6]/NET0131  ;
  assign n5596 = ~\u0_csr_r2_reg[3]/NET0131  & \u4_ps_cnt_reg[3]/NET0131  ;
  assign n5597 = ~n5595 & ~n5596 ;
  assign n5598 = n5594 & n5597 ;
  assign n5599 = n5591 & n5598 ;
  assign n5600 = n5584 & n5599 ;
  assign n5601 = ~\u0_csr_r2_reg[4]/NET0131  & ~\u0_csr_r2_reg[5]/NET0131  ;
  assign n5602 = ~\u0_csr_r2_reg[6]/NET0131  & ~\u0_csr_r2_reg[7]/NET0131  ;
  assign n5603 = n5601 & n5602 ;
  assign n5604 = ~\u0_csr_r2_reg[0]/NET0131  & ~\u0_csr_r2_reg[1]/NET0131  ;
  assign n5605 = ~\u0_csr_r2_reg[2]/NET0131  & ~\u0_csr_r2_reg[3]/NET0131  ;
  assign n5606 = n5604 & n5605 ;
  assign n5607 = n5603 & n5606 ;
  assign n5608 = n5600 & ~n5607 ;
  assign n5609 = \u4_ps_cnt_reg[0]/NET0131  & \u4_rfr_en_reg/NET0131  ;
  assign n5610 = \u4_ps_cnt_reg[1]/NET0131  & \u4_ps_cnt_reg[2]/NET0131  ;
  assign n5611 = n5609 & n5610 ;
  assign n5612 = \u4_ps_cnt_reg[3]/NET0131  & \u4_ps_cnt_reg[4]/NET0131  ;
  assign n5613 = n5611 & n5612 ;
  assign n5614 = \u4_ps_cnt_reg[3]/NET0131  & n5611 ;
  assign n5615 = ~\u4_ps_cnt_reg[4]/NET0131  & ~n5614 ;
  assign n5616 = ~n5613 & ~n5615 ;
  assign n5617 = ~n5608 & n5616 ;
  assign n5618 = \u4_rfr_ce_reg/NET0131  & \u4_rfr_cnt_reg[0]/NET0131  ;
  assign n5619 = \u4_rfr_cnt_reg[1]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5620 = ~n5618 & n5619 ;
  assign n5621 = ~\u4_rfr_cnt_reg[1]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5622 = n5618 & n5621 ;
  assign n5623 = ~n5620 & ~n5622 ;
  assign n5624 = ~\u5_state_reg[20]/NET0131  & n977 ;
  assign n5625 = ~\u5_state_reg[7]/NET0131  & n991 ;
  assign n5626 = n5624 & n5625 ;
  assign n5627 = n1056 & n5626 ;
  assign n5628 = n1065 & n5627 ;
  assign n5629 = ~\u5_state_reg[33]/NET0131  & ~\u5_state_reg[34]/NET0131  ;
  assign n5630 = \u5_state_reg[33]/NET0131  & \u5_state_reg[34]/NET0131  ;
  assign n5631 = ~\u5_state_reg[0]/NET0131  & ~\u5_state_reg[35]/NET0131  ;
  assign n5632 = ~n5630 & n5631 ;
  assign n5633 = ~n5629 & n5632 ;
  assign n5634 = n1057 & n3728 ;
  assign n5635 = n3726 & n5634 ;
  assign n5636 = n5633 & n5635 ;
  assign n5637 = n3704 & n5636 ;
  assign n5638 = n5628 & n5637 ;
  assign n5639 = n3724 & n5638 ;
  assign n5640 = ~\u0_init_req_reg/NET0131  & ~\u0_lmr_req_reg/NET0131  ;
  assign n5641 = ~\u4_rfr_req_reg/NET0131  & \u5_state_reg[35]/NET0131  ;
  assign n5642 = ~\u5_susp_req_r_reg/NET0131  & n5641 ;
  assign n5643 = n5640 & n5642 ;
  assign n5644 = n1898 & n5643 ;
  assign n5645 = ~n5639 & ~n5644 ;
  assign n5646 = ~\u4_rfr_ce_reg/NET0131  & ~\u4_rfr_cnt_reg[0]/NET0131  ;
  assign n5647 = ~\u5_rfr_ack_r_reg/NET0131  & ~n5618 ;
  assign n5648 = ~n5646 & n5647 ;
  assign n5649 = n4981 & n5618 ;
  assign n5650 = \u4_rfr_cnt_reg[2]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5651 = n5618 & n5619 ;
  assign n5652 = ~n5650 & ~n5651 ;
  assign n5653 = ~n5649 & ~n5652 ;
  assign n5654 = \u4_rfr_cnt_reg[3]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5655 = ~n5649 & n5654 ;
  assign n5656 = ~\u4_rfr_cnt_reg[3]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5657 = n5649 & n5656 ;
  assign n5658 = ~n5655 & ~n5657 ;
  assign n5659 = n4989 & n5649 ;
  assign n5660 = \u4_rfr_cnt_reg[4]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5661 = n5649 & n5654 ;
  assign n5662 = ~n5660 & ~n5661 ;
  assign n5663 = ~n5659 & ~n5662 ;
  assign n5664 = ~\u4_rfr_cnt_reg[5]/NET0131  & ~n5659 ;
  assign n5665 = \u4_rfr_cnt_reg[3]/NET0131  & \u4_rfr_cnt_reg[5]/NET0131  ;
  assign n5666 = \u4_rfr_cnt_reg[4]/NET0131  & n5665 ;
  assign n5667 = n5649 & n5666 ;
  assign n5668 = ~\u5_rfr_ack_r_reg/NET0131  & ~n5667 ;
  assign n5669 = ~n5664 & n5668 ;
  assign n5670 = \u4_rfr_cnt_reg[6]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5671 = ~n5667 & n5670 ;
  assign n5672 = ~\u4_rfr_cnt_reg[6]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5673 = n5667 & n5672 ;
  assign n5674 = ~n5671 & ~n5673 ;
  assign n5675 = \u4_rfr_cnt_reg[6]/NET0131  & \u4_rfr_cnt_reg[7]/NET0131  ;
  assign n5676 = n5667 & n5675 ;
  assign n5677 = \u4_rfr_cnt_reg[7]/NET0131  & ~\u5_rfr_ack_r_reg/NET0131  ;
  assign n5678 = n5667 & n5670 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5680 = ~n5676 & ~n5679 ;
  assign n5681 = \u5_cs_le_reg/P0001  & n1045 ;
  assign n5682 = \u0_wp_err_reg/NET0131  & wb_cyc_i_pad ;
  assign n5683 = ~n5681 & n5682 ;
  assign n5684 = \u0_u0_csc_reg[8]/P0001  & n4214 ;
  assign n5685 = n4199 & n5684 ;
  assign n5686 = \u0_u1_csc_reg[8]/P0001  & n4256 ;
  assign n5687 = n4241 & n5686 ;
  assign n5688 = ~n5685 & ~n5687 ;
  assign n5689 = \u5_cs_le_reg/P0001  & wb_we_i_pad ;
  assign n5690 = n1045 & n5689 ;
  assign n5691 = ~n5688 & n5690 ;
  assign n5692 = ~n5683 & ~n5691 ;
  assign n5693 = \u5_mc_adv_r1_reg/NET0131  & \u5_mc_le_reg/NET0131  ;
  assign n5694 = n1899 & ~n3258 ;
  assign n5695 = ~n1112 & ~n5694 ;
  assign n5696 = n1023 & n1111 ;
  assign n5697 = ~\u5_mc_le_reg/NET0131  & ~n5696 ;
  assign n5698 = n5695 & n5697 ;
  assign n5699 = ~n5693 & ~n5698 ;
  assign n5700 = ~n5114 & n5122 ;
  assign n5701 = n5122 & ~n5200 ;
  assign n5702 = n5204 & n5701 ;
  assign n5703 = ~n5700 & ~n5702 ;
  assign n5704 = ~n5114 & ~n5122 ;
  assign n5705 = ~n3647 & ~n5122 ;
  assign n5706 = n5176 & n5705 ;
  assign n5707 = ~n5704 & ~n5706 ;
  assign n5708 = n5703 & n5707 ;
  assign n5709 = \u5_cmd_asserted_reg/NET0131  & n1419 ;
  assign n5710 = n1096 & n5709 ;
  assign n5711 = n1078 & n5710 ;
  assign n5712 = ~\u5_ir_cnt_reg[0]/P0001  & n5711 ;
  assign n5713 = \u5_ir_cnt_reg[1]/P0001  & ~n5712 ;
  assign n5714 = ~\u5_ir_cnt_reg[0]/P0001  & ~\u5_ir_cnt_reg[1]/P0001  ;
  assign n5715 = n5711 & n5714 ;
  assign n5716 = ~\u5_state_reg[22]/NET0131  & ~n5715 ;
  assign n5717 = ~n5713 & n5716 ;
  assign n5718 = \u4_ps_cnt_reg[3]/NET0131  & \u4_ps_cnt_reg[5]/NET0131  ;
  assign n5719 = \u4_ps_cnt_reg[4]/NET0131  & n5718 ;
  assign n5720 = n5611 & n5719 ;
  assign n5721 = \u4_ps_cnt_reg[6]/NET0131  & n5720 ;
  assign n5722 = ~\u4_ps_cnt_reg[7]/NET0131  & ~n5721 ;
  assign n5723 = \u4_ps_cnt_reg[6]/NET0131  & \u4_ps_cnt_reg[7]/NET0131  ;
  assign n5724 = n5720 & n5723 ;
  assign n5725 = ~n5722 & ~n5724 ;
  assign n5726 = ~n5608 & n5725 ;
  assign n5727 = ~\u5_ir_cnt_reg[2]/P0001  & ~\u5_ir_cnt_reg[3]/P0001  ;
  assign n5728 = n5714 & n5727 ;
  assign n5729 = n5711 & n5728 ;
  assign n5730 = ~\u5_state_reg[22]/NET0131  & n5729 ;
  assign n5731 = ~\u5_ir_cnt_reg[2]/P0001  & n5714 ;
  assign n5732 = n5711 & n5731 ;
  assign n5733 = \u5_ir_cnt_reg[3]/P0001  & ~\u5_state_reg[22]/NET0131  ;
  assign n5734 = ~n5732 & n5733 ;
  assign n5735 = ~n5730 & ~n5734 ;
  assign n5736 = \u3_u0_wr_adr_reg[1]/NET0131  & ~n1043 ;
  assign n5737 = \u3_u0_wr_adr_reg[2]/NET0131  & ~n1043 ;
  assign n5738 = \u5_ir_cnt_reg[0]/P0001  & ~\u5_state_reg[22]/NET0131  ;
  assign n5739 = ~n5711 & n5738 ;
  assign n5740 = ~\u5_ir_cnt_reg[0]/P0001  & ~\u5_state_reg[22]/NET0131  ;
  assign n5741 = n5711 & n5740 ;
  assign n5742 = ~n5739 & ~n5741 ;
  assign n5743 = \u5_ir_cnt_reg[2]/P0001  & ~\u5_state_reg[22]/NET0131  ;
  assign n5744 = ~n5715 & n5743 ;
  assign n5745 = ~\u5_ir_cnt_reg[2]/P0001  & ~\u5_state_reg[22]/NET0131  ;
  assign n5746 = n5715 & n5745 ;
  assign n5747 = ~n5744 & ~n5746 ;
  assign n5748 = ~\u1_row_adr_reg[6]/P0001  & \u2_u1_b3_last_row_reg[6]/P0001  ;
  assign n5749 = \u1_row_adr_reg[7]/P0001  & ~\u2_u1_b3_last_row_reg[7]/P0001  ;
  assign n5750 = ~\u1_row_adr_reg[7]/P0001  & \u2_u1_b3_last_row_reg[7]/P0001  ;
  assign n5751 = ~n5749 & ~n5750 ;
  assign n5752 = ~n5748 & n5751 ;
  assign n5753 = \u1_row_adr_reg[0]/P0001  & ~\u2_u1_b3_last_row_reg[0]/P0001  ;
  assign n5754 = \u1_row_adr_reg[8]/P0001  & ~\u2_u1_b3_last_row_reg[8]/P0001  ;
  assign n5755 = ~n5753 & ~n5754 ;
  assign n5756 = ~\u1_row_adr_reg[11]/P0001  & \u2_u1_b3_last_row_reg[11]/P0001  ;
  assign n5757 = ~\u1_row_adr_reg[8]/P0001  & \u2_u1_b3_last_row_reg[8]/P0001  ;
  assign n5758 = ~n5756 & ~n5757 ;
  assign n5759 = n5755 & n5758 ;
  assign n5760 = ~\u1_row_adr_reg[1]/P0001  & \u2_u1_b3_last_row_reg[1]/P0001  ;
  assign n5761 = ~\u1_row_adr_reg[12]/P0001  & \u2_u1_b3_last_row_reg[12]/P0001  ;
  assign n5762 = ~n5760 & ~n5761 ;
  assign n5763 = \u1_row_adr_reg[1]/P0001  & ~\u2_u1_b3_last_row_reg[1]/P0001  ;
  assign n5764 = ~\u1_row_adr_reg[4]/P0001  & \u2_u1_b3_last_row_reg[4]/P0001  ;
  assign n5765 = ~n5763 & ~n5764 ;
  assign n5766 = n5762 & n5765 ;
  assign n5767 = n5759 & n5766 ;
  assign n5768 = n5752 & n5767 ;
  assign n5769 = \u1_row_adr_reg[11]/P0001  & ~\u2_u1_b3_last_row_reg[11]/P0001  ;
  assign n5770 = ~\u1_row_adr_reg[0]/P0001  & \u2_u1_b3_last_row_reg[0]/P0001  ;
  assign n5771 = ~n5769 & ~n5770 ;
  assign n5772 = \u1_row_adr_reg[2]/P0001  & ~\u2_u1_b3_last_row_reg[2]/P0001  ;
  assign n5773 = \u1_row_adr_reg[12]/P0001  & ~\u2_u1_b3_last_row_reg[12]/P0001  ;
  assign n5774 = ~n5772 & ~n5773 ;
  assign n5775 = n5771 & n5774 ;
  assign n5776 = ~\u1_row_adr_reg[10]/P0001  & ~\u2_u1_b3_last_row_reg[10]/P0001  ;
  assign n5777 = \u1_row_adr_reg[10]/P0001  & \u2_u1_b3_last_row_reg[10]/P0001  ;
  assign n5778 = ~n5776 & ~n5777 ;
  assign n5779 = \u1_row_adr_reg[3]/P0001  & ~\u2_u1_b3_last_row_reg[3]/P0001  ;
  assign n5780 = n3793 & ~n5779 ;
  assign n5781 = ~n5778 & n5780 ;
  assign n5782 = n5775 & n5781 ;
  assign n5783 = ~\u1_row_adr_reg[5]/P0001  & \u2_u1_b3_last_row_reg[5]/P0001  ;
  assign n5784 = ~\u1_row_adr_reg[9]/P0001  & \u2_u1_b3_last_row_reg[9]/P0001  ;
  assign n5785 = ~n5783 & ~n5784 ;
  assign n5786 = ~\u1_row_adr_reg[2]/P0001  & \u2_u1_b3_last_row_reg[2]/P0001  ;
  assign n5787 = \u1_row_adr_reg[4]/P0001  & ~\u2_u1_b3_last_row_reg[4]/P0001  ;
  assign n5788 = ~n5786 & ~n5787 ;
  assign n5789 = n5785 & n5788 ;
  assign n5790 = \u1_row_adr_reg[9]/P0001  & ~\u2_u1_b3_last_row_reg[9]/P0001  ;
  assign n5791 = \u1_row_adr_reg[5]/P0001  & ~\u2_u1_b3_last_row_reg[5]/P0001  ;
  assign n5792 = ~n5790 & ~n5791 ;
  assign n5793 = ~\u1_row_adr_reg[3]/P0001  & \u2_u1_b3_last_row_reg[3]/P0001  ;
  assign n5794 = \u1_row_adr_reg[6]/P0001  & ~\u2_u1_b3_last_row_reg[6]/P0001  ;
  assign n5795 = ~n5793 & ~n5794 ;
  assign n5796 = n5792 & n5795 ;
  assign n5797 = n5789 & n5796 ;
  assign n5798 = n5782 & n5797 ;
  assign n5799 = n5768 & n5798 ;
  assign n5800 = ~\u1_row_adr_reg[3]/P0001  & \u2_u1_b2_last_row_reg[3]/P0001  ;
  assign n5801 = \u1_row_adr_reg[3]/P0001  & ~\u2_u1_b2_last_row_reg[3]/P0001  ;
  assign n5802 = ~\u1_row_adr_reg[8]/P0001  & \u2_u1_b2_last_row_reg[8]/P0001  ;
  assign n5803 = ~n5801 & ~n5802 ;
  assign n5804 = ~n5800 & n5803 ;
  assign n5805 = ~\u1_row_adr_reg[4]/P0001  & \u2_u1_b2_last_row_reg[4]/P0001  ;
  assign n5806 = ~\u1_row_adr_reg[2]/P0001  & \u2_u1_b2_last_row_reg[2]/P0001  ;
  assign n5807 = ~n5805 & ~n5806 ;
  assign n5808 = \u1_row_adr_reg[8]/P0001  & ~\u2_u1_b2_last_row_reg[8]/P0001  ;
  assign n5809 = ~\u1_row_adr_reg[0]/P0001  & \u2_u1_b2_last_row_reg[0]/P0001  ;
  assign n5810 = ~n5808 & ~n5809 ;
  assign n5811 = n5807 & n5810 ;
  assign n5812 = ~\u1_row_adr_reg[7]/P0001  & \u2_u1_b2_last_row_reg[7]/P0001  ;
  assign n5813 = \u1_row_adr_reg[2]/P0001  & ~\u2_u1_b2_last_row_reg[2]/P0001  ;
  assign n5814 = ~n5812 & ~n5813 ;
  assign n5815 = \u1_row_adr_reg[7]/P0001  & ~\u2_u1_b2_last_row_reg[7]/P0001  ;
  assign n5816 = \u1_row_adr_reg[0]/P0001  & ~\u2_u1_b2_last_row_reg[0]/P0001  ;
  assign n5817 = ~n5815 & ~n5816 ;
  assign n5818 = n5814 & n5817 ;
  assign n5819 = n5811 & n5818 ;
  assign n5820 = n5804 & n5819 ;
  assign n5821 = \u1_row_adr_reg[1]/P0001  & ~\u2_u1_b2_last_row_reg[1]/P0001  ;
  assign n5822 = ~\u1_row_adr_reg[11]/P0001  & \u2_u1_b2_last_row_reg[11]/P0001  ;
  assign n5823 = ~n5821 & ~n5822 ;
  assign n5824 = \u1_row_adr_reg[11]/P0001  & ~\u2_u1_b2_last_row_reg[11]/P0001  ;
  assign n5825 = \u1_row_adr_reg[9]/P0001  & ~\u2_u1_b2_last_row_reg[9]/P0001  ;
  assign n5826 = ~n5824 & ~n5825 ;
  assign n5827 = n5823 & n5826 ;
  assign n5828 = \u1_row_adr_reg[12]/P0001  & ~\u2_u1_b2_last_row_reg[12]/P0001  ;
  assign n5829 = n3751 & ~n5828 ;
  assign n5830 = \u1_row_adr_reg[6]/P0001  & ~\u2_u1_b2_last_row_reg[6]/P0001  ;
  assign n5831 = \u1_row_adr_reg[5]/P0001  & ~\u2_u1_b2_last_row_reg[5]/P0001  ;
  assign n5832 = ~n5830 & ~n5831 ;
  assign n5833 = n5829 & n5832 ;
  assign n5834 = n5827 & n5833 ;
  assign n5835 = ~\u1_row_adr_reg[5]/P0001  & \u2_u1_b2_last_row_reg[5]/P0001  ;
  assign n5836 = ~\u1_row_adr_reg[9]/P0001  & \u2_u1_b2_last_row_reg[9]/P0001  ;
  assign n5837 = ~n5835 & ~n5836 ;
  assign n5838 = \u1_row_adr_reg[10]/P0001  & ~\u2_u1_b2_last_row_reg[10]/P0001  ;
  assign n5839 = \u1_row_adr_reg[4]/P0001  & ~\u2_u1_b2_last_row_reg[4]/P0001  ;
  assign n5840 = ~n5838 & ~n5839 ;
  assign n5841 = n5837 & n5840 ;
  assign n5842 = ~\u1_row_adr_reg[10]/P0001  & \u2_u1_b2_last_row_reg[10]/P0001  ;
  assign n5843 = ~\u1_row_adr_reg[1]/P0001  & \u2_u1_b2_last_row_reg[1]/P0001  ;
  assign n5844 = ~n5842 & ~n5843 ;
  assign n5845 = ~\u1_row_adr_reg[6]/P0001  & \u2_u1_b2_last_row_reg[6]/P0001  ;
  assign n5846 = ~\u1_row_adr_reg[12]/P0001  & \u2_u1_b2_last_row_reg[12]/P0001  ;
  assign n5847 = ~n5845 & ~n5846 ;
  assign n5848 = n5844 & n5847 ;
  assign n5849 = n5841 & n5848 ;
  assign n5850 = n5834 & n5849 ;
  assign n5851 = n5820 & n5850 ;
  assign n5852 = ~n5799 & ~n5851 ;
  assign n5853 = ~\u1_row_adr_reg[4]/P0001  & \u2_u1_b0_last_row_reg[4]/P0001  ;
  assign n5854 = \u1_row_adr_reg[5]/P0001  & ~\u2_u1_b0_last_row_reg[5]/P0001  ;
  assign n5855 = ~\u1_bank_adr_reg[0]/P0001  & ~\u1_bank_adr_reg[1]/P0001  ;
  assign n5856 = ~n5854 & n5855 ;
  assign n5857 = ~n5853 & n5856 ;
  assign n5858 = \u1_row_adr_reg[2]/P0001  & ~\u2_u1_b0_last_row_reg[2]/P0001  ;
  assign n5859 = \u1_row_adr_reg[9]/P0001  & ~\u2_u1_b0_last_row_reg[9]/P0001  ;
  assign n5860 = ~n5858 & ~n5859 ;
  assign n5861 = \u1_row_adr_reg[10]/P0001  & ~\u2_u1_b0_last_row_reg[10]/P0001  ;
  assign n5862 = \u1_row_adr_reg[1]/P0001  & ~\u2_u1_b0_last_row_reg[1]/P0001  ;
  assign n5863 = ~n5861 & ~n5862 ;
  assign n5864 = n5860 & n5863 ;
  assign n5865 = \u1_row_adr_reg[6]/P0001  & ~\u2_u1_b0_last_row_reg[6]/P0001  ;
  assign n5866 = \u1_row_adr_reg[11]/P0001  & ~\u2_u1_b0_last_row_reg[11]/P0001  ;
  assign n5867 = ~n5865 & ~n5866 ;
  assign n5868 = \u1_row_adr_reg[3]/P0001  & ~\u2_u1_b0_last_row_reg[3]/P0001  ;
  assign n5869 = ~\u1_row_adr_reg[9]/P0001  & \u2_u1_b0_last_row_reg[9]/P0001  ;
  assign n5870 = ~n5868 & ~n5869 ;
  assign n5871 = n5867 & n5870 ;
  assign n5872 = n5864 & n5871 ;
  assign n5873 = n5857 & n5872 ;
  assign n5874 = ~\u1_row_adr_reg[10]/P0001  & \u2_u1_b0_last_row_reg[10]/P0001  ;
  assign n5875 = \u1_row_adr_reg[12]/P0001  & ~\u2_u1_b0_last_row_reg[12]/P0001  ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = \u1_row_adr_reg[4]/P0001  & ~\u2_u1_b0_last_row_reg[4]/P0001  ;
  assign n5878 = ~\u1_row_adr_reg[8]/P0001  & \u2_u1_b0_last_row_reg[8]/P0001  ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = n5876 & n5879 ;
  assign n5881 = ~\u1_row_adr_reg[7]/P0001  & ~\u2_u1_b0_last_row_reg[7]/P0001  ;
  assign n5882 = \u1_row_adr_reg[7]/P0001  & \u2_u1_b0_last_row_reg[7]/P0001  ;
  assign n5883 = ~n5881 & ~n5882 ;
  assign n5884 = ~\u1_row_adr_reg[0]/P0001  & ~\u2_u1_b0_last_row_reg[0]/P0001  ;
  assign n5885 = \u1_row_adr_reg[0]/P0001  & \u2_u1_b0_last_row_reg[0]/P0001  ;
  assign n5886 = ~n5884 & ~n5885 ;
  assign n5887 = ~n5883 & ~n5886 ;
  assign n5888 = n5880 & n5887 ;
  assign n5889 = ~\u1_row_adr_reg[5]/P0001  & \u2_u1_b0_last_row_reg[5]/P0001  ;
  assign n5890 = ~\u1_row_adr_reg[11]/P0001  & \u2_u1_b0_last_row_reg[11]/P0001  ;
  assign n5891 = ~n5889 & ~n5890 ;
  assign n5892 = ~\u1_row_adr_reg[1]/P0001  & \u2_u1_b0_last_row_reg[1]/P0001  ;
  assign n5893 = ~\u1_row_adr_reg[2]/P0001  & \u2_u1_b0_last_row_reg[2]/P0001  ;
  assign n5894 = ~n5892 & ~n5893 ;
  assign n5895 = n5891 & n5894 ;
  assign n5896 = ~\u1_row_adr_reg[3]/P0001  & \u2_u1_b0_last_row_reg[3]/P0001  ;
  assign n5897 = ~\u1_row_adr_reg[12]/P0001  & \u2_u1_b0_last_row_reg[12]/P0001  ;
  assign n5898 = ~n5896 & ~n5897 ;
  assign n5899 = \u1_row_adr_reg[8]/P0001  & ~\u2_u1_b0_last_row_reg[8]/P0001  ;
  assign n5900 = ~\u1_row_adr_reg[6]/P0001  & \u2_u1_b0_last_row_reg[6]/P0001  ;
  assign n5901 = ~n5899 & ~n5900 ;
  assign n5902 = n5898 & n5901 ;
  assign n5903 = n5895 & n5902 ;
  assign n5904 = n5888 & n5903 ;
  assign n5905 = n5873 & n5904 ;
  assign n5906 = ~\u1_row_adr_reg[3]/P0001  & \u2_u1_b1_last_row_reg[3]/P0001  ;
  assign n5907 = \u1_row_adr_reg[12]/P0001  & ~\u2_u1_b1_last_row_reg[12]/P0001  ;
  assign n5908 = \u1_row_adr_reg[3]/P0001  & ~\u2_u1_b1_last_row_reg[3]/P0001  ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5910 = ~n5906 & n5909 ;
  assign n5911 = \u1_row_adr_reg[1]/P0001  & ~\u2_u1_b1_last_row_reg[1]/P0001  ;
  assign n5912 = ~\u1_row_adr_reg[6]/P0001  & \u2_u1_b1_last_row_reg[6]/P0001  ;
  assign n5913 = ~n5911 & ~n5912 ;
  assign n5914 = \u1_row_adr_reg[5]/P0001  & ~\u2_u1_b1_last_row_reg[5]/P0001  ;
  assign n5915 = ~\u1_row_adr_reg[12]/P0001  & \u2_u1_b1_last_row_reg[12]/P0001  ;
  assign n5916 = ~n5914 & ~n5915 ;
  assign n5917 = n5913 & n5916 ;
  assign n5918 = \u1_row_adr_reg[9]/P0001  & ~\u2_u1_b1_last_row_reg[9]/P0001  ;
  assign n5919 = ~\u1_row_adr_reg[5]/P0001  & \u2_u1_b1_last_row_reg[5]/P0001  ;
  assign n5920 = ~n5918 & ~n5919 ;
  assign n5921 = ~\u1_row_adr_reg[10]/P0001  & \u2_u1_b1_last_row_reg[10]/P0001  ;
  assign n5922 = \u1_row_adr_reg[6]/P0001  & ~\u2_u1_b1_last_row_reg[6]/P0001  ;
  assign n5923 = ~n5921 & ~n5922 ;
  assign n5924 = n5920 & n5923 ;
  assign n5925 = n5917 & n5924 ;
  assign n5926 = n5910 & n5925 ;
  assign n5927 = ~\u1_row_adr_reg[7]/P0001  & \u2_u1_b1_last_row_reg[7]/P0001  ;
  assign n5928 = ~\u1_row_adr_reg[11]/P0001  & \u2_u1_b1_last_row_reg[11]/P0001  ;
  assign n5929 = ~n5927 & ~n5928 ;
  assign n5930 = \u1_row_adr_reg[8]/P0001  & ~\u2_u1_b1_last_row_reg[8]/P0001  ;
  assign n5931 = \u1_row_adr_reg[10]/P0001  & ~\u2_u1_b1_last_row_reg[10]/P0001  ;
  assign n5932 = ~n5930 & ~n5931 ;
  assign n5933 = n5929 & n5932 ;
  assign n5934 = \u1_row_adr_reg[11]/P0001  & ~\u2_u1_b1_last_row_reg[11]/P0001  ;
  assign n5935 = n3684 & ~n5934 ;
  assign n5936 = \u1_row_adr_reg[2]/P0001  & ~\u2_u1_b1_last_row_reg[2]/P0001  ;
  assign n5937 = \u1_row_adr_reg[0]/P0001  & ~\u2_u1_b1_last_row_reg[0]/P0001  ;
  assign n5938 = ~n5936 & ~n5937 ;
  assign n5939 = n5935 & n5938 ;
  assign n5940 = n5933 & n5939 ;
  assign n5941 = ~\u1_row_adr_reg[1]/P0001  & \u2_u1_b1_last_row_reg[1]/P0001  ;
  assign n5942 = ~\u1_row_adr_reg[8]/P0001  & \u2_u1_b1_last_row_reg[8]/P0001  ;
  assign n5943 = ~n5941 & ~n5942 ;
  assign n5944 = ~\u1_row_adr_reg[9]/P0001  & \u2_u1_b1_last_row_reg[9]/P0001  ;
  assign n5945 = ~\u1_row_adr_reg[2]/P0001  & \u2_u1_b1_last_row_reg[2]/P0001  ;
  assign n5946 = ~n5944 & ~n5945 ;
  assign n5947 = n5943 & n5946 ;
  assign n5948 = \u1_row_adr_reg[4]/P0001  & ~\u2_u1_b1_last_row_reg[4]/P0001  ;
  assign n5949 = ~\u1_row_adr_reg[0]/P0001  & \u2_u1_b1_last_row_reg[0]/P0001  ;
  assign n5950 = ~n5948 & ~n5949 ;
  assign n5951 = \u1_row_adr_reg[7]/P0001  & ~\u2_u1_b1_last_row_reg[7]/P0001  ;
  assign n5952 = ~\u1_row_adr_reg[4]/P0001  & \u2_u1_b1_last_row_reg[4]/P0001  ;
  assign n5953 = ~n5951 & ~n5952 ;
  assign n5954 = n5950 & n5953 ;
  assign n5955 = n5947 & n5954 ;
  assign n5956 = n5940 & n5955 ;
  assign n5957 = n5926 & n5956 ;
  assign n5958 = ~n5905 & ~n5957 ;
  assign n5959 = n5852 & n5958 ;
  assign n5960 = ~n1919 & ~n5959 ;
  assign n5961 = \u1_row_adr_reg[5]/P0001  & ~\u2_u0_b2_last_row_reg[5]/P0001  ;
  assign n5962 = \u1_row_adr_reg[11]/P0001  & ~\u2_u0_b2_last_row_reg[11]/P0001  ;
  assign n5963 = ~\u1_row_adr_reg[11]/P0001  & \u2_u0_b2_last_row_reg[11]/P0001  ;
  assign n5964 = ~n5962 & ~n5963 ;
  assign n5965 = ~n5961 & n5964 ;
  assign n5966 = ~\u1_row_adr_reg[10]/P0001  & \u2_u0_b2_last_row_reg[10]/P0001  ;
  assign n5967 = \u1_row_adr_reg[9]/P0001  & ~\u2_u0_b2_last_row_reg[9]/P0001  ;
  assign n5968 = ~n5966 & ~n5967 ;
  assign n5969 = ~\u1_row_adr_reg[8]/P0001  & \u2_u0_b2_last_row_reg[8]/P0001  ;
  assign n5970 = \u1_row_adr_reg[8]/P0001  & ~\u2_u0_b2_last_row_reg[8]/P0001  ;
  assign n5971 = ~n5969 & ~n5970 ;
  assign n5972 = n5968 & n5971 ;
  assign n5973 = ~\u1_row_adr_reg[2]/P0001  & \u2_u0_b2_last_row_reg[2]/P0001  ;
  assign n5974 = ~\u1_row_adr_reg[1]/P0001  & \u2_u0_b2_last_row_reg[1]/P0001  ;
  assign n5975 = ~n5973 & ~n5974 ;
  assign n5976 = ~\u1_row_adr_reg[9]/P0001  & \u2_u0_b2_last_row_reg[9]/P0001  ;
  assign n5977 = \u1_row_adr_reg[3]/P0001  & ~\u2_u0_b2_last_row_reg[3]/P0001  ;
  assign n5978 = ~n5976 & ~n5977 ;
  assign n5979 = n5975 & n5978 ;
  assign n5980 = n5972 & n5979 ;
  assign n5981 = n5965 & n5980 ;
  assign n5982 = \u1_row_adr_reg[7]/P0001  & ~\u2_u0_b2_last_row_reg[7]/P0001  ;
  assign n5983 = n3751 & ~n5982 ;
  assign n5984 = \u1_row_adr_reg[6]/P0001  & ~\u2_u0_b2_last_row_reg[6]/P0001  ;
  assign n5985 = \u1_row_adr_reg[2]/P0001  & ~\u2_u0_b2_last_row_reg[2]/P0001  ;
  assign n5986 = ~n5984 & ~n5985 ;
  assign n5987 = n5983 & n5986 ;
  assign n5988 = ~\u1_row_adr_reg[4]/P0001  & ~\u2_u0_b2_last_row_reg[4]/P0001  ;
  assign n5989 = \u1_row_adr_reg[4]/P0001  & \u2_u0_b2_last_row_reg[4]/P0001  ;
  assign n5990 = ~n5988 & ~n5989 ;
  assign n5991 = ~\u1_row_adr_reg[0]/P0001  & ~\u2_u0_b2_last_row_reg[0]/P0001  ;
  assign n5992 = \u1_row_adr_reg[0]/P0001  & \u2_u0_b2_last_row_reg[0]/P0001  ;
  assign n5993 = ~n5991 & ~n5992 ;
  assign n5994 = ~n5990 & ~n5993 ;
  assign n5995 = n5987 & n5994 ;
  assign n5996 = \u1_row_adr_reg[12]/P0001  & ~\u2_u0_b2_last_row_reg[12]/P0001  ;
  assign n5997 = ~\u1_row_adr_reg[12]/P0001  & \u2_u0_b2_last_row_reg[12]/P0001  ;
  assign n5998 = ~n5996 & ~n5997 ;
  assign n5999 = ~\u1_row_adr_reg[5]/P0001  & \u2_u0_b2_last_row_reg[5]/P0001  ;
  assign n6000 = \u1_row_adr_reg[10]/P0001  & ~\u2_u0_b2_last_row_reg[10]/P0001  ;
  assign n6001 = ~n5999 & ~n6000 ;
  assign n6002 = n5998 & n6001 ;
  assign n6003 = ~\u1_row_adr_reg[6]/P0001  & \u2_u0_b2_last_row_reg[6]/P0001  ;
  assign n6004 = ~\u1_row_adr_reg[7]/P0001  & \u2_u0_b2_last_row_reg[7]/P0001  ;
  assign n6005 = ~n6003 & ~n6004 ;
  assign n6006 = ~\u1_row_adr_reg[3]/P0001  & \u2_u0_b2_last_row_reg[3]/P0001  ;
  assign n6007 = \u1_row_adr_reg[1]/P0001  & ~\u2_u0_b2_last_row_reg[1]/P0001  ;
  assign n6008 = ~n6006 & ~n6007 ;
  assign n6009 = n6005 & n6008 ;
  assign n6010 = n6002 & n6009 ;
  assign n6011 = n5995 & n6010 ;
  assign n6012 = n5981 & n6011 ;
  assign n6013 = \u1_row_adr_reg[3]/P0001  & ~\u2_u0_b1_last_row_reg[3]/P0001  ;
  assign n6014 = \u1_row_adr_reg[6]/P0001  & ~\u2_u0_b1_last_row_reg[6]/P0001  ;
  assign n6015 = ~\u1_row_adr_reg[12]/P0001  & \u2_u0_b1_last_row_reg[12]/P0001  ;
  assign n6016 = ~n6014 & ~n6015 ;
  assign n6017 = ~n6013 & n6016 ;
  assign n6018 = ~\u1_row_adr_reg[7]/P0001  & \u2_u0_b1_last_row_reg[7]/P0001  ;
  assign n6019 = \u1_row_adr_reg[1]/P0001  & ~\u2_u0_b1_last_row_reg[1]/P0001  ;
  assign n6020 = ~n6018 & ~n6019 ;
  assign n6021 = ~\u1_row_adr_reg[11]/P0001  & \u2_u0_b1_last_row_reg[11]/P0001  ;
  assign n6022 = \u1_row_adr_reg[11]/P0001  & ~\u2_u0_b1_last_row_reg[11]/P0001  ;
  assign n6023 = ~n6021 & ~n6022 ;
  assign n6024 = n6020 & n6023 ;
  assign n6025 = ~\u1_row_adr_reg[3]/P0001  & \u2_u0_b1_last_row_reg[3]/P0001  ;
  assign n6026 = \u1_row_adr_reg[8]/P0001  & ~\u2_u0_b1_last_row_reg[8]/P0001  ;
  assign n6027 = ~n6025 & ~n6026 ;
  assign n6028 = ~\u1_row_adr_reg[10]/P0001  & \u2_u0_b1_last_row_reg[10]/P0001  ;
  assign n6029 = ~\u1_row_adr_reg[0]/P0001  & \u2_u0_b1_last_row_reg[0]/P0001  ;
  assign n6030 = ~n6028 & ~n6029 ;
  assign n6031 = n6027 & n6030 ;
  assign n6032 = n6024 & n6031 ;
  assign n6033 = n6017 & n6032 ;
  assign n6034 = \u1_row_adr_reg[5]/P0001  & ~\u2_u0_b1_last_row_reg[5]/P0001  ;
  assign n6035 = ~\u1_row_adr_reg[9]/P0001  & \u2_u0_b1_last_row_reg[9]/P0001  ;
  assign n6036 = ~n6034 & ~n6035 ;
  assign n6037 = \u1_row_adr_reg[12]/P0001  & ~\u2_u0_b1_last_row_reg[12]/P0001  ;
  assign n6038 = ~\u1_row_adr_reg[6]/P0001  & \u2_u0_b1_last_row_reg[6]/P0001  ;
  assign n6039 = ~n6037 & ~n6038 ;
  assign n6040 = n6036 & n6039 ;
  assign n6041 = ~\u1_row_adr_reg[1]/P0001  & \u2_u0_b1_last_row_reg[1]/P0001  ;
  assign n6042 = n3684 & ~n6041 ;
  assign n6043 = \u1_row_adr_reg[9]/P0001  & ~\u2_u0_b1_last_row_reg[9]/P0001  ;
  assign n6044 = \u1_row_adr_reg[4]/P0001  & ~\u2_u0_b1_last_row_reg[4]/P0001  ;
  assign n6045 = ~n6043 & ~n6044 ;
  assign n6046 = n6042 & n6045 ;
  assign n6047 = n6040 & n6046 ;
  assign n6048 = \u1_row_adr_reg[10]/P0001  & ~\u2_u0_b1_last_row_reg[10]/P0001  ;
  assign n6049 = ~\u1_row_adr_reg[2]/P0001  & \u2_u0_b1_last_row_reg[2]/P0001  ;
  assign n6050 = ~n6048 & ~n6049 ;
  assign n6051 = ~\u1_row_adr_reg[8]/P0001  & \u2_u0_b1_last_row_reg[8]/P0001  ;
  assign n6052 = \u1_row_adr_reg[0]/P0001  & ~\u2_u0_b1_last_row_reg[0]/P0001  ;
  assign n6053 = ~n6051 & ~n6052 ;
  assign n6054 = n6050 & n6053 ;
  assign n6055 = \u1_row_adr_reg[7]/P0001  & ~\u2_u0_b1_last_row_reg[7]/P0001  ;
  assign n6056 = ~\u1_row_adr_reg[5]/P0001  & \u2_u0_b1_last_row_reg[5]/P0001  ;
  assign n6057 = ~n6055 & ~n6056 ;
  assign n6058 = ~\u1_row_adr_reg[4]/P0001  & \u2_u0_b1_last_row_reg[4]/P0001  ;
  assign n6059 = \u1_row_adr_reg[2]/P0001  & ~\u2_u0_b1_last_row_reg[2]/P0001  ;
  assign n6060 = ~n6058 & ~n6059 ;
  assign n6061 = n6057 & n6060 ;
  assign n6062 = n6054 & n6061 ;
  assign n6063 = n6047 & n6062 ;
  assign n6064 = n6033 & n6063 ;
  assign n6065 = ~n6012 & ~n6064 ;
  assign n6066 = ~\u1_row_adr_reg[12]/P0001  & \u2_u0_b0_last_row_reg[12]/P0001  ;
  assign n6067 = \u1_row_adr_reg[12]/P0001  & ~\u2_u0_b0_last_row_reg[12]/P0001  ;
  assign n6068 = \u1_row_adr_reg[5]/P0001  & ~\u2_u0_b0_last_row_reg[5]/P0001  ;
  assign n6069 = ~n6067 & ~n6068 ;
  assign n6070 = ~n6066 & n6069 ;
  assign n6071 = \u1_row_adr_reg[10]/P0001  & ~\u2_u0_b0_last_row_reg[10]/P0001  ;
  assign n6072 = \u1_row_adr_reg[11]/P0001  & ~\u2_u0_b0_last_row_reg[11]/P0001  ;
  assign n6073 = ~n6071 & ~n6072 ;
  assign n6074 = ~\u1_row_adr_reg[0]/P0001  & \u2_u0_b0_last_row_reg[0]/P0001  ;
  assign n6075 = ~\u1_row_adr_reg[6]/P0001  & \u2_u0_b0_last_row_reg[6]/P0001  ;
  assign n6076 = ~n6074 & ~n6075 ;
  assign n6077 = n6073 & n6076 ;
  assign n6078 = ~\u1_row_adr_reg[10]/P0001  & \u2_u0_b0_last_row_reg[10]/P0001  ;
  assign n6079 = \u1_row_adr_reg[6]/P0001  & ~\u2_u0_b0_last_row_reg[6]/P0001  ;
  assign n6080 = ~n6078 & ~n6079 ;
  assign n6081 = ~\u1_row_adr_reg[2]/P0001  & \u2_u0_b0_last_row_reg[2]/P0001  ;
  assign n6082 = ~\u1_row_adr_reg[9]/P0001  & \u2_u0_b0_last_row_reg[9]/P0001  ;
  assign n6083 = ~n6081 & ~n6082 ;
  assign n6084 = n6080 & n6083 ;
  assign n6085 = n6077 & n6084 ;
  assign n6086 = n6070 & n6085 ;
  assign n6087 = \u1_row_adr_reg[7]/P0001  & ~\u2_u0_b0_last_row_reg[7]/P0001  ;
  assign n6088 = \u1_row_adr_reg[1]/P0001  & ~\u2_u0_b0_last_row_reg[1]/P0001  ;
  assign n6089 = ~n6087 & ~n6088 ;
  assign n6090 = \u1_row_adr_reg[8]/P0001  & ~\u2_u0_b0_last_row_reg[8]/P0001  ;
  assign n6091 = ~\u1_row_adr_reg[11]/P0001  & \u2_u0_b0_last_row_reg[11]/P0001  ;
  assign n6092 = ~n6090 & ~n6091 ;
  assign n6093 = n6089 & n6092 ;
  assign n6094 = ~\u1_row_adr_reg[5]/P0001  & \u2_u0_b0_last_row_reg[5]/P0001  ;
  assign n6095 = n5855 & ~n6094 ;
  assign n6096 = ~\u1_row_adr_reg[8]/P0001  & \u2_u0_b0_last_row_reg[8]/P0001  ;
  assign n6097 = ~\u1_row_adr_reg[4]/P0001  & \u2_u0_b0_last_row_reg[4]/P0001  ;
  assign n6098 = ~n6096 & ~n6097 ;
  assign n6099 = n6095 & n6098 ;
  assign n6100 = n6093 & n6099 ;
  assign n6101 = ~\u1_row_adr_reg[3]/P0001  & \u2_u0_b0_last_row_reg[3]/P0001  ;
  assign n6102 = ~\u1_row_adr_reg[1]/P0001  & \u2_u0_b0_last_row_reg[1]/P0001  ;
  assign n6103 = ~n6101 & ~n6102 ;
  assign n6104 = \u1_row_adr_reg[0]/P0001  & ~\u2_u0_b0_last_row_reg[0]/P0001  ;
  assign n6105 = \u1_row_adr_reg[2]/P0001  & ~\u2_u0_b0_last_row_reg[2]/P0001  ;
  assign n6106 = ~n6104 & ~n6105 ;
  assign n6107 = n6103 & n6106 ;
  assign n6108 = \u1_row_adr_reg[3]/P0001  & ~\u2_u0_b0_last_row_reg[3]/P0001  ;
  assign n6109 = \u1_row_adr_reg[4]/P0001  & ~\u2_u0_b0_last_row_reg[4]/P0001  ;
  assign n6110 = ~n6108 & ~n6109 ;
  assign n6111 = \u1_row_adr_reg[9]/P0001  & ~\u2_u0_b0_last_row_reg[9]/P0001  ;
  assign n6112 = ~\u1_row_adr_reg[7]/P0001  & \u2_u0_b0_last_row_reg[7]/P0001  ;
  assign n6113 = ~n6111 & ~n6112 ;
  assign n6114 = n6110 & n6113 ;
  assign n6115 = n6107 & n6114 ;
  assign n6116 = n6100 & n6115 ;
  assign n6117 = n6086 & n6116 ;
  assign n6118 = ~\u1_row_adr_reg[0]/P0001  & \u2_u0_b3_last_row_reg[0]/P0001  ;
  assign n6119 = \u1_row_adr_reg[0]/P0001  & ~\u2_u0_b3_last_row_reg[0]/P0001  ;
  assign n6120 = \u1_row_adr_reg[11]/P0001  & ~\u2_u0_b3_last_row_reg[11]/P0001  ;
  assign n6121 = ~n6119 & ~n6120 ;
  assign n6122 = ~n6118 & n6121 ;
  assign n6123 = ~\u1_row_adr_reg[11]/P0001  & \u2_u0_b3_last_row_reg[11]/P0001  ;
  assign n6124 = \u1_row_adr_reg[7]/P0001  & ~\u2_u0_b3_last_row_reg[7]/P0001  ;
  assign n6125 = ~n6123 & ~n6124 ;
  assign n6126 = \u1_row_adr_reg[1]/P0001  & ~\u2_u0_b3_last_row_reg[1]/P0001  ;
  assign n6127 = ~\u1_row_adr_reg[12]/P0001  & \u2_u0_b3_last_row_reg[12]/P0001  ;
  assign n6128 = ~n6126 & ~n6127 ;
  assign n6129 = n6125 & n6128 ;
  assign n6130 = ~\u1_row_adr_reg[3]/P0001  & \u2_u0_b3_last_row_reg[3]/P0001  ;
  assign n6131 = \u1_row_adr_reg[10]/P0001  & ~\u2_u0_b3_last_row_reg[10]/P0001  ;
  assign n6132 = ~n6130 & ~n6131 ;
  assign n6133 = ~\u1_row_adr_reg[5]/P0001  & \u2_u0_b3_last_row_reg[5]/P0001  ;
  assign n6134 = ~\u1_row_adr_reg[9]/P0001  & \u2_u0_b3_last_row_reg[9]/P0001  ;
  assign n6135 = ~n6133 & ~n6134 ;
  assign n6136 = n6132 & n6135 ;
  assign n6137 = n6129 & n6136 ;
  assign n6138 = n6122 & n6137 ;
  assign n6139 = \u1_row_adr_reg[5]/P0001  & ~\u2_u0_b3_last_row_reg[5]/P0001  ;
  assign n6140 = ~\u1_row_adr_reg[10]/P0001  & \u2_u0_b3_last_row_reg[10]/P0001  ;
  assign n6141 = ~n6139 & ~n6140 ;
  assign n6142 = \u1_row_adr_reg[2]/P0001  & ~\u2_u0_b3_last_row_reg[2]/P0001  ;
  assign n6143 = ~\u1_row_adr_reg[8]/P0001  & \u2_u0_b3_last_row_reg[8]/P0001  ;
  assign n6144 = ~n6142 & ~n6143 ;
  assign n6145 = n6141 & n6144 ;
  assign n6146 = ~\u1_row_adr_reg[4]/P0001  & ~\u2_u0_b3_last_row_reg[4]/P0001  ;
  assign n6147 = \u1_row_adr_reg[4]/P0001  & \u2_u0_b3_last_row_reg[4]/P0001  ;
  assign n6148 = ~n6146 & ~n6147 ;
  assign n6149 = \u1_row_adr_reg[6]/P0001  & ~\u2_u0_b3_last_row_reg[6]/P0001  ;
  assign n6150 = n3793 & ~n6149 ;
  assign n6151 = ~n6148 & n6150 ;
  assign n6152 = n6145 & n6151 ;
  assign n6153 = \u1_row_adr_reg[3]/P0001  & ~\u2_u0_b3_last_row_reg[3]/P0001  ;
  assign n6154 = \u1_row_adr_reg[8]/P0001  & ~\u2_u0_b3_last_row_reg[8]/P0001  ;
  assign n6155 = ~n6153 & ~n6154 ;
  assign n6156 = ~\u1_row_adr_reg[2]/P0001  & \u2_u0_b3_last_row_reg[2]/P0001  ;
  assign n6157 = ~\u1_row_adr_reg[6]/P0001  & \u2_u0_b3_last_row_reg[6]/P0001  ;
  assign n6158 = ~n6156 & ~n6157 ;
  assign n6159 = n6155 & n6158 ;
  assign n6160 = ~\u1_row_adr_reg[7]/P0001  & \u2_u0_b3_last_row_reg[7]/P0001  ;
  assign n6161 = \u1_row_adr_reg[9]/P0001  & ~\u2_u0_b3_last_row_reg[9]/P0001  ;
  assign n6162 = ~n6160 & ~n6161 ;
  assign n6163 = ~\u1_row_adr_reg[1]/P0001  & \u2_u0_b3_last_row_reg[1]/P0001  ;
  assign n6164 = \u1_row_adr_reg[12]/P0001  & ~\u2_u0_b3_last_row_reg[12]/P0001  ;
  assign n6165 = ~n6163 & ~n6164 ;
  assign n6166 = n6162 & n6165 ;
  assign n6167 = n6159 & n6166 ;
  assign n6168 = n6152 & n6167 ;
  assign n6169 = n6138 & n6168 ;
  assign n6170 = ~n6117 & ~n6169 ;
  assign n6171 = n6065 & n6170 ;
  assign n6172 = n1840 & ~n6171 ;
  assign n6173 = ~n5960 & ~n6172 ;
  assign n6174 = n3398 & n3670 ;
  assign n6175 = ~n3372 & n6174 ;
  assign n6176 = ~n3381 & n6175 ;
  assign n6177 = n3678 & n6176 ;
  assign n6178 = \u5_cmd_asserted_reg/NET0131  & n1180 ;
  assign n6179 = \u5_susp_sel_r_reg/NET0131  & ~n6178 ;
  assign n6180 = n1924 & n1925 ;
  assign n6181 = n3858 & n6180 ;
  assign n6182 = n1308 & n6181 ;
  assign n6183 = ~n6179 & ~n6182 ;
  assign n6184 = \u0_u1_csc_reg[1]/NET0131  & n4259 ;
  assign n6185 = \u0_u0_csc_reg[1]/NET0131  & ~n4200 ;
  assign n6186 = n4214 & n6185 ;
  assign n6187 = n4199 & n6186 ;
  assign n6188 = ~n6184 & ~n6187 ;
  assign n6189 = \u0_u1_csc_reg[2]/NET0131  & n4259 ;
  assign n6190 = \u0_u0_csc_reg[2]/NET0131  & ~n4200 ;
  assign n6191 = n4214 & n6190 ;
  assign n6192 = n4199 & n6191 ;
  assign n6193 = ~n6189 & ~n6192 ;
  assign n6194 = \u0_u1_csc_reg[3]/NET0131  & n4259 ;
  assign n6195 = \u0_u0_csc_reg[3]/NET0131  & ~n4200 ;
  assign n6196 = n4214 & n6195 ;
  assign n6197 = n4199 & n6196 ;
  assign n6198 = ~n6194 & ~n6197 ;
  assign n6199 = ~\u4_ps_cnt_reg[3]/NET0131  & ~n5611 ;
  assign n6200 = ~n5614 & ~n6199 ;
  assign n6201 = ~n5608 & n6200 ;
  assign n6202 = ~\wb_addr_i[15]_pad  & ~n1546 ;
  assign n6203 = ~\u1_sram_addr_reg[13]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6204 = n1537 & n6203 ;
  assign n6205 = n1544 & n6204 ;
  assign n6206 = ~n1532 & ~n6205 ;
  assign n6207 = ~n6202 & n6206 ;
  assign n6208 = \u1_bank_adr_reg[0]/P0001  & n1537 ;
  assign n6209 = n1532 & n6208 ;
  assign n6210 = \u1_acs_addr_reg[13]/P0001  & ~n1537 ;
  assign n6211 = n1532 & n6210 ;
  assign n6212 = ~n6209 & ~n6211 ;
  assign n6213 = ~n6207 & n6212 ;
  assign n6214 = ~\wb_addr_i[16]_pad  & ~n1546 ;
  assign n6215 = ~\u1_sram_addr_reg[14]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6216 = n1537 & n6215 ;
  assign n6217 = n1544 & n6216 ;
  assign n6218 = ~n1532 & ~n6217 ;
  assign n6219 = ~n6214 & n6218 ;
  assign n6220 = \u1_bank_adr_reg[1]/P0001  & n1537 ;
  assign n6221 = n1532 & n6220 ;
  assign n6222 = \u1_acs_addr_reg[14]/P0001  & ~n1537 ;
  assign n6223 = n1532 & n6222 ;
  assign n6224 = ~n6221 & ~n6223 ;
  assign n6225 = ~n6219 & n6224 ;
  assign n6226 = \u1_col_adr_reg[9]/P0001  & n5550 ;
  assign n6227 = n4912 & ~n5550 ;
  assign n6228 = ~n5115 & n6227 ;
  assign n6229 = ~n6226 & ~n6228 ;
  assign n6230 = n5695 & ~n5696 ;
  assign n6231 = \u1_acs_addr_reg[16]/P0001  & ~n1537 ;
  assign n6232 = n1532 & n6231 ;
  assign n6233 = ~\wb_addr_i[18]_pad  & ~n1546 ;
  assign n6234 = ~\u1_sram_addr_reg[16]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6235 = n1537 & n6234 ;
  assign n6236 = n1544 & n6235 ;
  assign n6237 = ~n1532 & ~n6236 ;
  assign n6238 = ~n6233 & n6237 ;
  assign n6239 = ~n6232 & ~n6238 ;
  assign n6240 = \u1_acs_addr_reg[17]/P0001  & ~n1537 ;
  assign n6241 = n1532 & n6240 ;
  assign n6242 = ~\wb_addr_i[19]_pad  & ~n1546 ;
  assign n6243 = ~\u1_sram_addr_reg[17]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6244 = n1537 & n6243 ;
  assign n6245 = n1544 & n6244 ;
  assign n6246 = ~n1532 & ~n6245 ;
  assign n6247 = ~n6242 & n6246 ;
  assign n6248 = ~n6241 & ~n6247 ;
  assign n6249 = \u1_acs_addr_reg[18]/P0001  & ~n1537 ;
  assign n6250 = n1532 & n6249 ;
  assign n6251 = ~\wb_addr_i[20]_pad  & ~n1546 ;
  assign n6252 = ~\u1_sram_addr_reg[18]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6253 = n1537 & n6252 ;
  assign n6254 = n1544 & n6253 ;
  assign n6255 = ~n1532 & ~n6254 ;
  assign n6256 = ~n6251 & n6255 ;
  assign n6257 = ~n6250 & ~n6256 ;
  assign n6258 = \u1_acs_addr_reg[19]/P0001  & ~n1537 ;
  assign n6259 = n1532 & n6258 ;
  assign n6260 = ~\wb_addr_i[21]_pad  & ~n1546 ;
  assign n6261 = ~\u1_sram_addr_reg[19]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6262 = n1537 & n6261 ;
  assign n6263 = n1544 & n6262 ;
  assign n6264 = ~n1532 & ~n6263 ;
  assign n6265 = ~n6260 & n6264 ;
  assign n6266 = ~n6259 & ~n6265 ;
  assign n6267 = \u1_acs_addr_reg[21]/P0001  & ~n1537 ;
  assign n6268 = n1532 & n6267 ;
  assign n6269 = ~\wb_addr_i[23]_pad  & ~n1546 ;
  assign n6270 = ~\u1_sram_addr_reg[21]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6271 = n1537 & n6270 ;
  assign n6272 = n1544 & n6271 ;
  assign n6273 = ~n1532 & ~n6272 ;
  assign n6274 = ~n6269 & n6273 ;
  assign n6275 = ~n6268 & ~n6274 ;
  assign n6276 = \u1_acs_addr_reg[22]/P0001  & ~n1537 ;
  assign n6277 = n1532 & n6276 ;
  assign n6278 = ~\wb_addr_i[24]_pad  & ~n1546 ;
  assign n6279 = ~\u1_sram_addr_reg[22]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6280 = n1537 & n6279 ;
  assign n6281 = n1544 & n6280 ;
  assign n6282 = ~n1532 & ~n6281 ;
  assign n6283 = ~n6278 & n6282 ;
  assign n6284 = ~n6277 & ~n6283 ;
  assign n6285 = \u1_acs_addr_reg[23]/P0001  & ~n1537 ;
  assign n6286 = n1532 & n6285 ;
  assign n6287 = ~\wb_addr_i[25]_pad  & ~n1546 ;
  assign n6288 = ~\u1_sram_addr_reg[23]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6289 = n1537 & n6288 ;
  assign n6290 = n1544 & n6289 ;
  assign n6291 = ~n1532 & ~n6290 ;
  assign n6292 = ~n6287 & n6291 ;
  assign n6293 = ~n6286 & ~n6292 ;
  assign n6294 = \u1_acs_addr_reg[15]/P0001  & ~n1537 ;
  assign n6295 = n1532 & n6294 ;
  assign n6296 = ~\wb_addr_i[17]_pad  & ~n1546 ;
  assign n6297 = ~\u1_sram_addr_reg[15]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6298 = n1537 & n6297 ;
  assign n6299 = n1544 & n6298 ;
  assign n6300 = ~n1532 & ~n6299 ;
  assign n6301 = ~n6296 & n6300 ;
  assign n6302 = ~n6295 & ~n6301 ;
  assign n6303 = \u1_acs_addr_reg[20]/P0001  & ~n1537 ;
  assign n6304 = n1532 & n6303 ;
  assign n6305 = ~\wb_addr_i[22]_pad  & ~n1546 ;
  assign n6306 = ~\u1_sram_addr_reg[20]/P0001  & \u6_wr_hold_reg/NET0131  ;
  assign n6307 = n1537 & n6306 ;
  assign n6308 = n1544 & n6307 ;
  assign n6309 = ~n1532 & ~n6308 ;
  assign n6310 = ~n6305 & n6309 ;
  assign n6311 = ~n6304 & ~n6310 ;
  assign n6312 = \u1_acs_addr_reg[7]/P0001  & \u1_acs_addr_reg[8]/P0001  ;
  assign n6313 = n5146 & n6312 ;
  assign n6314 = ~\u1_acs_addr_reg[8]/P0001  & ~n5557 ;
  assign n6315 = ~n6313 & ~n6314 ;
  assign n6316 = \u4_ps_cnt_reg[1]/NET0131  & n5609 ;
  assign n6317 = ~\u4_ps_cnt_reg[2]/NET0131  & ~n6316 ;
  assign n6318 = ~n5611 & ~n6317 ;
  assign n6319 = ~n5608 & n6318 ;
  assign n6320 = ~\u4_ps_cnt_reg[5]/NET0131  & ~n5613 ;
  assign n6321 = ~n5720 & ~n6320 ;
  assign n6322 = ~n5608 & n6321 ;
  assign n6323 = ~\u4_ps_cnt_reg[6]/NET0131  & ~n5720 ;
  assign n6324 = ~n5721 & ~n6323 ;
  assign n6325 = ~n5608 & n6324 ;
  assign n6326 = ~\u4_ps_cnt_reg[0]/NET0131  & ~\u4_rfr_en_reg/NET0131  ;
  assign n6327 = ~n5609 & ~n6326 ;
  assign n6328 = ~n5608 & n6327 ;
  assign n6329 = ~\u4_ps_cnt_reg[1]/NET0131  & ~n5609 ;
  assign n6330 = ~n6316 & ~n6329 ;
  assign n6331 = ~n5608 & n6330 ;
  assign n6332 = \u0_init_req_reg/NET0131  & ~\u4_rfr_req_reg/NET0131  ;
  assign n6333 = n1309 & n6332 ;
  assign n6334 = n1308 & n6333 ;
  assign n6335 = \u1_acs_addr_reg[4]/P0001  & n5143 ;
  assign n6336 = ~\u1_acs_addr_reg[4]/P0001  & ~n5143 ;
  assign n6337 = ~n6335 & ~n6336 ;
  assign n6338 = \mem_ack_r_reg/P0001  & \u6_read_go_r1_reg/NET0131  ;
  assign n6339 = n1234 & n6338 ;
  assign n6340 = ~n1048 & n6339 ;
  assign n6341 = ~\u3_u0_rd_adr_reg[0]/NET0131  & n5380 ;
  assign n6342 = ~n6340 & n6341 ;
  assign n6343 = ~\u3_u0_rd_adr_reg[3]/NET0131  & n5380 ;
  assign n6344 = n6340 & n6343 ;
  assign n6345 = ~n6342 & ~n6344 ;
  assign n6346 = \u3_u0_rd_adr_reg[1]/NET0131  & n5380 ;
  assign n6347 = ~n6340 & n6346 ;
  assign n6348 = \u3_u0_rd_adr_reg[0]/NET0131  & n5380 ;
  assign n6349 = n6340 & n6348 ;
  assign n6350 = ~n6347 & ~n6349 ;
  assign n6351 = \u3_u0_rd_adr_reg[2]/NET0131  & n5380 ;
  assign n6352 = ~n6340 & n6351 ;
  assign n6353 = n6340 & n6346 ;
  assign n6354 = ~n6352 & ~n6353 ;
  assign n6355 = \u3_u0_rd_adr_reg[3]/NET0131  & n5380 ;
  assign n6356 = ~n6340 & n6355 ;
  assign n6357 = n6340 & n6351 ;
  assign n6358 = ~n6356 & ~n6357 ;
  assign n6359 = \u2_u0_bank2_open_reg/NET0131  & n3751 ;
  assign n6360 = \u2_u0_bank1_open_reg/NET0131  & n3684 ;
  assign n6361 = ~n6359 & ~n6360 ;
  assign n6362 = \u2_u0_bank3_open_reg/NET0131  & n3793 ;
  assign n6363 = \u2_u0_bank0_open_reg/NET0131  & n5855 ;
  assign n6364 = ~n6362 & ~n6363 ;
  assign n6365 = n6361 & n6364 ;
  assign n6366 = ~n1839 & ~n6365 ;
  assign n6367 = n1835 & n6366 ;
  assign n6368 = \u2_u1_bank2_open_reg/NET0131  & n3751 ;
  assign n6369 = \u2_u1_bank3_open_reg/NET0131  & n3793 ;
  assign n6370 = ~n6368 & ~n6369 ;
  assign n6371 = \u2_u1_bank0_open_reg/NET0131  & n5855 ;
  assign n6372 = \u2_u1_bank1_open_reg/NET0131  & n3684 ;
  assign n6373 = ~n6371 & ~n6372 ;
  assign n6374 = n6370 & n6373 ;
  assign n6375 = ~n1919 & ~n6374 ;
  assign n6376 = ~n6367 & ~n6375 ;
  assign n6377 = ~\u0_u0_addr_r_reg[5]/P0001  & ~\u0_u0_addr_r_reg[6]/P0001  ;
  assign n6378 = ~\u0_u0_addr_r_reg[3]/P0001  & n6377 ;
  assign n6379 = \u0_rf_we_reg/NET0131  & \u0_u0_addr_r_reg[4]/P0001  ;
  assign n6380 = ~\u0_u0_addr_r_reg[2]/P0001  & n6379 ;
  assign n6381 = n6378 & n6380 ;
  assign n6382 = ~\u0_u0_csc_reg[0]/NET0131  & ~n6381 ;
  assign n6383 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[0]_pad  ;
  assign n6384 = n6379 & n6383 ;
  assign n6385 = n6378 & n6384 ;
  assign n6386 = ~\u0_rst_r2_reg/NET0131  & ~n6385 ;
  assign n6387 = ~n6382 & n6386 ;
  assign n6388 = \poc_o[3]_pad  & \u0_rst_r2_reg/NET0131  ;
  assign n6389 = \poc_o[2]_pad  & \u0_rst_r2_reg/NET0131  ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = ~n6387 & n6390 ;
  assign n6392 = ~\u0_csc_reg[2]/NET0131  & ~\u0_csc_reg[3]/NET0131  ;
  assign n6393 = ~n2375 & n6392 ;
  assign n6394 = n2191 & n6392 ;
  assign n6395 = \u7_mc_data_ir_reg[2]/P0001  & n5304 ;
  assign n6396 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[26]/P0001  ;
  assign n6397 = ~n6395 & ~n6396 ;
  assign n6398 = \u7_mc_data_ir_reg[10]/P0001  & n5309 ;
  assign n6399 = n2191 & ~n6398 ;
  assign n6400 = n6397 & n6399 ;
  assign n6401 = ~n6394 & ~n6400 ;
  assign n6402 = ~n6393 & ~n6401 ;
  assign n6403 = ~\wb_addr_i[5]_pad  & ~\wb_addr_i[6]_pad  ;
  assign n6404 = ~\wb_addr_i[3]_pad  & n6403 ;
  assign n6405 = ~\wb_addr_i[2]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6406 = \u0_csr_r2_reg[2]/NET0131  & n6405 ;
  assign n6407 = n6404 & n6406 ;
  assign n6408 = ~\wb_addr_i[2]_pad  & \wb_addr_i[4]_pad  ;
  assign n6409 = \u0_u0_csc_reg[26]/P0001  & n6408 ;
  assign n6410 = n6404 & n6409 ;
  assign n6411 = \wb_addr_i[3]_pad  & n6403 ;
  assign n6412 = \wb_addr_i[2]_pad  & \wb_addr_i[4]_pad  ;
  assign n6413 = \u0_u1_tms_reg[26]/P0001  & n6412 ;
  assign n6414 = n6411 & n6413 ;
  assign n6415 = ~n6410 & ~n6414 ;
  assign n6416 = ~n6407 & n6415 ;
  assign n6417 = \u0_u1_csc_reg[26]/P0001  & n6408 ;
  assign n6418 = n6411 & n6417 ;
  assign n6419 = ~n2191 & ~n6418 ;
  assign n6420 = \wb_addr_i[2]_pad  & ~\wb_addr_i[3]_pad  ;
  assign n6421 = n6403 & n6420 ;
  assign n6422 = \u0_u0_tms_reg[26]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6423 = n6421 & n6422 ;
  assign n6424 = \poc_o[26]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6425 = n6421 & n6424 ;
  assign n6426 = ~n6423 & ~n6425 ;
  assign n6427 = n6419 & n6426 ;
  assign n6428 = n6416 & n6427 ;
  assign n6429 = ~n6402 & ~n6428 ;
  assign n6430 = \u7_mc_data_ir_reg[11]/P0001  & n5309 ;
  assign n6431 = \u7_mc_data_ir_reg[3]/P0001  & n5304 ;
  assign n6432 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[27]/P0001  ;
  assign n6433 = ~n6392 & ~n6432 ;
  assign n6434 = ~n6431 & n6433 ;
  assign n6435 = ~n6430 & n6434 ;
  assign n6436 = n2191 & n6435 ;
  assign n6437 = n2321 & n6394 ;
  assign n6438 = ~n6436 & ~n6437 ;
  assign n6439 = \u0_u1_csc_reg[27]/P0001  & n6408 ;
  assign n6440 = n6411 & n6439 ;
  assign n6441 = \u0_u0_csc_reg[27]/P0001  & n6408 ;
  assign n6442 = n6404 & n6441 ;
  assign n6443 = \u0_u1_tms_reg[27]/P0001  & n6412 ;
  assign n6444 = n6411 & n6443 ;
  assign n6445 = ~n6442 & ~n6444 ;
  assign n6446 = ~n6440 & n6445 ;
  assign n6447 = \u0_csr_r2_reg[3]/NET0131  & n6405 ;
  assign n6448 = n6404 & n6447 ;
  assign n6449 = ~n2191 & ~n6448 ;
  assign n6450 = \u0_u0_tms_reg[27]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6451 = n6421 & n6450 ;
  assign n6452 = \poc_o[27]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6453 = n6421 & n6452 ;
  assign n6454 = ~n6451 & ~n6453 ;
  assign n6455 = n6449 & n6454 ;
  assign n6456 = n6446 & n6455 ;
  assign n6457 = n6438 & ~n6456 ;
  assign n6458 = \u7_mc_data_ir_reg[12]/P0001  & n5309 ;
  assign n6459 = \u7_mc_data_ir_reg[4]/P0001  & n5304 ;
  assign n6460 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[28]/P0001  ;
  assign n6461 = ~n6392 & ~n6460 ;
  assign n6462 = ~n6459 & n6461 ;
  assign n6463 = ~n6458 & n6462 ;
  assign n6464 = n2191 & n6463 ;
  assign n6465 = n2335 & n6394 ;
  assign n6466 = ~n6464 & ~n6465 ;
  assign n6467 = \u0_u1_csc_reg[28]/P0001  & n6408 ;
  assign n6468 = n6411 & n6467 ;
  assign n6469 = \u0_u0_csc_reg[28]/P0001  & n6408 ;
  assign n6470 = n6404 & n6469 ;
  assign n6471 = \u0_u1_tms_reg[28]/P0001  & n6412 ;
  assign n6472 = n6411 & n6471 ;
  assign n6473 = ~n6470 & ~n6472 ;
  assign n6474 = ~n6468 & n6473 ;
  assign n6475 = \u0_csr_r2_reg[4]/NET0131  & n6405 ;
  assign n6476 = n6404 & n6475 ;
  assign n6477 = ~n2191 & ~n6476 ;
  assign n6478 = \u0_u0_tms_reg[28]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6479 = n6421 & n6478 ;
  assign n6480 = \poc_o[28]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6481 = n6421 & n6480 ;
  assign n6482 = ~n6479 & ~n6481 ;
  assign n6483 = n6477 & n6482 ;
  assign n6484 = n6474 & n6483 ;
  assign n6485 = n6466 & ~n6484 ;
  assign n6486 = \u7_mc_data_ir_reg[13]/P0001  & n5309 ;
  assign n6487 = \u7_mc_data_ir_reg[5]/P0001  & n5304 ;
  assign n6488 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[29]/P0001  ;
  assign n6489 = ~n6392 & ~n6488 ;
  assign n6490 = ~n6487 & n6489 ;
  assign n6491 = ~n6486 & n6490 ;
  assign n6492 = n2191 & n6491 ;
  assign n6493 = n2311 & n6394 ;
  assign n6494 = ~n6492 & ~n6493 ;
  assign n6495 = \u0_u1_csc_reg[29]/P0001  & n6408 ;
  assign n6496 = n6411 & n6495 ;
  assign n6497 = \u0_u0_csc_reg[29]/P0001  & n6408 ;
  assign n6498 = n6404 & n6497 ;
  assign n6499 = \u0_u1_tms_reg[29]/P0001  & n6412 ;
  assign n6500 = n6411 & n6499 ;
  assign n6501 = ~n6498 & ~n6500 ;
  assign n6502 = ~n6496 & n6501 ;
  assign n6503 = \u0_csr_r2_reg[5]/NET0131  & n6405 ;
  assign n6504 = n6404 & n6503 ;
  assign n6505 = ~n2191 & ~n6504 ;
  assign n6506 = \u0_u0_tms_reg[29]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6507 = n6421 & n6506 ;
  assign n6508 = \poc_o[29]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6509 = n6421 & n6508 ;
  assign n6510 = ~n6507 & ~n6509 ;
  assign n6511 = n6505 & n6510 ;
  assign n6512 = n6502 & n6511 ;
  assign n6513 = n6494 & ~n6512 ;
  assign n6514 = \u7_mc_data_ir_reg[15]/P0001  & n5309 ;
  assign n6515 = \u7_mc_data_ir_reg[7]/P0001  & n5304 ;
  assign n6516 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[31]/P0001  ;
  assign n6517 = ~n6392 & ~n6516 ;
  assign n6518 = ~n6515 & n6517 ;
  assign n6519 = ~n6514 & n6518 ;
  assign n6520 = n2191 & n6519 ;
  assign n6521 = n2358 & n6394 ;
  assign n6522 = ~n6520 & ~n6521 ;
  assign n6523 = \u0_u1_csc_reg[31]/P0001  & n6408 ;
  assign n6524 = n6411 & n6523 ;
  assign n6525 = \u0_u1_tms_reg[31]/P0001  & n6412 ;
  assign n6526 = n6411 & n6525 ;
  assign n6527 = \u0_csr_r2_reg[7]/NET0131  & n6405 ;
  assign n6528 = n6404 & n6527 ;
  assign n6529 = ~n6526 & ~n6528 ;
  assign n6530 = ~n6524 & n6529 ;
  assign n6531 = \u0_u0_csc_reg[31]/P0001  & n6408 ;
  assign n6532 = n6404 & n6531 ;
  assign n6533 = ~n2191 & ~n6532 ;
  assign n6534 = \u0_u0_tms_reg[31]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6535 = n6421 & n6534 ;
  assign n6536 = \poc_o[31]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6537 = n6421 & n6536 ;
  assign n6538 = ~n6535 & ~n6537 ;
  assign n6539 = n6533 & n6538 ;
  assign n6540 = n6530 & n6539 ;
  assign n6541 = n6522 & ~n6540 ;
  assign n6542 = ~\u0_u0_csc_reg[3]/NET0131  & \u0_u0_lmr_req_we_reg/NET0131  ;
  assign n6543 = n1836 & n6542 ;
  assign n6544 = \u0_u0_inited_reg/NET0131  & n6543 ;
  assign n6545 = \u0_lmr_ack_r_reg/P0001  & ~\u5_lmr_ack_reg/NET0131  ;
  assign n6546 = \u0_spec_req_cs_reg[0]/NET0131  & n6545 ;
  assign n6547 = \u0_u0_lmr_req_reg/NET0131  & ~n6546 ;
  assign n6548 = ~n6543 & n6547 ;
  assign n6549 = ~n6544 & ~n6548 ;
  assign n6550 = ~\u0_u1_csc_reg[3]/NET0131  & \u0_u1_lmr_req_we_reg/NET0131  ;
  assign n6551 = n1915 & n6550 ;
  assign n6552 = \u0_u1_inited_reg/NET0131  & n6551 ;
  assign n6553 = \u0_spec_req_cs_reg[1]/NET0131  & n6545 ;
  assign n6554 = \u0_u1_lmr_req_reg/NET0131  & ~n6553 ;
  assign n6555 = ~n6551 & n6554 ;
  assign n6556 = ~n6552 & ~n6555 ;
  assign n6557 = \u7_mc_data_ir_reg[14]/P0001  & n5309 ;
  assign n6558 = \u7_mc_data_ir_reg[6]/P0001  & n5304 ;
  assign n6559 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[30]/P0001  ;
  assign n6560 = ~n6392 & ~n6559 ;
  assign n6561 = ~n6558 & n6560 ;
  assign n6562 = ~n6557 & n6561 ;
  assign n6563 = n2191 & n6562 ;
  assign n6564 = n2304 & n6394 ;
  assign n6565 = ~n6563 & ~n6564 ;
  assign n6566 = \u0_u1_csc_reg[30]/P0001  & n6408 ;
  assign n6567 = n6411 & n6566 ;
  assign n6568 = \u0_u0_csc_reg[30]/P0001  & n6408 ;
  assign n6569 = n6404 & n6568 ;
  assign n6570 = \u0_u1_tms_reg[30]/P0001  & n6412 ;
  assign n6571 = n6411 & n6570 ;
  assign n6572 = ~n6569 & ~n6571 ;
  assign n6573 = ~n6567 & n6572 ;
  assign n6574 = \u0_csr_r2_reg[6]/NET0131  & n6405 ;
  assign n6575 = n6404 & n6574 ;
  assign n6576 = ~n2191 & ~n6575 ;
  assign n6577 = \u0_u0_tms_reg[30]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6578 = n6421 & n6577 ;
  assign n6579 = \poc_o[30]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6580 = n6421 & n6579 ;
  assign n6581 = ~n6578 & ~n6580 ;
  assign n6582 = n6576 & n6581 ;
  assign n6583 = n6573 & n6582 ;
  assign n6584 = n6565 & ~n6583 ;
  assign n6585 = \u7_mc_data_ir_reg[0]/P0001  & n5304 ;
  assign n6586 = \u7_mc_data_ir_reg[8]/P0001  & n5309 ;
  assign n6587 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[24]/P0001  ;
  assign n6588 = ~n6392 & ~n6587 ;
  assign n6589 = ~n6586 & n6588 ;
  assign n6590 = ~n6585 & n6589 ;
  assign n6591 = n2191 & n6590 ;
  assign n6592 = n2351 & n6394 ;
  assign n6593 = ~n6591 & ~n6592 ;
  assign n6594 = \u0_u1_csc_reg[24]/P0001  & n6408 ;
  assign n6595 = n6411 & n6594 ;
  assign n6596 = \u0_u0_csc_reg[24]/P0001  & n6408 ;
  assign n6597 = n6404 & n6596 ;
  assign n6598 = \u0_u1_tms_reg[24]/P0001  & n6412 ;
  assign n6599 = n6411 & n6598 ;
  assign n6600 = ~n6597 & ~n6599 ;
  assign n6601 = ~n6595 & n6600 ;
  assign n6602 = \u0_csr_r2_reg[0]/NET0131  & n6405 ;
  assign n6603 = n6404 & n6602 ;
  assign n6604 = ~n2191 & ~n6603 ;
  assign n6605 = \u0_u0_tms_reg[24]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6606 = n6421 & n6605 ;
  assign n6607 = \poc_o[24]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6608 = n6421 & n6607 ;
  assign n6609 = ~n6606 & ~n6608 ;
  assign n6610 = n6604 & n6609 ;
  assign n6611 = n6601 & n6610 ;
  assign n6612 = n6593 & ~n6611 ;
  assign n6613 = \u7_mc_data_ir_reg[1]/P0001  & n5304 ;
  assign n6614 = \u7_mc_data_ir_reg[9]/P0001  & n5309 ;
  assign n6615 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[25]/P0001  ;
  assign n6616 = ~n6392 & ~n6615 ;
  assign n6617 = ~n6614 & n6616 ;
  assign n6618 = ~n6613 & n6617 ;
  assign n6619 = n2191 & n6618 ;
  assign n6620 = n2328 & n6394 ;
  assign n6621 = ~n6619 & ~n6620 ;
  assign n6622 = \u0_u1_csc_reg[25]/P0001  & n6408 ;
  assign n6623 = n6411 & n6622 ;
  assign n6624 = \u0_u0_csc_reg[25]/P0001  & n6408 ;
  assign n6625 = n6404 & n6624 ;
  assign n6626 = \u0_u1_tms_reg[25]/P0001  & n6412 ;
  assign n6627 = n6411 & n6626 ;
  assign n6628 = ~n6625 & ~n6627 ;
  assign n6629 = ~n6623 & n6628 ;
  assign n6630 = \u0_csr_r2_reg[1]/NET0131  & n6405 ;
  assign n6631 = n6404 & n6630 ;
  assign n6632 = ~n2191 & ~n6631 ;
  assign n6633 = \u0_u0_tms_reg[25]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6634 = n6421 & n6633 ;
  assign n6635 = \poc_o[25]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6636 = n6421 & n6635 ;
  assign n6637 = ~n6634 & ~n6636 ;
  assign n6638 = n6632 & n6637 ;
  assign n6639 = n6629 & n6638 ;
  assign n6640 = n6621 & ~n6639 ;
  assign n6641 = ~n2562 & n6392 ;
  assign n6642 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[1]/P0001  ;
  assign n6643 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[1]/P0001  ;
  assign n6644 = ~n6642 & ~n6643 ;
  assign n6645 = ~n6392 & ~n6644 ;
  assign n6646 = n2191 & ~n6645 ;
  assign n6647 = ~n6641 & n6646 ;
  assign n6648 = \u0_u1_csc_reg[1]/NET0131  & n6408 ;
  assign n6649 = n6411 & n6648 ;
  assign n6650 = \u0_csc_mask_r_reg[1]/NET0131  & n6405 ;
  assign n6651 = n6411 & n6650 ;
  assign n6652 = ~n6649 & ~n6651 ;
  assign n6653 = \u0_u1_tms_reg[1]/P0001  & n6412 ;
  assign n6654 = n6411 & n6653 ;
  assign n6655 = mc_vpen_pad_o_pad & n6405 ;
  assign n6656 = n6404 & n6655 ;
  assign n6657 = ~n6654 & ~n6656 ;
  assign n6658 = n6652 & n6657 ;
  assign n6659 = \u0_u0_csc_reg[1]/NET0131  & n6408 ;
  assign n6660 = n6404 & n6659 ;
  assign n6661 = ~n2191 & ~n6660 ;
  assign n6662 = \poc_o[1]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6663 = n6421 & n6662 ;
  assign n6664 = \u0_u0_tms_reg[1]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6665 = n6421 & n6664 ;
  assign n6666 = ~n6663 & ~n6665 ;
  assign n6667 = n6661 & n6666 ;
  assign n6668 = n6658 & n6667 ;
  assign n6669 = ~n6647 & ~n6668 ;
  assign n6670 = ~n2545 & n6392 ;
  assign n6671 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[3]/P0001  ;
  assign n6672 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[3]/P0001  ;
  assign n6673 = ~n6671 & ~n6672 ;
  assign n6674 = ~n6392 & ~n6673 ;
  assign n6675 = n2191 & ~n6674 ;
  assign n6676 = ~n6670 & n6675 ;
  assign n6677 = \u0_csc_mask_r_reg[3]/NET0131  & n6405 ;
  assign n6678 = n6411 & n6677 ;
  assign n6679 = \u0_u0_csc_reg[3]/NET0131  & n6408 ;
  assign n6680 = n6404 & n6679 ;
  assign n6681 = ~n6678 & ~n6680 ;
  assign n6682 = \u0_u1_tms_reg[3]/P0001  & n6412 ;
  assign n6683 = n6411 & n6682 ;
  assign n6684 = \u0_csr_r_reg[3]/NET0131  & n6405 ;
  assign n6685 = n6404 & n6684 ;
  assign n6686 = ~n6683 & ~n6685 ;
  assign n6687 = n6681 & n6686 ;
  assign n6688 = \u0_u1_csc_reg[3]/NET0131  & n6408 ;
  assign n6689 = n6411 & n6688 ;
  assign n6690 = ~n2191 & ~n6689 ;
  assign n6691 = \poc_o[3]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6692 = n6421 & n6691 ;
  assign n6693 = \u0_u0_tms_reg[3]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6694 = n6421 & n6693 ;
  assign n6695 = ~n6692 & ~n6694 ;
  assign n6696 = n6690 & n6695 ;
  assign n6697 = n6687 & n6696 ;
  assign n6698 = ~n6676 & ~n6697 ;
  assign n6699 = ~n2538 & n6392 ;
  assign n6700 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[5]/P0001  ;
  assign n6701 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[5]/P0001  ;
  assign n6702 = ~n6700 & ~n6701 ;
  assign n6703 = ~n6392 & ~n6702 ;
  assign n6704 = n2191 & ~n6703 ;
  assign n6705 = ~n6699 & n6704 ;
  assign n6706 = \u0_csc_mask_r_reg[5]/NET0131  & n6405 ;
  assign n6707 = n6411 & n6706 ;
  assign n6708 = \u0_u1_tms_reg[5]/P0001  & n6412 ;
  assign n6709 = n6411 & n6708 ;
  assign n6710 = ~n6707 & ~n6709 ;
  assign n6711 = \u0_u1_csc_reg[5]/P0001  & n6408 ;
  assign n6712 = n6411 & n6711 ;
  assign n6713 = \u0_csr_r_reg[5]/NET0131  & n6405 ;
  assign n6714 = n6404 & n6713 ;
  assign n6715 = ~n6712 & ~n6714 ;
  assign n6716 = n6710 & n6715 ;
  assign n6717 = \u0_u0_csc_reg[5]/P0001  & n6408 ;
  assign n6718 = n6404 & n6717 ;
  assign n6719 = ~n2191 & ~n6718 ;
  assign n6720 = \u0_u0_tms_reg[5]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6721 = n6421 & n6720 ;
  assign n6722 = \poc_o[5]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6723 = n6421 & n6722 ;
  assign n6724 = ~n6721 & ~n6723 ;
  assign n6725 = n6719 & n6724 ;
  assign n6726 = n6716 & n6725 ;
  assign n6727 = ~n6705 & ~n6726 ;
  assign n6728 = ~n2218 & n6392 ;
  assign n6729 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[1]/P0001  ;
  assign n6730 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[9]/P0001  ;
  assign n6731 = ~n6729 & ~n6730 ;
  assign n6732 = ~n6392 & ~n6731 ;
  assign n6733 = n2191 & ~n6732 ;
  assign n6734 = ~n6728 & n6733 ;
  assign n6735 = \u0_u1_csc_reg[9]/P0001  & n6408 ;
  assign n6736 = n6411 & n6735 ;
  assign n6737 = \u0_u1_tms_reg[9]/P0001  & n6412 ;
  assign n6738 = n6411 & n6737 ;
  assign n6739 = ~n6736 & ~n6738 ;
  assign n6740 = \u0_u0_csc_reg[9]/P0001  & n6408 ;
  assign n6741 = n6404 & n6740 ;
  assign n6742 = \u0_csc_mask_r_reg[9]/NET0131  & n6405 ;
  assign n6743 = n6411 & n6742 ;
  assign n6744 = ~n6741 & ~n6743 ;
  assign n6745 = n6739 & n6744 ;
  assign n6746 = \u0_csr_r_reg[9]/NET0131  & n6405 ;
  assign n6747 = n6404 & n6746 ;
  assign n6748 = ~n2191 & ~n6747 ;
  assign n6749 = \u0_u0_tms_reg[9]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6750 = n6421 & n6749 ;
  assign n6751 = \poc_o[9]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6752 = n6421 & n6751 ;
  assign n6753 = ~n6750 & ~n6752 ;
  assign n6754 = n6748 & n6753 ;
  assign n6755 = n6745 & n6754 ;
  assign n6756 = ~n6734 & ~n6755 ;
  assign n6757 = ~n2522 & n6392 ;
  assign n6758 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[6]/P0001  ;
  assign n6759 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[6]/P0001  ;
  assign n6760 = ~n6758 & ~n6759 ;
  assign n6761 = ~n6392 & ~n6760 ;
  assign n6762 = n2191 & ~n6761 ;
  assign n6763 = ~n6757 & n6762 ;
  assign n6764 = \u0_u0_csc_reg[6]/P0001  & n6408 ;
  assign n6765 = n6404 & n6764 ;
  assign n6766 = \u0_u1_csc_reg[6]/P0001  & n6408 ;
  assign n6767 = n6411 & n6766 ;
  assign n6768 = ~n6765 & ~n6767 ;
  assign n6769 = \u0_csc_mask_r_reg[6]/NET0131  & n6405 ;
  assign n6770 = n6411 & n6769 ;
  assign n6771 = \u0_csr_r_reg[6]/NET0131  & n6405 ;
  assign n6772 = n6404 & n6771 ;
  assign n6773 = ~n6770 & ~n6772 ;
  assign n6774 = n6768 & n6773 ;
  assign n6775 = \u0_u1_tms_reg[6]/P0001  & n6412 ;
  assign n6776 = n6411 & n6775 ;
  assign n6777 = ~n2191 & ~n6776 ;
  assign n6778 = \u0_u0_tms_reg[6]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6779 = n6421 & n6778 ;
  assign n6780 = \poc_o[6]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6781 = n6421 & n6780 ;
  assign n6782 = ~n6779 & ~n6781 ;
  assign n6783 = n6777 & n6782 ;
  assign n6784 = n6774 & n6783 ;
  assign n6785 = ~n6763 & ~n6784 ;
  assign n6786 = ~n2508 & n6392 ;
  assign n6787 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[4]/P0001  ;
  assign n6788 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[4]/P0001  ;
  assign n6789 = ~n6787 & ~n6788 ;
  assign n6790 = ~n6392 & ~n6789 ;
  assign n6791 = n2191 & ~n6790 ;
  assign n6792 = ~n6786 & n6791 ;
  assign n6793 = \u0_u0_csc_reg[4]/P0001  & n6408 ;
  assign n6794 = n6404 & n6793 ;
  assign n6795 = \u0_u1_csc_reg[4]/P0001  & n6408 ;
  assign n6796 = n6411 & n6795 ;
  assign n6797 = ~n6794 & ~n6796 ;
  assign n6798 = \u0_csc_mask_r_reg[4]/NET0131  & n6405 ;
  assign n6799 = n6411 & n6798 ;
  assign n6800 = \u0_csr_r_reg[4]/NET0131  & n6405 ;
  assign n6801 = n6404 & n6800 ;
  assign n6802 = ~n6799 & ~n6801 ;
  assign n6803 = n6797 & n6802 ;
  assign n6804 = \u0_u1_tms_reg[4]/P0001  & n6412 ;
  assign n6805 = n6411 & n6804 ;
  assign n6806 = ~n2191 & ~n6805 ;
  assign n6807 = \u0_u0_tms_reg[4]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6808 = n6421 & n6807 ;
  assign n6809 = \poc_o[4]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6810 = n6421 & n6809 ;
  assign n6811 = ~n6808 & ~n6810 ;
  assign n6812 = n6806 & n6811 ;
  assign n6813 = n6803 & n6812 ;
  assign n6814 = ~n6792 & ~n6813 ;
  assign n6815 = \u5_tmr2_done_reg/NET0131  & n1385 ;
  assign n6816 = n1384 & n6815 ;
  assign n6817 = n1122 & n6816 ;
  assign n6818 = \u5_state_reg[45]/NET0131  & ~n2739 ;
  assign n6819 = ~n2736 & n6818 ;
  assign n6820 = ~n2734 & n6819 ;
  assign n6821 = n3723 & n5634 ;
  assign n6822 = n3727 & n6821 ;
  assign n6823 = n5628 & n6822 ;
  assign n6824 = n964 & n1007 ;
  assign n6825 = n1069 & n1356 ;
  assign n6826 = n6824 & n6825 ;
  assign n6827 = n1051 & n6826 ;
  assign n6828 = n6823 & n6827 ;
  assign n6829 = ~n6820 & ~n6828 ;
  assign n6830 = ~\u1_acs_addr_reg[10]/P0001  & ~n5149 ;
  assign n6831 = ~n5152 & ~n6830 ;
  assign n6832 = \u0_init_ack_r_reg/P0001  & ~\u5_state_reg[26]/NET0131  ;
  assign n6833 = \u0_spec_req_cs_reg[0]/NET0131  & n6832 ;
  assign n6834 = n983 & n6833 ;
  assign n6835 = \u0_u0_init_req_reg/NET0131  & ~n6834 ;
  assign n6836 = \u0_u0_init_req_we_reg/NET0131  & ~\u0_u0_inited_reg/NET0131  ;
  assign n6837 = n1838 & n6836 ;
  assign n6838 = ~n6835 & ~n6837 ;
  assign n6839 = \u0_spec_req_cs_reg[1]/NET0131  & n6832 ;
  assign n6840 = n983 & n6839 ;
  assign n6841 = \u0_u1_init_req_reg/NET0131  & ~n6840 ;
  assign n6842 = \u0_u1_init_req_we_reg/NET0131  & ~\u0_u1_inited_reg/NET0131  ;
  assign n6843 = n1917 & n6842 ;
  assign n6844 = ~n6841 & ~n6843 ;
  assign n6845 = \u5_tmr2_done_reg/NET0131  & n1297 ;
  assign n6846 = n1296 & n6845 ;
  assign n6847 = n1292 & n6846 ;
  assign n6848 = \u3_byte2_reg[0]/P0001  & n5304 ;
  assign n6849 = \u7_mc_data_ir_reg[0]/P0001  & n5309 ;
  assign n6850 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[16]/P0001  ;
  assign n6851 = ~n6392 & ~n6850 ;
  assign n6852 = ~n6849 & n6851 ;
  assign n6853 = ~n6848 & n6852 ;
  assign n6854 = n2191 & n6853 ;
  assign n6855 = n2445 & n6394 ;
  assign n6856 = ~n6854 & ~n6855 ;
  assign n6857 = \u0_u1_csc_reg[16]/P0001  & n6408 ;
  assign n6858 = n6411 & n6857 ;
  assign n6859 = ~n2191 & ~n6858 ;
  assign n6860 = \u0_u1_tms_reg[16]/P0001  & n6412 ;
  assign n6861 = n6411 & n6860 ;
  assign n6862 = \u0_u0_csc_reg[16]/P0001  & n6408 ;
  assign n6863 = n6404 & n6862 ;
  assign n6864 = ~n6861 & ~n6863 ;
  assign n6865 = n6859 & n6864 ;
  assign n6866 = ~\poc_o[16]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6867 = ~\u0_u0_tms_reg[16]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6868 = ~n6866 & ~n6867 ;
  assign n6869 = n6421 & n6868 ;
  assign n6870 = n6865 & ~n6869 ;
  assign n6871 = n6856 & ~n6870 ;
  assign n6872 = \u3_byte2_reg[1]/P0001  & n5304 ;
  assign n6873 = \u7_mc_data_ir_reg[1]/P0001  & n5309 ;
  assign n6874 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[17]/P0001  ;
  assign n6875 = ~n6392 & ~n6874 ;
  assign n6876 = ~n6873 & n6875 ;
  assign n6877 = ~n6872 & n6876 ;
  assign n6878 = n2191 & n6877 ;
  assign n6879 = n2405 & n6394 ;
  assign n6880 = ~n6878 & ~n6879 ;
  assign n6881 = \u0_u1_csc_reg[17]/P0001  & n6408 ;
  assign n6882 = n6411 & n6881 ;
  assign n6883 = ~n2191 & ~n6882 ;
  assign n6884 = \u0_u1_tms_reg[17]/P0001  & n6412 ;
  assign n6885 = n6411 & n6884 ;
  assign n6886 = \u0_u0_csc_reg[17]/P0001  & n6408 ;
  assign n6887 = n6404 & n6886 ;
  assign n6888 = ~n6885 & ~n6887 ;
  assign n6889 = n6883 & n6888 ;
  assign n6890 = ~\poc_o[17]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6891 = ~\u0_u0_tms_reg[17]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6892 = ~n6890 & ~n6891 ;
  assign n6893 = n6421 & n6892 ;
  assign n6894 = n6889 & ~n6893 ;
  assign n6895 = n6880 & ~n6894 ;
  assign n6896 = \u3_byte2_reg[2]/P0001  & n5304 ;
  assign n6897 = \u7_mc_data_ir_reg[2]/P0001  & n5309 ;
  assign n6898 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[18]/P0001  ;
  assign n6899 = ~n6392 & ~n6898 ;
  assign n6900 = ~n6897 & n6899 ;
  assign n6901 = ~n6896 & n6900 ;
  assign n6902 = n2191 & n6901 ;
  assign n6903 = n2469 & n6394 ;
  assign n6904 = ~n6902 & ~n6903 ;
  assign n6905 = \u0_u1_csc_reg[18]/P0001  & n6408 ;
  assign n6906 = n6411 & n6905 ;
  assign n6907 = ~n2191 & ~n6906 ;
  assign n6908 = \u0_u1_tms_reg[18]/P0001  & n6412 ;
  assign n6909 = n6411 & n6908 ;
  assign n6910 = \u0_u0_csc_reg[18]/P0001  & n6408 ;
  assign n6911 = n6404 & n6910 ;
  assign n6912 = ~n6909 & ~n6911 ;
  assign n6913 = n6907 & n6912 ;
  assign n6914 = ~\poc_o[18]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6915 = ~\u0_u0_tms_reg[18]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6916 = ~n6914 & ~n6915 ;
  assign n6917 = n6421 & n6916 ;
  assign n6918 = n6913 & ~n6917 ;
  assign n6919 = n6904 & ~n6918 ;
  assign n6920 = \u3_byte2_reg[3]/P0001  & n5304 ;
  assign n6921 = \u7_mc_data_ir_reg[3]/P0001  & n5309 ;
  assign n6922 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[19]/P0001  ;
  assign n6923 = ~n6392 & ~n6922 ;
  assign n6924 = ~n6921 & n6923 ;
  assign n6925 = ~n6920 & n6924 ;
  assign n6926 = n2191 & n6925 ;
  assign n6927 = n2422 & n6394 ;
  assign n6928 = ~n6926 & ~n6927 ;
  assign n6929 = \u0_u1_csc_reg[19]/P0001  & n6408 ;
  assign n6930 = n6411 & n6929 ;
  assign n6931 = ~n2191 & ~n6930 ;
  assign n6932 = \u0_u1_tms_reg[19]/P0001  & n6412 ;
  assign n6933 = n6411 & n6932 ;
  assign n6934 = \u0_u0_csc_reg[19]/P0001  & n6408 ;
  assign n6935 = n6404 & n6934 ;
  assign n6936 = ~n6933 & ~n6935 ;
  assign n6937 = n6931 & n6936 ;
  assign n6938 = ~\poc_o[19]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6939 = ~\u0_u0_tms_reg[19]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6940 = ~n6938 & ~n6939 ;
  assign n6941 = n6421 & n6940 ;
  assign n6942 = n6937 & ~n6941 ;
  assign n6943 = n6928 & ~n6942 ;
  assign n6944 = \u3_byte2_reg[4]/P0001  & n5304 ;
  assign n6945 = \u7_mc_data_ir_reg[4]/P0001  & n5309 ;
  assign n6946 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[20]/P0001  ;
  assign n6947 = ~n6392 & ~n6946 ;
  assign n6948 = ~n6945 & n6947 ;
  assign n6949 = ~n6944 & n6948 ;
  assign n6950 = n2191 & n6949 ;
  assign n6951 = n2429 & n6394 ;
  assign n6952 = ~n6950 & ~n6951 ;
  assign n6953 = \u0_u1_csc_reg[20]/P0001  & n6408 ;
  assign n6954 = n6411 & n6953 ;
  assign n6955 = ~n2191 & ~n6954 ;
  assign n6956 = \u0_u1_tms_reg[20]/P0001  & n6412 ;
  assign n6957 = n6411 & n6956 ;
  assign n6958 = \u0_u0_csc_reg[20]/P0001  & n6408 ;
  assign n6959 = n6404 & n6958 ;
  assign n6960 = ~n6957 & ~n6959 ;
  assign n6961 = n6955 & n6960 ;
  assign n6962 = ~\poc_o[20]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6963 = ~\u0_u0_tms_reg[20]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = n6421 & n6964 ;
  assign n6966 = n6961 & ~n6965 ;
  assign n6967 = n6952 & ~n6966 ;
  assign n6968 = \u3_byte2_reg[6]/P0001  & n5304 ;
  assign n6969 = \u7_mc_data_ir_reg[6]/P0001  & n5309 ;
  assign n6970 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[22]/P0001  ;
  assign n6971 = ~n6392 & ~n6970 ;
  assign n6972 = ~n6969 & n6971 ;
  assign n6973 = ~n6968 & n6972 ;
  assign n6974 = n2191 & n6973 ;
  assign n6975 = n2415 & n6394 ;
  assign n6976 = ~n6974 & ~n6975 ;
  assign n6977 = \u0_u1_csc_reg[22]/P0001  & n6408 ;
  assign n6978 = n6411 & n6977 ;
  assign n6979 = ~n2191 & ~n6978 ;
  assign n6980 = \u0_u1_tms_reg[22]/P0001  & n6412 ;
  assign n6981 = n6411 & n6980 ;
  assign n6982 = \u0_u0_csc_reg[22]/P0001  & n6408 ;
  assign n6983 = n6404 & n6982 ;
  assign n6984 = ~n6981 & ~n6983 ;
  assign n6985 = n6979 & n6984 ;
  assign n6986 = ~\poc_o[22]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n6987 = ~\u0_u0_tms_reg[22]/P0001  & \wb_addr_i[4]_pad  ;
  assign n6988 = ~n6986 & ~n6987 ;
  assign n6989 = n6421 & n6988 ;
  assign n6990 = n6985 & ~n6989 ;
  assign n6991 = n6976 & ~n6990 ;
  assign n6992 = \u3_byte2_reg[7]/P0001  & n5304 ;
  assign n6993 = \u7_mc_data_ir_reg[7]/P0001  & n5309 ;
  assign n6994 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[23]/P0001  ;
  assign n6995 = ~n6392 & ~n6994 ;
  assign n6996 = ~n6993 & n6995 ;
  assign n6997 = ~n6992 & n6996 ;
  assign n6998 = n2191 & n6997 ;
  assign n6999 = n2452 & n6394 ;
  assign n7000 = ~n6998 & ~n6999 ;
  assign n7001 = \u0_u1_csc_reg[23]/P0001  & n6408 ;
  assign n7002 = n6411 & n7001 ;
  assign n7003 = ~n2191 & ~n7002 ;
  assign n7004 = \u0_u1_tms_reg[23]/P0001  & n6412 ;
  assign n7005 = n6411 & n7004 ;
  assign n7006 = \u0_u0_csc_reg[23]/P0001  & n6408 ;
  assign n7007 = n6404 & n7006 ;
  assign n7008 = ~n7005 & ~n7007 ;
  assign n7009 = n7003 & n7008 ;
  assign n7010 = ~\poc_o[23]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7011 = ~\u0_u0_tms_reg[23]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7012 = ~n7010 & ~n7011 ;
  assign n7013 = n6421 & n7012 ;
  assign n7014 = n7009 & ~n7013 ;
  assign n7015 = n7000 & ~n7014 ;
  assign n7016 = \u3_byte2_reg[5]/P0001  & n5304 ;
  assign n7017 = \u7_mc_data_ir_reg[5]/P0001  & n5309 ;
  assign n7018 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[21]/P0001  ;
  assign n7019 = ~n6392 & ~n7018 ;
  assign n7020 = ~n7017 & n7019 ;
  assign n7021 = ~n7016 & n7020 ;
  assign n7022 = n2191 & n7021 ;
  assign n7023 = n2398 & n6394 ;
  assign n7024 = ~n7022 & ~n7023 ;
  assign n7025 = \u0_u1_csc_reg[21]/P0001  & n6408 ;
  assign n7026 = n6411 & n7025 ;
  assign n7027 = ~n2191 & ~n7026 ;
  assign n7028 = \u0_u1_tms_reg[21]/P0001  & n6412 ;
  assign n7029 = n6411 & n7028 ;
  assign n7030 = \u0_u0_csc_reg[21]/P0001  & n6408 ;
  assign n7031 = n6404 & n7030 ;
  assign n7032 = ~n7029 & ~n7031 ;
  assign n7033 = n7027 & n7032 ;
  assign n7034 = ~\poc_o[21]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7035 = ~\u0_u0_tms_reg[21]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7036 = ~n7034 & ~n7035 ;
  assign n7037 = n6421 & n7036 ;
  assign n7038 = n7033 & ~n7037 ;
  assign n7039 = n7024 & ~n7038 ;
  assign n7040 = ~n2235 & n6392 ;
  assign n7041 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[3]/P0001  ;
  assign n7042 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[11]/P0001  ;
  assign n7043 = ~n7041 & ~n7042 ;
  assign n7044 = ~n6392 & ~n7043 ;
  assign n7045 = n2191 & ~n7044 ;
  assign n7046 = ~n7040 & n7045 ;
  assign n7047 = \u0_u1_csc_reg[11]/P0001  & n6408 ;
  assign n7048 = n6411 & n7047 ;
  assign n7049 = ~n2191 & ~n7048 ;
  assign n7050 = \u0_u1_tms_reg[11]/P0001  & n6412 ;
  assign n7051 = n6411 & n7050 ;
  assign n7052 = \u0_u0_csc_reg[11]/P0001  & n6408 ;
  assign n7053 = n6404 & n7052 ;
  assign n7054 = ~n7051 & ~n7053 ;
  assign n7055 = n7049 & n7054 ;
  assign n7056 = ~\poc_o[11]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7057 = ~\u0_u0_tms_reg[11]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7058 = ~n7056 & ~n7057 ;
  assign n7059 = n6421 & n7058 ;
  assign n7060 = n7055 & ~n7059 ;
  assign n7061 = ~n7046 & ~n7060 ;
  assign n7062 = ~n2242 & n6392 ;
  assign n7063 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[4]/P0001  ;
  assign n7064 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[12]/P0001  ;
  assign n7065 = ~n7063 & ~n7064 ;
  assign n7066 = ~n6392 & ~n7065 ;
  assign n7067 = n2191 & ~n7066 ;
  assign n7068 = ~n7062 & n7067 ;
  assign n7069 = \u0_u1_csc_reg[12]/P0001  & n6408 ;
  assign n7070 = n6411 & n7069 ;
  assign n7071 = ~n2191 & ~n7070 ;
  assign n7072 = \u0_u1_tms_reg[12]/P0001  & n6412 ;
  assign n7073 = n6411 & n7072 ;
  assign n7074 = \u0_u0_csc_reg[12]/P0001  & n6408 ;
  assign n7075 = n6404 & n7074 ;
  assign n7076 = ~n7073 & ~n7075 ;
  assign n7077 = n7071 & n7076 ;
  assign n7078 = ~\poc_o[12]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7079 = ~\u0_u0_tms_reg[12]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7080 = ~n7078 & ~n7079 ;
  assign n7081 = n6421 & n7080 ;
  assign n7082 = n7077 & ~n7081 ;
  assign n7083 = ~n7068 & ~n7082 ;
  assign n7084 = ~n2228 & n6392 ;
  assign n7085 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[6]/P0001  ;
  assign n7086 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[14]/P0001  ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7088 = ~n6392 & ~n7087 ;
  assign n7089 = n2191 & ~n7088 ;
  assign n7090 = ~n7084 & n7089 ;
  assign n7091 = \u0_u1_csc_reg[14]/P0001  & n6408 ;
  assign n7092 = n6411 & n7091 ;
  assign n7093 = ~n2191 & ~n7092 ;
  assign n7094 = \u0_u1_tms_reg[14]/P0001  & n6412 ;
  assign n7095 = n6411 & n7094 ;
  assign n7096 = \u0_u0_csc_reg[14]/P0001  & n6408 ;
  assign n7097 = n6404 & n7096 ;
  assign n7098 = ~n7095 & ~n7097 ;
  assign n7099 = n7093 & n7098 ;
  assign n7100 = ~\poc_o[14]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7101 = ~\u0_u0_tms_reg[14]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7102 = ~n7100 & ~n7101 ;
  assign n7103 = n6421 & n7102 ;
  assign n7104 = n7099 & ~n7103 ;
  assign n7105 = ~n7090 & ~n7104 ;
  assign n7106 = ~n2265 & n6392 ;
  assign n7107 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[7]/P0001  ;
  assign n7108 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[15]/P0001  ;
  assign n7109 = ~n7107 & ~n7108 ;
  assign n7110 = ~n6392 & ~n7109 ;
  assign n7111 = n2191 & ~n7110 ;
  assign n7112 = ~n7106 & n7111 ;
  assign n7113 = \u0_u1_csc_reg[15]/P0001  & n6408 ;
  assign n7114 = n6411 & n7113 ;
  assign n7115 = ~n2191 & ~n7114 ;
  assign n7116 = \u0_u1_tms_reg[15]/P0001  & n6412 ;
  assign n7117 = n6411 & n7116 ;
  assign n7118 = \u0_u0_csc_reg[15]/P0001  & n6408 ;
  assign n7119 = n6404 & n7118 ;
  assign n7120 = ~n7117 & ~n7119 ;
  assign n7121 = n7115 & n7120 ;
  assign n7122 = ~\poc_o[15]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7123 = ~\u0_u0_tms_reg[15]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7124 = ~n7122 & ~n7123 ;
  assign n7125 = n6421 & n7124 ;
  assign n7126 = n7121 & ~n7125 ;
  assign n7127 = ~n7112 & ~n7126 ;
  assign n7128 = ~n2211 & n6392 ;
  assign n7129 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[5]/P0001  ;
  assign n7130 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[13]/P0001  ;
  assign n7131 = ~n7129 & ~n7130 ;
  assign n7132 = ~n6392 & ~n7131 ;
  assign n7133 = n2191 & ~n7132 ;
  assign n7134 = ~n7128 & n7133 ;
  assign n7135 = \u0_u1_csc_reg[13]/P0001  & n6408 ;
  assign n7136 = n6411 & n7135 ;
  assign n7137 = ~n2191 & ~n7136 ;
  assign n7138 = \u0_u1_tms_reg[13]/P0001  & n6412 ;
  assign n7139 = n6411 & n7138 ;
  assign n7140 = \u0_u0_csc_reg[13]/P0001  & n6408 ;
  assign n7141 = n6404 & n7140 ;
  assign n7142 = ~n7139 & ~n7141 ;
  assign n7143 = n7137 & n7142 ;
  assign n7144 = ~\poc_o[13]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7145 = ~\u0_u0_tms_reg[13]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7146 = ~n7144 & ~n7145 ;
  assign n7147 = n6421 & n7146 ;
  assign n7148 = n7143 & ~n7147 ;
  assign n7149 = ~n7134 & ~n7148 ;
  assign n7150 = ~\u0_u0_csc_reg[1]/NET0131  & ~n6381 ;
  assign n7151 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[1]_pad  ;
  assign n7152 = n6379 & n7151 ;
  assign n7153 = n6378 & n7152 ;
  assign n7154 = ~\u0_rst_r2_reg/NET0131  & ~n7153 ;
  assign n7155 = ~n7150 & n7154 ;
  assign n7156 = ~n6389 & ~n7155 ;
  assign n7157 = ~\u0_u0_csc_reg[2]/NET0131  & ~n6381 ;
  assign n7158 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[2]_pad  ;
  assign n7159 = n6379 & n7158 ;
  assign n7160 = n6378 & n7159 ;
  assign n7161 = ~\u0_rst_r2_reg/NET0131  & ~n7160 ;
  assign n7162 = ~n7157 & n7161 ;
  assign n7163 = ~n6388 & ~n7162 ;
  assign n7164 = \u1_acs_addr_reg[4]/P0001  & \u1_acs_addr_reg[5]/P0001  ;
  assign n7165 = n5143 & n7164 ;
  assign n7166 = ~\u1_acs_addr_reg[6]/P0001  & ~n7165 ;
  assign n7167 = ~n5146 & ~n7166 ;
  assign n7168 = ~n2491 & n6392 ;
  assign n7169 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[0]/P0001  ;
  assign n7170 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[0]/P0001  ;
  assign n7171 = ~n7169 & ~n7170 ;
  assign n7172 = ~n6392 & ~n7171 ;
  assign n7173 = n2191 & ~n7172 ;
  assign n7174 = ~n7168 & n7173 ;
  assign n7175 = \u0_u0_csc_reg[0]/NET0131  & n6408 ;
  assign n7176 = n6404 & n7175 ;
  assign n7177 = \u0_csc_mask_r_reg[0]/NET0131  & n6405 ;
  assign n7178 = n6411 & n7177 ;
  assign n7179 = ~n7176 & ~n7178 ;
  assign n7180 = \u0_u1_csc_reg[0]/NET0131  & n6408 ;
  assign n7181 = n6411 & n7180 ;
  assign n7182 = \u0_csr_r_reg[0]/P0001  & n6405 ;
  assign n7183 = n6404 & n7182 ;
  assign n7184 = ~n7181 & ~n7183 ;
  assign n7185 = n7179 & n7184 ;
  assign n7186 = \u0_u1_tms_reg[0]/P0001  & n6412 ;
  assign n7187 = n6411 & n7186 ;
  assign n7188 = ~n2191 & ~n7187 ;
  assign n7189 = \u0_u0_tms_reg[0]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7190 = n6421 & n7189 ;
  assign n7191 = \poc_o[0]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7192 = n6421 & n7191 ;
  assign n7193 = ~n7190 & ~n7192 ;
  assign n7194 = n7188 & n7193 ;
  assign n7195 = n7185 & n7194 ;
  assign n7196 = ~n7174 & ~n7195 ;
  assign n7197 = ~n2282 & n6392 ;
  assign n7198 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[2]/P0001  ;
  assign n7199 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[10]/P0001  ;
  assign n7200 = ~n7198 & ~n7199 ;
  assign n7201 = ~n6392 & ~n7200 ;
  assign n7202 = n2191 & ~n7201 ;
  assign n7203 = ~n7197 & n7202 ;
  assign n7204 = \u0_u0_csc_reg[10]/P0001  & n6408 ;
  assign n7205 = n6404 & n7204 ;
  assign n7206 = \u0_csr_r_reg[10]/NET0131  & n6405 ;
  assign n7207 = n6404 & n7206 ;
  assign n7208 = ~n7205 & ~n7207 ;
  assign n7209 = \u0_u1_csc_reg[10]/P0001  & n6408 ;
  assign n7210 = n6411 & n7209 ;
  assign n7211 = \u0_csc_mask_r_reg[10]/NET0131  & n6405 ;
  assign n7212 = n6411 & n7211 ;
  assign n7213 = ~n7210 & ~n7212 ;
  assign n7214 = n7208 & n7213 ;
  assign n7215 = \u0_u1_tms_reg[10]/P0001  & n6412 ;
  assign n7216 = n6411 & n7215 ;
  assign n7217 = ~n2191 & ~n7216 ;
  assign n7218 = \u0_u0_tms_reg[10]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7219 = n6421 & n7218 ;
  assign n7220 = \poc_o[10]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7221 = n6421 & n7220 ;
  assign n7222 = ~n7219 & ~n7221 ;
  assign n7223 = n7217 & n7222 ;
  assign n7224 = n7214 & n7223 ;
  assign n7225 = ~n7203 & ~n7224 ;
  assign n7226 = ~n2498 & n6392 ;
  assign n7227 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[2]/P0001  ;
  assign n7228 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[2]/P0001  ;
  assign n7229 = ~n7227 & ~n7228 ;
  assign n7230 = ~n6392 & ~n7229 ;
  assign n7231 = n2191 & ~n7230 ;
  assign n7232 = ~n7226 & n7231 ;
  assign n7233 = \u0_csr_r_reg[2]/NET0131  & n6405 ;
  assign n7234 = n6404 & n7233 ;
  assign n7235 = \u0_u0_csc_reg[2]/NET0131  & n6408 ;
  assign n7236 = n6404 & n7235 ;
  assign n7237 = ~n7234 & ~n7236 ;
  assign n7238 = \u0_u1_tms_reg[2]/P0001  & n6412 ;
  assign n7239 = n6411 & n7238 ;
  assign n7240 = \u0_csc_mask_r_reg[2]/NET0131  & n6405 ;
  assign n7241 = n6411 & n7240 ;
  assign n7242 = ~n7239 & ~n7241 ;
  assign n7243 = n7237 & n7242 ;
  assign n7244 = \u0_u1_csc_reg[2]/NET0131  & n6408 ;
  assign n7245 = n6411 & n7244 ;
  assign n7246 = ~n2191 & ~n7245 ;
  assign n7247 = \u0_u0_tms_reg[2]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7248 = n6421 & n7247 ;
  assign n7249 = \poc_o[2]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7250 = n6421 & n7249 ;
  assign n7251 = ~n7248 & ~n7250 ;
  assign n7252 = n7246 & n7251 ;
  assign n7253 = n7243 & n7252 ;
  assign n7254 = ~n7232 & ~n7253 ;
  assign n7255 = ~n2515 & n6392 ;
  assign n7256 = ~\u0_csc_reg[5]/NET0131  & \u3_byte0_reg[7]/P0001  ;
  assign n7257 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[7]/P0001  ;
  assign n7258 = ~n7256 & ~n7257 ;
  assign n7259 = ~n6392 & ~n7258 ;
  assign n7260 = n2191 & ~n7259 ;
  assign n7261 = ~n7255 & n7260 ;
  assign n7262 = \u0_u0_csc_reg[7]/P0001  & n6408 ;
  assign n7263 = n6404 & n7262 ;
  assign n7264 = \u0_csc_mask_r_reg[7]/NET0131  & n6405 ;
  assign n7265 = n6411 & n7264 ;
  assign n7266 = ~n7263 & ~n7265 ;
  assign n7267 = \u0_u1_csc_reg[7]/P0001  & n6408 ;
  assign n7268 = n6411 & n7267 ;
  assign n7269 = \u0_csr_r_reg[7]/NET0131  & n6405 ;
  assign n7270 = n6404 & n7269 ;
  assign n7271 = ~n7268 & ~n7270 ;
  assign n7272 = n7266 & n7271 ;
  assign n7273 = \u0_u1_tms_reg[7]/P0001  & n6412 ;
  assign n7274 = n6411 & n7273 ;
  assign n7275 = ~n2191 & ~n7274 ;
  assign n7276 = \u0_u0_tms_reg[7]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7277 = n6421 & n7276 ;
  assign n7278 = \poc_o[7]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7279 = n6421 & n7278 ;
  assign n7280 = ~n7277 & ~n7279 ;
  assign n7281 = n7275 & n7280 ;
  assign n7282 = n7272 & n7281 ;
  assign n7283 = ~n7261 & ~n7282 ;
  assign n7284 = ~n2258 & n6392 ;
  assign n7285 = ~\u0_csc_reg[5]/NET0131  & \u3_byte1_reg[0]/P0001  ;
  assign n7286 = \u0_csc_reg[5]/NET0131  & \u7_mc_data_ir_reg[8]/P0001  ;
  assign n7287 = ~n7285 & ~n7286 ;
  assign n7288 = ~n6392 & ~n7287 ;
  assign n7289 = n2191 & ~n7288 ;
  assign n7290 = ~n7284 & n7289 ;
  assign n7291 = \u0_u0_csc_reg[8]/P0001  & n6408 ;
  assign n7292 = n6404 & n7291 ;
  assign n7293 = \u0_csr_r_reg[8]/NET0131  & n6405 ;
  assign n7294 = n6404 & n7293 ;
  assign n7295 = ~n7292 & ~n7294 ;
  assign n7296 = \u0_u1_csc_reg[8]/P0001  & n6408 ;
  assign n7297 = n6411 & n7296 ;
  assign n7298 = \u0_csc_mask_r_reg[8]/NET0131  & n6405 ;
  assign n7299 = n6411 & n7298 ;
  assign n7300 = ~n7297 & ~n7299 ;
  assign n7301 = n7295 & n7300 ;
  assign n7302 = \u0_u1_tms_reg[8]/P0001  & n6412 ;
  assign n7303 = n6411 & n7302 ;
  assign n7304 = ~n2191 & ~n7303 ;
  assign n7305 = \u0_u0_tms_reg[8]/P0001  & \wb_addr_i[4]_pad  ;
  assign n7306 = n6421 & n7305 ;
  assign n7307 = \poc_o[8]_pad  & ~\wb_addr_i[4]_pad  ;
  assign n7308 = n6421 & n7307 ;
  assign n7309 = ~n7306 & ~n7308 ;
  assign n7310 = n7304 & n7309 ;
  assign n7311 = n7301 & n7310 ;
  assign n7312 = ~n7290 & ~n7311 ;
  assign n7313 = ~\u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[5]_pad  ;
  assign n7314 = n6379 & n7313 ;
  assign n7315 = n6378 & n7314 ;
  assign n7316 = ~\u0_rst_r2_reg/NET0131  & n7315 ;
  assign n7317 = ~\u0_rst_r2_reg/NET0131  & \u0_u0_csc_reg[5]/P0001  ;
  assign n7318 = ~n6381 & n7317 ;
  assign n7319 = ~n7316 & ~n7318 ;
  assign n7320 = \poc_o[1]_pad  & \u0_rst_r2_reg/NET0131  ;
  assign n7321 = n7319 & ~n7320 ;
  assign n7322 = ~\u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[4]_pad  ;
  assign n7323 = n6379 & n7322 ;
  assign n7324 = n6378 & n7323 ;
  assign n7325 = ~\u0_rst_r2_reg/NET0131  & n7324 ;
  assign n7326 = ~\u0_rst_r2_reg/NET0131  & \u0_u0_csc_reg[4]/P0001  ;
  assign n7327 = ~n6381 & n7326 ;
  assign n7328 = ~n7325 & ~n7327 ;
  assign n7329 = \poc_o[0]_pad  & \u0_rst_r2_reg/NET0131  ;
  assign n7330 = n7328 & ~n7329 ;
  assign n7331 = \u5_state_reg[45]/NET0131  & ~n2733 ;
  assign n7332 = ~n2730 & n7331 ;
  assign n7333 = n2740 & n7332 ;
  assign n7334 = ~\u0_u0_csc_reg[11]/P0001  & ~n6381 ;
  assign n7335 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[11]_pad  ;
  assign n7336 = n6379 & n7335 ;
  assign n7337 = n6378 & n7336 ;
  assign n7338 = ~\u0_rst_r2_reg/NET0131  & ~n7337 ;
  assign n7339 = ~n7334 & n7338 ;
  assign n7340 = ~\u0_u0_csc_reg[12]/P0001  & ~n6381 ;
  assign n7341 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[12]_pad  ;
  assign n7342 = n6379 & n7341 ;
  assign n7343 = n6378 & n7342 ;
  assign n7344 = ~\u0_rst_r2_reg/NET0131  & ~n7343 ;
  assign n7345 = ~n7340 & n7344 ;
  assign n7346 = \u0_u0_addr_r_reg[3]/P0001  & n6377 ;
  assign n7347 = \u0_u0_addr_r_reg[2]/P0001  & n6379 ;
  assign n7348 = n7346 & n7347 ;
  assign n7349 = ~\u0_u1_tms_reg[19]/P0001  & ~n7348 ;
  assign n7350 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[19]_pad  ;
  assign n7351 = n6379 & n7350 ;
  assign n7352 = n7346 & n7351 ;
  assign n7353 = ~\u0_rst_r2_reg/NET0131  & ~n7352 ;
  assign n7354 = ~n7349 & n7353 ;
  assign n7355 = ~\u0_u0_csc_reg[13]/P0001  & ~n6381 ;
  assign n7356 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[13]_pad  ;
  assign n7357 = n6379 & n7356 ;
  assign n7358 = n6378 & n7357 ;
  assign n7359 = ~\u0_rst_r2_reg/NET0131  & ~n7358 ;
  assign n7360 = ~n7355 & n7359 ;
  assign n7361 = ~\u0_u0_csc_reg[14]/P0001  & ~n6381 ;
  assign n7362 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[14]_pad  ;
  assign n7363 = n6379 & n7362 ;
  assign n7364 = n6378 & n7363 ;
  assign n7365 = ~\u0_rst_r2_reg/NET0131  & ~n7364 ;
  assign n7366 = ~n7361 & n7365 ;
  assign n7367 = ~\u0_u0_csc_reg[16]/P0001  & ~n6381 ;
  assign n7368 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[16]_pad  ;
  assign n7369 = n6379 & n7368 ;
  assign n7370 = n6378 & n7369 ;
  assign n7371 = ~\u0_rst_r2_reg/NET0131  & ~n7370 ;
  assign n7372 = ~n7367 & n7371 ;
  assign n7373 = ~\u0_u0_csc_reg[17]/P0001  & ~n6381 ;
  assign n7374 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[17]_pad  ;
  assign n7375 = n6379 & n7374 ;
  assign n7376 = n6378 & n7375 ;
  assign n7377 = ~\u0_rst_r2_reg/NET0131  & ~n7376 ;
  assign n7378 = ~n7373 & n7377 ;
  assign n7379 = ~\u0_u0_csc_reg[20]/P0001  & ~n6381 ;
  assign n7380 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[20]_pad  ;
  assign n7381 = n6379 & n7380 ;
  assign n7382 = n6378 & n7381 ;
  assign n7383 = ~\u0_rst_r2_reg/NET0131  & ~n7382 ;
  assign n7384 = ~n7379 & n7383 ;
  assign n7385 = ~\u0_u0_csc_reg[21]/P0001  & ~n6381 ;
  assign n7386 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[21]_pad  ;
  assign n7387 = n6379 & n7386 ;
  assign n7388 = n6378 & n7387 ;
  assign n7389 = ~\u0_rst_r2_reg/NET0131  & ~n7388 ;
  assign n7390 = ~n7385 & n7389 ;
  assign n7391 = ~\u0_u0_csc_reg[22]/P0001  & ~n6381 ;
  assign n7392 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[22]_pad  ;
  assign n7393 = n6379 & n7392 ;
  assign n7394 = n6378 & n7393 ;
  assign n7395 = ~\u0_rst_r2_reg/NET0131  & ~n7394 ;
  assign n7396 = ~n7391 & n7395 ;
  assign n7397 = ~\u0_u0_csc_reg[24]/P0001  & ~n6381 ;
  assign n7398 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[24]_pad  ;
  assign n7399 = n6379 & n7398 ;
  assign n7400 = n6378 & n7399 ;
  assign n7401 = ~\u0_rst_r2_reg/NET0131  & ~n7400 ;
  assign n7402 = ~n7397 & n7401 ;
  assign n7403 = ~\u0_u0_csc_reg[26]/P0001  & ~n6381 ;
  assign n7404 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[26]_pad  ;
  assign n7405 = n6379 & n7404 ;
  assign n7406 = n6378 & n7405 ;
  assign n7407 = ~\u0_rst_r2_reg/NET0131  & ~n7406 ;
  assign n7408 = ~n7403 & n7407 ;
  assign n7409 = ~\u0_u0_csc_reg[27]/P0001  & ~n6381 ;
  assign n7410 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[27]_pad  ;
  assign n7411 = n6379 & n7410 ;
  assign n7412 = n6378 & n7411 ;
  assign n7413 = ~\u0_rst_r2_reg/NET0131  & ~n7412 ;
  assign n7414 = ~n7409 & n7413 ;
  assign n7415 = ~\u0_u0_csc_reg[28]/P0001  & ~n6381 ;
  assign n7416 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[28]_pad  ;
  assign n7417 = n6379 & n7416 ;
  assign n7418 = n6378 & n7417 ;
  assign n7419 = ~\u0_rst_r2_reg/NET0131  & ~n7418 ;
  assign n7420 = ~n7415 & n7419 ;
  assign n7421 = ~\u0_u1_tms_reg[23]/P0001  & ~n7348 ;
  assign n7422 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[23]_pad  ;
  assign n7423 = n6379 & n7422 ;
  assign n7424 = n7346 & n7423 ;
  assign n7425 = ~\u0_rst_r2_reg/NET0131  & ~n7424 ;
  assign n7426 = ~n7421 & n7425 ;
  assign n7427 = ~\u0_u0_csc_reg[30]/P0001  & ~n6381 ;
  assign n7428 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[30]_pad  ;
  assign n7429 = n6379 & n7428 ;
  assign n7430 = n6378 & n7429 ;
  assign n7431 = ~\u0_rst_r2_reg/NET0131  & ~n7430 ;
  assign n7432 = ~n7427 & n7431 ;
  assign n7433 = ~\u0_u0_csc_reg[3]/NET0131  & ~n6381 ;
  assign n7434 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[3]_pad  ;
  assign n7435 = n6379 & n7434 ;
  assign n7436 = n6378 & n7435 ;
  assign n7437 = ~\u0_rst_r2_reg/NET0131  & ~n7436 ;
  assign n7438 = ~n7433 & n7437 ;
  assign n7439 = ~\u0_u0_csc_reg[25]/P0001  & ~n6381 ;
  assign n7440 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[25]_pad  ;
  assign n7441 = n6379 & n7440 ;
  assign n7442 = n6378 & n7441 ;
  assign n7443 = ~\u0_rst_r2_reg/NET0131  & ~n7442 ;
  assign n7444 = ~n7439 & n7443 ;
  assign n7445 = ~\u0_u1_tms_reg[17]/P0001  & ~n7348 ;
  assign n7446 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[17]_pad  ;
  assign n7447 = n6379 & n7446 ;
  assign n7448 = n7346 & n7447 ;
  assign n7449 = ~\u0_rst_r2_reg/NET0131  & ~n7448 ;
  assign n7450 = ~n7445 & n7449 ;
  assign n7451 = ~\u0_u1_tms_reg[16]/P0001  & ~n7348 ;
  assign n7452 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[16]_pad  ;
  assign n7453 = n6379 & n7452 ;
  assign n7454 = n7346 & n7453 ;
  assign n7455 = ~\u0_rst_r2_reg/NET0131  & ~n7454 ;
  assign n7456 = ~n7451 & n7455 ;
  assign n7457 = n6378 & n7347 ;
  assign n7458 = \u0_u0_tms_reg[0]/P0001  & ~n7457 ;
  assign n7459 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[0]_pad  ;
  assign n7460 = n6379 & n7459 ;
  assign n7461 = n6378 & n7460 ;
  assign n7462 = ~\u0_rst_r2_reg/NET0131  & ~n7461 ;
  assign n7463 = ~n7458 & n7462 ;
  assign n7464 = \u0_u0_tms_reg[10]/P0001  & ~n7457 ;
  assign n7465 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[10]_pad  ;
  assign n7466 = n6379 & n7465 ;
  assign n7467 = n6378 & n7466 ;
  assign n7468 = ~\u0_rst_r2_reg/NET0131  & ~n7467 ;
  assign n7469 = ~n7464 & n7468 ;
  assign n7470 = \u0_u0_tms_reg[11]/P0001  & ~n7457 ;
  assign n7471 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[11]_pad  ;
  assign n7472 = n6379 & n7471 ;
  assign n7473 = n6378 & n7472 ;
  assign n7474 = ~\u0_rst_r2_reg/NET0131  & ~n7473 ;
  assign n7475 = ~n7470 & n7474 ;
  assign n7476 = \u0_u0_tms_reg[12]/P0001  & ~n7457 ;
  assign n7477 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[12]_pad  ;
  assign n7478 = n6379 & n7477 ;
  assign n7479 = n6378 & n7478 ;
  assign n7480 = ~\u0_rst_r2_reg/NET0131  & ~n7479 ;
  assign n7481 = ~n7476 & n7480 ;
  assign n7482 = \u0_u0_tms_reg[14]/P0001  & ~n7457 ;
  assign n7483 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[14]_pad  ;
  assign n7484 = n6379 & n7483 ;
  assign n7485 = n6378 & n7484 ;
  assign n7486 = ~\u0_rst_r2_reg/NET0131  & ~n7485 ;
  assign n7487 = ~n7482 & n7486 ;
  assign n7488 = \u0_u0_tms_reg[13]/P0001  & ~n7457 ;
  assign n7489 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[13]_pad  ;
  assign n7490 = n6379 & n7489 ;
  assign n7491 = n6378 & n7490 ;
  assign n7492 = ~\u0_rst_r2_reg/NET0131  & ~n7491 ;
  assign n7493 = ~n7488 & n7492 ;
  assign n7494 = \u0_u0_tms_reg[15]/P0001  & ~n7457 ;
  assign n7495 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[15]_pad  ;
  assign n7496 = n6379 & n7495 ;
  assign n7497 = n6378 & n7496 ;
  assign n7498 = ~\u0_rst_r2_reg/NET0131  & ~n7497 ;
  assign n7499 = ~n7494 & n7498 ;
  assign n7500 = \u0_u0_tms_reg[16]/P0001  & ~n7457 ;
  assign n7501 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[16]_pad  ;
  assign n7502 = n6379 & n7501 ;
  assign n7503 = n6378 & n7502 ;
  assign n7504 = ~\u0_rst_r2_reg/NET0131  & ~n7503 ;
  assign n7505 = ~n7500 & n7504 ;
  assign n7506 = \u0_u0_tms_reg[17]/P0001  & ~n7457 ;
  assign n7507 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[17]_pad  ;
  assign n7508 = n6379 & n7507 ;
  assign n7509 = n6378 & n7508 ;
  assign n7510 = ~\u0_rst_r2_reg/NET0131  & ~n7509 ;
  assign n7511 = ~n7506 & n7510 ;
  assign n7512 = \u0_u0_tms_reg[18]/P0001  & ~n7457 ;
  assign n7513 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[18]_pad  ;
  assign n7514 = n6379 & n7513 ;
  assign n7515 = n6378 & n7514 ;
  assign n7516 = ~\u0_rst_r2_reg/NET0131  & ~n7515 ;
  assign n7517 = ~n7512 & n7516 ;
  assign n7518 = \u0_u0_tms_reg[19]/P0001  & ~n7457 ;
  assign n7519 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[19]_pad  ;
  assign n7520 = n6379 & n7519 ;
  assign n7521 = n6378 & n7520 ;
  assign n7522 = ~\u0_rst_r2_reg/NET0131  & ~n7521 ;
  assign n7523 = ~n7518 & n7522 ;
  assign n7524 = \u0_u0_tms_reg[1]/P0001  & ~n7457 ;
  assign n7525 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[1]_pad  ;
  assign n7526 = n6379 & n7525 ;
  assign n7527 = n6378 & n7526 ;
  assign n7528 = ~\u0_rst_r2_reg/NET0131  & ~n7527 ;
  assign n7529 = ~n7524 & n7528 ;
  assign n7530 = \u0_u0_tms_reg[21]/P0001  & ~n7457 ;
  assign n7531 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[21]_pad  ;
  assign n7532 = n6379 & n7531 ;
  assign n7533 = n6378 & n7532 ;
  assign n7534 = ~\u0_rst_r2_reg/NET0131  & ~n7533 ;
  assign n7535 = ~n7530 & n7534 ;
  assign n7536 = \u0_u0_tms_reg[22]/P0001  & ~n7457 ;
  assign n7537 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[22]_pad  ;
  assign n7538 = n6379 & n7537 ;
  assign n7539 = n6378 & n7538 ;
  assign n7540 = ~\u0_rst_r2_reg/NET0131  & ~n7539 ;
  assign n7541 = ~n7536 & n7540 ;
  assign n7542 = \u0_u0_tms_reg[23]/P0001  & ~n7457 ;
  assign n7543 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[23]_pad  ;
  assign n7544 = n6379 & n7543 ;
  assign n7545 = n6378 & n7544 ;
  assign n7546 = ~\u0_rst_r2_reg/NET0131  & ~n7545 ;
  assign n7547 = ~n7542 & n7546 ;
  assign n7548 = \u0_u0_tms_reg[24]/P0001  & ~n7457 ;
  assign n7549 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[24]_pad  ;
  assign n7550 = n6379 & n7549 ;
  assign n7551 = n6378 & n7550 ;
  assign n7552 = ~\u0_rst_r2_reg/NET0131  & ~n7551 ;
  assign n7553 = ~n7548 & n7552 ;
  assign n7554 = \u0_u0_tms_reg[25]/P0001  & ~n7457 ;
  assign n7555 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[25]_pad  ;
  assign n7556 = n6379 & n7555 ;
  assign n7557 = n6378 & n7556 ;
  assign n7558 = ~\u0_rst_r2_reg/NET0131  & ~n7557 ;
  assign n7559 = ~n7554 & n7558 ;
  assign n7560 = \u0_u0_tms_reg[26]/P0001  & ~n7457 ;
  assign n7561 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[26]_pad  ;
  assign n7562 = n6379 & n7561 ;
  assign n7563 = n6378 & n7562 ;
  assign n7564 = ~\u0_rst_r2_reg/NET0131  & ~n7563 ;
  assign n7565 = ~n7560 & n7564 ;
  assign n7566 = \u0_u0_tms_reg[27]/P0001  & ~n7457 ;
  assign n7567 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[27]_pad  ;
  assign n7568 = n6379 & n7567 ;
  assign n7569 = n6378 & n7568 ;
  assign n7570 = ~\u0_rst_r2_reg/NET0131  & ~n7569 ;
  assign n7571 = ~n7566 & n7570 ;
  assign n7572 = ~\u0_u1_tms_reg[22]/P0001  & ~n7348 ;
  assign n7573 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[22]_pad  ;
  assign n7574 = n6379 & n7573 ;
  assign n7575 = n7346 & n7574 ;
  assign n7576 = ~\u0_rst_r2_reg/NET0131  & ~n7575 ;
  assign n7577 = ~n7572 & n7576 ;
  assign n7578 = \u0_u0_tms_reg[28]/P0001  & ~n7457 ;
  assign n7579 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[28]_pad  ;
  assign n7580 = n6379 & n7579 ;
  assign n7581 = n6378 & n7580 ;
  assign n7582 = ~\u0_rst_r2_reg/NET0131  & ~n7581 ;
  assign n7583 = ~n7578 & n7582 ;
  assign n7584 = \u0_u0_tms_reg[29]/P0001  & ~n7457 ;
  assign n7585 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[29]_pad  ;
  assign n7586 = n6379 & n7585 ;
  assign n7587 = n6378 & n7586 ;
  assign n7588 = ~\u0_rst_r2_reg/NET0131  & ~n7587 ;
  assign n7589 = ~n7584 & n7588 ;
  assign n7590 = \u0_u0_tms_reg[2]/P0001  & ~n7457 ;
  assign n7591 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[2]_pad  ;
  assign n7592 = n6379 & n7591 ;
  assign n7593 = n6378 & n7592 ;
  assign n7594 = ~\u0_rst_r2_reg/NET0131  & ~n7593 ;
  assign n7595 = ~n7590 & n7594 ;
  assign n7596 = ~\u0_u0_csc_reg[15]/P0001  & ~n6381 ;
  assign n7597 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[15]_pad  ;
  assign n7598 = n6379 & n7597 ;
  assign n7599 = n6378 & n7598 ;
  assign n7600 = ~\u0_rst_r2_reg/NET0131  & ~n7599 ;
  assign n7601 = ~n7596 & n7600 ;
  assign n7602 = \u0_u0_tms_reg[30]/P0001  & ~n7457 ;
  assign n7603 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[30]_pad  ;
  assign n7604 = n6379 & n7603 ;
  assign n7605 = n6378 & n7604 ;
  assign n7606 = ~\u0_rst_r2_reg/NET0131  & ~n7605 ;
  assign n7607 = ~n7602 & n7606 ;
  assign n7608 = \u0_u0_tms_reg[3]/P0001  & ~n7457 ;
  assign n7609 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[3]_pad  ;
  assign n7610 = n6379 & n7609 ;
  assign n7611 = n6378 & n7610 ;
  assign n7612 = ~\u0_rst_r2_reg/NET0131  & ~n7611 ;
  assign n7613 = ~n7608 & n7612 ;
  assign n7614 = \u0_u0_tms_reg[4]/P0001  & ~n7457 ;
  assign n7615 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[4]_pad  ;
  assign n7616 = n6379 & n7615 ;
  assign n7617 = n6378 & n7616 ;
  assign n7618 = ~\u0_rst_r2_reg/NET0131  & ~n7617 ;
  assign n7619 = ~n7614 & n7618 ;
  assign n7620 = \u0_u0_tms_reg[5]/P0001  & ~n7457 ;
  assign n7621 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[5]_pad  ;
  assign n7622 = n6379 & n7621 ;
  assign n7623 = n6378 & n7622 ;
  assign n7624 = ~\u0_rst_r2_reg/NET0131  & ~n7623 ;
  assign n7625 = ~n7620 & n7624 ;
  assign n7626 = \u0_u0_tms_reg[6]/P0001  & ~n7457 ;
  assign n7627 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[6]_pad  ;
  assign n7628 = n6379 & n7627 ;
  assign n7629 = n6378 & n7628 ;
  assign n7630 = ~\u0_rst_r2_reg/NET0131  & ~n7629 ;
  assign n7631 = ~n7626 & n7630 ;
  assign n7632 = \u0_u0_tms_reg[7]/P0001  & ~n7457 ;
  assign n7633 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[7]_pad  ;
  assign n7634 = n6379 & n7633 ;
  assign n7635 = n6378 & n7634 ;
  assign n7636 = ~\u0_rst_r2_reg/NET0131  & ~n7635 ;
  assign n7637 = ~n7632 & n7636 ;
  assign n7638 = \u0_u0_tms_reg[8]/P0001  & ~n7457 ;
  assign n7639 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[8]_pad  ;
  assign n7640 = n6379 & n7639 ;
  assign n7641 = n6378 & n7640 ;
  assign n7642 = ~\u0_rst_r2_reg/NET0131  & ~n7641 ;
  assign n7643 = ~n7638 & n7642 ;
  assign n7644 = \u0_u0_tms_reg[9]/P0001  & ~n7457 ;
  assign n7645 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[9]_pad  ;
  assign n7646 = n6379 & n7645 ;
  assign n7647 = n6378 & n7646 ;
  assign n7648 = ~\u0_rst_r2_reg/NET0131  & ~n7647 ;
  assign n7649 = ~n7644 & n7648 ;
  assign n7650 = n6380 & n7346 ;
  assign n7651 = ~\u0_u1_csc_reg[0]/NET0131  & ~n7650 ;
  assign n7652 = n6384 & n7346 ;
  assign n7653 = ~\u0_rst_r2_reg/NET0131  & ~n7652 ;
  assign n7654 = ~n7651 & n7653 ;
  assign n7655 = ~\u0_u1_csc_reg[10]/P0001  & ~n7650 ;
  assign n7656 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[10]_pad  ;
  assign n7657 = n6379 & n7656 ;
  assign n7658 = n7346 & n7657 ;
  assign n7659 = ~\u0_rst_r2_reg/NET0131  & ~n7658 ;
  assign n7660 = ~n7655 & n7659 ;
  assign n7661 = ~\u0_u1_csc_reg[11]/P0001  & ~n7650 ;
  assign n7662 = n7336 & n7346 ;
  assign n7663 = ~\u0_rst_r2_reg/NET0131  & ~n7662 ;
  assign n7664 = ~n7661 & n7663 ;
  assign n7665 = ~\u0_u1_csc_reg[12]/P0001  & ~n7650 ;
  assign n7666 = n7342 & n7346 ;
  assign n7667 = ~\u0_rst_r2_reg/NET0131  & ~n7666 ;
  assign n7668 = ~n7665 & n7667 ;
  assign n7669 = ~\u0_u1_csc_reg[13]/P0001  & ~n7650 ;
  assign n7670 = n7346 & n7357 ;
  assign n7671 = ~\u0_rst_r2_reg/NET0131  & ~n7670 ;
  assign n7672 = ~n7669 & n7671 ;
  assign n7673 = ~\u0_u1_csc_reg[14]/P0001  & ~n7650 ;
  assign n7674 = n7346 & n7363 ;
  assign n7675 = ~\u0_rst_r2_reg/NET0131  & ~n7674 ;
  assign n7676 = ~n7673 & n7675 ;
  assign n7677 = ~\u0_u1_csc_reg[15]/P0001  & ~n7650 ;
  assign n7678 = n7346 & n7598 ;
  assign n7679 = ~\u0_rst_r2_reg/NET0131  & ~n7678 ;
  assign n7680 = ~n7677 & n7679 ;
  assign n7681 = ~\u0_u1_csc_reg[17]/P0001  & ~n7650 ;
  assign n7682 = n7346 & n7375 ;
  assign n7683 = ~\u0_rst_r2_reg/NET0131  & ~n7682 ;
  assign n7684 = ~n7681 & n7683 ;
  assign n7685 = ~\u0_u1_csc_reg[18]/P0001  & ~n7650 ;
  assign n7686 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[18]_pad  ;
  assign n7687 = n6379 & n7686 ;
  assign n7688 = n7346 & n7687 ;
  assign n7689 = ~\u0_rst_r2_reg/NET0131  & ~n7688 ;
  assign n7690 = ~n7685 & n7689 ;
  assign n7691 = ~\u0_u1_csc_reg[19]/P0001  & ~n7650 ;
  assign n7692 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[19]_pad  ;
  assign n7693 = n6379 & n7692 ;
  assign n7694 = n7346 & n7693 ;
  assign n7695 = ~\u0_rst_r2_reg/NET0131  & ~n7694 ;
  assign n7696 = ~n7691 & n7695 ;
  assign n7697 = ~\u0_u1_csc_reg[1]/NET0131  & ~n7650 ;
  assign n7698 = n7152 & n7346 ;
  assign n7699 = ~\u0_rst_r2_reg/NET0131  & ~n7698 ;
  assign n7700 = ~n7697 & n7699 ;
  assign n7701 = ~\u0_u1_csc_reg[20]/P0001  & ~n7650 ;
  assign n7702 = n7346 & n7381 ;
  assign n7703 = ~\u0_rst_r2_reg/NET0131  & ~n7702 ;
  assign n7704 = ~n7701 & n7703 ;
  assign n7705 = ~\u0_u0_csc_reg[29]/P0001  & ~n6381 ;
  assign n7706 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[29]_pad  ;
  assign n7707 = n6379 & n7706 ;
  assign n7708 = n6378 & n7707 ;
  assign n7709 = ~\u0_rst_r2_reg/NET0131  & ~n7708 ;
  assign n7710 = ~n7705 & n7709 ;
  assign n7711 = ~\u0_u1_csc_reg[22]/P0001  & ~n7650 ;
  assign n7712 = n7346 & n7393 ;
  assign n7713 = ~\u0_rst_r2_reg/NET0131  & ~n7712 ;
  assign n7714 = ~n7711 & n7713 ;
  assign n7715 = ~\u0_u1_csc_reg[23]/P0001  & ~n7650 ;
  assign n7716 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[23]_pad  ;
  assign n7717 = n6379 & n7716 ;
  assign n7718 = n7346 & n7717 ;
  assign n7719 = ~\u0_rst_r2_reg/NET0131  & ~n7718 ;
  assign n7720 = ~n7715 & n7719 ;
  assign n7721 = ~\u0_u1_csc_reg[21]/P0001  & ~n7650 ;
  assign n7722 = n7346 & n7387 ;
  assign n7723 = ~\u0_rst_r2_reg/NET0131  & ~n7722 ;
  assign n7724 = ~n7721 & n7723 ;
  assign n7725 = ~\u0_u1_csc_reg[24]/P0001  & ~n7650 ;
  assign n7726 = n7346 & n7399 ;
  assign n7727 = ~\u0_rst_r2_reg/NET0131  & ~n7726 ;
  assign n7728 = ~n7725 & n7727 ;
  assign n7729 = ~\u0_u1_csc_reg[25]/P0001  & ~n7650 ;
  assign n7730 = n7346 & n7441 ;
  assign n7731 = ~\u0_rst_r2_reg/NET0131  & ~n7730 ;
  assign n7732 = ~n7729 & n7731 ;
  assign n7733 = ~\u0_u1_csc_reg[26]/P0001  & ~n7650 ;
  assign n7734 = n7346 & n7405 ;
  assign n7735 = ~\u0_rst_r2_reg/NET0131  & ~n7734 ;
  assign n7736 = ~n7733 & n7735 ;
  assign n7737 = ~\u0_u1_csc_reg[27]/P0001  & ~n7650 ;
  assign n7738 = n7346 & n7411 ;
  assign n7739 = ~\u0_rst_r2_reg/NET0131  & ~n7738 ;
  assign n7740 = ~n7737 & n7739 ;
  assign n7741 = ~\u0_u1_csc_reg[28]/P0001  & ~n7650 ;
  assign n7742 = n7346 & n7417 ;
  assign n7743 = ~\u0_rst_r2_reg/NET0131  & ~n7742 ;
  assign n7744 = ~n7741 & n7743 ;
  assign n7745 = ~\u0_u0_csc_reg[7]/P0001  & ~n6381 ;
  assign n7746 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[7]_pad  ;
  assign n7747 = n6379 & n7746 ;
  assign n7748 = n6378 & n7747 ;
  assign n7749 = ~\u0_rst_r2_reg/NET0131  & ~n7748 ;
  assign n7750 = ~n7745 & n7749 ;
  assign n7751 = ~\u0_u1_csc_reg[29]/P0001  & ~n7650 ;
  assign n7752 = n7346 & n7707 ;
  assign n7753 = ~\u0_rst_r2_reg/NET0131  & ~n7752 ;
  assign n7754 = ~n7751 & n7753 ;
  assign n7755 = ~\u0_u1_csc_reg[2]/NET0131  & ~n7650 ;
  assign n7756 = n7159 & n7346 ;
  assign n7757 = ~\u0_rst_r2_reg/NET0131  & ~n7756 ;
  assign n7758 = ~n7755 & n7757 ;
  assign n7759 = ~\u0_u1_csc_reg[30]/P0001  & ~n7650 ;
  assign n7760 = n7346 & n7429 ;
  assign n7761 = ~\u0_rst_r2_reg/NET0131  & ~n7760 ;
  assign n7762 = ~n7759 & n7761 ;
  assign n7763 = ~\u0_u1_csc_reg[31]/P0001  & ~n7650 ;
  assign n7764 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[31]_pad  ;
  assign n7765 = n6379 & n7764 ;
  assign n7766 = n7346 & n7765 ;
  assign n7767 = ~\u0_rst_r2_reg/NET0131  & ~n7766 ;
  assign n7768 = ~n7763 & n7767 ;
  assign n7769 = ~\u0_u1_csc_reg[4]/P0001  & ~n7650 ;
  assign n7770 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[4]_pad  ;
  assign n7771 = n6379 & n7770 ;
  assign n7772 = n7346 & n7771 ;
  assign n7773 = ~\u0_rst_r2_reg/NET0131  & ~n7772 ;
  assign n7774 = ~n7769 & n7773 ;
  assign n7775 = ~\u0_u1_csc_reg[3]/NET0131  & ~n7650 ;
  assign n7776 = n7346 & n7435 ;
  assign n7777 = ~\u0_rst_r2_reg/NET0131  & ~n7776 ;
  assign n7778 = ~n7775 & n7777 ;
  assign n7779 = ~\u0_u1_csc_reg[5]/P0001  & ~n7650 ;
  assign n7780 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[5]_pad  ;
  assign n7781 = n6379 & n7780 ;
  assign n7782 = n7346 & n7781 ;
  assign n7783 = ~\u0_rst_r2_reg/NET0131  & ~n7782 ;
  assign n7784 = ~n7779 & n7783 ;
  assign n7785 = ~\u0_u1_csc_reg[6]/P0001  & ~n7650 ;
  assign n7786 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[6]_pad  ;
  assign n7787 = n6379 & n7786 ;
  assign n7788 = n7346 & n7787 ;
  assign n7789 = ~\u0_rst_r2_reg/NET0131  & ~n7788 ;
  assign n7790 = ~n7785 & n7789 ;
  assign n7791 = ~\u0_u0_csc_reg[8]/P0001  & ~n6381 ;
  assign n7792 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[8]_pad  ;
  assign n7793 = n6379 & n7792 ;
  assign n7794 = n6378 & n7793 ;
  assign n7795 = ~\u0_rst_r2_reg/NET0131  & ~n7794 ;
  assign n7796 = ~n7791 & n7795 ;
  assign n7797 = ~\u0_u1_csc_reg[8]/P0001  & ~n7650 ;
  assign n7798 = n7346 & n7793 ;
  assign n7799 = ~\u0_rst_r2_reg/NET0131  & ~n7798 ;
  assign n7800 = ~n7797 & n7799 ;
  assign n7801 = ~\u0_u1_csc_reg[7]/P0001  & ~n7650 ;
  assign n7802 = n7346 & n7747 ;
  assign n7803 = ~\u0_rst_r2_reg/NET0131  & ~n7802 ;
  assign n7804 = ~n7801 & n7803 ;
  assign n7805 = ~\u0_u1_csc_reg[9]/P0001  & ~n7650 ;
  assign n7806 = ~\u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[9]_pad  ;
  assign n7807 = n6379 & n7806 ;
  assign n7808 = n7346 & n7807 ;
  assign n7809 = ~\u0_rst_r2_reg/NET0131  & ~n7808 ;
  assign n7810 = ~n7805 & n7809 ;
  assign n7811 = ~\u0_u1_tms_reg[0]/P0001  & ~n7348 ;
  assign n7812 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[0]_pad  ;
  assign n7813 = n6379 & n7812 ;
  assign n7814 = n7346 & n7813 ;
  assign n7815 = ~\u0_rst_r2_reg/NET0131  & ~n7814 ;
  assign n7816 = ~n7811 & n7815 ;
  assign n7817 = ~\u0_u1_tms_reg[30]/P0001  & ~n7348 ;
  assign n7818 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[30]_pad  ;
  assign n7819 = n6379 & n7818 ;
  assign n7820 = n7346 & n7819 ;
  assign n7821 = ~\u0_rst_r2_reg/NET0131  & ~n7820 ;
  assign n7822 = ~n7817 & n7821 ;
  assign n7823 = ~\u0_u1_tms_reg[10]/P0001  & ~n7348 ;
  assign n7824 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[10]_pad  ;
  assign n7825 = n6379 & n7824 ;
  assign n7826 = n7346 & n7825 ;
  assign n7827 = ~\u0_rst_r2_reg/NET0131  & ~n7826 ;
  assign n7828 = ~n7823 & n7827 ;
  assign n7829 = ~\u0_u1_tms_reg[11]/P0001  & ~n7348 ;
  assign n7830 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[11]_pad  ;
  assign n7831 = n6379 & n7830 ;
  assign n7832 = n7346 & n7831 ;
  assign n7833 = ~\u0_rst_r2_reg/NET0131  & ~n7832 ;
  assign n7834 = ~n7829 & n7833 ;
  assign n7835 = ~\u0_u1_tms_reg[12]/P0001  & ~n7348 ;
  assign n7836 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[12]_pad  ;
  assign n7837 = n6379 & n7836 ;
  assign n7838 = n7346 & n7837 ;
  assign n7839 = ~\u0_rst_r2_reg/NET0131  & ~n7838 ;
  assign n7840 = ~n7835 & n7839 ;
  assign n7841 = ~\u0_u1_tms_reg[13]/P0001  & ~n7348 ;
  assign n7842 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[13]_pad  ;
  assign n7843 = n6379 & n7842 ;
  assign n7844 = n7346 & n7843 ;
  assign n7845 = ~\u0_rst_r2_reg/NET0131  & ~n7844 ;
  assign n7846 = ~n7841 & n7845 ;
  assign n7847 = ~\u0_u1_tms_reg[14]/P0001  & ~n7348 ;
  assign n7848 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[14]_pad  ;
  assign n7849 = n6379 & n7848 ;
  assign n7850 = n7346 & n7849 ;
  assign n7851 = ~\u0_rst_r2_reg/NET0131  & ~n7850 ;
  assign n7852 = ~n7847 & n7851 ;
  assign n7853 = ~\u0_u1_tms_reg[15]/P0001  & ~n7348 ;
  assign n7854 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[15]_pad  ;
  assign n7855 = n6379 & n7854 ;
  assign n7856 = n7346 & n7855 ;
  assign n7857 = ~\u0_rst_r2_reg/NET0131  & ~n7856 ;
  assign n7858 = ~n7853 & n7857 ;
  assign n7859 = ~\u0_u1_tms_reg[18]/P0001  & ~n7348 ;
  assign n7860 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[18]_pad  ;
  assign n7861 = n6379 & n7860 ;
  assign n7862 = n7346 & n7861 ;
  assign n7863 = ~\u0_rst_r2_reg/NET0131  & ~n7862 ;
  assign n7864 = ~n7859 & n7863 ;
  assign n7865 = ~\u0_u1_tms_reg[20]/P0001  & ~n7348 ;
  assign n7866 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[20]_pad  ;
  assign n7867 = n6379 & n7866 ;
  assign n7868 = n7346 & n7867 ;
  assign n7869 = ~\u0_rst_r2_reg/NET0131  & ~n7868 ;
  assign n7870 = ~n7865 & n7869 ;
  assign n7871 = ~\u0_u1_tms_reg[21]/P0001  & ~n7348 ;
  assign n7872 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[21]_pad  ;
  assign n7873 = n6379 & n7872 ;
  assign n7874 = n7346 & n7873 ;
  assign n7875 = ~\u0_rst_r2_reg/NET0131  & ~n7874 ;
  assign n7876 = ~n7871 & n7875 ;
  assign n7877 = ~\u0_u1_tms_reg[24]/P0001  & ~n7348 ;
  assign n7878 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[24]_pad  ;
  assign n7879 = n6379 & n7878 ;
  assign n7880 = n7346 & n7879 ;
  assign n7881 = ~\u0_rst_r2_reg/NET0131  & ~n7880 ;
  assign n7882 = ~n7877 & n7881 ;
  assign n7883 = ~\u0_u1_tms_reg[25]/P0001  & ~n7348 ;
  assign n7884 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[25]_pad  ;
  assign n7885 = n6379 & n7884 ;
  assign n7886 = n7346 & n7885 ;
  assign n7887 = ~\u0_rst_r2_reg/NET0131  & ~n7886 ;
  assign n7888 = ~n7883 & n7887 ;
  assign n7889 = ~\u0_u1_tms_reg[27]/P0001  & ~n7348 ;
  assign n7890 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[27]_pad  ;
  assign n7891 = n6379 & n7890 ;
  assign n7892 = n7346 & n7891 ;
  assign n7893 = ~\u0_rst_r2_reg/NET0131  & ~n7892 ;
  assign n7894 = ~n7889 & n7893 ;
  assign n7895 = ~\u0_u1_tms_reg[2]/P0001  & ~n7348 ;
  assign n7896 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[2]_pad  ;
  assign n7897 = n6379 & n7896 ;
  assign n7898 = n7346 & n7897 ;
  assign n7899 = ~\u0_rst_r2_reg/NET0131  & ~n7898 ;
  assign n7900 = ~n7895 & n7899 ;
  assign n7901 = ~\u0_u1_tms_reg[31]/P0001  & ~n7348 ;
  assign n7902 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[31]_pad  ;
  assign n7903 = n6379 & n7902 ;
  assign n7904 = n7346 & n7903 ;
  assign n7905 = ~\u0_rst_r2_reg/NET0131  & ~n7904 ;
  assign n7906 = ~n7901 & n7905 ;
  assign n7907 = ~\u0_u0_csc_reg[23]/P0001  & ~n6381 ;
  assign n7908 = n6378 & n7717 ;
  assign n7909 = ~\u0_rst_r2_reg/NET0131  & ~n7908 ;
  assign n7910 = ~n7907 & n7909 ;
  assign n7911 = ~\u0_u1_tms_reg[3]/P0001  & ~n7348 ;
  assign n7912 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[3]_pad  ;
  assign n7913 = n6379 & n7912 ;
  assign n7914 = n7346 & n7913 ;
  assign n7915 = ~\u0_rst_r2_reg/NET0131  & ~n7914 ;
  assign n7916 = ~n7911 & n7915 ;
  assign n7917 = ~\u0_u1_tms_reg[5]/P0001  & ~n7348 ;
  assign n7918 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[5]_pad  ;
  assign n7919 = n6379 & n7918 ;
  assign n7920 = n7346 & n7919 ;
  assign n7921 = ~\u0_rst_r2_reg/NET0131  & ~n7920 ;
  assign n7922 = ~n7917 & n7921 ;
  assign n7923 = ~\u0_u1_tms_reg[8]/P0001  & ~n7348 ;
  assign n7924 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[8]_pad  ;
  assign n7925 = n6379 & n7924 ;
  assign n7926 = n7346 & n7925 ;
  assign n7927 = ~\u0_rst_r2_reg/NET0131  & ~n7926 ;
  assign n7928 = ~n7923 & n7927 ;
  assign n7929 = ~\u0_u1_tms_reg[9]/P0001  & ~n7348 ;
  assign n7930 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[9]_pad  ;
  assign n7931 = n6379 & n7930 ;
  assign n7932 = n7346 & n7931 ;
  assign n7933 = ~\u0_rst_r2_reg/NET0131  & ~n7932 ;
  assign n7934 = ~n7929 & n7933 ;
  assign n7935 = \u0_u0_tms_reg[20]/P0001  & ~n7457 ;
  assign n7936 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[20]_pad  ;
  assign n7937 = n6379 & n7936 ;
  assign n7938 = n6378 & n7937 ;
  assign n7939 = ~\u0_rst_r2_reg/NET0131  & ~n7938 ;
  assign n7940 = ~n7935 & n7939 ;
  assign n7941 = ~\u0_u1_tms_reg[1]/P0001  & ~n7348 ;
  assign n7942 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[1]_pad  ;
  assign n7943 = n6379 & n7942 ;
  assign n7944 = n7346 & n7943 ;
  assign n7945 = ~\u0_rst_r2_reg/NET0131  & ~n7944 ;
  assign n7946 = ~n7941 & n7945 ;
  assign n7947 = ~\u0_u1_tms_reg[6]/P0001  & ~n7348 ;
  assign n7948 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[6]_pad  ;
  assign n7949 = n6379 & n7948 ;
  assign n7950 = n7346 & n7949 ;
  assign n7951 = ~\u0_rst_r2_reg/NET0131  & ~n7950 ;
  assign n7952 = ~n7947 & n7951 ;
  assign n7953 = ~\u0_u1_tms_reg[29]/P0001  & ~n7348 ;
  assign n7954 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[29]_pad  ;
  assign n7955 = n6379 & n7954 ;
  assign n7956 = n7346 & n7955 ;
  assign n7957 = ~\u0_rst_r2_reg/NET0131  & ~n7956 ;
  assign n7958 = ~n7953 & n7957 ;
  assign n7959 = ~\u0_u1_tms_reg[28]/P0001  & ~n7348 ;
  assign n7960 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[28]_pad  ;
  assign n7961 = n6379 & n7960 ;
  assign n7962 = n7346 & n7961 ;
  assign n7963 = ~\u0_rst_r2_reg/NET0131  & ~n7962 ;
  assign n7964 = ~n7959 & n7963 ;
  assign n7965 = ~\u0_u1_tms_reg[4]/P0001  & ~n7348 ;
  assign n7966 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[4]_pad  ;
  assign n7967 = n6379 & n7966 ;
  assign n7968 = n7346 & n7967 ;
  assign n7969 = ~\u0_rst_r2_reg/NET0131  & ~n7968 ;
  assign n7970 = ~n7965 & n7969 ;
  assign n7971 = ~\u0_u0_csc_reg[10]/P0001  & ~n6381 ;
  assign n7972 = n6378 & n7657 ;
  assign n7973 = ~\u0_rst_r2_reg/NET0131  & ~n7972 ;
  assign n7974 = ~n7971 & n7973 ;
  assign n7975 = ~\u0_u1_tms_reg[26]/P0001  & ~n7348 ;
  assign n7976 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[26]_pad  ;
  assign n7977 = n6379 & n7976 ;
  assign n7978 = n7346 & n7977 ;
  assign n7979 = ~\u0_rst_r2_reg/NET0131  & ~n7978 ;
  assign n7980 = ~n7975 & n7979 ;
  assign n7981 = ~\u0_u1_csc_reg[16]/P0001  & ~n7650 ;
  assign n7982 = n7346 & n7369 ;
  assign n7983 = ~\u0_rst_r2_reg/NET0131  & ~n7982 ;
  assign n7984 = ~n7981 & n7983 ;
  assign n7985 = ~\u0_u0_csc_reg[18]/P0001  & ~n6381 ;
  assign n7986 = n6378 & n7687 ;
  assign n7987 = ~\u0_rst_r2_reg/NET0131  & ~n7986 ;
  assign n7988 = ~n7985 & n7987 ;
  assign n7989 = ~\u0_u0_csc_reg[31]/P0001  & ~n6381 ;
  assign n7990 = n6378 & n7765 ;
  assign n7991 = ~\u0_rst_r2_reg/NET0131  & ~n7990 ;
  assign n7992 = ~n7989 & n7991 ;
  assign n7993 = \u0_u0_tms_reg[31]/P0001  & ~n7457 ;
  assign n7994 = \u0_u0_addr_r_reg[2]/P0001  & \wb_data_i[31]_pad  ;
  assign n7995 = n6379 & n7994 ;
  assign n7996 = n6378 & n7995 ;
  assign n7997 = ~\u0_rst_r2_reg/NET0131  & ~n7996 ;
  assign n7998 = ~n7993 & n7997 ;
  assign n7999 = ~\u0_u1_tms_reg[7]/P0001  & ~n7348 ;
  assign n8000 = \u0_u0_addr_r_reg[2]/P0001  & ~\wb_data_i[7]_pad  ;
  assign n8001 = n6379 & n8000 ;
  assign n8002 = n7346 & n8001 ;
  assign n8003 = ~\u0_rst_r2_reg/NET0131  & ~n8002 ;
  assign n8004 = ~n7999 & n8003 ;
  assign n8005 = ~\u0_u0_csc_reg[19]/P0001  & ~n6381 ;
  assign n8006 = n6378 & n7693 ;
  assign n8007 = ~\u0_rst_r2_reg/NET0131  & ~n8006 ;
  assign n8008 = ~n8005 & n8007 ;
  assign n8009 = ~\u0_u0_csc_reg[6]/P0001  & ~n6381 ;
  assign n8010 = n6378 & n7787 ;
  assign n8011 = ~\u0_rst_r2_reg/NET0131  & ~n8010 ;
  assign n8012 = ~n8009 & n8011 ;
  assign n8013 = ~\u0_u0_csc_reg[9]/P0001  & ~n6381 ;
  assign n8014 = n6378 & n7807 ;
  assign n8015 = ~\u0_rst_r2_reg/NET0131  & ~n8014 ;
  assign n8016 = ~n8013 & n8015 ;
  assign n8017 = \u1_acs_addr_reg[2]/P0001  & n5141 ;
  assign n8018 = ~\u1_acs_addr_reg[3]/P0001  & ~n8017 ;
  assign n8019 = ~n5143 & ~n8018 ;
  assign n8020 = ~\u0_u1_inited_reg/NET0131  & ~n6840 ;
  assign n8021 = ~\u0_u0_inited_reg/NET0131  & ~n6834 ;
  assign n8022 = n983 & n6832 ;
  assign n8023 = ~n5640 & ~n6545 ;
  assign n8024 = ~n8022 & n8023 ;
  assign n8025 = ~n1048 & n1234 ;
  assign n8026 = n1231 & n2191 ;
  assign n8027 = ~\u6_read_go_r_reg/NET0131  & ~n8026 ;
  assign n8028 = n8025 & ~n8027 ;
  assign n8029 = ~n3350 & ~n3352 ;
  assign n8030 = ~\u1_acs_addr_reg[9]/P0001  & ~n6313 ;
  assign n8031 = ~n5149 & ~n8030 ;
  assign n8032 = \wb_data_i[11]_pad  & ~\wb_data_i[13]_pad  ;
  assign n8033 = ~\wb_data_i[11]_pad  & \wb_data_i[13]_pad  ;
  assign n8034 = ~n8032 & ~n8033 ;
  assign n8035 = ~\wb_data_i[15]_pad  & ~\wb_data_i[8]_pad  ;
  assign n8036 = \wb_data_i[15]_pad  & \wb_data_i[8]_pad  ;
  assign n8037 = ~n8035 & ~n8036 ;
  assign n8038 = \wb_data_i[9]_pad  & n8037 ;
  assign n8039 = ~\wb_data_i[9]_pad  & ~n8037 ;
  assign n8040 = ~n8038 & ~n8039 ;
  assign n8041 = \wb_data_i[10]_pad  & ~\wb_data_i[12]_pad  ;
  assign n8042 = ~\wb_data_i[10]_pad  & \wb_data_i[12]_pad  ;
  assign n8043 = ~n8041 & ~n8042 ;
  assign n8044 = \wb_data_i[14]_pad  & n8043 ;
  assign n8045 = ~\wb_data_i[14]_pad  & ~n8043 ;
  assign n8046 = ~n8044 & ~n8045 ;
  assign n8047 = n8040 & ~n8046 ;
  assign n8048 = ~n8040 & n8046 ;
  assign n8049 = ~n8047 & ~n8048 ;
  assign n8050 = n8034 & n8049 ;
  assign n8051 = ~n8034 & ~n8049 ;
  assign n8052 = ~n8050 & ~n8051 ;
  assign n8053 = \wb_data_i[1]_pad  & ~\wb_data_i[6]_pad  ;
  assign n8054 = ~\wb_data_i[1]_pad  & \wb_data_i[6]_pad  ;
  assign n8055 = ~n8053 & ~n8054 ;
  assign n8056 = ~\wb_data_i[2]_pad  & ~\wb_data_i[4]_pad  ;
  assign n8057 = \wb_data_i[2]_pad  & \wb_data_i[4]_pad  ;
  assign n8058 = ~n8056 & ~n8057 ;
  assign n8059 = \wb_data_i[5]_pad  & n8058 ;
  assign n8060 = ~\wb_data_i[5]_pad  & ~n8058 ;
  assign n8061 = ~n8059 & ~n8060 ;
  assign n8062 = \wb_data_i[0]_pad  & ~\wb_data_i[7]_pad  ;
  assign n8063 = ~\wb_data_i[0]_pad  & \wb_data_i[7]_pad  ;
  assign n8064 = ~n8062 & ~n8063 ;
  assign n8065 = \wb_data_i[3]_pad  & n8064 ;
  assign n8066 = ~\wb_data_i[3]_pad  & ~n8064 ;
  assign n8067 = ~n8065 & ~n8066 ;
  assign n8068 = n8061 & ~n8067 ;
  assign n8069 = ~n8061 & n8067 ;
  assign n8070 = ~n8068 & ~n8069 ;
  assign n8071 = n8055 & n8070 ;
  assign n8072 = ~n8055 & ~n8070 ;
  assign n8073 = ~n8071 & ~n8072 ;
  assign n8074 = \wb_data_i[27]_pad  & ~\wb_data_i[29]_pad  ;
  assign n8075 = ~\wb_data_i[27]_pad  & \wb_data_i[29]_pad  ;
  assign n8076 = ~n8074 & ~n8075 ;
  assign n8077 = ~\wb_data_i[24]_pad  & ~\wb_data_i[31]_pad  ;
  assign n8078 = \wb_data_i[24]_pad  & \wb_data_i[31]_pad  ;
  assign n8079 = ~n8077 & ~n8078 ;
  assign n8080 = \wb_data_i[30]_pad  & n8079 ;
  assign n8081 = ~\wb_data_i[30]_pad  & ~n8079 ;
  assign n8082 = ~n8080 & ~n8081 ;
  assign n8083 = \wb_data_i[26]_pad  & ~\wb_data_i[28]_pad  ;
  assign n8084 = ~\wb_data_i[26]_pad  & \wb_data_i[28]_pad  ;
  assign n8085 = ~n8083 & ~n8084 ;
  assign n8086 = \wb_data_i[25]_pad  & n8085 ;
  assign n8087 = ~\wb_data_i[25]_pad  & ~n8085 ;
  assign n8088 = ~n8086 & ~n8087 ;
  assign n8089 = n8082 & ~n8088 ;
  assign n8090 = ~n8082 & n8088 ;
  assign n8091 = ~n8089 & ~n8090 ;
  assign n8092 = n8076 & n8091 ;
  assign n8093 = ~n8076 & ~n8091 ;
  assign n8094 = ~n8092 & ~n8093 ;
  assign n8095 = \wb_data_i[17]_pad  & ~\wb_data_i[22]_pad  ;
  assign n8096 = ~\wb_data_i[17]_pad  & \wb_data_i[22]_pad  ;
  assign n8097 = ~n8095 & ~n8096 ;
  assign n8098 = ~\wb_data_i[16]_pad  & ~\wb_data_i[23]_pad  ;
  assign n8099 = \wb_data_i[16]_pad  & \wb_data_i[23]_pad  ;
  assign n8100 = ~n8098 & ~n8099 ;
  assign n8101 = \wb_data_i[21]_pad  & n8100 ;
  assign n8102 = ~\wb_data_i[21]_pad  & ~n8100 ;
  assign n8103 = ~n8101 & ~n8102 ;
  assign n8104 = \wb_data_i[18]_pad  & ~\wb_data_i[20]_pad  ;
  assign n8105 = ~\wb_data_i[18]_pad  & \wb_data_i[20]_pad  ;
  assign n8106 = ~n8104 & ~n8105 ;
  assign n8107 = \wb_data_i[19]_pad  & n8106 ;
  assign n8108 = ~\wb_data_i[19]_pad  & ~n8106 ;
  assign n8109 = ~n8107 & ~n8108 ;
  assign n8110 = n8103 & ~n8109 ;
  assign n8111 = ~n8103 & n8109 ;
  assign n8112 = ~n8110 & ~n8111 ;
  assign n8113 = n8097 & n8112 ;
  assign n8114 = ~n8097 & ~n8112 ;
  assign n8115 = ~n8113 & ~n8114 ;
  assign n8116 = \u6_write_go_r_reg/NET0131  & wb_cyc_i_pad ;
  assign n8117 = wb_cyc_i_pad & n2165 ;
  assign n8118 = n2191 & n8117 ;
  assign n8119 = ~n8116 & ~n8118 ;
  assign n8120 = ~\u0_init_req_reg/NET0131  & ~\u0_u1_lmr_req_reg/NET0131  ;
  assign n8121 = \u0_init_req_reg/NET0131  & ~\u0_u1_init_req_reg/NET0131  ;
  assign n8122 = ~n8120 & ~n8121 ;
  assign n8123 = \u0_sreq_cs_le_reg/NET0131  & ~n8122 ;
  assign n8124 = ~\u0_spec_req_cs_reg[1]/NET0131  & ~\u0_sreq_cs_le_reg/NET0131  ;
  assign n8125 = \u0_init_req_reg/NET0131  & ~\u0_u0_init_req_reg/NET0131  ;
  assign n8126 = ~\u0_init_req_reg/NET0131  & ~\u0_u0_lmr_req_reg/NET0131  ;
  assign n8127 = \u0_sreq_cs_le_reg/NET0131  & ~n8126 ;
  assign n8128 = ~n8125 & n8127 ;
  assign n8129 = ~n8124 & ~n8128 ;
  assign n8130 = ~n8123 & n8129 ;
  assign n8131 = ~\u1_acs_addr_reg[2]/P0001  & ~n5141 ;
  assign n8132 = ~n8017 & ~n8131 ;
  assign n8133 = ~\u1_acs_addr_reg[5]/P0001  & ~n6335 ;
  assign n8134 = ~n7165 & ~n8133 ;
  assign n8135 = ~suspended_o_pad & ~\u0_csr_r_reg[2]/NET0131  ;
  assign n8136 = ~\u0_rf_we_reg/NET0131  & wb_we_i_pad ;
  assign n8137 = n1045 & n8136 ;
  assign n8138 = n2589 & n8137 ;
  assign n8139 = \u5_lookup_ready1_reg/NET0131  & n1045 ;
  assign n8140 = \u0_rf_we_reg/NET0131  & ~\u0_u0_addr_r_reg[2]/P0001  ;
  assign n8141 = ~\u0_u0_addr_r_reg[4]/P0001  & n8140 ;
  assign n8142 = n6378 & n8141 ;
  assign n8143 = n7346 & n8141 ;
  assign n8144 = \u0_spec_req_cs_reg[0]/NET0131  & ~\u0_sreq_cs_le_reg/NET0131  ;
  assign n8145 = ~n8128 & ~n8144 ;
  assign n8146 = ~\mem_ack_r_reg/P0001  & ~\u0_csc_reg[1]/NET0131  ;
  assign n8147 = n6392 & n8146 ;
  assign n8148 = ~\u5_state_reg[26]/NET0131  & n983 ;
  assign n8149 = ~n1838 & ~n1917 ;
  assign n8150 = \u6_wr_hold_reg/NET0131  & ~n1045 ;
  assign n8151 = ~n1046 & ~n8150 ;
  assign n8152 = ~\u1_acs_addr_reg[0]/P0001  & ~\u1_acs_addr_reg[1]/P0001  ;
  assign n8153 = ~n5141 & ~n8152 ;
  assign n8154 = \u6_rmw_en_reg/NET0131  & wb_cyc_i_pad ;
  assign n8155 = ~wb_ack_o_pad & ~n8154 ;
  assign n8156 = \u5_cmd_asserted_reg/NET0131  & ~\u5_mc_le_reg/NET0131  ;
  assign n8157 = \u5_cmd_asserted2_reg/NET0131  & \u5_mc_le_reg/NET0131  ;
  assign n8158 = ~n8156 & ~n8157 ;
  assign n8159 = ~\u0_u0_lmr_req_reg/NET0131  & ~\u0_u1_lmr_req_reg/NET0131  ;
  assign n8160 = ~\u0_u0_init_req_reg/NET0131  & ~\u0_u1_init_req_reg/NET0131  ;
  assign n8161 = ~\u5_state_reg[1]/NET0131  & ~\u5_state_reg[54]/NET0131  ;
  assign n8162 = \u5_state_reg[1]/NET0131  & \u5_state_reg[54]/NET0131  ;
  assign n8163 = ~n8161 & ~n8162 ;
  assign n8164 = ~n1144 & ~n1320 ;
  assign n8165 = ~\u5_state_reg[0]/NET0131  & n1007 ;
  assign n8166 = ~n8164 & n8165 ;
  assign n8167 = n1052 & n8166 ;
  assign n8168 = ~n1069 & ~n8167 ;
  assign n8169 = ~\u5_state_reg[46]/NET0131  & ~n1378 ;
  assign n8170 = ~n1390 & n8169 ;
  assign n8171 = ~\u5_state_reg[49]/NET0131  & n969 ;
  assign n8172 = \u5_state_reg[46]/NET0131  & ~n1383 ;
  assign n8173 = n8171 & ~n8172 ;
  assign n8174 = ~n8170 & n8173 ;
  assign n8175 = n1306 & n8174 ;
  assign n8176 = n1380 & n8175 ;
  assign n8177 = ~n1108 & ~n1345 ;
  assign n8178 = n1011 & ~n8177 ;
  assign n8179 = ~n1150 & ~n1360 ;
  assign n8180 = n1007 & ~n8179 ;
  assign n8181 = n1294 & n8180 ;
  assign n8182 = ~n8178 & ~n8181 ;
  assign n8183 = n1028 & n1383 ;
  assign n8184 = n3701 & n8183 ;
  assign n8185 = n1380 & n8184 ;
  assign n8186 = ~n8182 & n8185 ;
  assign n8187 = ~n8176 & ~n8186 ;
  assign n8188 = ~n1357 & n1379 ;
  assign n8189 = ~n1385 & ~n1393 ;
  assign n8190 = n961 & ~n8189 ;
  assign n8191 = ~n8188 & ~n8190 ;
  assign n8192 = n971 & n1029 ;
  assign n8193 = n1011 & n1383 ;
  assign n8194 = n8192 & n8193 ;
  assign n8195 = ~n8191 & n8194 ;
  assign n8196 = ~n8167 & ~n8195 ;
  assign n8197 = n8187 & n8196 ;
  assign n8198 = ~n8168 & ~n8197 ;
  assign n8199 = n6822 & ~n8163 ;
  assign n8200 = n5628 & n8199 ;
  assign n8201 = n8198 & n8200 ;
  assign n8202 = ~n8163 & ~n8201 ;
  assign n8203 = ~\u5_state_reg[1]/NET0131  & n1897 ;
  assign n8204 = ~n1966 & n8203 ;
  assign n8205 = ~n1954 & n8204 ;
  assign n8206 = ~\u4_rfr_req_reg/NET0131  & ~\u5_state_reg[54]/NET0131  ;
  assign n8207 = n1905 & n8206 ;
  assign n8208 = n1998 & n8207 ;
  assign n8209 = ~n8201 & ~n8208 ;
  assign n8210 = ~n8205 & n8209 ;
  assign n8211 = ~n8202 & ~n8210 ;
  assign n8212 = ~\u5_cmd_asserted_reg/NET0131  & ~\u5_state_reg[10]/NET0131  ;
  assign n8213 = n1184 & ~n8212 ;
  assign n8214 = ~\u5_tmr_done_reg/NET0131  & n1138 ;
  assign n8215 = n1036 & n8214 ;
  assign n8216 = ~n8213 & ~n8215 ;
  assign n8217 = \u5_tmr_done_reg/NET0131  & n1331 ;
  assign n8218 = ~\u5_cmd_asserted_reg/NET0131  & n1135 ;
  assign n8219 = ~n8217 & ~n8218 ;
  assign n8220 = ~\u5_tmr_done_reg/NET0131  & n1373 ;
  assign n8221 = ~n5711 & ~n8220 ;
  assign n8222 = ~\u5_cmd_asserted_reg/NET0131  & n1455 ;
  assign n8223 = n1096 & n8222 ;
  assign n8224 = n1078 & n8223 ;
  assign n8225 = ~n1171 & ~n8224 ;
  assign n8226 = \u5_state_reg[26]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n8227 = ~n3336 & ~n8226 ;
  assign n8228 = n1373 & ~n8227 ;
  assign n8229 = ~\u5_cmd_asserted_reg/NET0131  & n1265 ;
  assign n8230 = ~n8228 & ~n8229 ;
  assign n8231 = ~\u5_state_reg[38]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n8232 = \u5_tmr2_done_reg/NET0131  & ~n2739 ;
  assign n8233 = ~n2736 & n8232 ;
  assign n8234 = ~n8231 & ~n8233 ;
  assign n8235 = n1323 & n8234 ;
  assign n8236 = n1532 & ~n1537 ;
  assign n8237 = ~n1904 & n8236 ;
  assign n8238 = n1922 & n8237 ;
  assign n8239 = \u5_state_reg[36]/NET0131  & n1922 ;
  assign n8240 = ~n2809 & n8239 ;
  assign n8241 = ~n8238 & ~n8240 ;
  assign n8242 = \u5_state_reg[36]/NET0131  & ~n2811 ;
  assign n8243 = ~n1922 & n8242 ;
  assign n8244 = n8241 & ~n8243 ;
  assign n8245 = n1929 & ~n8244 ;
  assign n8246 = ~\u5_cmd_asserted_reg/NET0131  & n1249 ;
  assign n8247 = n1248 & n8246 ;
  assign n8248 = \u5_state_reg[13]/NET0131  & ~n3158 ;
  assign n8249 = ~n1431 & ~n8248 ;
  assign n8250 = n1193 & ~n8249 ;
  assign n8251 = ~n1238 & ~n8250 ;
  assign n8252 = ~n8247 & n8251 ;
  assign n8253 = n3858 & n5395 ;
  assign n8254 = n1308 & n8253 ;
  assign n8255 = ~\u5_cmd_asserted_reg/NET0131  & n1453 ;
  assign n8256 = ~n8254 & ~n8255 ;
  assign n8257 = ~\u5_cmd_asserted_reg/NET0131  & ~\u5_state_reg[28]/NET0131  ;
  assign n8258 = n1462 & ~n8257 ;
  assign n8259 = \u5_state_reg[28]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n8260 = ~n3124 & n8259 ;
  assign n8261 = ~n8258 & ~n8260 ;
  assign n8262 = ~\u5_cmd_asserted_reg/NET0131  & ~\u5_state_reg[30]/NET0131  ;
  assign n8263 = n1135 & ~n8262 ;
  assign n8264 = ~\u5_resume_req_r_reg/NET0131  & n1104 ;
  assign n8265 = ~n8263 & ~n8264 ;
  assign n8266 = n1929 & ~n2810 ;
  assign n8267 = ~\u5_state_reg[33]/NET0131  & ~n2812 ;
  assign n8268 = n8266 & ~n8267 ;
  assign n8269 = ~\u5_cmd_asserted_reg/NET0131  & n1462 ;
  assign n8270 = ~n6182 & ~n8269 ;
  assign n8271 = \u5_state_reg[32]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n8272 = ~n3559 & n8271 ;
  assign n8273 = ~n1327 & ~n8272 ;
  assign n8274 = n1309 & n1995 ;
  assign n8275 = n1308 & n8274 ;
  assign n8276 = ~\u5_cmd_asserted_reg/NET0131  & n1465 ;
  assign n8277 = n1032 & n8276 ;
  assign n8278 = ~n2004 & ~n8277 ;
  assign n8279 = ~n8275 & n8278 ;
  assign n8280 = ~\u2_row_same_reg/P0001  & ~n3176 ;
  assign n8281 = n3172 & n8280 ;
  assign n8282 = n1922 & n8281 ;
  assign n8283 = \u5_state_reg[4]/NET0131  & n1922 ;
  assign n8284 = ~n2809 & n8283 ;
  assign n8285 = ~n8282 & ~n8284 ;
  assign n8286 = \u5_state_reg[4]/NET0131  & ~n2811 ;
  assign n8287 = ~n1922 & n8286 ;
  assign n8288 = n8278 & ~n8287 ;
  assign n8289 = n8285 & n8288 ;
  assign n8290 = ~n8279 & ~n8289 ;
  assign n8291 = ~\u5_cmd_asserted_reg/NET0131  & ~\u5_state_reg[23]/NET0131  ;
  assign n8292 = n1455 & ~n8291 ;
  assign n8293 = n1096 & n8292 ;
  assign n8294 = n1078 & n8293 ;
  assign n8295 = \u5_state_reg[23]/NET0131  & ~\u5_tmr_done_reg/NET0131  ;
  assign n8296 = ~n3559 & n8295 ;
  assign n8297 = ~n8294 & ~n8296 ;
  assign n8298 = \u6_write_go_r1_reg/NET0131  & wb_cyc_i_pad ;
  assign n8299 = ~n1231 & n8298 ;
  assign n8300 = \u5_state_reg[44]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n8301 = ~n1882 & n8300 ;
  assign n8302 = ~n1395 & ~n8301 ;
  assign n8303 = ~n1898 & ~n2189 ;
  assign n8304 = \u6_read_go_r1_reg/NET0131  & wb_cyc_i_pad ;
  assign n8305 = ~\u5_state_reg[39]/NET0131  & ~\u5_tmr2_done_reg/NET0131  ;
  assign n8306 = n1415 & ~n8305 ;
  assign n8307 = n968 & n8306 ;
  assign n8308 = n1088 & n8307 ;
  assign n8309 = n960 & n1353 ;
  assign n8310 = n964 & n8309 ;
  assign n8311 = n1122 & n8310 ;
  assign n8312 = ~n8308 & ~n8311 ;
  assign n8313 = \u5_tmr2_done_reg/NET0131  & ~n1147 ;
  assign n8314 = ~n1941 & ~n8313 ;
  assign n8315 = \u5_tmr2_done_reg/NET0131  & ~n2821 ;
  assign n8316 = ~n2820 & n8315 ;
  assign n8317 = n1281 & ~n8316 ;
  assign n8318 = n2158 & ~n8317 ;
  assign n8319 = ~n3688 & n5855 ;
  assign n8320 = n1840 & n8319 ;
  assign n8321 = ~n1839 & n5855 ;
  assign n8322 = n1835 & n8321 ;
  assign n8323 = ~n3743 & n8322 ;
  assign n8324 = \u2_u0_bank0_open_reg/NET0131  & ~n8323 ;
  assign n8325 = ~\u5_rfr_ack_r_reg/NET0131  & n8324 ;
  assign n8326 = ~n3736 & n8325 ;
  assign n8327 = ~n8320 & ~n8326 ;
  assign n8328 = ~n1919 & n8319 ;
  assign n8329 = n3763 & n5855 ;
  assign n8330 = \u2_u1_bank0_open_reg/NET0131  & ~n8329 ;
  assign n8331 = ~\u5_rfr_ack_r_reg/NET0131  & n8330 ;
  assign n8332 = ~n3762 & n8331 ;
  assign n8333 = ~n8328 & ~n8332 ;
  assign n8334 = ~n1512 & ~n1513 ;
  assign n8335 = ~\u5_cmd_asserted_reg/NET0131  & n1316 ;
  assign n8336 = n1254 & n8335 ;
  assign n8337 = \u5_tmr_done_reg/NET0131  & n1255 ;
  assign n8338 = n1254 & n8337 ;
  assign n8339 = ~n8336 & ~n8338 ;
  assign n8340 = ~n1260 & ~n1889 ;
  assign n8341 = ~\u5_state_reg[12]/NET0131  & ~n1966 ;
  assign n8342 = ~n1954 & n8341 ;
  assign n8343 = n1094 & ~n8342 ;
  assign n8344 = n3295 & n8343 ;
  assign n8345 = \u5_state_reg[12]/NET0131  & ~n2698 ;
  assign n8346 = ~n2700 & ~n8345 ;
  assign n8347 = ~\u5_mem_ack_r_reg/NET0131  & ~n2700 ;
  assign n8348 = ~n1899 & n8347 ;
  assign n8349 = ~n8346 & ~n8348 ;
  assign n8350 = n1413 & n8349 ;
  assign n8351 = ~n8344 & ~n8350 ;
  assign n8352 = n967 & n971 ;
  assign n8353 = n1088 & n8352 ;
  assign n8354 = ~n1089 & ~n1408 ;
  assign n8355 = ~\u7_mc_br_r_reg/P0001  & ~n1089 ;
  assign n8356 = ~n8354 & ~n8355 ;
  assign n8357 = n8353 & n8356 ;
  assign n8358 = n1400 & n2168 ;
  assign n8359 = n1143 & n1899 ;
  assign n8360 = ~n8358 & ~n8359 ;
  assign n8361 = n1897 & ~n8360 ;
  assign n8362 = \u3_u0_wr_adr_reg[0]/NET0131  & n5380 ;
  assign n8363 = ~n1043 & n8362 ;
  assign n8364 = \u3_u0_wr_adr_reg[1]/NET0131  & n5380 ;
  assign n8365 = n1043 & n8364 ;
  assign n8366 = ~n8363 & ~n8365 ;
  assign n8367 = \u3_u0_wr_adr_reg[0]/NET0131  & ~n1043 ;
  assign n8368 = \u7_mc_dqm_r_reg[0]/P0001  & ~n1045 ;
  assign n8369 = \wb_sel_i[0]_pad  & n1045 ;
  assign n8370 = ~n8368 & ~n8369 ;
  assign n8371 = \u7_mc_dqm_r_reg[1]/P0001  & ~n1045 ;
  assign n8372 = \wb_sel_i[1]_pad  & n1045 ;
  assign n8373 = ~n8371 & ~n8372 ;
  assign n8374 = \u7_mc_dqm_r_reg[2]/P0001  & ~n1045 ;
  assign n8375 = \wb_sel_i[2]_pad  & n1045 ;
  assign n8376 = ~n8374 & ~n8375 ;
  assign n8377 = \u7_mc_dqm_r_reg[3]/P0001  & ~n1045 ;
  assign n8378 = \wb_sel_i[3]_pad  & n1045 ;
  assign n8379 = ~n8377 & ~n8378 ;
  assign n8380 = \u5_cmd_del_reg[0]/NET0131  & \u5_wr_cycle_reg/NET0131  ;
  assign n8381 = \u5_wr_cycle_reg/NET0131  & ~n8380 ;
  assign n8382 = ~n1985 & ~n8380 ;
  assign n8383 = n2018 & n8382 ;
  assign n8384 = ~n8381 & ~n8383 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g22/_0_  = n1044 ;
  assign \g23/_0_  = ~n1043 ;
  assign \g25_dup61718/_2_  = n1048 ;
  assign \g43466/_0_  = ~n1557 ;
  assign \g43467/_0_  = ~n1580 ;
  assign \g43468/_0_  = ~n1600 ;
  assign \g43469/_0_  = ~n1620 ;
  assign \g43470/_0_  = ~n1643 ;
  assign \g43471/_0_  = ~n1666 ;
  assign \g43472/_0_  = ~n1689 ;
  assign \g43473/_0_  = ~n1712 ;
  assign \g43474/_0_  = ~n1735 ;
  assign \g43475/_0_  = ~n1758 ;
  assign \g43476/_0_  = ~n1781 ;
  assign \g43477/_0_  = ~n1804 ;
  assign \g43478/_0_  = ~n1827 ;
  assign \g43512/_0_  = ~n1982 ;
  assign \g43513/_0_  = ~n1983 ;
  assign \g43544/_3_  = ~n2019 ;
  assign \g43545/_0_  = n2024 ;
  assign \g43554/_0_  = n2145 ;
  assign \g43555/_0_  = ~n2592 ;
  assign \g43557/_0_  = ~n2593 ;
  assign \g43558/_0_  = n2659 ;
  assign \g43571/_2_  = ~n2718 ;
  assign \g43632/_0_  = n2760 ;
  assign \g43633/_0_  = n2775 ;
  assign \g43635/_0_  = ~n2790 ;
  assign \g43636/_0_  = ~n2798 ;
  assign \g43637/_0_  = n2803 ;
  assign \g43638/_0_  = ~n2829 ;
  assign \g43639/_0_  = ~n2843 ;
  assign \g43640/_0_  = n2855 ;
  assign \g43642/_0_  = n1337 ;
  assign \g43662/_0_  = ~n2860 ;
  assign \g43663/_0_  = ~n2863 ;
  assign \g43664/_0_  = ~n2866 ;
  assign \g43665/_0_  = ~n2869 ;
  assign \g43668/_0_  = ~n2912 ;
  assign \g43670/_0_  = ~n2929 ;
  assign \g43671/_0_  = ~n2936 ;
  assign \g43673/_0_  = ~n3003 ;
  assign \g43674/_0_  = n3063 ;
  assign \g43692/_0_  = n3067 ;
  assign \g43695/_0_  = n3073 ;
  assign \g43696/_0_  = ~n3076 ;
  assign \g43697/_0_  = n3086 ;
  assign \g43698/_0_  = n3102 ;
  assign \g43700/_0_  = n3120 ;
  assign \g43701/_0_  = ~n3127 ;
  assign \g43703/_0_  = n3142 ;
  assign \g43705/_0_  = n3155 ;
  assign \g43707/_0_  = ~n3163 ;
  assign \g43708/_0_  = n3187 ;
  assign \g43710/_0_  = ~n3196 ;
  assign \g43717/_0_  = ~n3202 ;
  assign \g43719/_0_  = ~n3204 ;
  assign \g43720/_0_  = n3208 ;
  assign \g43721/_0_  = n3227 ;
  assign \g43722/_1_  = ~n3233 ;
  assign \g43723/_0_  = ~n3244 ;
  assign \g43725/_0_  = ~n3251 ;
  assign \g43729/_0_  = n3252 ;
  assign \g43731/_0_  = ~n3259 ;
  assign \g43734/_0_  = ~n3268 ;
  assign \g43735/_0_  = ~n3276 ;
  assign \g43737/_0_  = ~n3277 ;
  assign \g43744/_0_  = ~n3282 ;
  assign \g43747/_0_  = ~n3287 ;
  assign \g43760/_2_  = ~n3291 ;
  assign \g43770/_1_  = ~n3307 ;
  assign \g43775/_2_  = ~n3312 ;
  assign \g43780/_2_  = ~n3330 ;
  assign \g43786/_0_  = n3332 ;
  assign \g43787/_1_  = ~n3346 ;
  assign \g43847/_0_  = ~n3359 ;
  assign \g43848/_1_  = ~n3364 ;
  assign \g43858/_1_  = ~n3371 ;
  assign \g43891/_3_  = n3421 ;
  assign \g43895/_0_  = n3457 ;
  assign \g43934/_0_  = n3483 ;
  assign \g43936/_3_  = ~n3510 ;
  assign \g43954/_3_  = ~n3524 ;
  assign \g43961/_0_  = ~n3558 ;
  assign \g44016/_1_  = n3561 ;
  assign \g44067/_0_  = ~n3579 ;
  assign \g44094/_0_  = ~n3596 ;
  assign \g44096/_0_  = n3617 ;
  assign \g44104/_0_  = ~n3640 ;
  assign \g44122/_0_  = n3657 ;
  assign \g44172/_0_  = ~n3521 ;
  assign \g44209/_0_  = ~n3683 ;
  assign \g44219/_0_  = ~n3750 ;
  assign \g44220/_0_  = ~n3760 ;
  assign \g44222/_0_  = ~n3768 ;
  assign \g44223/_0_  = ~n3774 ;
  assign \g44241/_2_  = n3792 ;
  assign \g44252/_0_  = ~n3802 ;
  assign \g44253/_0_  = ~n3808 ;
  assign \g44255/_2_  = ~n3822 ;
  assign \g44263/_2_  = ~n3842 ;
  assign \g44470/_0_  = ~n3856 ;
  assign \g44538/_0_  = ~n3900 ;
  assign \g44539/_0_  = ~n3910 ;
  assign \g44540/_0_  = ~n3920 ;
  assign \g44541/_0_  = ~n3930 ;
  assign \g44542/_0_  = ~n3940 ;
  assign \g44543/_0_  = ~n3950 ;
  assign \g44544/_0_  = ~n3960 ;
  assign \g44545/_0_  = ~n3970 ;
  assign \g44546/_0_  = ~n3980 ;
  assign \g44547/_0_  = ~n3990 ;
  assign \g44548/_0_  = ~n4000 ;
  assign \g44549/_0_  = ~n4010 ;
  assign \g44550/_0_  = ~n4020 ;
  assign \g44551/_0_  = ~n4030 ;
  assign \g44552/_0_  = ~n4040 ;
  assign \g44553/_0_  = ~n4050 ;
  assign \g44554/_0_  = ~n4060 ;
  assign \g44555/_0_  = ~n4070 ;
  assign \g44556/_0_  = ~n4080 ;
  assign \g44557/_0_  = ~n4090 ;
  assign \g44558/_0_  = ~n4100 ;
  assign \g44559/_0_  = ~n4110 ;
  assign \g44560/_0_  = ~n4120 ;
  assign \g44561/_0_  = ~n4130 ;
  assign \g44562/_0_  = ~n4140 ;
  assign \g44563/_0_  = ~n4150 ;
  assign \g44564/_0_  = ~n4160 ;
  assign \g44565/_0_  = ~n4170 ;
  assign \g44566/_0_  = ~n4267 ;
  assign \g44567/_0_  = ~n4279 ;
  assign \g44568/_0_  = ~n4291 ;
  assign \g44569/_0_  = ~n4303 ;
  assign \g44570/_0_  = ~n4315 ;
  assign \g44571/_0_  = ~n4327 ;
  assign \g44572/_0_  = ~n4339 ;
  assign \g44573/_0_  = ~n4351 ;
  assign \g44574/_0_  = ~n4363 ;
  assign \g44575/_0_  = ~n4375 ;
  assign \g44576/_0_  = ~n4387 ;
  assign \g44577/_0_  = ~n4399 ;
  assign \g44578/_0_  = ~n4411 ;
  assign \g44579/_0_  = ~n4423 ;
  assign \g44580/_0_  = ~n4435 ;
  assign \g44581/_0_  = ~n4447 ;
  assign \g44582/_0_  = ~n4459 ;
  assign \g44583/_0_  = ~n4471 ;
  assign \g44584/_0_  = ~n4483 ;
  assign \g44585/_0_  = ~n4495 ;
  assign \g44586/_0_  = ~n4507 ;
  assign \g44588/_0_  = ~n4519 ;
  assign \g44589/_0_  = ~n4531 ;
  assign \g44590/_0_  = ~n4543 ;
  assign \g44591/_0_  = ~n4555 ;
  assign \g44592/_0_  = ~n4567 ;
  assign \g44593/_0_  = ~n4579 ;
  assign \g44594/_0_  = ~n4591 ;
  assign \g44595/_0_  = ~n4609 ;
  assign \g44596/_0_  = ~n4626 ;
  assign \g44636/_2_  = ~n4644 ;
  assign \g44646/_0_  = ~n4654 ;
  assign \g44647/_0_  = ~n4663 ;
  assign \g44648/_0_  = ~n4672 ;
  assign \g44649/_0_  = ~n4681 ;
  assign \g44650/_0_  = ~n4690 ;
  assign \g44651/_0_  = ~n4699 ;
  assign \g44652/_0_  = ~n4707 ;
  assign \g44653/_0_  = ~n4715 ;
  assign \g44654/_0_  = ~n4723 ;
  assign \g44655/_0_  = ~n4731 ;
  assign \g44656/_0_  = ~n4739 ;
  assign \g44657/_0_  = ~n4747 ;
  assign \g44665/_0_  = ~n4751 ;
  assign \g44666/_0_  = ~n4760 ;
  assign \g44667/_0_  = ~n4769 ;
  assign \g44668/_0_  = ~n4778 ;
  assign \g44752/_0_  = ~n4793 ;
  assign \g44753/_0_  = ~n4803 ;
  assign \g44873/_0_  = ~n1472 ;
  assign \g44939/_0_  = ~n4816 ;
  assign \g44942/_0_  = ~n4824 ;
  assign \g44945/_0_  = ~n4833 ;
  assign \g45023/_2_  = ~n4848 ;
  assign \g45090/_0_  = n4645 ;
  assign \g45141/_0_  = n4857 ;
  assign \g45147/_3_  = ~n4868 ;
  assign \g45155/_0_  = ~n4882 ;
  assign \g45190/_0_  = n4884 ;
  assign \g45195/_2_  = ~n4900 ;
  assign \g45199/_2_  = ~n4919 ;
  assign \g45201/_2_  = ~n4932 ;
  assign \g45324/_0_  = ~n4947 ;
  assign \g45334/_2_  = ~n4968 ;
  assign \g45336/_0_  = ~n4866 ;
  assign \g45388/_0_  = ~n4975 ;
  assign \g45391/_0_  = n4995 ;
  assign \g45413/_2_  = ~n5011 ;
  assign \g45530/_0_  = ~n5024 ;
  assign \g45532/_0_  = n5037 ;
  assign \g45533/_0_  = n5052 ;
  assign \g45534/_0_  = n5065 ;
  assign \g45739/_2_  = ~n5086 ;
  assign \g45743/_2_  = ~n5107 ;
  assign \g45767/_0_  = n5140 ;
  assign \g45782/_0_  = n5154 ;
  assign \g45830/_3_  = ~n5184 ;
  assign \g45834/_3_  = ~n5210 ;
  assign \g45835/_3_  = ~n5220 ;
  assign \g45836/_3_  = ~n5234 ;
  assign \g45837/_3_  = ~n5243 ;
  assign \g45839/_3_  = ~n5252 ;
  assign \g45840/_3_  = ~n5261 ;
  assign \g45841/_3_  = ~n5270 ;
  assign \g45842/_3_  = ~n5279 ;
  assign \g45843/_3_  = ~n5287 ;
  assign \g45844/_3_  = n5292 ;
  assign \g45845/_3_  = ~n5295 ;
  assign \g46191/_0_  = ~n5297 ;
  assign \g46193/_3_  = ~n5303 ;
  assign \g46256/_3_  = n5316 ;
  assign \g46257/_3_  = n5325 ;
  assign \g46258/_3_  = n5334 ;
  assign \g46259/_3_  = n5343 ;
  assign \g46260/_3_  = n5352 ;
  assign \g46261/_3_  = n5361 ;
  assign \g46262/_3_  = n5370 ;
  assign \g46263/_3_  = n5379 ;
  assign \g46278/_0_  = n5385 ;
  assign \g46292/_0_  = ~n5390 ;
  assign \g46293/_0_  = ~n5394 ;
  assign \g46312/_0_  = ~n5403 ;
  assign \g46367/_2_  = ~n5424 ;
  assign \g46370/_2_  = ~n5437 ;
  assign \g46380/_2_  = ~n5458 ;
  assign \g46386/_2_  = ~n5475 ;
  assign \g46388/_2_  = ~n5494 ;
  assign \g46392/_2_  = ~n5511 ;
  assign \g46395/_2_  = ~n5528 ;
  assign \g46399/_2_  = ~n5541 ;
  assign \g46420/_0_  = n5543 ;
  assign \g46446/_0_  = ~n5547 ;
  assign \g46493/_0_  = ~n5556 ;
  assign \g46510/_0_  = n5559 ;
  assign \g46669/_2_  = n5569 ;
  assign \g46691/_0_  = n5617 ;
  assign \g46708/_0_  = ~n5623 ;
  assign \g46721/_00_  = ~n5645 ;
  assign \g46776/_0_  = n5648 ;
  assign \g46777/_0_  = n5653 ;
  assign \g46778/_0_  = ~n5658 ;
  assign \g46779/_0_  = n5663 ;
  assign \g46780/_0_  = n5669 ;
  assign \g46782/_0_  = ~n5674 ;
  assign \g46784/_0_  = n5680 ;
  assign \g46932/_0_  = ~n5692 ;
  assign \g47112/_0_  = ~n5699 ;
  assign \g47124/_0_  = n5708 ;
  assign \g47265/_0_  = ~n5717 ;
  assign \g47270/_0_  = n5726 ;
  assign \g47275/_0_  = ~n5735 ;
  assign \g47300/_1_  = n5736 ;
  assign \g47305/_1_  = n5737 ;
  assign \g47338/_0_  = ~n5742 ;
  assign \g47339/_0_  = ~n5747 ;
  assign \g47352/_0_  = ~n6173 ;
  assign \g47699/_3_  = n6177 ;
  assign \g47711/_0_  = ~n6183 ;
  assign \g47719/_3_  = ~n6188 ;
  assign \g47721/_3_  = ~n6193 ;
  assign \g47723/_3_  = ~n6198 ;
  assign \g47853/_0_  = n6201 ;
  assign \g48094/_0_  = ~n6213 ;
  assign \g48095/_0_  = ~n6225 ;
  assign \g48177/_2_  = ~n6229 ;
  assign \g48194/_0_  = ~n6230 ;
  assign \g48369/_2_  = ~n6239 ;
  assign \g48371/_2_  = ~n6248 ;
  assign \g48373/_2_  = ~n6257 ;
  assign \g48375/_2_  = ~n6266 ;
  assign \g48377/_2_  = ~n6275 ;
  assign \g48379/_2_  = ~n6284 ;
  assign \g48381/_2_  = ~n6293 ;
  assign \g48383/_2_  = ~n6302 ;
  assign \g48385/_2_  = ~n6311 ;
  assign \g48535/_0_  = n6315 ;
  assign \g48569/_0_  = n6319 ;
  assign \g48570/_0_  = n6322 ;
  assign \g48571/_0_  = n6325 ;
  assign \g48836/_0_  = n6328 ;
  assign \g48843/_0_  = n6331 ;
  assign \g49187/_3_  = n5151 ;
  assign \g49375/_2_  = n6334 ;
  assign \g49633/_0_  = n6337 ;
  assign \g49788/_1_  = n3769 ;
  assign \g49800/_1_  = n3761 ;
  assign \g49802/_1_  = n3803 ;
  assign \g49806/_1_  = n3690 ;
  assign \g49853/_1_  = n3795 ;
  assign \g49883/_0_  = n6345 ;
  assign \g49884/_0_  = ~n6350 ;
  assign \g49885/_0_  = ~n6354 ;
  assign \g49886/_0_  = ~n6358 ;
  assign \g49976/_1_  = n3753 ;
  assign \g50038/_0_  = ~n6376 ;
  assign \g50082/_0_  = ~n6391 ;
  assign \g50083/_0_  = n5608 ;
  assign \g50167/_3_  = n6429 ;
  assign \g50168/_3_  = n6457 ;
  assign \g50169/_3_  = n6485 ;
  assign \g50170/_3_  = n6513 ;
  assign \g50171/_3_  = n6541 ;
  assign \g50177/_0_  = ~n6549 ;
  assign \g50190/_0_  = ~n6556 ;
  assign \g50236/_0_  = n4216 ;
  assign \g50251/_3_  = n6584 ;
  assign \g50256/_0_  = n4258 ;
  assign \g50318/_3_  = n6612 ;
  assign \g50319/_3_  = n6640 ;
  assign \g50350/_3_  = n6669 ;
  assign \g50351/_3_  = n6698 ;
  assign \g50352/_3_  = n6727 ;
  assign \g50353/_3_  = n6756 ;
  assign \g50354/_3_  = n6785 ;
  assign \g50355/_3_  = n6814 ;
  assign \g50361/_2_  = n6817 ;
  assign \g50366/_0_  = ~n6829 ;
  assign \g50393/_0_  = n6831 ;
  assign \g50552/_1_  = n2042 ;
  assign \g51108/_0_  = ~n6838 ;
  assign \g51160/_0_  = ~n6844 ;
  assign \g51290/_1_  = n6847 ;
  assign \g51327/_3_  = n6871 ;
  assign \g51328/_3_  = n6895 ;
  assign \g51329/_3_  = n6919 ;
  assign \g51330/_3_  = n6943 ;
  assign \g51331/_3_  = n6967 ;
  assign \g51332/_3_  = n6991 ;
  assign \g51333/_3_  = n7015 ;
  assign \g51334/_3_  = n7039 ;
  assign \g51339/_3_  = n7061 ;
  assign \g51340/_3_  = n7083 ;
  assign \g51341/_3_  = n7105 ;
  assign \g51342/_3_  = n7127 ;
  assign \g51343/_3_  = n7149 ;
  assign \g51346/_0_  = ~n7156 ;
  assign \g51347/_0_  = ~n7163 ;
  assign \g51348/_0_  = n7167 ;
  assign \g51381/_3_  = n7196 ;
  assign \g51382/_3_  = n7225 ;
  assign \g51383/_3_  = n7254 ;
  assign \g51386/_3_  = n7283 ;
  assign \g51387/_3_  = n7312 ;
  assign \g51405/_3_  = ~n7321 ;
  assign \g51410/_3_  = ~n7330 ;
  assign \g51883/_0_  = n7333 ;
  assign \g51916/_0_  = n5600 ;
  assign \g51947/_0_  = n7339 ;
  assign \g51948/_0_  = n7345 ;
  assign \g51949/_0_  = n7354 ;
  assign \g51950/_0_  = n7360 ;
  assign \g51951/_0_  = n7366 ;
  assign \g51952/_0_  = n7372 ;
  assign \g51953/_0_  = n7378 ;
  assign \g51954/_0_  = n7384 ;
  assign \g51955/_0_  = n7390 ;
  assign \g51956/_0_  = n7396 ;
  assign \g51957/_0_  = n7402 ;
  assign \g51958/_0_  = n7408 ;
  assign \g51959/_0_  = n7414 ;
  assign \g51960/_0_  = n7420 ;
  assign \g51961/_0_  = n7426 ;
  assign \g51962/_0_  = n7432 ;
  assign \g51963/_0_  = n7438 ;
  assign \g51964/_0_  = n7444 ;
  assign \g51965/_0_  = n7450 ;
  assign \g51967/_0_  = n7456 ;
  assign \g51968/_0_  = ~n7463 ;
  assign \g51969/_0_  = ~n7469 ;
  assign \g51970/_0_  = ~n7475 ;
  assign \g51971/_0_  = ~n7481 ;
  assign \g51972/_0_  = ~n7487 ;
  assign \g51973/_0_  = ~n7493 ;
  assign \g51974/_0_  = ~n7499 ;
  assign \g51975/_0_  = ~n7505 ;
  assign \g51976/_0_  = ~n7511 ;
  assign \g51977/_0_  = ~n7517 ;
  assign \g51978/_0_  = ~n7523 ;
  assign \g51979/_0_  = ~n7529 ;
  assign \g51980/_0_  = ~n7535 ;
  assign \g51981/_0_  = ~n7541 ;
  assign \g51982/_0_  = ~n7547 ;
  assign \g51983/_0_  = ~n7553 ;
  assign \g51984/_0_  = ~n7559 ;
  assign \g51985/_0_  = ~n7565 ;
  assign \g51986/_0_  = ~n7571 ;
  assign \g51987/_0_  = n7577 ;
  assign \g51988/_0_  = ~n7583 ;
  assign \g51989/_0_  = ~n7589 ;
  assign \g51990/_0_  = ~n7595 ;
  assign \g51991/_0_  = n7601 ;
  assign \g51992/_0_  = ~n7607 ;
  assign \g51993/_0_  = ~n7613 ;
  assign \g51994/_0_  = ~n7619 ;
  assign \g51995/_0_  = ~n7625 ;
  assign \g51996/_0_  = ~n7631 ;
  assign \g51997/_0_  = ~n7637 ;
  assign \g51998/_0_  = ~n7643 ;
  assign \g51999/_0_  = ~n7649 ;
  assign \g52000/_0_  = n7654 ;
  assign \g52001/_0_  = n7660 ;
  assign \g52002/_0_  = n7664 ;
  assign \g52003/_0_  = n7668 ;
  assign \g52004/_0_  = n7672 ;
  assign \g52005/_0_  = n7676 ;
  assign \g52006/_0_  = n7680 ;
  assign \g52007/_0_  = n7684 ;
  assign \g52008/_0_  = n7690 ;
  assign \g52009/_0_  = n7696 ;
  assign \g52010/_0_  = n7700 ;
  assign \g52011/_0_  = n7704 ;
  assign \g52012/_0_  = n7710 ;
  assign \g52013/_0_  = n7714 ;
  assign \g52014/_0_  = n7720 ;
  assign \g52015/_0_  = n7724 ;
  assign \g52016/_0_  = n7728 ;
  assign \g52017/_0_  = n7732 ;
  assign \g52018/_0_  = n7736 ;
  assign \g52019/_0_  = n7740 ;
  assign \g52020/_0_  = n7744 ;
  assign \g52021/_0_  = n7750 ;
  assign \g52022/_0_  = n7754 ;
  assign \g52023/_0_  = n7758 ;
  assign \g52024/_0_  = n7762 ;
  assign \g52025/_0_  = n7768 ;
  assign \g52026/_0_  = n7774 ;
  assign \g52027/_0_  = n7778 ;
  assign \g52028/_0_  = n7784 ;
  assign \g52029/_0_  = n7790 ;
  assign \g52030/_0_  = n7796 ;
  assign \g52031/_0_  = n7800 ;
  assign \g52032/_0_  = n7804 ;
  assign \g52033/_0_  = n7810 ;
  assign \g52034/_0_  = n7816 ;
  assign \g52035/_0_  = n7822 ;
  assign \g52036/_0_  = n7828 ;
  assign \g52037/_0_  = n7834 ;
  assign \g52038/_0_  = n7840 ;
  assign \g52039/_0_  = n7846 ;
  assign \g52040/_0_  = n7852 ;
  assign \g52041/_0_  = n7858 ;
  assign \g52042/_0_  = n7864 ;
  assign \g52043/_0_  = n7870 ;
  assign \g52044/_0_  = n7876 ;
  assign \g52045/_0_  = n7882 ;
  assign \g52046/_0_  = n7888 ;
  assign \g52047/_0_  = n7894 ;
  assign \g52049/_0_  = n7900 ;
  assign \g52050/_0_  = n7906 ;
  assign \g52051/_0_  = n7910 ;
  assign \g52052/_0_  = n7916 ;
  assign \g52053/_0_  = n7922 ;
  assign \g52054/_0_  = n7928 ;
  assign \g52055/_0_  = n7934 ;
  assign \g52056/_0_  = ~n7940 ;
  assign \g52057/_0_  = n7946 ;
  assign \g52058/_0_  = n7952 ;
  assign \g52061/_0_  = n7958 ;
  assign \g52065/_0_  = n7964 ;
  assign \g52066/_0_  = n7970 ;
  assign \g52067/_0_  = n7974 ;
  assign \g52068/_0_  = n7980 ;
  assign \g52069/_0_  = n7984 ;
  assign \g52070/_0_  = n7988 ;
  assign \g52071/_0_  = n7992 ;
  assign \g52073/_0_  = ~n7998 ;
  assign \g52074/_0_  = n8004 ;
  assign \g52075/_0_  = n8008 ;
  assign \g52082/_0_  = n8012 ;
  assign \g52083/_0_  = n8016 ;
  assign \g52158/_0_  = n8019 ;
  assign \g52201/_0_  = ~n8020 ;
  assign \g52202/_0_  = ~n8021 ;
  assign \g52346/_0_  = n2069 ;
  assign \g52351/_0_  = ~n8024 ;
  assign \g52390/_0_  = n8028 ;
  assign \g52847/_0_  = ~n8029 ;
  assign \g52854/_0_  = n8031 ;
  assign \g52968/_0_  = ~n8052 ;
  assign \g52969/_0_  = ~n8073 ;
  assign \g52970/_0_  = ~n8094 ;
  assign \g52971/_0_  = ~n8115 ;
  assign \g52984/_0_  = ~n8119 ;
  assign \g52994/_0_  = n5728 ;
  assign \g53019/_0_  = n7457 ;
  assign \g53030/_0_  = n7348 ;
  assign \g53094/_1_  = n6381 ;
  assign \g53106/_0_  = n7650 ;
  assign \g53150/_0_  = n8130 ;
  assign \g53256/_0_  = n8132 ;
  assign \g53297/_0_  = n8134 ;
  assign \g53345/_0_  = n8135 ;
  assign \g53359/_0_  = n8138 ;
  assign \g53375/_0_  = n8139 ;
  assign \g53474/_1__syn_2  = n8142 ;
  assign \g53475/_2_  = n8143 ;
  assign \g53593/_0_  = ~n8145 ;
  assign \g53643/_1_  = ~n8147 ;
  assign \g53655/_0_  = ~n8148 ;
  assign \g53710/_0_  = ~n8149 ;
  assign \g53786/_0_  = ~n8151 ;
  assign \g53837/_0_  = n8153 ;
  assign \g53888/_1_  = n5681 ;
  assign \g53909/_0_  = ~n1062 ;
  assign \g54253/_2_  = ~n8155 ;
  assign \g54394/_3_  = ~n5550 ;
  assign \g54413/_0_  = ~n8158 ;
  assign \g55420/_0_  = ~n8159 ;
  assign \g55587/_0_  = ~n8160 ;
  assign \g55852/_0_  = ~\u5_mc_le_reg/NET0131  ;
  assign \g57020/_0_  = ~\u1_acs_addr_reg[0]/P0001  ;
  assign \g59450/_0_  = ~n8211 ;
  assign \g59488/_2_  = ~n1511 ;
  assign \g59752/_0_  = ~n8216 ;
  assign \g59786/_0_  = ~n8219 ;
  assign \g59854/_0_  = ~n8221 ;
  assign \g59878/_0_  = ~n8225 ;
  assign \g59902/_0_  = ~n8230 ;
  assign \g59924/_0_  = n8235 ;
  assign \g59947/_0_  = n8245 ;
  assign \g59972/_0_  = ~n8252 ;
  assign \g59996/_0_  = ~n8256 ;
  assign \g60017/_0_  = ~n8261 ;
  assign \g60040/_0_  = ~n8265 ;
  assign \g60064/_0_  = n8268 ;
  assign \g60095/_0_  = ~n8270 ;
  assign \g60119/_0_  = ~n8273 ;
  assign \g60145/_1_  = n8290 ;
  assign \g60165/_0_  = ~n8297 ;
  assign \g60407/_2_  = n1895 ;
  assign \g60408/_0_  = n8299 ;
  assign \g60613/_2_  = ~n8302 ;
  assign \g60649/_0_  = n8303 ;
  assign \g60771/_0_  = n8304 ;
  assign \g60908/_1_  = ~n8312 ;
  assign \g60911/_0_  = n8314 ;
  assign \g60977/_0_  = ~n3889 ;
  assign \g61/_0_  = n1084 ;
  assign \g61002/_0_  = ~n8318 ;
  assign \g61308/_0_  = ~n8327 ;
  assign \g61312/_1_  = n8320 ;
  assign \g61314/_0_  = ~n8333 ;
  assign \g61319/_1_  = n8328 ;
  assign \g61342/_1_  = ~n8334 ;
  assign \g61360/_0_  = ~n8339 ;
  assign \g61377/_0_  = ~n8340 ;
  assign \g61423/_1_  = n1899 ;
  assign \g61426/_0_  = n1898 ;
  assign \g61479/_1_  = ~n8351 ;
  assign \g61523/_1_  = n8357 ;
  assign \g61558/_1_  = n3411 ;
  assign \g61652/_0_  = n8361 ;
  assign \g61866/_0_  = ~n8366 ;
  assign \g61868/_1_  = n8367 ;
  assign \g61887/_0_  = ~n1966 ;
  assign \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3  = ~n8370 ;
  assign \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3  = ~n8373 ;
  assign \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3  = ~n8376 ;
  assign \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3  = ~n8379 ;
  assign \u7_mc_we__reg/_05_  = n8384 ;
endmodule
