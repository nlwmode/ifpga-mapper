module top (\B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] , \B[8] , \B[9] , \B[10] , \M[0] , \M[1] , \M[2] , \M[3] , \E[0] , \E[1] , \E[2] );
	input \B[0]  ;
	input \B[1]  ;
	input \B[2]  ;
	input \B[3]  ;
	input \B[4]  ;
	input \B[5]  ;
	input \B[6]  ;
	input \B[7]  ;
	input \B[8]  ;
	input \B[9]  ;
	input \B[10]  ;
	output \M[0]  ;
	output \M[1]  ;
	output \M[2]  ;
	output \M[3]  ;
	output \E[0]  ;
	output \E[1]  ;
	output \E[2]  ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w14_ ;
	wire _w13_ ;
	wire _w12_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\B[6] ,
		\B[7] ,
		_w12_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\B[10] ,
		_w12_,
		_w13_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\B[5] ,
		\B[6] ,
		_w14_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\B[9] ,
		_w14_,
		_w15_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\B[4] ,
		\B[7] ,
		_w16_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\B[2] ,
		\B[7] ,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\B[1] ,
		\B[5] ,
		_w18_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w17_,
		_w18_,
		_w19_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w16_,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\B[3] ,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\B[3] ,
		\B[4] ,
		_w22_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\B[7] ,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w21_,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\B[8] ,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\B[4] ,
		\B[8] ,
		_w26_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\B[5] ,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\B[6] ,
		\B[7] ,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\B[1] ,
		\B[4] ,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w26_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\B[0] ,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		\B[0] ,
		_w29_,
		_w32_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		_w28_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w31_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\B[4] ,
		\B[8] ,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\B[5] ,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w34_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w27_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w25_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\B[9] ,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\B[5] ,
		\B[6] ,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\B[3] ,
		\B[4] ,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\B[1] ,
		\B[2] ,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w16_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w35_,
		_w42_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\B[7] ,
		\B[8] ,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		\B[1] ,
		\B[2] ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\B[9] ,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		_w46_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		_w41_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w15_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w40_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\B[10] ,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\B[2] ,
		\B[3] ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\B[2] ,
		\B[3] ,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\B[8] ,
		\B[9] ,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w56_,
		_w57_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\B[10] ,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\B[7] ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\B[8] ,
		\B[10] ,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\B[9] ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w62_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\B[6] ,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w13_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w55_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\B[6] ,
		\B[7] ,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\B[9] ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w63_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\B[4] ,
		_w28_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\B[4] ,
		_w58_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\B[1] ,
		\B[2] ,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\B[7] ,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\B[3] ,
		_w72_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w73_,
		_w75_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\B[4] ,
		\B[9] ,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		\B[7] ,
		\B[9] ,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\B[6] ,
		_w58_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w79_,
		_w80_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w81_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w78_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\B[5] ,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\B[9] ,
		_w26_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w80_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\B[6] ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\B[7] ,
		_w42_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w58_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\B[8] ,
		\B[9] ,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w17_,
		_w79_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\B[1] ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\B[4] ,
		\B[7] ,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\B[0] ,
		_w74_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\B[0] ,
		\B[2] ,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		_w94_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w95_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w91_,
		_w93_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w98_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\B[6] ,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w80_,
		_w90_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\B[5] ,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w85_,
		_w88_,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w104_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\B[10] ,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\B[6] ,
		\B[9] ,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\B[2] ,
		_w42_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w108_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		\B[4] ,
		_w108_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\B[3] ,
		\B[5] ,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\B[6] ,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w111_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\B[2] ,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\B[1] ,
		_w41_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w111_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\B[3] ,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w110_,
		_w115_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\B[7] ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\B[10] ,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\B[8] ,
		_w69_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w71_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w107_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\B[0] ,
		\B[6] ,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w22_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\B[3] ,
		\B[4] ,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\B[5] ,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w128_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\B[1] ,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\B[4] ,
		\B[6] ,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\B[0] ,
		\B[1] ,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		_w42_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w133_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\B[5] ,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w132_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\B[2] ,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\B[3] ,
		\B[6] ,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		\B[2] ,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w112_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\B[4] ,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w139_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\B[7] ,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\B[5] ,
		\B[6] ,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w42_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\B[2] ,
		_w14_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w116_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		_w42_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w147_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w145_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		\B[8] ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\B[4] ,
		\B[5] ,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w17_,
		_w140_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w28_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		_w154_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w69_,
		_w154_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w153_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\B[9] ,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w94_,
		_w146_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w12_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\B[8] ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w161_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\B[10] ,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\B[5] ,
		\B[8] ,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\B[9] ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w63_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		_w69_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\B[5] ,
		\B[7] ,
		_w171_
	);
	LUT2 #(
		.INIT('h2)
	) name160 (
		\B[8] ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\B[10] ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name162 (
		\B[9] ,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w170_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w166_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		\B[9] ,
		\B[10] ,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		\B[5] ,
		_w47_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w133_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\B[7] ,
		_w146_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\B[2] ,
		_w35_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w180_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w179_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		\B[3] ,
		_w177_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		_w183_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\B[8] ,
		_w180_,
		_w186_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		\B[9] ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\B[5] ,
		_w74_,
		_w188_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\B[7] ,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w89_,
		_w146_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\B[5] ,
		\B[6] ,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w134_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w162_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		_w57_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		\B[4] ,
		_w112_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\B[6] ,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w191_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w195_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\B[8] ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\B[3] ,
		\B[8] ,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w56_,
		_w154_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		_w70_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w187_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		_w200_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\B[10] ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w109_,
		_w146_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		_w47_,
		_w192_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w208_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w56_,
		_w186_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w57_,
		_w134_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w178_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w211_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\B[4] ,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		_w177_,
		_w210_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w47_,
		_w177_,
		_w218_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w208_,
		_w218_,
		_w219_
	);
	assign \M[0]  = _w68_ ;
	assign \M[1]  = _w126_ ;
	assign \M[2]  = _w176_ ;
	assign \M[3]  = _w185_ ;
	assign \E[0]  = _w207_ ;
	assign \E[1]  = _w217_ ;
	assign \E[2]  = _w219_ ;
endmodule;