module top( ADS_n_pad , \Address[0]_pad  , \Address[10]_pad  , \Address[11]_pad  , \Address[12]_pad  , \Address[13]_pad  , \Address[14]_pad  , \Address[15]_pad  , \Address[16]_pad  , \Address[17]_pad  , \Address[18]_pad  , \Address[19]_pad  , \Address[1]_pad  , \Address[20]_pad  , \Address[21]_pad  , \Address[22]_pad  , \Address[23]_pad  , \Address[24]_pad  , \Address[25]_pad  , \Address[26]_pad  , \Address[27]_pad  , \Address[28]_pad  , \Address[29]_pad  , \Address[2]_pad  , \Address[3]_pad  , \Address[4]_pad  , \Address[5]_pad  , \Address[6]_pad  , \Address[7]_pad  , \Address[8]_pad  , \Address[9]_pad  , \BE_n[0]_pad  , \BE_n[1]_pad  , \BE_n[2]_pad  , \BE_n[3]_pad  , \BS16_n_pad  , \ByteEnable_reg[0]/NET0131  , \ByteEnable_reg[1]/NET0131  , \ByteEnable_reg[2]/NET0131  , \ByteEnable_reg[3]/NET0131  , \CodeFetch_reg/NET0131  , D_C_n_pad , \DataWidth_reg[0]/NET0131  , \DataWidth_reg[1]/NET0131  , \Datai[0]_pad  , \Datai[10]_pad  , \Datai[11]_pad  , \Datai[12]_pad  , \Datai[13]_pad  , \Datai[14]_pad  , \Datai[15]_pad  , \Datai[16]_pad  , \Datai[17]_pad  , \Datai[18]_pad  , \Datai[19]_pad  , \Datai[1]_pad  , \Datai[20]_pad  , \Datai[21]_pad  , \Datai[22]_pad  , \Datai[23]_pad  , \Datai[24]_pad  , \Datai[25]_pad  , \Datai[26]_pad  , \Datai[27]_pad  , \Datai[28]_pad  , \Datai[29]_pad  , \Datai[2]_pad  , \Datai[30]_pad  , \Datai[31]_pad  , \Datai[3]_pad  , \Datai[4]_pad  , \Datai[5]_pad  , \Datai[6]_pad  , \Datai[7]_pad  , \Datai[8]_pad  , \Datai[9]_pad  , \Datao[0]_pad  , \Datao[10]_pad  , \Datao[11]_pad  , \Datao[12]_pad  , \Datao[13]_pad  , \Datao[14]_pad  , \Datao[15]_pad  , \Datao[16]_pad  , \Datao[17]_pad  , \Datao[18]_pad  , \Datao[19]_pad  , \Datao[1]_pad  , \Datao[20]_pad  , \Datao[21]_pad  , \Datao[22]_pad  , \Datao[23]_pad  , \Datao[24]_pad  , \Datao[25]_pad  , \Datao[26]_pad  , \Datao[27]_pad  , \Datao[28]_pad  , \Datao[29]_pad  , \Datao[2]_pad  , \Datao[30]_pad  , \Datao[3]_pad  , \Datao[4]_pad  , \Datao[5]_pad  , \Datao[6]_pad  , \Datao[7]_pad  , \Datao[8]_pad  , \Datao[9]_pad  , \EAX_reg[0]/NET0131  , \EAX_reg[10]/NET0131  , \EAX_reg[11]/NET0131  , \EAX_reg[12]/NET0131  , \EAX_reg[13]/NET0131  , \EAX_reg[14]/NET0131  , \EAX_reg[15]/NET0131  , \EAX_reg[16]/NET0131  , \EAX_reg[17]/NET0131  , \EAX_reg[18]/NET0131  , \EAX_reg[19]/NET0131  , \EAX_reg[1]/NET0131  , \EAX_reg[20]/NET0131  , \EAX_reg[21]/NET0131  , \EAX_reg[22]/NET0131  , \EAX_reg[23]/NET0131  , \EAX_reg[24]/NET0131  , \EAX_reg[25]/NET0131  , \EAX_reg[26]/NET0131  , \EAX_reg[27]/NET0131  , \EAX_reg[28]/NET0131  , \EAX_reg[29]/NET0131  , \EAX_reg[2]/NET0131  , \EAX_reg[30]/NET0131  , \EAX_reg[31]/NET0131  , \EAX_reg[3]/NET0131  , \EAX_reg[4]/NET0131  , \EAX_reg[5]/NET0131  , \EAX_reg[6]/NET0131  , \EAX_reg[7]/NET0131  , \EAX_reg[8]/NET0131  , \EAX_reg[9]/NET0131  , \EBX_reg[0]/NET0131  , \EBX_reg[10]/NET0131  , \EBX_reg[11]/NET0131  , \EBX_reg[12]/NET0131  , \EBX_reg[13]/NET0131  , \EBX_reg[14]/NET0131  , \EBX_reg[15]/NET0131  , \EBX_reg[16]/NET0131  , \EBX_reg[17]/NET0131  , \EBX_reg[18]/NET0131  , \EBX_reg[19]/NET0131  , \EBX_reg[1]/NET0131  , \EBX_reg[20]/NET0131  , \EBX_reg[21]/NET0131  , \EBX_reg[22]/NET0131  , \EBX_reg[23]/NET0131  , \EBX_reg[24]/NET0131  , \EBX_reg[25]/NET0131  , \EBX_reg[26]/NET0131  , \EBX_reg[27]/NET0131  , \EBX_reg[28]/NET0131  , \EBX_reg[29]/NET0131  , \EBX_reg[2]/NET0131  , \EBX_reg[30]/NET0131  , \EBX_reg[31]/NET0131  , \EBX_reg[3]/NET0131  , \EBX_reg[4]/NET0131  , \EBX_reg[5]/NET0131  , \EBX_reg[6]/NET0131  , \EBX_reg[7]/NET0131  , \EBX_reg[8]/NET0131  , \EBX_reg[9]/NET0131  , \Flush_reg/NET0131  , HOLD_pad , \InstAddrPointer_reg[0]/NET0131  , \InstAddrPointer_reg[10]/NET0131  , \InstAddrPointer_reg[11]/NET0131  , \InstAddrPointer_reg[12]/NET0131  , \InstAddrPointer_reg[13]/NET0131  , \InstAddrPointer_reg[14]/NET0131  , \InstAddrPointer_reg[15]/NET0131  , \InstAddrPointer_reg[16]/NET0131  , \InstAddrPointer_reg[17]/NET0131  , \InstAddrPointer_reg[18]/NET0131  , \InstAddrPointer_reg[19]/NET0131  , \InstAddrPointer_reg[1]/NET0131  , \InstAddrPointer_reg[20]/NET0131  , \InstAddrPointer_reg[21]/NET0131  , \InstAddrPointer_reg[22]/NET0131  , \InstAddrPointer_reg[23]/NET0131  , \InstAddrPointer_reg[24]/NET0131  , \InstAddrPointer_reg[25]/NET0131  , \InstAddrPointer_reg[26]/NET0131  , \InstAddrPointer_reg[27]/NET0131  , \InstAddrPointer_reg[28]/NET0131  , \InstAddrPointer_reg[29]/NET0131  , \InstAddrPointer_reg[2]/NET0131  , \InstAddrPointer_reg[30]/NET0131  , \InstAddrPointer_reg[31]/NET0131  , \InstAddrPointer_reg[3]/NET0131  , \InstAddrPointer_reg[4]/NET0131  , \InstAddrPointer_reg[5]/NET0131  , \InstAddrPointer_reg[6]/NET0131  , \InstAddrPointer_reg[7]/NET0131  , \InstAddrPointer_reg[8]/NET0131  , \InstAddrPointer_reg[9]/NET0131  , \InstQueueRd_Addr_reg[0]/NET0131  , \InstQueueRd_Addr_reg[1]/NET0131  , \InstQueueRd_Addr_reg[2]/NET0131  , \InstQueueRd_Addr_reg[3]/NET0131  , \InstQueueWr_Addr_reg[0]/NET0131  , \InstQueueWr_Addr_reg[1]/NET0131  , \InstQueueWr_Addr_reg[2]/NET0131  , \InstQueueWr_Addr_reg[3]/NET0131  , \InstQueue_reg[0][0]/NET0131  , \InstQueue_reg[0][1]/NET0131  , \InstQueue_reg[0][2]/NET0131  , \InstQueue_reg[0][3]/NET0131  , \InstQueue_reg[0][4]/NET0131  , \InstQueue_reg[0][5]/NET0131  , \InstQueue_reg[0][6]/NET0131  , \InstQueue_reg[0][7]/NET0131  , \InstQueue_reg[10][0]/NET0131  , \InstQueue_reg[10][1]/NET0131  , \InstQueue_reg[10][2]/NET0131  , \InstQueue_reg[10][3]/NET0131  , \InstQueue_reg[10][4]/NET0131  , \InstQueue_reg[10][5]/NET0131  , \InstQueue_reg[10][6]/NET0131  , \InstQueue_reg[10][7]/NET0131  , \InstQueue_reg[11][0]/NET0131  , \InstQueue_reg[11][1]/NET0131  , \InstQueue_reg[11][2]/NET0131  , \InstQueue_reg[11][3]/NET0131  , \InstQueue_reg[11][4]/NET0131  , \InstQueue_reg[11][5]/NET0131  , \InstQueue_reg[11][6]/NET0131  , \InstQueue_reg[11][7]/NET0131  , \InstQueue_reg[12][0]/NET0131  , \InstQueue_reg[12][1]/NET0131  , \InstQueue_reg[12][2]/NET0131  , \InstQueue_reg[12][3]/NET0131  , \InstQueue_reg[12][4]/NET0131  , \InstQueue_reg[12][5]/NET0131  , \InstQueue_reg[12][6]/NET0131  , \InstQueue_reg[12][7]/NET0131  , \InstQueue_reg[13][0]/NET0131  , \InstQueue_reg[13][1]/NET0131  , \InstQueue_reg[13][2]/NET0131  , \InstQueue_reg[13][3]/NET0131  , \InstQueue_reg[13][4]/NET0131  , \InstQueue_reg[13][5]/NET0131  , \InstQueue_reg[13][6]/NET0131  , \InstQueue_reg[13][7]/NET0131  , \InstQueue_reg[14][0]/NET0131  , \InstQueue_reg[14][1]/NET0131  , \InstQueue_reg[14][2]/NET0131  , \InstQueue_reg[14][3]/NET0131  , \InstQueue_reg[14][4]/NET0131  , \InstQueue_reg[14][5]/NET0131  , \InstQueue_reg[14][6]/NET0131  , \InstQueue_reg[14][7]/NET0131  , \InstQueue_reg[15][0]/NET0131  , \InstQueue_reg[15][1]/NET0131  , \InstQueue_reg[15][2]/NET0131  , \InstQueue_reg[15][3]/NET0131  , \InstQueue_reg[15][4]/NET0131  , \InstQueue_reg[15][5]/NET0131  , \InstQueue_reg[15][6]/NET0131  , \InstQueue_reg[15][7]/NET0131  , \InstQueue_reg[1][0]/NET0131  , \InstQueue_reg[1][1]/NET0131  , \InstQueue_reg[1][2]/NET0131  , \InstQueue_reg[1][3]/NET0131  , \InstQueue_reg[1][4]/NET0131  , \InstQueue_reg[1][5]/NET0131  , \InstQueue_reg[1][6]/NET0131  , \InstQueue_reg[1][7]/NET0131  , \InstQueue_reg[2][0]/NET0131  , \InstQueue_reg[2][1]/NET0131  , \InstQueue_reg[2][2]/NET0131  , \InstQueue_reg[2][3]/NET0131  , \InstQueue_reg[2][4]/NET0131  , \InstQueue_reg[2][5]/NET0131  , \InstQueue_reg[2][6]/NET0131  , \InstQueue_reg[2][7]/NET0131  , \InstQueue_reg[3][0]/NET0131  , \InstQueue_reg[3][1]/NET0131  , \InstQueue_reg[3][2]/NET0131  , \InstQueue_reg[3][3]/NET0131  , \InstQueue_reg[3][4]/NET0131  , \InstQueue_reg[3][5]/NET0131  , \InstQueue_reg[3][6]/NET0131  , \InstQueue_reg[3][7]/NET0131  , \InstQueue_reg[4][0]/NET0131  , \InstQueue_reg[4][1]/NET0131  , \InstQueue_reg[4][2]/NET0131  , \InstQueue_reg[4][3]/NET0131  , \InstQueue_reg[4][4]/NET0131  , \InstQueue_reg[4][5]/NET0131  , \InstQueue_reg[4][6]/NET0131  , \InstQueue_reg[4][7]/NET0131  , \InstQueue_reg[5][0]/NET0131  , \InstQueue_reg[5][1]/NET0131  , \InstQueue_reg[5][2]/NET0131  , \InstQueue_reg[5][3]/NET0131  , \InstQueue_reg[5][4]/NET0131  , \InstQueue_reg[5][5]/NET0131  , \InstQueue_reg[5][6]/NET0131  , \InstQueue_reg[5][7]/NET0131  , \InstQueue_reg[6][0]/NET0131  , \InstQueue_reg[6][1]/NET0131  , \InstQueue_reg[6][2]/NET0131  , \InstQueue_reg[6][3]/NET0131  , \InstQueue_reg[6][4]/NET0131  , \InstQueue_reg[6][5]/NET0131  , \InstQueue_reg[6][6]/NET0131  , \InstQueue_reg[6][7]/NET0131  , \InstQueue_reg[7][0]/NET0131  , \InstQueue_reg[7][1]/NET0131  , \InstQueue_reg[7][2]/NET0131  , \InstQueue_reg[7][3]/NET0131  , \InstQueue_reg[7][4]/NET0131  , \InstQueue_reg[7][5]/NET0131  , \InstQueue_reg[7][6]/NET0131  , \InstQueue_reg[7][7]/NET0131  , \InstQueue_reg[8][0]/NET0131  , \InstQueue_reg[8][1]/NET0131  , \InstQueue_reg[8][2]/NET0131  , \InstQueue_reg[8][3]/NET0131  , \InstQueue_reg[8][4]/NET0131  , \InstQueue_reg[8][5]/NET0131  , \InstQueue_reg[8][6]/NET0131  , \InstQueue_reg[8][7]/NET0131  , \InstQueue_reg[9][0]/NET0131  , \InstQueue_reg[9][1]/NET0131  , \InstQueue_reg[9][2]/NET0131  , \InstQueue_reg[9][3]/NET0131  , \InstQueue_reg[9][4]/NET0131  , \InstQueue_reg[9][5]/NET0131  , \InstQueue_reg[9][6]/NET0131  , \InstQueue_reg[9][7]/NET0131  , M_IO_n_pad , \MemoryFetch_reg/NET0131  , \More_reg/NET0131  , NA_n_pad , \PhyAddrPointer_reg[0]/NET0131  , \PhyAddrPointer_reg[10]/NET0131  , \PhyAddrPointer_reg[11]/NET0131  , \PhyAddrPointer_reg[12]/NET0131  , \PhyAddrPointer_reg[13]/NET0131  , \PhyAddrPointer_reg[14]/NET0131  , \PhyAddrPointer_reg[15]/NET0131  , \PhyAddrPointer_reg[16]/NET0131  , \PhyAddrPointer_reg[17]/NET0131  , \PhyAddrPointer_reg[18]/NET0131  , \PhyAddrPointer_reg[19]/NET0131  , \PhyAddrPointer_reg[1]/NET0131  , \PhyAddrPointer_reg[20]/NET0131  , \PhyAddrPointer_reg[21]/NET0131  , \PhyAddrPointer_reg[22]/NET0131  , \PhyAddrPointer_reg[23]/NET0131  , \PhyAddrPointer_reg[24]/NET0131  , \PhyAddrPointer_reg[25]/NET0131  , \PhyAddrPointer_reg[26]/NET0131  , \PhyAddrPointer_reg[27]/NET0131  , \PhyAddrPointer_reg[28]/NET0131  , \PhyAddrPointer_reg[29]/NET0131  , \PhyAddrPointer_reg[2]/NET0131  , \PhyAddrPointer_reg[30]/NET0131  , \PhyAddrPointer_reg[31]/NET0131  , \PhyAddrPointer_reg[3]/NET0131  , \PhyAddrPointer_reg[4]/NET0131  , \PhyAddrPointer_reg[5]/NET0131  , \PhyAddrPointer_reg[6]/NET0131  , \PhyAddrPointer_reg[7]/NET0131  , \PhyAddrPointer_reg[8]/NET0131  , \PhyAddrPointer_reg[9]/NET0131  , READY_n_pad , \ReadRequest_reg/NET0131  , \RequestPending_reg/NET0131  , \State2_reg[0]/NET0131  , \State2_reg[1]/NET0131  , \State2_reg[2]/NET0131  , \State2_reg[3]/NET0131  , \State_reg[0]/NET0131  , \State_reg[1]/NET0131  , \State_reg[2]/NET0131  , W_R_n_pad , \lWord_reg[0]/NET0131  , \lWord_reg[10]/NET0131  , \lWord_reg[11]/NET0131  , \lWord_reg[12]/NET0131  , \lWord_reg[13]/NET0131  , \lWord_reg[14]/NET0131  , \lWord_reg[15]/NET0131  , \lWord_reg[1]/NET0131  , \lWord_reg[2]/NET0131  , \lWord_reg[3]/NET0131  , \lWord_reg[4]/NET0131  , \lWord_reg[5]/NET0131  , \lWord_reg[6]/NET0131  , \lWord_reg[7]/NET0131  , \lWord_reg[8]/NET0131  , \lWord_reg[9]/NET0131  , \rEIP_reg[0]/NET0131  , \rEIP_reg[10]/NET0131  , \rEIP_reg[11]/NET0131  , \rEIP_reg[12]/NET0131  , \rEIP_reg[13]/NET0131  , \rEIP_reg[14]/NET0131  , \rEIP_reg[15]/NET0131  , \rEIP_reg[16]/NET0131  , \rEIP_reg[17]/NET0131  , \rEIP_reg[18]/NET0131  , \rEIP_reg[19]/NET0131  , \rEIP_reg[1]/NET0131  , \rEIP_reg[20]/NET0131  , \rEIP_reg[21]/NET0131  , \rEIP_reg[22]/NET0131  , \rEIP_reg[23]/NET0131  , \rEIP_reg[24]/NET0131  , \rEIP_reg[25]/NET0131  , \rEIP_reg[26]/NET0131  , \rEIP_reg[27]/NET0131  , \rEIP_reg[28]/NET0131  , \rEIP_reg[29]/NET0131  , \rEIP_reg[2]/NET0131  , \rEIP_reg[30]/NET0131  , \rEIP_reg[31]/NET0131  , \rEIP_reg[3]/NET0131  , \rEIP_reg[4]/NET0131  , \rEIP_reg[5]/NET0131  , \rEIP_reg[6]/NET0131  , \rEIP_reg[7]/NET0131  , \rEIP_reg[8]/NET0131  , \rEIP_reg[9]/NET0131  , \uWord_reg[0]/NET0131  , \uWord_reg[10]/NET0131  , \uWord_reg[11]/NET0131  , \uWord_reg[12]/NET0131  , \uWord_reg[13]/NET0131  , \uWord_reg[14]/NET0131  , \uWord_reg[1]/NET0131  , \uWord_reg[2]/NET0131  , \uWord_reg[3]/NET0131  , \uWord_reg[4]/NET0131  , \uWord_reg[5]/NET0131  , \uWord_reg[6]/NET0131  , \uWord_reg[7]/NET0131  , \uWord_reg[8]/NET0131  , \uWord_reg[9]/NET0131  , \_al_n0  , \_al_n1  , \g47406/_2_  , \g47407/_2_  , \g47411/_0_  , \g47413/_0_  , \g47424/_0_  , \g47434/_0_  , \g47437/_0_  , \g47447/_2_  , \g47448/_0_  , \g47451/_0_  , \g47452/_0_  , \g47453/_0_  , \g47465/_2_  , \g47466/_0_  , \g47467/_0_  , \g47471/_0_  , \g47485/_0_  , \g47486/_0_  , \g47487/_2_  , \g47488/_0_  , \g47489/_2_  , \g47491/_0_  , \g47494/_0_  , \g47510/_0_  , \g47511/_0_  , \g47512/_0_  , \g47515/_0_  , \g47516/_0_  , \g47517/_2_  , \g47524/_0_  , \g47525/_0_  , \g47550/_0_  , \g47551/_2_  , \g47552/_0_  , \g47554/_0_  , \g47555/_0_  , \g47556/_0_  , \g47558/_0_  , \g47563/_0_  , \g47564/_0_  , \g47565/_0_  , \g47584/_0_  , \g47592/_0_  , \g47597/_0_  , \g47598/_0_  , \g47601/_0_  , \g47602/_0_  , \g47603/_0_  , \g47604/_0_  , \g47606/_0_  , \g47630/_0_  , \g47636/_0_  , \g47641/_0_  , \g47642/_0_  , \g47643/_0_  , \g47644/_0_  , \g47645/_0_  , \g47646/_0_  , \g47648/_0_  , \g47679/_0_  , \g47680/_0_  , \g47681/_0_  , \g47683/_0_  , \g47687/_0_  , \g47690/_0_  , \g47746/_0_  , \g47747/_0_  , \g47754/_0_  , \g47756/_0_  , \g47804/_0_  , \g47805/_0_  , \g47806/_0_  , \g47807/_0_  , \g47809/_0_  , \g47810/_0_  , \g47812/_0_  , \g47813/_0_  , \g47814/_0_  , \g47815/_0_  , \g47816/_0_  , \g47817/_0_  , \g47818/_0_  , \g47819/_0_  , \g47820/_0_  , \g47821/_0_  , \g47836/_0_  , \g47848/_0_  , \g47851/_0_  , \g47852/_0_  , \g47943/_0_  , \g47944/_0_  , \g47945/_0_  , \g47946/_0_  , \g47947/_0_  , \g47949/_0_  , \g47950/_0_  , \g47952/_0_  , \g47953/_0_  , \g47954/_0_  , \g47955/_0_  , \g47956/_0_  , \g47957/_0_  , \g47958/_0_  , \g47959/_0_  , \g47960/_0_  , \g47999/_0_  , \g48/_0_  , \g48005/_0_  , \g48006/_0_  , \g48007/_0_  , \g48008/_0_  , \g48009/_0_  , \g48010/_0_  , \g48011/_0_  , \g48012/_0_  , \g48013/_0_  , \g48014/_0_  , \g48015/_0_  , \g48057/_0_  , \g48058/_0_  , \g48059/_0_  , \g48060/_0_  , \g48061/_0_  , \g48062/_0_  , \g48063/_0_  , \g48064/_0_  , \g48066/_0_  , \g48067/_0_  , \g48068/_0_  , \g48069/_0_  , \g48070/_0_  , \g48071/_0_  , \g48073/_0_  , \g48074/_0_  , \g48075/_0_  , \g48076/_0_  , \g48077/_0_  , \g48078/_0_  , \g48079/_0_  , \g48080/_0_  , \g48081/_0_  , \g48082/_0_  , \g48084/_0_  , \g48085/_0_  , \g48086/_0_  , \g48087/_0_  , \g48089/_0_  , \g48090/_0_  , \g48091/_0_  , \g48093/_0_  , \g48094/_0_  , \g48119/_0_  , \g48120/_0_  , \g48121/_0_  , \g48122/_0_  , \g48123/_0_  , \g48124/_0_  , \g48125/_0_  , \g48126/_0_  , \g48127/_0_  , \g48128/_0_  , \g48129/_0_  , \g48130/_0_  , \g48131/_0_  , \g48132/_0_  , \g48133/_0_  , \g48134/_0_  , \g48135/_0_  , \g48136/_0_  , \g48137/_0_  , \g48138/_0_  , \g48140/_0_  , \g48144/_0_  , \g48145/_0_  , \g48146/_0_  , \g48147/_0_  , \g48148/_0_  , \g48150/_0_  , \g48151/_0_  , \g48152/_0_  , \g48153/_0_  , \g48154/_0_  , \g48176/_0_  , \g48189/_0_  , \g48192/_0_  , \g48193/_0_  , \g48194/_0_  , \g48195/_0_  , \g48196/_0_  , \g48197/_0_  , \g48198/_0_  , \g48199/_0_  , \g48200/_0_  , \g48263/_0_  , \g48265/_0_  , \g48273/_0_  , \g48313/_0_  , \g48318/_0_  , \g48319/_0_  , \g48321/_0_  , \g48323/_0_  , \g48324/_0_  , \g48325/_0_  , \g48326/_0_  , \g48327/_0_  , \g48328/_0_  , \g48329/_0_  , \g48330/_0_  , \g48331/_0_  , \g48332/_0_  , \g48333/_0_  , \g48472/_0_  , \g48519/_0_  , \g48520/_0_  , \g48521/_0_  , \g48522/_0_  , \g48523/_0_  , \g48524/_0_  , \g48525/_0_  , \g48527/_0_  , \g48529/_0_  , \g48530/_0_  , \g48531/_0_  , \g48532/_0_  , \g48533/_0_  , \g48534/_0_  , \g48535/_0_  , \g48536/_0_  , \g48537/_0_  , \g48538/_0_  , \g48539/_0_  , \g48540/_0_  , \g48541/_0_  , \g48542/_0_  , \g48543/_0_  , \g48545/_0_  , \g48546/_0_  , \g48547/_0_  , \g48639/_0_  , \g48642/_0_  , \g48645/_0_  , \g48648/_0_  , \g48652/_0_  , \g48655/_0_  , \g48658/_0_  , \g48661/_0_  , \g48664/_0_  , \g48667/_0_  , \g48670/_0_  , \g48673/_0_  , \g48678/_0_  , \g48681/_0_  , \g48684/_0_  , \g48688/_0_  , \g48793/_0_  , \g48812/_0_  , \g48813/_0_  , \g48814/_0_  , \g48824/_0_  , \g48825/_0_  , \g48826/_0_  , \g48827/_0_  , \g48828/_0_  , \g48829/_0_  , \g48830/_0_  , \g48831/_0_  , \g48833/_0_  , \g48834/_0_  , \g48835/_0_  , \g48836/_0_  , \g48837/_0_  , \g48838/_0_  , \g48839/_0_  , \g48840/_0_  , \g48841/_0_  , \g48842/_0_  , \g48843/_0_  , \g48844/_0_  , \g48845/_0_  , \g48846/_0_  , \g48847/_0_  , \g48848/_0_  , \g48908/_0_  , \g48909/_0_  , \g48910/_0_  , \g48912/_0_  , \g48913/_0_  , \g48915/_0_  , \g48917/_0_  , \g48932/_0_  , \g48933/_0_  , \g48935/_0_  , \g48937/_0_  , \g48938/_0_  , \g48939/_0_  , \g48940/_0_  , \g48942/_0_  , \g48945/_0_  , \g48971/_0_  , \g49007/_0_  , \g49047/_0_  , \g49048/_0_  , \g49050/_0_  , \g49182/_0_  , \g49280/_0_  , \g49332/_0_  , \g49335/_0_  , \g49336/_0_  , \g49337/_0_  , \g49338/_0_  , \g49339/_0_  , \g49340/_0_  , \g49341/_0_  , \g49342/_0_  , \g49343/_0_  , \g49344/_0_  , \g49345/_0_  , \g49346/_0_  , \g49347/_0_  , \g49348/_0_  , \g49349/_0_  , \g49356/_0_  , \g49375/_0_  , \g49396/_0_  , \g49397/_0_  , \g49400/_0_  , \g49404/_0_  , \g49406/_0_  , \g49414/_0_  , \g49422/_0_  , \g49426/_0_  , \g49430/_0_  , \g49434/_0_  , \g49437/_0_  , \g49440/_0_  , \g49441/_0_  , \g49444/_0_  , \g49448/_0_  , \g49451/_0_  , \g49455/_0_  , \g49456/_0_  , \g49460/_0_  , \g49466/_0_  , \g49563/_0_  , \g49592/_0_  , \g49915/_0_  , \g49941/_0_  , \g50023/_0_  , \g50026/_0_  , \g50029/_0_  , \g50031/_0_  , \g50033/_0_  , \g50035/_0_  , \g50037/_0_  , \g50040/_0_  , \g50050/_0_  , \g50056/_0_  , \g50059/_0_  , \g50065/_0_  , \g50067/_0_  , \g50150/_0_  , \g50283/_0_  , \g50284/_0_  , \g50501/_0_  , \g50594/_0_  , \g50807/_0_  , \g50866/_0_  , \g50875/_0_  , \g51449/_0_  , \g51510/_0_  , \g51534/_0_  , \g52310/_0_  , \g53066/_0_  , \g53087/_0_  , \g53151/_0_  , \g53608/_0_  , \g53634/_0_  , \g54053/_0_  , \g54091/_0_  , \g54103/_0_  , \g54268/_0_  , \g54277/_0_  , \g54287/_0_  , \g54294/_0_  , \g54449/_0_  , \g54453/_0_  , \g54484/_0_  , \g54528/_0_  , \g54582/_0_  , \g55448/_0_  , \g55693/_1_  , \g55874/_0_  , \g56203/_0_  , \g56303/_0_  , \g56329/_0_  , \g56336/_0_  , \g56345/_0_  , \g56367/_0_  , \g56411/_0_  , \g56529/_0_  , \g56858/_0_  , \g60443/_1_  , \g63395/_0_  , \g63442/_0_  , \g63595/_0_  , \g63996/_0_  , \g64048/_0_  , \g64071/_0_  , \g64085/_0_  , \g64096/_0_  , \g64119/_0_  , \g64216/_0_  , \g64513/_0_  , \g64566/_0_  , \g64694/_0_  , \g64913/_0_  );
  input ADS_n_pad ;
  input \Address[0]_pad  ;
  input \Address[10]_pad  ;
  input \Address[11]_pad  ;
  input \Address[12]_pad  ;
  input \Address[13]_pad  ;
  input \Address[14]_pad  ;
  input \Address[15]_pad  ;
  input \Address[16]_pad  ;
  input \Address[17]_pad  ;
  input \Address[18]_pad  ;
  input \Address[19]_pad  ;
  input \Address[1]_pad  ;
  input \Address[20]_pad  ;
  input \Address[21]_pad  ;
  input \Address[22]_pad  ;
  input \Address[23]_pad  ;
  input \Address[24]_pad  ;
  input \Address[25]_pad  ;
  input \Address[26]_pad  ;
  input \Address[27]_pad  ;
  input \Address[28]_pad  ;
  input \Address[29]_pad  ;
  input \Address[2]_pad  ;
  input \Address[3]_pad  ;
  input \Address[4]_pad  ;
  input \Address[5]_pad  ;
  input \Address[6]_pad  ;
  input \Address[7]_pad  ;
  input \Address[8]_pad  ;
  input \Address[9]_pad  ;
  input \BE_n[0]_pad  ;
  input \BE_n[1]_pad  ;
  input \BE_n[2]_pad  ;
  input \BE_n[3]_pad  ;
  input \BS16_n_pad  ;
  input \ByteEnable_reg[0]/NET0131  ;
  input \ByteEnable_reg[1]/NET0131  ;
  input \ByteEnable_reg[2]/NET0131  ;
  input \ByteEnable_reg[3]/NET0131  ;
  input \CodeFetch_reg/NET0131  ;
  input D_C_n_pad ;
  input \DataWidth_reg[0]/NET0131  ;
  input \DataWidth_reg[1]/NET0131  ;
  input \Datai[0]_pad  ;
  input \Datai[10]_pad  ;
  input \Datai[11]_pad  ;
  input \Datai[12]_pad  ;
  input \Datai[13]_pad  ;
  input \Datai[14]_pad  ;
  input \Datai[15]_pad  ;
  input \Datai[16]_pad  ;
  input \Datai[17]_pad  ;
  input \Datai[18]_pad  ;
  input \Datai[19]_pad  ;
  input \Datai[1]_pad  ;
  input \Datai[20]_pad  ;
  input \Datai[21]_pad  ;
  input \Datai[22]_pad  ;
  input \Datai[23]_pad  ;
  input \Datai[24]_pad  ;
  input \Datai[25]_pad  ;
  input \Datai[26]_pad  ;
  input \Datai[27]_pad  ;
  input \Datai[28]_pad  ;
  input \Datai[29]_pad  ;
  input \Datai[2]_pad  ;
  input \Datai[30]_pad  ;
  input \Datai[31]_pad  ;
  input \Datai[3]_pad  ;
  input \Datai[4]_pad  ;
  input \Datai[5]_pad  ;
  input \Datai[6]_pad  ;
  input \Datai[7]_pad  ;
  input \Datai[8]_pad  ;
  input \Datai[9]_pad  ;
  input \Datao[0]_pad  ;
  input \Datao[10]_pad  ;
  input \Datao[11]_pad  ;
  input \Datao[12]_pad  ;
  input \Datao[13]_pad  ;
  input \Datao[14]_pad  ;
  input \Datao[15]_pad  ;
  input \Datao[16]_pad  ;
  input \Datao[17]_pad  ;
  input \Datao[18]_pad  ;
  input \Datao[19]_pad  ;
  input \Datao[1]_pad  ;
  input \Datao[20]_pad  ;
  input \Datao[21]_pad  ;
  input \Datao[22]_pad  ;
  input \Datao[23]_pad  ;
  input \Datao[24]_pad  ;
  input \Datao[25]_pad  ;
  input \Datao[26]_pad  ;
  input \Datao[27]_pad  ;
  input \Datao[28]_pad  ;
  input \Datao[29]_pad  ;
  input \Datao[2]_pad  ;
  input \Datao[30]_pad  ;
  input \Datao[3]_pad  ;
  input \Datao[4]_pad  ;
  input \Datao[5]_pad  ;
  input \Datao[6]_pad  ;
  input \Datao[7]_pad  ;
  input \Datao[8]_pad  ;
  input \Datao[9]_pad  ;
  input \EAX_reg[0]/NET0131  ;
  input \EAX_reg[10]/NET0131  ;
  input \EAX_reg[11]/NET0131  ;
  input \EAX_reg[12]/NET0131  ;
  input \EAX_reg[13]/NET0131  ;
  input \EAX_reg[14]/NET0131  ;
  input \EAX_reg[15]/NET0131  ;
  input \EAX_reg[16]/NET0131  ;
  input \EAX_reg[17]/NET0131  ;
  input \EAX_reg[18]/NET0131  ;
  input \EAX_reg[19]/NET0131  ;
  input \EAX_reg[1]/NET0131  ;
  input \EAX_reg[20]/NET0131  ;
  input \EAX_reg[21]/NET0131  ;
  input \EAX_reg[22]/NET0131  ;
  input \EAX_reg[23]/NET0131  ;
  input \EAX_reg[24]/NET0131  ;
  input \EAX_reg[25]/NET0131  ;
  input \EAX_reg[26]/NET0131  ;
  input \EAX_reg[27]/NET0131  ;
  input \EAX_reg[28]/NET0131  ;
  input \EAX_reg[29]/NET0131  ;
  input \EAX_reg[2]/NET0131  ;
  input \EAX_reg[30]/NET0131  ;
  input \EAX_reg[31]/NET0131  ;
  input \EAX_reg[3]/NET0131  ;
  input \EAX_reg[4]/NET0131  ;
  input \EAX_reg[5]/NET0131  ;
  input \EAX_reg[6]/NET0131  ;
  input \EAX_reg[7]/NET0131  ;
  input \EAX_reg[8]/NET0131  ;
  input \EAX_reg[9]/NET0131  ;
  input \EBX_reg[0]/NET0131  ;
  input \EBX_reg[10]/NET0131  ;
  input \EBX_reg[11]/NET0131  ;
  input \EBX_reg[12]/NET0131  ;
  input \EBX_reg[13]/NET0131  ;
  input \EBX_reg[14]/NET0131  ;
  input \EBX_reg[15]/NET0131  ;
  input \EBX_reg[16]/NET0131  ;
  input \EBX_reg[17]/NET0131  ;
  input \EBX_reg[18]/NET0131  ;
  input \EBX_reg[19]/NET0131  ;
  input \EBX_reg[1]/NET0131  ;
  input \EBX_reg[20]/NET0131  ;
  input \EBX_reg[21]/NET0131  ;
  input \EBX_reg[22]/NET0131  ;
  input \EBX_reg[23]/NET0131  ;
  input \EBX_reg[24]/NET0131  ;
  input \EBX_reg[25]/NET0131  ;
  input \EBX_reg[26]/NET0131  ;
  input \EBX_reg[27]/NET0131  ;
  input \EBX_reg[28]/NET0131  ;
  input \EBX_reg[29]/NET0131  ;
  input \EBX_reg[2]/NET0131  ;
  input \EBX_reg[30]/NET0131  ;
  input \EBX_reg[31]/NET0131  ;
  input \EBX_reg[3]/NET0131  ;
  input \EBX_reg[4]/NET0131  ;
  input \EBX_reg[5]/NET0131  ;
  input \EBX_reg[6]/NET0131  ;
  input \EBX_reg[7]/NET0131  ;
  input \EBX_reg[8]/NET0131  ;
  input \EBX_reg[9]/NET0131  ;
  input \Flush_reg/NET0131  ;
  input HOLD_pad ;
  input \InstAddrPointer_reg[0]/NET0131  ;
  input \InstAddrPointer_reg[10]/NET0131  ;
  input \InstAddrPointer_reg[11]/NET0131  ;
  input \InstAddrPointer_reg[12]/NET0131  ;
  input \InstAddrPointer_reg[13]/NET0131  ;
  input \InstAddrPointer_reg[14]/NET0131  ;
  input \InstAddrPointer_reg[15]/NET0131  ;
  input \InstAddrPointer_reg[16]/NET0131  ;
  input \InstAddrPointer_reg[17]/NET0131  ;
  input \InstAddrPointer_reg[18]/NET0131  ;
  input \InstAddrPointer_reg[19]/NET0131  ;
  input \InstAddrPointer_reg[1]/NET0131  ;
  input \InstAddrPointer_reg[20]/NET0131  ;
  input \InstAddrPointer_reg[21]/NET0131  ;
  input \InstAddrPointer_reg[22]/NET0131  ;
  input \InstAddrPointer_reg[23]/NET0131  ;
  input \InstAddrPointer_reg[24]/NET0131  ;
  input \InstAddrPointer_reg[25]/NET0131  ;
  input \InstAddrPointer_reg[26]/NET0131  ;
  input \InstAddrPointer_reg[27]/NET0131  ;
  input \InstAddrPointer_reg[28]/NET0131  ;
  input \InstAddrPointer_reg[29]/NET0131  ;
  input \InstAddrPointer_reg[2]/NET0131  ;
  input \InstAddrPointer_reg[30]/NET0131  ;
  input \InstAddrPointer_reg[31]/NET0131  ;
  input \InstAddrPointer_reg[3]/NET0131  ;
  input \InstAddrPointer_reg[4]/NET0131  ;
  input \InstAddrPointer_reg[5]/NET0131  ;
  input \InstAddrPointer_reg[6]/NET0131  ;
  input \InstAddrPointer_reg[7]/NET0131  ;
  input \InstAddrPointer_reg[8]/NET0131  ;
  input \InstAddrPointer_reg[9]/NET0131  ;
  input \InstQueueRd_Addr_reg[0]/NET0131  ;
  input \InstQueueRd_Addr_reg[1]/NET0131  ;
  input \InstQueueRd_Addr_reg[2]/NET0131  ;
  input \InstQueueRd_Addr_reg[3]/NET0131  ;
  input \InstQueueWr_Addr_reg[0]/NET0131  ;
  input \InstQueueWr_Addr_reg[1]/NET0131  ;
  input \InstQueueWr_Addr_reg[2]/NET0131  ;
  input \InstQueueWr_Addr_reg[3]/NET0131  ;
  input \InstQueue_reg[0][0]/NET0131  ;
  input \InstQueue_reg[0][1]/NET0131  ;
  input \InstQueue_reg[0][2]/NET0131  ;
  input \InstQueue_reg[0][3]/NET0131  ;
  input \InstQueue_reg[0][4]/NET0131  ;
  input \InstQueue_reg[0][5]/NET0131  ;
  input \InstQueue_reg[0][6]/NET0131  ;
  input \InstQueue_reg[0][7]/NET0131  ;
  input \InstQueue_reg[10][0]/NET0131  ;
  input \InstQueue_reg[10][1]/NET0131  ;
  input \InstQueue_reg[10][2]/NET0131  ;
  input \InstQueue_reg[10][3]/NET0131  ;
  input \InstQueue_reg[10][4]/NET0131  ;
  input \InstQueue_reg[10][5]/NET0131  ;
  input \InstQueue_reg[10][6]/NET0131  ;
  input \InstQueue_reg[10][7]/NET0131  ;
  input \InstQueue_reg[11][0]/NET0131  ;
  input \InstQueue_reg[11][1]/NET0131  ;
  input \InstQueue_reg[11][2]/NET0131  ;
  input \InstQueue_reg[11][3]/NET0131  ;
  input \InstQueue_reg[11][4]/NET0131  ;
  input \InstQueue_reg[11][5]/NET0131  ;
  input \InstQueue_reg[11][6]/NET0131  ;
  input \InstQueue_reg[11][7]/NET0131  ;
  input \InstQueue_reg[12][0]/NET0131  ;
  input \InstQueue_reg[12][1]/NET0131  ;
  input \InstQueue_reg[12][2]/NET0131  ;
  input \InstQueue_reg[12][3]/NET0131  ;
  input \InstQueue_reg[12][4]/NET0131  ;
  input \InstQueue_reg[12][5]/NET0131  ;
  input \InstQueue_reg[12][6]/NET0131  ;
  input \InstQueue_reg[12][7]/NET0131  ;
  input \InstQueue_reg[13][0]/NET0131  ;
  input \InstQueue_reg[13][1]/NET0131  ;
  input \InstQueue_reg[13][2]/NET0131  ;
  input \InstQueue_reg[13][3]/NET0131  ;
  input \InstQueue_reg[13][4]/NET0131  ;
  input \InstQueue_reg[13][5]/NET0131  ;
  input \InstQueue_reg[13][6]/NET0131  ;
  input \InstQueue_reg[13][7]/NET0131  ;
  input \InstQueue_reg[14][0]/NET0131  ;
  input \InstQueue_reg[14][1]/NET0131  ;
  input \InstQueue_reg[14][2]/NET0131  ;
  input \InstQueue_reg[14][3]/NET0131  ;
  input \InstQueue_reg[14][4]/NET0131  ;
  input \InstQueue_reg[14][5]/NET0131  ;
  input \InstQueue_reg[14][6]/NET0131  ;
  input \InstQueue_reg[14][7]/NET0131  ;
  input \InstQueue_reg[15][0]/NET0131  ;
  input \InstQueue_reg[15][1]/NET0131  ;
  input \InstQueue_reg[15][2]/NET0131  ;
  input \InstQueue_reg[15][3]/NET0131  ;
  input \InstQueue_reg[15][4]/NET0131  ;
  input \InstQueue_reg[15][5]/NET0131  ;
  input \InstQueue_reg[15][6]/NET0131  ;
  input \InstQueue_reg[15][7]/NET0131  ;
  input \InstQueue_reg[1][0]/NET0131  ;
  input \InstQueue_reg[1][1]/NET0131  ;
  input \InstQueue_reg[1][2]/NET0131  ;
  input \InstQueue_reg[1][3]/NET0131  ;
  input \InstQueue_reg[1][4]/NET0131  ;
  input \InstQueue_reg[1][5]/NET0131  ;
  input \InstQueue_reg[1][6]/NET0131  ;
  input \InstQueue_reg[1][7]/NET0131  ;
  input \InstQueue_reg[2][0]/NET0131  ;
  input \InstQueue_reg[2][1]/NET0131  ;
  input \InstQueue_reg[2][2]/NET0131  ;
  input \InstQueue_reg[2][3]/NET0131  ;
  input \InstQueue_reg[2][4]/NET0131  ;
  input \InstQueue_reg[2][5]/NET0131  ;
  input \InstQueue_reg[2][6]/NET0131  ;
  input \InstQueue_reg[2][7]/NET0131  ;
  input \InstQueue_reg[3][0]/NET0131  ;
  input \InstQueue_reg[3][1]/NET0131  ;
  input \InstQueue_reg[3][2]/NET0131  ;
  input \InstQueue_reg[3][3]/NET0131  ;
  input \InstQueue_reg[3][4]/NET0131  ;
  input \InstQueue_reg[3][5]/NET0131  ;
  input \InstQueue_reg[3][6]/NET0131  ;
  input \InstQueue_reg[3][7]/NET0131  ;
  input \InstQueue_reg[4][0]/NET0131  ;
  input \InstQueue_reg[4][1]/NET0131  ;
  input \InstQueue_reg[4][2]/NET0131  ;
  input \InstQueue_reg[4][3]/NET0131  ;
  input \InstQueue_reg[4][4]/NET0131  ;
  input \InstQueue_reg[4][5]/NET0131  ;
  input \InstQueue_reg[4][6]/NET0131  ;
  input \InstQueue_reg[4][7]/NET0131  ;
  input \InstQueue_reg[5][0]/NET0131  ;
  input \InstQueue_reg[5][1]/NET0131  ;
  input \InstQueue_reg[5][2]/NET0131  ;
  input \InstQueue_reg[5][3]/NET0131  ;
  input \InstQueue_reg[5][4]/NET0131  ;
  input \InstQueue_reg[5][5]/NET0131  ;
  input \InstQueue_reg[5][6]/NET0131  ;
  input \InstQueue_reg[5][7]/NET0131  ;
  input \InstQueue_reg[6][0]/NET0131  ;
  input \InstQueue_reg[6][1]/NET0131  ;
  input \InstQueue_reg[6][2]/NET0131  ;
  input \InstQueue_reg[6][3]/NET0131  ;
  input \InstQueue_reg[6][4]/NET0131  ;
  input \InstQueue_reg[6][5]/NET0131  ;
  input \InstQueue_reg[6][6]/NET0131  ;
  input \InstQueue_reg[6][7]/NET0131  ;
  input \InstQueue_reg[7][0]/NET0131  ;
  input \InstQueue_reg[7][1]/NET0131  ;
  input \InstQueue_reg[7][2]/NET0131  ;
  input \InstQueue_reg[7][3]/NET0131  ;
  input \InstQueue_reg[7][4]/NET0131  ;
  input \InstQueue_reg[7][5]/NET0131  ;
  input \InstQueue_reg[7][6]/NET0131  ;
  input \InstQueue_reg[7][7]/NET0131  ;
  input \InstQueue_reg[8][0]/NET0131  ;
  input \InstQueue_reg[8][1]/NET0131  ;
  input \InstQueue_reg[8][2]/NET0131  ;
  input \InstQueue_reg[8][3]/NET0131  ;
  input \InstQueue_reg[8][4]/NET0131  ;
  input \InstQueue_reg[8][5]/NET0131  ;
  input \InstQueue_reg[8][6]/NET0131  ;
  input \InstQueue_reg[8][7]/NET0131  ;
  input \InstQueue_reg[9][0]/NET0131  ;
  input \InstQueue_reg[9][1]/NET0131  ;
  input \InstQueue_reg[9][2]/NET0131  ;
  input \InstQueue_reg[9][3]/NET0131  ;
  input \InstQueue_reg[9][4]/NET0131  ;
  input \InstQueue_reg[9][5]/NET0131  ;
  input \InstQueue_reg[9][6]/NET0131  ;
  input \InstQueue_reg[9][7]/NET0131  ;
  input M_IO_n_pad ;
  input \MemoryFetch_reg/NET0131  ;
  input \More_reg/NET0131  ;
  input NA_n_pad ;
  input \PhyAddrPointer_reg[0]/NET0131  ;
  input \PhyAddrPointer_reg[10]/NET0131  ;
  input \PhyAddrPointer_reg[11]/NET0131  ;
  input \PhyAddrPointer_reg[12]/NET0131  ;
  input \PhyAddrPointer_reg[13]/NET0131  ;
  input \PhyAddrPointer_reg[14]/NET0131  ;
  input \PhyAddrPointer_reg[15]/NET0131  ;
  input \PhyAddrPointer_reg[16]/NET0131  ;
  input \PhyAddrPointer_reg[17]/NET0131  ;
  input \PhyAddrPointer_reg[18]/NET0131  ;
  input \PhyAddrPointer_reg[19]/NET0131  ;
  input \PhyAddrPointer_reg[1]/NET0131  ;
  input \PhyAddrPointer_reg[20]/NET0131  ;
  input \PhyAddrPointer_reg[21]/NET0131  ;
  input \PhyAddrPointer_reg[22]/NET0131  ;
  input \PhyAddrPointer_reg[23]/NET0131  ;
  input \PhyAddrPointer_reg[24]/NET0131  ;
  input \PhyAddrPointer_reg[25]/NET0131  ;
  input \PhyAddrPointer_reg[26]/NET0131  ;
  input \PhyAddrPointer_reg[27]/NET0131  ;
  input \PhyAddrPointer_reg[28]/NET0131  ;
  input \PhyAddrPointer_reg[29]/NET0131  ;
  input \PhyAddrPointer_reg[2]/NET0131  ;
  input \PhyAddrPointer_reg[30]/NET0131  ;
  input \PhyAddrPointer_reg[31]/NET0131  ;
  input \PhyAddrPointer_reg[3]/NET0131  ;
  input \PhyAddrPointer_reg[4]/NET0131  ;
  input \PhyAddrPointer_reg[5]/NET0131  ;
  input \PhyAddrPointer_reg[6]/NET0131  ;
  input \PhyAddrPointer_reg[7]/NET0131  ;
  input \PhyAddrPointer_reg[8]/NET0131  ;
  input \PhyAddrPointer_reg[9]/NET0131  ;
  input READY_n_pad ;
  input \ReadRequest_reg/NET0131  ;
  input \RequestPending_reg/NET0131  ;
  input \State2_reg[0]/NET0131  ;
  input \State2_reg[1]/NET0131  ;
  input \State2_reg[2]/NET0131  ;
  input \State2_reg[3]/NET0131  ;
  input \State_reg[0]/NET0131  ;
  input \State_reg[1]/NET0131  ;
  input \State_reg[2]/NET0131  ;
  input W_R_n_pad ;
  input \lWord_reg[0]/NET0131  ;
  input \lWord_reg[10]/NET0131  ;
  input \lWord_reg[11]/NET0131  ;
  input \lWord_reg[12]/NET0131  ;
  input \lWord_reg[13]/NET0131  ;
  input \lWord_reg[14]/NET0131  ;
  input \lWord_reg[15]/NET0131  ;
  input \lWord_reg[1]/NET0131  ;
  input \lWord_reg[2]/NET0131  ;
  input \lWord_reg[3]/NET0131  ;
  input \lWord_reg[4]/NET0131  ;
  input \lWord_reg[5]/NET0131  ;
  input \lWord_reg[6]/NET0131  ;
  input \lWord_reg[7]/NET0131  ;
  input \lWord_reg[8]/NET0131  ;
  input \lWord_reg[9]/NET0131  ;
  input \rEIP_reg[0]/NET0131  ;
  input \rEIP_reg[10]/NET0131  ;
  input \rEIP_reg[11]/NET0131  ;
  input \rEIP_reg[12]/NET0131  ;
  input \rEIP_reg[13]/NET0131  ;
  input \rEIP_reg[14]/NET0131  ;
  input \rEIP_reg[15]/NET0131  ;
  input \rEIP_reg[16]/NET0131  ;
  input \rEIP_reg[17]/NET0131  ;
  input \rEIP_reg[18]/NET0131  ;
  input \rEIP_reg[19]/NET0131  ;
  input \rEIP_reg[1]/NET0131  ;
  input \rEIP_reg[20]/NET0131  ;
  input \rEIP_reg[21]/NET0131  ;
  input \rEIP_reg[22]/NET0131  ;
  input \rEIP_reg[23]/NET0131  ;
  input \rEIP_reg[24]/NET0131  ;
  input \rEIP_reg[25]/NET0131  ;
  input \rEIP_reg[26]/NET0131  ;
  input \rEIP_reg[27]/NET0131  ;
  input \rEIP_reg[28]/NET0131  ;
  input \rEIP_reg[29]/NET0131  ;
  input \rEIP_reg[2]/NET0131  ;
  input \rEIP_reg[30]/NET0131  ;
  input \rEIP_reg[31]/NET0131  ;
  input \rEIP_reg[3]/NET0131  ;
  input \rEIP_reg[4]/NET0131  ;
  input \rEIP_reg[5]/NET0131  ;
  input \rEIP_reg[6]/NET0131  ;
  input \rEIP_reg[7]/NET0131  ;
  input \rEIP_reg[8]/NET0131  ;
  input \rEIP_reg[9]/NET0131  ;
  input \uWord_reg[0]/NET0131  ;
  input \uWord_reg[10]/NET0131  ;
  input \uWord_reg[11]/NET0131  ;
  input \uWord_reg[12]/NET0131  ;
  input \uWord_reg[13]/NET0131  ;
  input \uWord_reg[14]/NET0131  ;
  input \uWord_reg[1]/NET0131  ;
  input \uWord_reg[2]/NET0131  ;
  input \uWord_reg[3]/NET0131  ;
  input \uWord_reg[4]/NET0131  ;
  input \uWord_reg[5]/NET0131  ;
  input \uWord_reg[6]/NET0131  ;
  input \uWord_reg[7]/NET0131  ;
  input \uWord_reg[8]/NET0131  ;
  input \uWord_reg[9]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g47406/_2_  ;
  output \g47407/_2_  ;
  output \g47411/_0_  ;
  output \g47413/_0_  ;
  output \g47424/_0_  ;
  output \g47434/_0_  ;
  output \g47437/_0_  ;
  output \g47447/_2_  ;
  output \g47448/_0_  ;
  output \g47451/_0_  ;
  output \g47452/_0_  ;
  output \g47453/_0_  ;
  output \g47465/_2_  ;
  output \g47466/_0_  ;
  output \g47467/_0_  ;
  output \g47471/_0_  ;
  output \g47485/_0_  ;
  output \g47486/_0_  ;
  output \g47487/_2_  ;
  output \g47488/_0_  ;
  output \g47489/_2_  ;
  output \g47491/_0_  ;
  output \g47494/_0_  ;
  output \g47510/_0_  ;
  output \g47511/_0_  ;
  output \g47512/_0_  ;
  output \g47515/_0_  ;
  output \g47516/_0_  ;
  output \g47517/_2_  ;
  output \g47524/_0_  ;
  output \g47525/_0_  ;
  output \g47550/_0_  ;
  output \g47551/_2_  ;
  output \g47552/_0_  ;
  output \g47554/_0_  ;
  output \g47555/_0_  ;
  output \g47556/_0_  ;
  output \g47558/_0_  ;
  output \g47563/_0_  ;
  output \g47564/_0_  ;
  output \g47565/_0_  ;
  output \g47584/_0_  ;
  output \g47592/_0_  ;
  output \g47597/_0_  ;
  output \g47598/_0_  ;
  output \g47601/_0_  ;
  output \g47602/_0_  ;
  output \g47603/_0_  ;
  output \g47604/_0_  ;
  output \g47606/_0_  ;
  output \g47630/_0_  ;
  output \g47636/_0_  ;
  output \g47641/_0_  ;
  output \g47642/_0_  ;
  output \g47643/_0_  ;
  output \g47644/_0_  ;
  output \g47645/_0_  ;
  output \g47646/_0_  ;
  output \g47648/_0_  ;
  output \g47679/_0_  ;
  output \g47680/_0_  ;
  output \g47681/_0_  ;
  output \g47683/_0_  ;
  output \g47687/_0_  ;
  output \g47690/_0_  ;
  output \g47746/_0_  ;
  output \g47747/_0_  ;
  output \g47754/_0_  ;
  output \g47756/_0_  ;
  output \g47804/_0_  ;
  output \g47805/_0_  ;
  output \g47806/_0_  ;
  output \g47807/_0_  ;
  output \g47809/_0_  ;
  output \g47810/_0_  ;
  output \g47812/_0_  ;
  output \g47813/_0_  ;
  output \g47814/_0_  ;
  output \g47815/_0_  ;
  output \g47816/_0_  ;
  output \g47817/_0_  ;
  output \g47818/_0_  ;
  output \g47819/_0_  ;
  output \g47820/_0_  ;
  output \g47821/_0_  ;
  output \g47836/_0_  ;
  output \g47848/_0_  ;
  output \g47851/_0_  ;
  output \g47852/_0_  ;
  output \g47943/_0_  ;
  output \g47944/_0_  ;
  output \g47945/_0_  ;
  output \g47946/_0_  ;
  output \g47947/_0_  ;
  output \g47949/_0_  ;
  output \g47950/_0_  ;
  output \g47952/_0_  ;
  output \g47953/_0_  ;
  output \g47954/_0_  ;
  output \g47955/_0_  ;
  output \g47956/_0_  ;
  output \g47957/_0_  ;
  output \g47958/_0_  ;
  output \g47959/_0_  ;
  output \g47960/_0_  ;
  output \g47999/_0_  ;
  output \g48/_0_  ;
  output \g48005/_0_  ;
  output \g48006/_0_  ;
  output \g48007/_0_  ;
  output \g48008/_0_  ;
  output \g48009/_0_  ;
  output \g48010/_0_  ;
  output \g48011/_0_  ;
  output \g48012/_0_  ;
  output \g48013/_0_  ;
  output \g48014/_0_  ;
  output \g48015/_0_  ;
  output \g48057/_0_  ;
  output \g48058/_0_  ;
  output \g48059/_0_  ;
  output \g48060/_0_  ;
  output \g48061/_0_  ;
  output \g48062/_0_  ;
  output \g48063/_0_  ;
  output \g48064/_0_  ;
  output \g48066/_0_  ;
  output \g48067/_0_  ;
  output \g48068/_0_  ;
  output \g48069/_0_  ;
  output \g48070/_0_  ;
  output \g48071/_0_  ;
  output \g48073/_0_  ;
  output \g48074/_0_  ;
  output \g48075/_0_  ;
  output \g48076/_0_  ;
  output \g48077/_0_  ;
  output \g48078/_0_  ;
  output \g48079/_0_  ;
  output \g48080/_0_  ;
  output \g48081/_0_  ;
  output \g48082/_0_  ;
  output \g48084/_0_  ;
  output \g48085/_0_  ;
  output \g48086/_0_  ;
  output \g48087/_0_  ;
  output \g48089/_0_  ;
  output \g48090/_0_  ;
  output \g48091/_0_  ;
  output \g48093/_0_  ;
  output \g48094/_0_  ;
  output \g48119/_0_  ;
  output \g48120/_0_  ;
  output \g48121/_0_  ;
  output \g48122/_0_  ;
  output \g48123/_0_  ;
  output \g48124/_0_  ;
  output \g48125/_0_  ;
  output \g48126/_0_  ;
  output \g48127/_0_  ;
  output \g48128/_0_  ;
  output \g48129/_0_  ;
  output \g48130/_0_  ;
  output \g48131/_0_  ;
  output \g48132/_0_  ;
  output \g48133/_0_  ;
  output \g48134/_0_  ;
  output \g48135/_0_  ;
  output \g48136/_0_  ;
  output \g48137/_0_  ;
  output \g48138/_0_  ;
  output \g48140/_0_  ;
  output \g48144/_0_  ;
  output \g48145/_0_  ;
  output \g48146/_0_  ;
  output \g48147/_0_  ;
  output \g48148/_0_  ;
  output \g48150/_0_  ;
  output \g48151/_0_  ;
  output \g48152/_0_  ;
  output \g48153/_0_  ;
  output \g48154/_0_  ;
  output \g48176/_0_  ;
  output \g48189/_0_  ;
  output \g48192/_0_  ;
  output \g48193/_0_  ;
  output \g48194/_0_  ;
  output \g48195/_0_  ;
  output \g48196/_0_  ;
  output \g48197/_0_  ;
  output \g48198/_0_  ;
  output \g48199/_0_  ;
  output \g48200/_0_  ;
  output \g48263/_0_  ;
  output \g48265/_0_  ;
  output \g48273/_0_  ;
  output \g48313/_0_  ;
  output \g48318/_0_  ;
  output \g48319/_0_  ;
  output \g48321/_0_  ;
  output \g48323/_0_  ;
  output \g48324/_0_  ;
  output \g48325/_0_  ;
  output \g48326/_0_  ;
  output \g48327/_0_  ;
  output \g48328/_0_  ;
  output \g48329/_0_  ;
  output \g48330/_0_  ;
  output \g48331/_0_  ;
  output \g48332/_0_  ;
  output \g48333/_0_  ;
  output \g48472/_0_  ;
  output \g48519/_0_  ;
  output \g48520/_0_  ;
  output \g48521/_0_  ;
  output \g48522/_0_  ;
  output \g48523/_0_  ;
  output \g48524/_0_  ;
  output \g48525/_0_  ;
  output \g48527/_0_  ;
  output \g48529/_0_  ;
  output \g48530/_0_  ;
  output \g48531/_0_  ;
  output \g48532/_0_  ;
  output \g48533/_0_  ;
  output \g48534/_0_  ;
  output \g48535/_0_  ;
  output \g48536/_0_  ;
  output \g48537/_0_  ;
  output \g48538/_0_  ;
  output \g48539/_0_  ;
  output \g48540/_0_  ;
  output \g48541/_0_  ;
  output \g48542/_0_  ;
  output \g48543/_0_  ;
  output \g48545/_0_  ;
  output \g48546/_0_  ;
  output \g48547/_0_  ;
  output \g48639/_0_  ;
  output \g48642/_0_  ;
  output \g48645/_0_  ;
  output \g48648/_0_  ;
  output \g48652/_0_  ;
  output \g48655/_0_  ;
  output \g48658/_0_  ;
  output \g48661/_0_  ;
  output \g48664/_0_  ;
  output \g48667/_0_  ;
  output \g48670/_0_  ;
  output \g48673/_0_  ;
  output \g48678/_0_  ;
  output \g48681/_0_  ;
  output \g48684/_0_  ;
  output \g48688/_0_  ;
  output \g48793/_0_  ;
  output \g48812/_0_  ;
  output \g48813/_0_  ;
  output \g48814/_0_  ;
  output \g48824/_0_  ;
  output \g48825/_0_  ;
  output \g48826/_0_  ;
  output \g48827/_0_  ;
  output \g48828/_0_  ;
  output \g48829/_0_  ;
  output \g48830/_0_  ;
  output \g48831/_0_  ;
  output \g48833/_0_  ;
  output \g48834/_0_  ;
  output \g48835/_0_  ;
  output \g48836/_0_  ;
  output \g48837/_0_  ;
  output \g48838/_0_  ;
  output \g48839/_0_  ;
  output \g48840/_0_  ;
  output \g48841/_0_  ;
  output \g48842/_0_  ;
  output \g48843/_0_  ;
  output \g48844/_0_  ;
  output \g48845/_0_  ;
  output \g48846/_0_  ;
  output \g48847/_0_  ;
  output \g48848/_0_  ;
  output \g48908/_0_  ;
  output \g48909/_0_  ;
  output \g48910/_0_  ;
  output \g48912/_0_  ;
  output \g48913/_0_  ;
  output \g48915/_0_  ;
  output \g48917/_0_  ;
  output \g48932/_0_  ;
  output \g48933/_0_  ;
  output \g48935/_0_  ;
  output \g48937/_0_  ;
  output \g48938/_0_  ;
  output \g48939/_0_  ;
  output \g48940/_0_  ;
  output \g48942/_0_  ;
  output \g48945/_0_  ;
  output \g48971/_0_  ;
  output \g49007/_0_  ;
  output \g49047/_0_  ;
  output \g49048/_0_  ;
  output \g49050/_0_  ;
  output \g49182/_0_  ;
  output \g49280/_0_  ;
  output \g49332/_0_  ;
  output \g49335/_0_  ;
  output \g49336/_0_  ;
  output \g49337/_0_  ;
  output \g49338/_0_  ;
  output \g49339/_0_  ;
  output \g49340/_0_  ;
  output \g49341/_0_  ;
  output \g49342/_0_  ;
  output \g49343/_0_  ;
  output \g49344/_0_  ;
  output \g49345/_0_  ;
  output \g49346/_0_  ;
  output \g49347/_0_  ;
  output \g49348/_0_  ;
  output \g49349/_0_  ;
  output \g49356/_0_  ;
  output \g49375/_0_  ;
  output \g49396/_0_  ;
  output \g49397/_0_  ;
  output \g49400/_0_  ;
  output \g49404/_0_  ;
  output \g49406/_0_  ;
  output \g49414/_0_  ;
  output \g49422/_0_  ;
  output \g49426/_0_  ;
  output \g49430/_0_  ;
  output \g49434/_0_  ;
  output \g49437/_0_  ;
  output \g49440/_0_  ;
  output \g49441/_0_  ;
  output \g49444/_0_  ;
  output \g49448/_0_  ;
  output \g49451/_0_  ;
  output \g49455/_0_  ;
  output \g49456/_0_  ;
  output \g49460/_0_  ;
  output \g49466/_0_  ;
  output \g49563/_0_  ;
  output \g49592/_0_  ;
  output \g49915/_0_  ;
  output \g49941/_0_  ;
  output \g50023/_0_  ;
  output \g50026/_0_  ;
  output \g50029/_0_  ;
  output \g50031/_0_  ;
  output \g50033/_0_  ;
  output \g50035/_0_  ;
  output \g50037/_0_  ;
  output \g50040/_0_  ;
  output \g50050/_0_  ;
  output \g50056/_0_  ;
  output \g50059/_0_  ;
  output \g50065/_0_  ;
  output \g50067/_0_  ;
  output \g50150/_0_  ;
  output \g50283/_0_  ;
  output \g50284/_0_  ;
  output \g50501/_0_  ;
  output \g50594/_0_  ;
  output \g50807/_0_  ;
  output \g50866/_0_  ;
  output \g50875/_0_  ;
  output \g51449/_0_  ;
  output \g51510/_0_  ;
  output \g51534/_0_  ;
  output \g52310/_0_  ;
  output \g53066/_0_  ;
  output \g53087/_0_  ;
  output \g53151/_0_  ;
  output \g53608/_0_  ;
  output \g53634/_0_  ;
  output \g54053/_0_  ;
  output \g54091/_0_  ;
  output \g54103/_0_  ;
  output \g54268/_0_  ;
  output \g54277/_0_  ;
  output \g54287/_0_  ;
  output \g54294/_0_  ;
  output \g54449/_0_  ;
  output \g54453/_0_  ;
  output \g54484/_0_  ;
  output \g54528/_0_  ;
  output \g54582/_0_  ;
  output \g55448/_0_  ;
  output \g55693/_1_  ;
  output \g55874/_0_  ;
  output \g56203/_0_  ;
  output \g56303/_0_  ;
  output \g56329/_0_  ;
  output \g56336/_0_  ;
  output \g56345/_0_  ;
  output \g56367/_0_  ;
  output \g56411/_0_  ;
  output \g56529/_0_  ;
  output \g56858/_0_  ;
  output \g60443/_1_  ;
  output \g63395/_0_  ;
  output \g63442/_0_  ;
  output \g63595/_0_  ;
  output \g63996/_0_  ;
  output \g64048/_0_  ;
  output \g64071/_0_  ;
  output \g64085/_0_  ;
  output \g64096/_0_  ;
  output \g64119/_0_  ;
  output \g64216/_0_  ;
  output \g64513/_0_  ;
  output \g64566/_0_  ;
  output \g64694/_0_  ;
  output \g64913/_0_  ;
  wire n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 ;
  assign n452 = \InstQueueRd_Addr_reg[2]/NET0131  & ~\InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n457 = ~\InstQueueRd_Addr_reg[0]/NET0131  & \InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n482 = n452 & n457 ;
  assign n546 = \InstQueue_reg[6][2]/NET0131  & n482 ;
  assign n453 = \InstQueueRd_Addr_reg[0]/NET0131  & \InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n464 = \InstQueueRd_Addr_reg[2]/NET0131  & \InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n522 = n453 & n464 ;
  assign n547 = \InstQueue_reg[15][2]/NET0131  & n522 ;
  assign n560 = ~n546 & ~n547 ;
  assign n463 = \InstQueueRd_Addr_reg[0]/NET0131  & ~\InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n490 = n452 & n463 ;
  assign n548 = \InstQueue_reg[5][2]/NET0131  & n490 ;
  assign n460 = ~\InstQueueRd_Addr_reg[2]/NET0131  & \InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n492 = n453 & n460 ;
  assign n549 = \InstQueue_reg[11][2]/NET0131  & n492 ;
  assign n561 = ~n548 & ~n549 ;
  assign n568 = n560 & n561 ;
  assign n456 = ~\InstQueueRd_Addr_reg[2]/NET0131  & ~\InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n476 = n453 & n456 ;
  assign n542 = \InstQueue_reg[3][2]/NET0131  & n476 ;
  assign n465 = n463 & n464 ;
  assign n543 = \InstQueue_reg[13][2]/NET0131  & n465 ;
  assign n558 = ~n542 & ~n543 ;
  assign n467 = ~\InstQueueRd_Addr_reg[0]/NET0131  & ~\InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n486 = n460 & n467 ;
  assign n544 = \InstQueue_reg[8][2]/NET0131  & n486 ;
  assign n474 = n456 & n467 ;
  assign n545 = \InstQueue_reg[0][2]/NET0131  & n474 ;
  assign n559 = ~n544 & ~n545 ;
  assign n569 = n558 & n559 ;
  assign n570 = n568 & n569 ;
  assign n484 = n460 & n463 ;
  assign n554 = \InstQueue_reg[9][2]/NET0131  & n484 ;
  assign n472 = n452 & n467 ;
  assign n555 = \InstQueue_reg[4][2]/NET0131  & n472 ;
  assign n564 = ~n554 & ~n555 ;
  assign n454 = n452 & n453 ;
  assign n556 = \InstQueue_reg[7][2]/NET0131  & n454 ;
  assign n461 = n457 & n460 ;
  assign n557 = \InstQueue_reg[10][2]/NET0131  & n461 ;
  assign n565 = ~n556 & ~n557 ;
  assign n566 = n564 & n565 ;
  assign n488 = n456 & n463 ;
  assign n550 = \InstQueue_reg[1][2]/NET0131  & n488 ;
  assign n458 = n456 & n457 ;
  assign n551 = \InstQueue_reg[2][2]/NET0131  & n458 ;
  assign n562 = ~n550 & ~n551 ;
  assign n470 = n457 & n464 ;
  assign n552 = \InstQueue_reg[14][2]/NET0131  & n470 ;
  assign n468 = n464 & n467 ;
  assign n553 = \InstQueue_reg[12][2]/NET0131  & n468 ;
  assign n563 = ~n552 & ~n553 ;
  assign n567 = n562 & n563 ;
  assign n571 = n566 & n567 ;
  assign n572 = n570 & n571 ;
  assign n478 = \InstQueueRd_Addr_reg[1]/NET0131  & \InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n479 = \InstQueueRd_Addr_reg[3]/NET0131  & n478 ;
  assign n577 = \InstQueueRd_Addr_reg[0]/NET0131  & \InstQueue_reg[15][1]/NET0131  ;
  assign n578 = n479 & n577 ;
  assign n579 = \InstQueue_reg[7][1]/NET0131  & n454 ;
  assign n592 = ~n578 & ~n579 ;
  assign n580 = \InstQueue_reg[9][1]/NET0131  & n484 ;
  assign n581 = \InstQueue_reg[3][1]/NET0131  & n476 ;
  assign n593 = ~n580 & ~n581 ;
  assign n600 = n592 & n593 ;
  assign n573 = \InstQueue_reg[6][1]/NET0131  & n482 ;
  assign n574 = \InstQueue_reg[4][1]/NET0131  & n472 ;
  assign n590 = ~n573 & ~n574 ;
  assign n575 = \InstQueue_reg[0][1]/NET0131  & n474 ;
  assign n576 = \InstQueue_reg[8][1]/NET0131  & n486 ;
  assign n591 = ~n575 & ~n576 ;
  assign n601 = n590 & n591 ;
  assign n602 = n600 & n601 ;
  assign n586 = \InstQueue_reg[2][1]/NET0131  & n458 ;
  assign n587 = \InstQueue_reg[12][1]/NET0131  & n468 ;
  assign n596 = ~n586 & ~n587 ;
  assign n588 = \InstQueue_reg[14][1]/NET0131  & n470 ;
  assign n589 = \InstQueue_reg[11][1]/NET0131  & n492 ;
  assign n597 = ~n588 & ~n589 ;
  assign n598 = n596 & n597 ;
  assign n582 = \InstQueue_reg[13][1]/NET0131  & n465 ;
  assign n583 = \InstQueue_reg[10][1]/NET0131  & n461 ;
  assign n594 = ~n582 & ~n583 ;
  assign n584 = \InstQueue_reg[1][1]/NET0131  & n488 ;
  assign n585 = \InstQueue_reg[5][1]/NET0131  & n490 ;
  assign n595 = ~n584 & ~n585 ;
  assign n599 = n594 & n595 ;
  assign n603 = n598 & n599 ;
  assign n604 = n602 & n603 ;
  assign n737 = n572 & n604 ;
  assign n469 = \InstQueue_reg[12][0]/NET0131  & n468 ;
  assign n471 = \InstQueue_reg[14][0]/NET0131  & n470 ;
  assign n496 = ~n469 & ~n471 ;
  assign n473 = \InstQueue_reg[4][0]/NET0131  & n472 ;
  assign n475 = \InstQueue_reg[0][0]/NET0131  & n474 ;
  assign n497 = ~n473 & ~n475 ;
  assign n504 = n496 & n497 ;
  assign n455 = \InstQueue_reg[7][0]/NET0131  & n454 ;
  assign n459 = \InstQueue_reg[2][0]/NET0131  & n458 ;
  assign n494 = ~n455 & ~n459 ;
  assign n462 = \InstQueue_reg[10][0]/NET0131  & n461 ;
  assign n466 = \InstQueue_reg[13][0]/NET0131  & n465 ;
  assign n495 = ~n462 & ~n466 ;
  assign n505 = n494 & n495 ;
  assign n506 = n504 & n505 ;
  assign n487 = \InstQueue_reg[8][0]/NET0131  & n486 ;
  assign n489 = \InstQueue_reg[1][0]/NET0131  & n488 ;
  assign n500 = ~n487 & ~n489 ;
  assign n491 = \InstQueue_reg[5][0]/NET0131  & n490 ;
  assign n493 = \InstQueue_reg[11][0]/NET0131  & n492 ;
  assign n501 = ~n491 & ~n493 ;
  assign n502 = n500 & n501 ;
  assign n477 = \InstQueue_reg[3][0]/NET0131  & n476 ;
  assign n480 = \InstQueueRd_Addr_reg[0]/NET0131  & \InstQueue_reg[15][0]/NET0131  ;
  assign n481 = n479 & n480 ;
  assign n498 = ~n477 & ~n481 ;
  assign n483 = \InstQueue_reg[6][0]/NET0131  & n482 ;
  assign n485 = \InstQueue_reg[9][0]/NET0131  & n484 ;
  assign n499 = ~n483 & ~n485 ;
  assign n503 = n498 & n499 ;
  assign n507 = n502 & n503 ;
  assign n508 = n506 & n507 ;
  assign n513 = \InstQueue_reg[4][3]/NET0131  & n472 ;
  assign n514 = \InstQueue_reg[1][3]/NET0131  & n488 ;
  assign n528 = ~n513 & ~n514 ;
  assign n515 = \InstQueue_reg[13][3]/NET0131  & n465 ;
  assign n516 = \InstQueue_reg[10][3]/NET0131  & n461 ;
  assign n529 = ~n515 & ~n516 ;
  assign n536 = n528 & n529 ;
  assign n509 = \InstQueue_reg[3][3]/NET0131  & n476 ;
  assign n510 = \InstQueue_reg[8][3]/NET0131  & n486 ;
  assign n526 = ~n509 & ~n510 ;
  assign n511 = \InstQueue_reg[5][3]/NET0131  & n490 ;
  assign n512 = \InstQueue_reg[12][3]/NET0131  & n468 ;
  assign n527 = ~n511 & ~n512 ;
  assign n537 = n526 & n527 ;
  assign n538 = n536 & n537 ;
  assign n521 = \InstQueue_reg[2][3]/NET0131  & n458 ;
  assign n523 = \InstQueue_reg[15][3]/NET0131  & n522 ;
  assign n532 = ~n521 & ~n523 ;
  assign n524 = \InstQueue_reg[6][3]/NET0131  & n482 ;
  assign n525 = \InstQueue_reg[0][3]/NET0131  & n474 ;
  assign n533 = ~n524 & ~n525 ;
  assign n534 = n532 & n533 ;
  assign n517 = \InstQueue_reg[14][3]/NET0131  & n470 ;
  assign n518 = \InstQueue_reg[9][3]/NET0131  & n484 ;
  assign n530 = ~n517 & ~n518 ;
  assign n519 = \InstQueue_reg[7][3]/NET0131  & n454 ;
  assign n520 = \InstQueue_reg[11][3]/NET0131  & n492 ;
  assign n531 = ~n519 & ~n520 ;
  assign n535 = n530 & n531 ;
  assign n539 = n534 & n535 ;
  assign n540 = n538 & n539 ;
  assign n776 = n508 & n540 ;
  assign n786 = n737 & n776 ;
  assign n705 = \InstQueue_reg[13][6]/NET0131  & n465 ;
  assign n706 = \InstQueue_reg[1][6]/NET0131  & n488 ;
  assign n719 = ~n705 & ~n706 ;
  assign n707 = \InstQueue_reg[0][6]/NET0131  & n474 ;
  assign n708 = \InstQueue_reg[9][6]/NET0131  & n484 ;
  assign n720 = ~n707 & ~n708 ;
  assign n727 = n719 & n720 ;
  assign n701 = \InstQueue_reg[3][6]/NET0131  & n476 ;
  assign n702 = \InstQueue_reg[8][6]/NET0131  & n486 ;
  assign n717 = ~n701 & ~n702 ;
  assign n703 = \InstQueue_reg[15][6]/NET0131  & n522 ;
  assign n704 = \InstQueue_reg[5][6]/NET0131  & n490 ;
  assign n718 = ~n703 & ~n704 ;
  assign n728 = n717 & n718 ;
  assign n729 = n727 & n728 ;
  assign n713 = \InstQueue_reg[2][6]/NET0131  & n458 ;
  assign n714 = \InstQueue_reg[7][6]/NET0131  & n454 ;
  assign n723 = ~n713 & ~n714 ;
  assign n715 = \InstQueue_reg[12][6]/NET0131  & n468 ;
  assign n716 = \InstQueue_reg[10][6]/NET0131  & n461 ;
  assign n724 = ~n715 & ~n716 ;
  assign n725 = n723 & n724 ;
  assign n709 = \InstQueue_reg[14][6]/NET0131  & n470 ;
  assign n710 = \InstQueue_reg[6][6]/NET0131  & n482 ;
  assign n721 = ~n709 & ~n710 ;
  assign n711 = \InstQueue_reg[4][6]/NET0131  & n472 ;
  assign n712 = \InstQueue_reg[11][6]/NET0131  & n492 ;
  assign n722 = ~n711 & ~n712 ;
  assign n726 = n721 & n722 ;
  assign n730 = n725 & n726 ;
  assign n731 = n729 & n730 ;
  assign n611 = \InstQueue_reg[0][5]/NET0131  & n474 ;
  assign n612 = \InstQueue_reg[1][5]/NET0131  & n488 ;
  assign n625 = ~n611 & ~n612 ;
  assign n613 = \InstQueue_reg[4][5]/NET0131  & n472 ;
  assign n614 = \InstQueue_reg[6][5]/NET0131  & n482 ;
  assign n626 = ~n613 & ~n614 ;
  assign n633 = n625 & n626 ;
  assign n607 = \InstQueue_reg[3][5]/NET0131  & n476 ;
  assign n608 = \InstQueue_reg[11][5]/NET0131  & n492 ;
  assign n623 = ~n607 & ~n608 ;
  assign n609 = \InstQueue_reg[15][5]/NET0131  & n522 ;
  assign n610 = \InstQueue_reg[5][5]/NET0131  & n490 ;
  assign n624 = ~n609 & ~n610 ;
  assign n634 = n623 & n624 ;
  assign n635 = n633 & n634 ;
  assign n619 = \InstQueue_reg[2][5]/NET0131  & n458 ;
  assign n620 = \InstQueue_reg[13][5]/NET0131  & n465 ;
  assign n629 = ~n619 & ~n620 ;
  assign n621 = \InstQueue_reg[12][5]/NET0131  & n468 ;
  assign n622 = \InstQueue_reg[10][5]/NET0131  & n461 ;
  assign n630 = ~n621 & ~n622 ;
  assign n631 = n629 & n630 ;
  assign n615 = \InstQueue_reg[14][5]/NET0131  & n470 ;
  assign n616 = \InstQueue_reg[9][5]/NET0131  & n484 ;
  assign n627 = ~n615 & ~n616 ;
  assign n617 = \InstQueue_reg[8][5]/NET0131  & n486 ;
  assign n618 = \InstQueue_reg[7][5]/NET0131  & n454 ;
  assign n628 = ~n617 & ~n618 ;
  assign n632 = n627 & n628 ;
  assign n636 = n631 & n632 ;
  assign n637 = n635 & n636 ;
  assign n673 = \InstQueueRd_Addr_reg[0]/NET0131  & \InstQueue_reg[15][7]/NET0131  ;
  assign n674 = n479 & n673 ;
  assign n675 = \InstQueue_reg[4][7]/NET0131  & n472 ;
  assign n688 = ~n674 & ~n675 ;
  assign n676 = \InstQueue_reg[0][7]/NET0131  & n474 ;
  assign n677 = \InstQueue_reg[14][7]/NET0131  & n470 ;
  assign n689 = ~n676 & ~n677 ;
  assign n696 = n688 & n689 ;
  assign n669 = \InstQueue_reg[12][7]/NET0131  & n468 ;
  assign n670 = \InstQueue_reg[13][7]/NET0131  & n465 ;
  assign n686 = ~n669 & ~n670 ;
  assign n671 = \InstQueue_reg[5][7]/NET0131  & n490 ;
  assign n672 = \InstQueue_reg[11][7]/NET0131  & n492 ;
  assign n687 = ~n671 & ~n672 ;
  assign n697 = n686 & n687 ;
  assign n698 = n696 & n697 ;
  assign n682 = \InstQueue_reg[6][7]/NET0131  & n482 ;
  assign n683 = \InstQueue_reg[1][7]/NET0131  & n488 ;
  assign n692 = ~n682 & ~n683 ;
  assign n684 = \InstQueue_reg[9][7]/NET0131  & n484 ;
  assign n685 = \InstQueue_reg[8][7]/NET0131  & n486 ;
  assign n693 = ~n684 & ~n685 ;
  assign n694 = n692 & n693 ;
  assign n678 = \InstQueue_reg[3][7]/NET0131  & n476 ;
  assign n679 = \InstQueue_reg[7][7]/NET0131  & n454 ;
  assign n690 = ~n678 & ~n679 ;
  assign n680 = \InstQueue_reg[10][7]/NET0131  & n461 ;
  assign n681 = \InstQueue_reg[2][7]/NET0131  & n458 ;
  assign n691 = ~n680 & ~n681 ;
  assign n695 = n690 & n691 ;
  assign n699 = n694 & n695 ;
  assign n700 = n698 & n699 ;
  assign n780 = n637 & ~n700 ;
  assign n787 = ~n731 & n780 ;
  assign n788 = n786 & n787 ;
  assign n741 = ~\InstQueueRd_Addr_reg[3]/NET0131  & \InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n742 = ~\InstQueueRd_Addr_reg[2]/NET0131  & \InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n743 = \InstQueueRd_Addr_reg[2]/NET0131  & ~\InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n744 = ~\InstQueueRd_Addr_reg[1]/NET0131  & \InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n745 = \InstQueueRd_Addr_reg[1]/NET0131  & ~\InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n746 = \InstQueueRd_Addr_reg[0]/NET0131  & ~\InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n747 = ~n745 & ~n746 ;
  assign n748 = ~n744 & ~n747 ;
  assign n749 = ~n743 & ~n748 ;
  assign n750 = ~n742 & ~n749 ;
  assign n751 = n741 & ~n750 ;
  assign n752 = \InstQueueRd_Addr_reg[3]/NET0131  & ~\InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n753 = ~n750 & ~n752 ;
  assign n754 = ~n741 & ~n753 ;
  assign n755 = ~n742 & ~n743 ;
  assign n756 = n748 & ~n755 ;
  assign n757 = ~n748 & n755 ;
  assign n758 = ~n756 & ~n757 ;
  assign n759 = ~n754 & n758 ;
  assign n760 = ~n751 & ~n759 ;
  assign n762 = ~n744 & n747 ;
  assign n830 = ~n744 & ~n745 ;
  assign n831 = n746 & ~n830 ;
  assign n832 = ~n762 & ~n831 ;
  assign n833 = ~n754 & n832 ;
  assign n834 = n760 & ~n833 ;
  assign n541 = ~n508 & ~n540 ;
  assign n605 = n572 & ~n604 ;
  assign n606 = n541 & n605 ;
  assign n642 = \InstQueue_reg[0][4]/NET0131  & n474 ;
  assign n643 = \InstQueue_reg[2][4]/NET0131  & n458 ;
  assign n656 = ~n642 & ~n643 ;
  assign n644 = \InstQueue_reg[12][4]/NET0131  & n468 ;
  assign n645 = \InstQueue_reg[4][4]/NET0131  & n472 ;
  assign n657 = ~n644 & ~n645 ;
  assign n664 = n656 & n657 ;
  assign n638 = \InstQueue_reg[14][4]/NET0131  & n470 ;
  assign n639 = \InstQueue_reg[10][4]/NET0131  & n461 ;
  assign n654 = ~n638 & ~n639 ;
  assign n640 = \InstQueue_reg[11][4]/NET0131  & n492 ;
  assign n641 = \InstQueue_reg[5][4]/NET0131  & n490 ;
  assign n655 = ~n640 & ~n641 ;
  assign n665 = n654 & n655 ;
  assign n666 = n664 & n665 ;
  assign n650 = \InstQueue_reg[1][4]/NET0131  & n488 ;
  assign n651 = \InstQueue_reg[7][4]/NET0131  & n454 ;
  assign n660 = ~n650 & ~n651 ;
  assign n652 = \InstQueue_reg[9][4]/NET0131  & n484 ;
  assign n653 = \InstQueue_reg[15][4]/NET0131  & n522 ;
  assign n661 = ~n652 & ~n653 ;
  assign n662 = n660 & n661 ;
  assign n646 = \InstQueue_reg[3][4]/NET0131  & n476 ;
  assign n647 = \InstQueue_reg[6][4]/NET0131  & n482 ;
  assign n658 = ~n646 & ~n647 ;
  assign n648 = \InstQueue_reg[13][4]/NET0131  & n465 ;
  assign n649 = \InstQueue_reg[8][4]/NET0131  & n486 ;
  assign n659 = ~n648 & ~n649 ;
  assign n663 = n658 & n659 ;
  assign n667 = n662 & n663 ;
  assign n668 = n666 & n667 ;
  assign n779 = n668 & n731 ;
  assign n781 = n779 & n780 ;
  assign n782 = n606 & n781 ;
  assign n767 = n668 & ~n731 ;
  assign n768 = ~n637 & ~n700 ;
  assign n769 = n767 & n768 ;
  assign n777 = ~n572 & n776 ;
  assign n778 = n769 & n777 ;
  assign n840 = n604 & n778 ;
  assign n841 = ~n782 & ~n840 ;
  assign n842 = ~n834 & ~n841 ;
  assign n770 = n541 & n737 ;
  assign n783 = n770 & n781 ;
  assign n804 = ~n604 & n777 ;
  assign n835 = n769 & n804 ;
  assign n836 = ~n783 & ~n835 ;
  assign n824 = ~\State_reg[0]/NET0131  & \State_reg[1]/NET0131  ;
  assign n825 = ~\State_reg[2]/NET0131  & n824 ;
  assign n826 = ~\State_reg[0]/NET0131  & ~\State_reg[1]/NET0131  ;
  assign n827 = \State_reg[2]/NET0131  & n826 ;
  assign n828 = ~n825 & ~n827 ;
  assign n856 = ~n828 & ~n834 ;
  assign n857 = ~n836 & n856 ;
  assign n858 = ~n842 & ~n857 ;
  assign n872 = ~READY_n_pad & ~n858 ;
  assign n873 = ~n788 & ~n872 ;
  assign n874 = ~n478 & ~n858 ;
  assign n875 = n873 & ~n874 ;
  assign n876 = ~\InstQueueRd_Addr_reg[3]/NET0131  & ~n478 ;
  assign n877 = ~n479 & ~n876 ;
  assign n878 = ~n875 & n877 ;
  assign n732 = ~n668 & ~n700 ;
  assign n733 = n731 & n732 ;
  assign n734 = ~n637 & n733 ;
  assign n735 = n606 & n734 ;
  assign n736 = n508 & ~n540 ;
  assign n738 = n736 & n737 ;
  assign n739 = n734 & n738 ;
  assign n740 = ~n735 & ~n739 ;
  assign n771 = n769 & n770 ;
  assign n772 = n605 & n769 ;
  assign n773 = n541 & n772 ;
  assign n774 = ~n771 & ~n773 ;
  assign n775 = n740 & n774 ;
  assign n859 = READY_n_pad & ~n858 ;
  assign n860 = n834 & ~n841 ;
  assign n861 = n836 & ~n860 ;
  assign n862 = ~n856 & ~n861 ;
  assign n863 = ~n859 & ~n862 ;
  assign n864 = n775 & n863 ;
  assign n865 = \InstQueueRd_Addr_reg[3]/NET0131  & ~n864 ;
  assign n784 = ~n778 & ~n782 ;
  assign n785 = ~n783 & n784 ;
  assign n789 = n785 & ~n788 ;
  assign n790 = n775 & n789 ;
  assign n791 = n700 & n767 ;
  assign n792 = n637 & n791 ;
  assign n793 = ~n733 & ~n792 ;
  assign n794 = n786 & ~n793 ;
  assign n795 = ~n508 & n540 ;
  assign n796 = n605 & n795 ;
  assign n797 = n792 & n796 ;
  assign n799 = n604 & n637 ;
  assign n800 = n700 & n799 ;
  assign n798 = n540 & ~n572 ;
  assign n801 = n779 & n798 ;
  assign n802 = n800 & n801 ;
  assign n807 = ~n797 & ~n802 ;
  assign n803 = n736 & n772 ;
  assign n805 = ~n637 & n791 ;
  assign n806 = n804 & n805 ;
  assign n808 = ~n803 & ~n806 ;
  assign n809 = n807 & n808 ;
  assign n810 = ~n794 & n809 ;
  assign n811 = ~n790 & n810 ;
  assign n866 = \InstQueueRd_Addr_reg[2]/NET0131  & n453 ;
  assign n867 = \InstQueueRd_Addr_reg[3]/NET0131  & ~n866 ;
  assign n868 = ~n454 & ~n867 ;
  assign n869 = ~n811 & ~n868 ;
  assign n761 = ~\InstQueueRd_Addr_reg[0]/NET0131  & \InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n763 = ~n761 & n762 ;
  assign n764 = ~n751 & n763 ;
  assign n765 = ~n760 & ~n764 ;
  assign n766 = ~n740 & n765 ;
  assign n870 = ~\InstQueueRd_Addr_reg[2]/NET0131  & ~n453 ;
  assign n871 = n766 & ~n870 ;
  assign n879 = ~n869 & ~n871 ;
  assign n880 = ~n865 & n879 ;
  assign n881 = ~n878 & n880 ;
  assign n882 = \InstQueueWr_Addr_reg[3]/NET0131  & n881 ;
  assign n812 = ~n766 & n811 ;
  assign n813 = ~\InstQueueRd_Addr_reg[0]/NET0131  & n812 ;
  assign n814 = ~n740 & ~n765 ;
  assign n815 = n774 & ~n814 ;
  assign n816 = \InstQueueRd_Addr_reg[0]/NET0131  & n789 ;
  assign n817 = n815 & n816 ;
  assign n818 = ~n813 & ~n817 ;
  assign n819 = \InstQueueWr_Addr_reg[0]/NET0131  & ~n818 ;
  assign n821 = ~\InstQueueWr_Addr_reg[1]/NET0131  & ~n819 ;
  assign n829 = ~READY_n_pad & ~n828 ;
  assign n837 = ~n834 & ~n836 ;
  assign n838 = n829 & n837 ;
  assign n839 = ~n788 & ~n838 ;
  assign n843 = ~READY_n_pad & n842 ;
  assign n844 = n839 & ~n843 ;
  assign n845 = ~\InstQueueRd_Addr_reg[1]/NET0131  & ~n844 ;
  assign n822 = ~n457 & ~n463 ;
  assign n823 = ~n812 & ~n822 ;
  assign n846 = ~READY_n_pad & ~n834 ;
  assign n847 = ~n841 & ~n846 ;
  assign n848 = n829 & ~n834 ;
  assign n849 = ~n836 & ~n848 ;
  assign n850 = ~n847 & ~n849 ;
  assign n851 = n815 & n850 ;
  assign n852 = \InstQueueRd_Addr_reg[1]/NET0131  & ~n851 ;
  assign n853 = ~n823 & ~n852 ;
  assign n854 = ~n845 & n853 ;
  assign n855 = ~n821 & n854 ;
  assign n820 = \InstQueueWr_Addr_reg[1]/NET0131  & n819 ;
  assign n885 = ~\InstQueueRd_Addr_reg[1]/NET0131  & ~\InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n886 = ~n478 & ~n885 ;
  assign n887 = ~n873 & n886 ;
  assign n883 = ~n866 & ~n870 ;
  assign n889 = ~n811 & n883 ;
  assign n884 = n766 & ~n883 ;
  assign n888 = \InstQueueRd_Addr_reg[2]/NET0131  & ~n851 ;
  assign n890 = ~n884 & ~n888 ;
  assign n891 = ~n889 & n890 ;
  assign n892 = ~n887 & n891 ;
  assign n893 = \InstQueueWr_Addr_reg[2]/NET0131  & n892 ;
  assign n894 = ~n820 & ~n893 ;
  assign n895 = ~n855 & n894 ;
  assign n896 = ~n882 & n895 ;
  assign n917 = ~\InstQueueWr_Addr_reg[2]/NET0131  & ~n892 ;
  assign n918 = ~n882 & n917 ;
  assign n897 = \InstQueueWr_Addr_reg[3]/NET0131  & n892 ;
  assign n898 = ~n881 & ~n897 ;
  assign n900 = READY_n_pad & n842 ;
  assign n901 = ~n829 & n837 ;
  assign n902 = ~n900 & ~n901 ;
  assign n903 = \Flush_reg/NET0131  & ~n902 ;
  assign n899 = n765 & n771 ;
  assign n904 = ~n761 & ~n830 ;
  assign n905 = n833 & ~n904 ;
  assign n906 = n760 & ~n905 ;
  assign n907 = n773 & ~n906 ;
  assign n908 = ~n899 & ~n907 ;
  assign n909 = ~n903 & n908 ;
  assign n913 = ~\More_reg/NET0131  & ~n834 ;
  assign n914 = ~n850 & ~n913 ;
  assign n910 = n773 & n906 ;
  assign n911 = ~n765 & n771 ;
  assign n912 = ~n814 & ~n911 ;
  assign n915 = ~n910 & n912 ;
  assign n916 = ~n914 & n915 ;
  assign n919 = n909 & n916 ;
  assign n920 = ~n898 & n919 ;
  assign n921 = ~n918 & n920 ;
  assign n922 = ~n896 & n921 ;
  assign n923 = n783 & ~n834 ;
  assign n924 = ~\DataWidth_reg[1]/NET0131  & n829 ;
  assign n925 = n923 & n924 ;
  assign n926 = n922 & ~n925 ;
  assign n927 = \State2_reg[0]/NET0131  & ~\State2_reg[3]/NET0131  ;
  assign n928 = \State2_reg[2]/NET0131  & n927 ;
  assign n929 = ~\State2_reg[1]/NET0131  & n928 ;
  assign n930 = ~n926 & n929 ;
  assign n939 = ~\State2_reg[2]/NET0131  & n927 ;
  assign n931 = ~\State2_reg[0]/NET0131  & ~\State2_reg[3]/NET0131  ;
  assign n940 = \State2_reg[2]/NET0131  & n931 ;
  assign n941 = ~n939 & ~n940 ;
  assign n942 = READY_n_pad & \State2_reg[1]/NET0131  ;
  assign n943 = ~n941 & n942 ;
  assign n932 = \State2_reg[1]/NET0131  & ~\State2_reg[2]/NET0131  ;
  assign n933 = n931 & n932 ;
  assign n934 = ~\DataWidth_reg[1]/NET0131  & n933 ;
  assign n935 = ~\State2_reg[1]/NET0131  & ~\State2_reg[2]/NET0131  ;
  assign n936 = \State2_reg[0]/NET0131  & n935 ;
  assign n937 = ~\State2_reg[3]/NET0131  & n936 ;
  assign n938 = ~READY_n_pad & n937 ;
  assign n944 = ~n934 & ~n938 ;
  assign n945 = ~n943 & n944 ;
  assign n946 = ~n930 & n945 ;
  assign n947 = n922 & n925 ;
  assign n948 = n929 & ~n947 ;
  assign n949 = \State2_reg[1]/NET0131  & \State2_reg[2]/NET0131  ;
  assign n955 = ~\State2_reg[3]/NET0131  & n949 ;
  assign n956 = \State2_reg[0]/NET0131  & n955 ;
  assign n957 = ~\Flush_reg/NET0131  & \InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n958 = \InstQueueRd_Addr_reg[3]/NET0131  & ~n467 ;
  assign n959 = n957 & n958 ;
  assign n960 = n956 & ~n959 ;
  assign n954 = READY_n_pad & n939 ;
  assign n950 = READY_n_pad & n949 ;
  assign n951 = n931 & ~n950 ;
  assign n952 = \State2_reg[3]/NET0131  & n935 ;
  assign n953 = \State2_reg[0]/NET0131  & n952 ;
  assign n961 = ~n951 & ~n953 ;
  assign n962 = ~n954 & n961 ;
  assign n963 = ~n960 & n962 ;
  assign n964 = ~n948 & n963 ;
  assign n965 = ~\State2_reg[0]/NET0131  & n952 ;
  assign n966 = ~n956 & ~n965 ;
  assign n967 = \State2_reg[1]/NET0131  & n939 ;
  assign n968 = ~READY_n_pad & n967 ;
  assign n969 = \DataWidth_reg[1]/NET0131  & n933 ;
  assign n970 = ~n929 & ~n940 ;
  assign n971 = ~n969 & n970 ;
  assign n972 = ~n968 & n971 ;
  assign n973 = \InstAddrPointer_reg[30]/NET0131  & n906 ;
  assign n1325 = \InstAddrPointer_reg[17]/NET0131  & \InstAddrPointer_reg[18]/NET0131  ;
  assign n1326 = \InstAddrPointer_reg[19]/NET0131  & n1325 ;
  assign n981 = \InstAddrPointer_reg[6]/NET0131  & \InstAddrPointer_reg[7]/NET0131  ;
  assign n974 = \InstAddrPointer_reg[1]/NET0131  & \InstAddrPointer_reg[2]/NET0131  ;
  assign n975 = \InstAddrPointer_reg[3]/NET0131  & n974 ;
  assign n976 = \InstAddrPointer_reg[4]/NET0131  & n975 ;
  assign n1291 = \InstAddrPointer_reg[5]/NET0131  & n976 ;
  assign n1292 = n981 & n1291 ;
  assign n1293 = \InstAddrPointer_reg[8]/NET0131  & \InstAddrPointer_reg[9]/NET0131  ;
  assign n1294 = \InstAddrPointer_reg[10]/NET0131  & n1293 ;
  assign n1295 = n1292 & n1294 ;
  assign n1296 = \InstAddrPointer_reg[11]/NET0131  & \InstAddrPointer_reg[12]/NET0131  ;
  assign n1297 = \InstAddrPointer_reg[13]/NET0131  & n1296 ;
  assign n1298 = n1295 & n1297 ;
  assign n1327 = \InstAddrPointer_reg[14]/NET0131  & \InstAddrPointer_reg[15]/NET0131  ;
  assign n1328 = \InstAddrPointer_reg[16]/NET0131  & n1327 ;
  assign n1329 = n1298 & n1328 ;
  assign n1330 = n1326 & n1329 ;
  assign n1362 = \InstAddrPointer_reg[21]/NET0131  & \InstAddrPointer_reg[22]/NET0131  ;
  assign n1365 = \InstAddrPointer_reg[23]/NET0131  & n1362 ;
  assign n1366 = \InstAddrPointer_reg[20]/NET0131  & n1365 ;
  assign n1488 = n1330 & n1366 ;
  assign n1489 = \InstAddrPointer_reg[24]/NET0131  & n1488 ;
  assign n1490 = \InstAddrPointer_reg[25]/NET0131  & n1489 ;
  assign n1386 = \InstAddrPointer_reg[26]/NET0131  & \InstAddrPointer_reg[27]/NET0131  ;
  assign n1505 = \InstAddrPointer_reg[28]/NET0131  & n1386 ;
  assign n1506 = n1490 & n1505 ;
  assign n1507 = \InstAddrPointer_reg[29]/NET0131  & n1506 ;
  assign n1513 = ~\InstAddrPointer_reg[30]/NET0131  & ~n1507 ;
  assign n1514 = \InstAddrPointer_reg[30]/NET0131  & n1507 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1094 = \InstQueue_reg[12][4]/NET0131  & n492 ;
  assign n1095 = \InstQueue_reg[3][4]/NET0131  & n458 ;
  assign n1113 = ~n1094 & ~n1095 ;
  assign n1096 = \InstQueue_reg[8][4]/NET0131  & n454 ;
  assign n1097 = \InstQueue_reg[9][4]/NET0131  & n486 ;
  assign n1114 = ~n1096 & ~n1097 ;
  assign n1118 = n1113 & n1114 ;
  assign n1090 = \InstQueue_reg[4][4]/NET0131  & n476 ;
  assign n1091 = \InstQueue_reg[2][4]/NET0131  & n488 ;
  assign n1111 = ~n1090 & ~n1091 ;
  assign n1092 = \InstQueue_reg[7][4]/NET0131  & n482 ;
  assign n1093 = \InstQueue_reg[10][4]/NET0131  & n484 ;
  assign n1112 = ~n1092 & ~n1093 ;
  assign n1119 = n1111 & n1112 ;
  assign n1120 = n1118 & n1119 ;
  assign n1016 = ~\InstQueueRd_Addr_reg[0]/NET0131  & n478 ;
  assign n1098 = \InstQueue_reg[15][4]/NET0131  & n1016 ;
  assign n1099 = ~n868 & n1098 ;
  assign n1100 = \InstQueue_reg[11][4]/NET0131  & n461 ;
  assign n1101 = \InstQueue_reg[5][4]/NET0131  & n472 ;
  assign n1115 = ~n1100 & ~n1101 ;
  assign n1102 = \InstQueue_reg[6][4]/NET0131  & n490 ;
  assign n1103 = \InstQueue_reg[14][4]/NET0131  & n465 ;
  assign n1116 = ~n1102 & ~n1103 ;
  assign n1117 = n1115 & n1116 ;
  assign n1121 = ~n1099 & n1117 ;
  assign n1104 = \InstQueue_reg[1][4]/NET0131  & n467 ;
  assign n1105 = \InstQueue_reg[0][4]/NET0131  & n453 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = ~n883 & ~n1106 ;
  assign n1108 = n868 & n1107 ;
  assign n1019 = \InstQueueRd_Addr_reg[3]/NET0131  & n883 ;
  assign n1109 = \InstQueue_reg[13][4]/NET0131  & n467 ;
  assign n1110 = n1019 & n1109 ;
  assign n1122 = ~n1108 & ~n1110 ;
  assign n1123 = n1121 & n1122 ;
  assign n1124 = n1120 & n1123 ;
  assign n1408 = ~\InstAddrPointer_reg[4]/NET0131  & ~n975 ;
  assign n1409 = ~n976 & ~n1408 ;
  assign n1410 = n1124 & ~n1409 ;
  assign n1170 = \InstQueue_reg[8][2]/NET0131  & n454 ;
  assign n1171 = \InstQueue_reg[13][2]/NET0131  & n468 ;
  assign n1185 = ~n1170 & ~n1171 ;
  assign n1172 = \InstQueue_reg[0][2]/NET0131  & n522 ;
  assign n1173 = \InstQueue_reg[14][2]/NET0131  & n465 ;
  assign n1186 = ~n1172 & ~n1173 ;
  assign n1192 = n1185 & n1186 ;
  assign n1166 = \InstQueue_reg[5][2]/NET0131  & n472 ;
  assign n1167 = \InstQueue_reg[6][2]/NET0131  & n490 ;
  assign n1183 = ~n1166 & ~n1167 ;
  assign n1168 = \InstQueue_reg[12][2]/NET0131  & n492 ;
  assign n1169 = \InstQueue_reg[9][2]/NET0131  & n486 ;
  assign n1184 = ~n1168 & ~n1169 ;
  assign n1193 = n1183 & n1184 ;
  assign n1194 = n1192 & n1193 ;
  assign n1181 = \InstQueue_reg[7][2]/NET0131  & n1016 ;
  assign n1182 = n868 & n1181 ;
  assign n1180 = \InstQueue_reg[2][2]/NET0131  & n488 ;
  assign n1178 = \InstQueue_reg[10][2]/NET0131  & n484 ;
  assign n1179 = \InstQueue_reg[3][2]/NET0131  & n458 ;
  assign n1189 = ~n1178 & ~n1179 ;
  assign n1190 = ~n1180 & n1189 ;
  assign n1174 = \InstQueue_reg[1][2]/NET0131  & n474 ;
  assign n1175 = \InstQueue_reg[4][2]/NET0131  & n476 ;
  assign n1187 = ~n1174 & ~n1175 ;
  assign n1176 = \InstQueue_reg[11][2]/NET0131  & n461 ;
  assign n1177 = \InstQueue_reg[15][2]/NET0131  & n470 ;
  assign n1188 = ~n1176 & ~n1177 ;
  assign n1191 = n1187 & n1188 ;
  assign n1195 = n1190 & n1191 ;
  assign n1196 = ~n1182 & n1195 ;
  assign n1197 = n1194 & n1196 ;
  assign n1411 = ~\InstAddrPointer_reg[1]/NET0131  & ~\InstAddrPointer_reg[2]/NET0131  ;
  assign n1412 = ~n974 & ~n1411 ;
  assign n1413 = n1197 & ~n1412 ;
  assign n1135 = \InstQueue_reg[14][3]/NET0131  & n465 ;
  assign n1136 = \InstQueue_reg[8][3]/NET0131  & n454 ;
  assign n1150 = ~n1135 & ~n1136 ;
  assign n1137 = \InstQueue_reg[9][3]/NET0131  & n486 ;
  assign n1138 = \InstQueue_reg[12][3]/NET0131  & n492 ;
  assign n1151 = ~n1137 & ~n1138 ;
  assign n1157 = n1150 & n1151 ;
  assign n1131 = \InstQueue_reg[1][3]/NET0131  & n474 ;
  assign n1132 = \InstQueue_reg[3][3]/NET0131  & n458 ;
  assign n1148 = ~n1131 & ~n1132 ;
  assign n1133 = \InstQueue_reg[6][3]/NET0131  & n490 ;
  assign n1134 = \InstQueue_reg[13][3]/NET0131  & n468 ;
  assign n1149 = ~n1133 & ~n1134 ;
  assign n1158 = n1148 & n1149 ;
  assign n1159 = n1157 & n1158 ;
  assign n1146 = \InstQueue_reg[7][3]/NET0131  & n1016 ;
  assign n1147 = n868 & n1146 ;
  assign n1145 = \InstQueue_reg[0][3]/NET0131  & n522 ;
  assign n1143 = \InstQueue_reg[15][3]/NET0131  & n470 ;
  assign n1144 = \InstQueue_reg[11][3]/NET0131  & n461 ;
  assign n1154 = ~n1143 & ~n1144 ;
  assign n1155 = ~n1145 & n1154 ;
  assign n1139 = \InstQueue_reg[2][3]/NET0131  & n488 ;
  assign n1140 = \InstQueue_reg[4][3]/NET0131  & n476 ;
  assign n1152 = ~n1139 & ~n1140 ;
  assign n1141 = \InstQueue_reg[5][3]/NET0131  & n472 ;
  assign n1142 = \InstQueue_reg[10][3]/NET0131  & n484 ;
  assign n1153 = ~n1141 & ~n1142 ;
  assign n1156 = n1152 & n1153 ;
  assign n1160 = n1155 & n1156 ;
  assign n1161 = ~n1147 & n1160 ;
  assign n1162 = n1159 & n1161 ;
  assign n1414 = ~\InstAddrPointer_reg[3]/NET0131  & ~n974 ;
  assign n1415 = ~n975 & ~n1414 ;
  assign n1416 = n1162 & ~n1415 ;
  assign n1417 = ~n1413 & ~n1416 ;
  assign n1418 = ~n1197 & n1412 ;
  assign n1206 = \InstQueue_reg[6][1]/NET0131  & n490 ;
  assign n1207 = \InstQueue_reg[13][1]/NET0131  & n468 ;
  assign n1220 = ~n1206 & ~n1207 ;
  assign n1208 = \InstQueue_reg[0][1]/NET0131  & n522 ;
  assign n1209 = \InstQueue_reg[11][1]/NET0131  & n461 ;
  assign n1221 = ~n1208 & ~n1209 ;
  assign n1228 = n1220 & n1221 ;
  assign n1202 = \InstQueue_reg[9][1]/NET0131  & n486 ;
  assign n1203 = \InstQueue_reg[12][1]/NET0131  & n492 ;
  assign n1218 = ~n1202 & ~n1203 ;
  assign n1204 = \InstQueue_reg[4][1]/NET0131  & n476 ;
  assign n1205 = \InstQueue_reg[1][1]/NET0131  & n474 ;
  assign n1219 = ~n1204 & ~n1205 ;
  assign n1229 = n1218 & n1219 ;
  assign n1230 = n1228 & n1229 ;
  assign n1214 = \InstQueue_reg[8][1]/NET0131  & n454 ;
  assign n1215 = \InstQueue_reg[3][1]/NET0131  & n458 ;
  assign n1224 = ~n1214 & ~n1215 ;
  assign n1216 = \InstQueue_reg[14][1]/NET0131  & n465 ;
  assign n1217 = \InstQueue_reg[5][1]/NET0131  & n472 ;
  assign n1225 = ~n1216 & ~n1217 ;
  assign n1226 = n1224 & n1225 ;
  assign n1210 = \InstQueue_reg[15][1]/NET0131  & n470 ;
  assign n1211 = \InstQueue_reg[2][1]/NET0131  & n488 ;
  assign n1222 = ~n1210 & ~n1211 ;
  assign n1212 = \InstQueue_reg[7][1]/NET0131  & n482 ;
  assign n1213 = \InstQueue_reg[10][1]/NET0131  & n484 ;
  assign n1223 = ~n1212 & ~n1213 ;
  assign n1227 = n1222 & n1223 ;
  assign n1231 = n1226 & n1227 ;
  assign n1232 = n1230 & n1231 ;
  assign n1236 = ~\InstAddrPointer_reg[1]/NET0131  & ~n1232 ;
  assign n1419 = \InstAddrPointer_reg[1]/NET0131  & n1232 ;
  assign n1241 = \InstQueue_reg[1][0]/NET0131  & n474 ;
  assign n1242 = \InstQueue_reg[11][0]/NET0131  & n461 ;
  assign n1255 = ~n1241 & ~n1242 ;
  assign n1243 = \InstQueue_reg[6][0]/NET0131  & n490 ;
  assign n1244 = \InstQueue_reg[0][0]/NET0131  & n522 ;
  assign n1256 = ~n1243 & ~n1244 ;
  assign n1263 = n1255 & n1256 ;
  assign n1237 = \InstQueue_reg[9][0]/NET0131  & n486 ;
  assign n1238 = \InstQueue_reg[12][0]/NET0131  & n492 ;
  assign n1253 = ~n1237 & ~n1238 ;
  assign n1239 = \InstQueue_reg[4][0]/NET0131  & n476 ;
  assign n1240 = \InstQueue_reg[14][0]/NET0131  & n465 ;
  assign n1254 = ~n1239 & ~n1240 ;
  assign n1264 = n1253 & n1254 ;
  assign n1265 = n1263 & n1264 ;
  assign n1249 = \InstQueue_reg[8][0]/NET0131  & n454 ;
  assign n1250 = \InstQueue_reg[3][0]/NET0131  & n458 ;
  assign n1259 = ~n1249 & ~n1250 ;
  assign n1251 = \InstQueue_reg[13][0]/NET0131  & n468 ;
  assign n1252 = \InstQueue_reg[5][0]/NET0131  & n472 ;
  assign n1260 = ~n1251 & ~n1252 ;
  assign n1261 = n1259 & n1260 ;
  assign n1245 = \InstQueue_reg[15][0]/NET0131  & n470 ;
  assign n1246 = \InstQueue_reg[2][0]/NET0131  & n488 ;
  assign n1257 = ~n1245 & ~n1246 ;
  assign n1247 = \InstQueue_reg[7][0]/NET0131  & n482 ;
  assign n1248 = \InstQueue_reg[10][0]/NET0131  & n484 ;
  assign n1258 = ~n1247 & ~n1248 ;
  assign n1262 = n1257 & n1258 ;
  assign n1266 = n1261 & n1262 ;
  assign n1267 = n1265 & n1266 ;
  assign n1420 = \InstAddrPointer_reg[0]/NET0131  & ~n1267 ;
  assign n1421 = ~n1419 & n1420 ;
  assign n1422 = ~n1236 & ~n1421 ;
  assign n1423 = ~n1418 & n1422 ;
  assign n1424 = n1417 & ~n1423 ;
  assign n1425 = ~n1124 & n1409 ;
  assign n1426 = ~n1162 & n1415 ;
  assign n1427 = ~n1425 & ~n1426 ;
  assign n1428 = ~n1424 & n1427 ;
  assign n1429 = ~n1410 & ~n1428 ;
  assign n988 = \InstQueue_reg[1][7]/NET0131  & n474 ;
  assign n989 = \InstQueue_reg[8][7]/NET0131  & n454 ;
  assign n1002 = ~n988 & ~n989 ;
  assign n990 = \InstQueue_reg[14][7]/NET0131  & n465 ;
  assign n991 = \InstQueue_reg[7][7]/NET0131  & n482 ;
  assign n1003 = ~n990 & ~n991 ;
  assign n1010 = n1002 & n1003 ;
  assign n984 = \InstQueue_reg[10][7]/NET0131  & n484 ;
  assign n985 = \InstQueue_reg[4][7]/NET0131  & n476 ;
  assign n1000 = ~n984 & ~n985 ;
  assign n986 = \InstQueue_reg[12][7]/NET0131  & n492 ;
  assign n987 = \InstQueue_reg[3][7]/NET0131  & n458 ;
  assign n1001 = ~n986 & ~n987 ;
  assign n1011 = n1000 & n1001 ;
  assign n1012 = n1010 & n1011 ;
  assign n996 = \InstQueue_reg[11][7]/NET0131  & n461 ;
  assign n997 = \InstQueue_reg[0][7]/NET0131  & n522 ;
  assign n1006 = ~n996 & ~n997 ;
  assign n998 = \InstQueue_reg[15][7]/NET0131  & n470 ;
  assign n999 = \InstQueue_reg[6][7]/NET0131  & n490 ;
  assign n1007 = ~n998 & ~n999 ;
  assign n1008 = n1006 & n1007 ;
  assign n992 = \InstQueue_reg[2][7]/NET0131  & n488 ;
  assign n993 = \InstQueue_reg[5][7]/NET0131  & n472 ;
  assign n1004 = ~n992 & ~n993 ;
  assign n994 = \InstQueue_reg[9][7]/NET0131  & n486 ;
  assign n995 = \InstQueue_reg[13][7]/NET0131  & n468 ;
  assign n1005 = ~n994 & ~n995 ;
  assign n1009 = n1004 & n1005 ;
  assign n1013 = n1008 & n1009 ;
  assign n1014 = n1012 & n1013 ;
  assign n1430 = \InstAddrPointer_reg[6]/NET0131  & n1291 ;
  assign n1431 = ~\InstAddrPointer_reg[7]/NET0131  & ~n1430 ;
  assign n1432 = ~n1292 & ~n1431 ;
  assign n1433 = n1014 & ~n1432 ;
  assign n1434 = \InstAddrPointer_reg[8]/NET0131  & n1292 ;
  assign n1435 = ~\InstAddrPointer_reg[8]/NET0131  & ~n1292 ;
  assign n1436 = ~n1434 & ~n1435 ;
  assign n1437 = ~n1433 & n1436 ;
  assign n1022 = \InstQueue_reg[0][6]/NET0131  & n522 ;
  assign n1023 = \InstQueue_reg[14][6]/NET0131  & n465 ;
  assign n1036 = ~n1022 & ~n1023 ;
  assign n1024 = \InstQueue_reg[8][6]/NET0131  & n454 ;
  assign n1025 = \InstQueue_reg[9][6]/NET0131  & n486 ;
  assign n1037 = ~n1024 & ~n1025 ;
  assign n1026 = \InstQueue_reg[6][6]/NET0131  & n490 ;
  assign n1027 = \InstQueue_reg[15][6]/NET0131  & n470 ;
  assign n1038 = ~n1026 & ~n1027 ;
  assign n1045 = n1037 & n1038 ;
  assign n1046 = n1036 & n1045 ;
  assign n1032 = \InstQueue_reg[11][6]/NET0131  & n461 ;
  assign n1033 = \InstQueue_reg[10][6]/NET0131  & n484 ;
  assign n1041 = ~n1032 & ~n1033 ;
  assign n1034 = \InstQueue_reg[2][6]/NET0131  & n488 ;
  assign n1035 = \InstQueue_reg[12][6]/NET0131  & n492 ;
  assign n1042 = ~n1034 & ~n1035 ;
  assign n1043 = n1041 & n1042 ;
  assign n1028 = \InstQueue_reg[3][6]/NET0131  & n458 ;
  assign n1029 = \InstQueue_reg[1][6]/NET0131  & n474 ;
  assign n1039 = ~n1028 & ~n1029 ;
  assign n1030 = \InstQueue_reg[4][6]/NET0131  & n476 ;
  assign n1031 = \InstQueue_reg[5][6]/NET0131  & n472 ;
  assign n1040 = ~n1030 & ~n1031 ;
  assign n1044 = n1039 & n1040 ;
  assign n1047 = n1043 & n1044 ;
  assign n1017 = \InstQueue_reg[7][6]/NET0131  & n1016 ;
  assign n1018 = n868 & n1017 ;
  assign n1020 = \InstQueue_reg[13][6]/NET0131  & n467 ;
  assign n1021 = n1019 & n1020 ;
  assign n1048 = ~n1018 & ~n1021 ;
  assign n1049 = n1047 & n1048 ;
  assign n1050 = n1046 & n1049 ;
  assign n1438 = ~\InstAddrPointer_reg[6]/NET0131  & ~n1291 ;
  assign n1439 = ~n1430 & ~n1438 ;
  assign n1440 = n1050 & ~n1439 ;
  assign n1062 = \InstQueue_reg[8][5]/NET0131  & n454 ;
  assign n1063 = \InstQueue_reg[0][5]/NET0131  & n522 ;
  assign n1076 = ~n1062 & ~n1063 ;
  assign n1064 = \InstQueue_reg[4][5]/NET0131  & n476 ;
  assign n1065 = \InstQueue_reg[10][5]/NET0131  & n484 ;
  assign n1077 = ~n1064 & ~n1065 ;
  assign n1084 = n1076 & n1077 ;
  assign n1058 = \InstQueue_reg[7][5]/NET0131  & n482 ;
  assign n1059 = \InstQueue_reg[12][5]/NET0131  & n492 ;
  assign n1074 = ~n1058 & ~n1059 ;
  assign n1060 = \InstQueue_reg[9][5]/NET0131  & n486 ;
  assign n1061 = \InstQueue_reg[6][5]/NET0131  & n490 ;
  assign n1075 = ~n1060 & ~n1061 ;
  assign n1085 = n1074 & n1075 ;
  assign n1086 = n1084 & n1085 ;
  assign n1070 = \InstQueue_reg[1][5]/NET0131  & n474 ;
  assign n1071 = \InstQueue_reg[11][5]/NET0131  & n461 ;
  assign n1080 = ~n1070 & ~n1071 ;
  assign n1072 = \InstQueue_reg[3][5]/NET0131  & n458 ;
  assign n1073 = \InstQueue_reg[5][5]/NET0131  & n472 ;
  assign n1081 = ~n1072 & ~n1073 ;
  assign n1082 = n1080 & n1081 ;
  assign n1066 = \InstQueue_reg[2][5]/NET0131  & n488 ;
  assign n1067 = \InstQueue_reg[14][5]/NET0131  & n465 ;
  assign n1078 = ~n1066 & ~n1067 ;
  assign n1068 = \InstQueue_reg[13][5]/NET0131  & n468 ;
  assign n1069 = \InstQueue_reg[15][5]/NET0131  & n470 ;
  assign n1079 = ~n1068 & ~n1069 ;
  assign n1083 = n1078 & n1079 ;
  assign n1087 = n1082 & n1083 ;
  assign n1088 = n1086 & n1087 ;
  assign n1441 = ~\InstAddrPointer_reg[5]/NET0131  & ~n976 ;
  assign n1442 = ~n1291 & ~n1441 ;
  assign n1443 = n1088 & ~n1442 ;
  assign n1444 = ~n1440 & ~n1443 ;
  assign n1445 = n1437 & n1444 ;
  assign n1446 = n1429 & n1445 ;
  assign n1447 = ~n1014 & n1432 ;
  assign n1448 = ~n1050 & n1439 ;
  assign n1449 = ~n1088 & n1442 ;
  assign n1450 = ~n1440 & n1449 ;
  assign n1451 = ~n1448 & ~n1450 ;
  assign n1452 = ~n1447 & n1451 ;
  assign n1453 = n1437 & ~n1452 ;
  assign n1454 = ~n1446 & ~n1453 ;
  assign n1331 = \InstAddrPointer_reg[20]/NET0131  & n1330 ;
  assign n1455 = ~\InstAddrPointer_reg[20]/NET0131  & ~n1330 ;
  assign n1456 = ~n1331 & ~n1455 ;
  assign n1347 = \InstAddrPointer_reg[17]/NET0131  & n1329 ;
  assign n1348 = \InstAddrPointer_reg[18]/NET0131  & n1347 ;
  assign n1466 = ~\InstAddrPointer_reg[18]/NET0131  & ~n1347 ;
  assign n1467 = ~n1348 & ~n1466 ;
  assign n1468 = \InstAddrPointer_reg[14]/NET0131  & n1298 ;
  assign n1469 = ~\InstAddrPointer_reg[15]/NET0131  & ~n1468 ;
  assign n1470 = n1298 & n1327 ;
  assign n1471 = ~n1469 & ~n1470 ;
  assign n1472 = \InstAddrPointer_reg[16]/NET0131  & n1471 ;
  assign n1473 = \InstAddrPointer_reg[17]/NET0131  & n1472 ;
  assign n1474 = n1467 & n1473 ;
  assign n1464 = ~\InstAddrPointer_reg[19]/NET0131  & ~n1348 ;
  assign n1465 = ~n1330 & ~n1464 ;
  assign n1457 = \InstAddrPointer_reg[10]/NET0131  & \InstAddrPointer_reg[11]/NET0131  ;
  assign n1303 = n1295 & n1296 ;
  assign n1458 = \InstAddrPointer_reg[11]/NET0131  & n1295 ;
  assign n1459 = ~\InstAddrPointer_reg[12]/NET0131  & ~n1458 ;
  assign n1460 = ~n1303 & ~n1459 ;
  assign n1461 = \InstAddrPointer_reg[13]/NET0131  & \InstAddrPointer_reg[14]/NET0131  ;
  assign n1462 = n1460 & n1461 ;
  assign n1463 = n1457 & n1462 ;
  assign n1475 = ~\InstAddrPointer_reg[9]/NET0131  & ~n1434 ;
  assign n1476 = n1292 & n1293 ;
  assign n1477 = ~n1475 & ~n1476 ;
  assign n1478 = n1463 & n1477 ;
  assign n1479 = n1465 & n1478 ;
  assign n1480 = n1474 & n1479 ;
  assign n1481 = n1456 & n1480 ;
  assign n1482 = ~n1454 & n1481 ;
  assign n1483 = \InstAddrPointer_reg[21]/NET0131  & n1331 ;
  assign n1484 = ~\InstAddrPointer_reg[21]/NET0131  & ~n1331 ;
  assign n1485 = ~n1483 & ~n1484 ;
  assign n1486 = \InstAddrPointer_reg[22]/NET0131  & n1485 ;
  assign n1487 = n1482 & n1486 ;
  assign n1491 = n1386 & n1490 ;
  assign n1370 = \InstAddrPointer_reg[23]/NET0131  & \InstAddrPointer_reg[24]/NET0131  ;
  assign n1378 = \InstAddrPointer_reg[25]/NET0131  & n1370 ;
  assign n1383 = \InstAddrPointer_reg[26]/NET0131  & n1378 ;
  assign n1492 = n1331 & n1362 ;
  assign n1493 = n1383 & n1492 ;
  assign n1494 = ~\InstAddrPointer_reg[27]/NET0131  & ~n1493 ;
  assign n1495 = ~n1491 & ~n1494 ;
  assign n1496 = ~\InstAddrPointer_reg[24]/NET0131  & ~n1488 ;
  assign n1497 = ~n1489 & ~n1496 ;
  assign n1498 = \InstAddrPointer_reg[25]/NET0131  & n1497 ;
  assign n1499 = \InstAddrPointer_reg[26]/NET0131  & n1498 ;
  assign n1500 = n1495 & n1499 ;
  assign n1501 = ~\InstAddrPointer_reg[23]/NET0131  & ~n1492 ;
  assign n1502 = ~n1488 & ~n1501 ;
  assign n1503 = \InstAddrPointer_reg[28]/NET0131  & n1502 ;
  assign n1504 = n1500 & n1503 ;
  assign n1508 = ~\InstAddrPointer_reg[29]/NET0131  & ~n1506 ;
  assign n1509 = ~n1507 & ~n1508 ;
  assign n1510 = n1504 & n1509 ;
  assign n1516 = n1487 & n1510 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1511 = \InstAddrPointer_reg[30]/NET0131  & n1510 ;
  assign n1512 = n1487 & n1511 ;
  assign n1518 = n1014 & ~n1512 ;
  assign n1519 = ~n1517 & n1518 ;
  assign n977 = \InstAddrPointer_reg[0]/NET0131  & n976 ;
  assign n978 = \InstAddrPointer_reg[5]/NET0131  & n977 ;
  assign n979 = \InstAddrPointer_reg[6]/NET0131  & n978 ;
  assign n980 = ~\InstAddrPointer_reg[7]/NET0131  & ~n979 ;
  assign n982 = n978 & n981 ;
  assign n983 = ~n980 & ~n982 ;
  assign n1015 = ~n983 & n1014 ;
  assign n1051 = ~\InstAddrPointer_reg[6]/NET0131  & ~n978 ;
  assign n1052 = ~n979 & ~n1051 ;
  assign n1053 = n1050 & ~n1052 ;
  assign n1054 = ~n1015 & ~n1053 ;
  assign n1055 = ~n1050 & n1052 ;
  assign n1125 = \InstAddrPointer_reg[0]/NET0131  & \InstAddrPointer_reg[1]/NET0131  ;
  assign n1126 = \InstAddrPointer_reg[2]/NET0131  & n1125 ;
  assign n1127 = \InstAddrPointer_reg[3]/NET0131  & n1126 ;
  assign n1163 = ~\InstAddrPointer_reg[3]/NET0131  & ~n1126 ;
  assign n1164 = ~n1127 & ~n1163 ;
  assign n1165 = n1162 & ~n1164 ;
  assign n1198 = ~\InstAddrPointer_reg[2]/NET0131  & ~n1125 ;
  assign n1199 = ~n1126 & ~n1198 ;
  assign n1200 = n1197 & ~n1199 ;
  assign n1201 = ~n1165 & ~n1200 ;
  assign n1233 = ~\InstAddrPointer_reg[0]/NET0131  & ~\InstAddrPointer_reg[1]/NET0131  ;
  assign n1234 = ~n1125 & ~n1233 ;
  assign n1235 = n1232 & ~n1234 ;
  assign n1268 = \InstAddrPointer_reg[0]/NET0131  & n1267 ;
  assign n1269 = ~n1236 & n1268 ;
  assign n1270 = ~n1235 & ~n1269 ;
  assign n1271 = n1201 & n1270 ;
  assign n1272 = ~n1162 & n1164 ;
  assign n1273 = ~n1197 & n1199 ;
  assign n1274 = ~n1165 & n1273 ;
  assign n1275 = ~n1272 & ~n1274 ;
  assign n1276 = ~n1271 & n1275 ;
  assign n1056 = ~\InstAddrPointer_reg[5]/NET0131  & ~n977 ;
  assign n1057 = ~n978 & ~n1056 ;
  assign n1089 = ~n1057 & n1088 ;
  assign n1128 = ~\InstAddrPointer_reg[4]/NET0131  & ~n1127 ;
  assign n1129 = ~n977 & ~n1128 ;
  assign n1130 = n1124 & ~n1129 ;
  assign n1277 = ~n1089 & ~n1130 ;
  assign n1278 = ~n1276 & n1277 ;
  assign n1279 = n1057 & ~n1088 ;
  assign n1280 = ~n1124 & n1129 ;
  assign n1281 = ~n1089 & n1280 ;
  assign n1282 = ~n1279 & ~n1281 ;
  assign n1283 = ~n1278 & n1282 ;
  assign n1284 = ~n1055 & n1283 ;
  assign n1285 = n1054 & ~n1284 ;
  assign n1304 = \InstAddrPointer_reg[0]/NET0131  & n1303 ;
  assign n1308 = n982 & n1293 ;
  assign n1309 = \InstAddrPointer_reg[10]/NET0131  & n1308 ;
  assign n1310 = \InstAddrPointer_reg[11]/NET0131  & n1309 ;
  assign n1311 = ~\InstAddrPointer_reg[12]/NET0131  & ~n1310 ;
  assign n1312 = ~n1304 & ~n1311 ;
  assign n1287 = \InstAddrPointer_reg[8]/NET0131  & n982 ;
  assign n1313 = ~\InstAddrPointer_reg[9]/NET0131  & ~n1287 ;
  assign n1314 = ~n1308 & ~n1313 ;
  assign n1315 = ~\InstAddrPointer_reg[10]/NET0131  & ~n1308 ;
  assign n1316 = ~n1309 & ~n1315 ;
  assign n1317 = ~n1314 & ~n1316 ;
  assign n1318 = ~\InstAddrPointer_reg[11]/NET0131  & ~n1309 ;
  assign n1319 = ~n1310 & ~n1318 ;
  assign n1320 = n1317 & ~n1319 ;
  assign n1321 = ~n1312 & n1320 ;
  assign n1286 = ~\InstAddrPointer_reg[8]/NET0131  & ~n982 ;
  assign n1288 = ~n1286 & ~n1287 ;
  assign n1289 = n983 & ~n1014 ;
  assign n1290 = ~n1288 & ~n1289 ;
  assign n1299 = \InstAddrPointer_reg[0]/NET0131  & n1298 ;
  assign n1300 = ~\InstAddrPointer_reg[14]/NET0131  & ~n1299 ;
  assign n1301 = \InstAddrPointer_reg[14]/NET0131  & n1299 ;
  assign n1302 = ~n1300 & ~n1301 ;
  assign n1305 = ~\InstAddrPointer_reg[13]/NET0131  & ~n1304 ;
  assign n1306 = ~n1299 & ~n1305 ;
  assign n1307 = ~n1302 & ~n1306 ;
  assign n1322 = n1290 & n1307 ;
  assign n1323 = n1321 & n1322 ;
  assign n1324 = ~n1285 & n1323 ;
  assign n1332 = \InstAddrPointer_reg[0]/NET0131  & n1331 ;
  assign n1333 = ~\InstAddrPointer_reg[21]/NET0131  & ~n1332 ;
  assign n1334 = \InstAddrPointer_reg[21]/NET0131  & n1332 ;
  assign n1335 = ~n1333 & ~n1334 ;
  assign n1336 = \InstAddrPointer_reg[0]/NET0131  & n1330 ;
  assign n1337 = ~\InstAddrPointer_reg[20]/NET0131  & ~n1336 ;
  assign n1338 = ~n1332 & ~n1337 ;
  assign n1339 = ~n1335 & ~n1338 ;
  assign n1340 = ~\InstAddrPointer_reg[15]/NET0131  & ~n1301 ;
  assign n1341 = n1299 & n1327 ;
  assign n1342 = ~n1340 & ~n1341 ;
  assign n1343 = ~\InstAddrPointer_reg[16]/NET0131  & ~n1341 ;
  assign n1344 = n1299 & n1328 ;
  assign n1345 = ~n1343 & ~n1344 ;
  assign n1346 = ~n1342 & ~n1345 ;
  assign n1349 = \InstAddrPointer_reg[0]/NET0131  & n1348 ;
  assign n1350 = ~\InstAddrPointer_reg[19]/NET0131  & ~n1349 ;
  assign n1351 = ~n1336 & ~n1350 ;
  assign n1352 = ~\InstAddrPointer_reg[17]/NET0131  & ~n1344 ;
  assign n1353 = \InstAddrPointer_reg[0]/NET0131  & n1347 ;
  assign n1354 = ~n1352 & ~n1353 ;
  assign n1355 = ~\InstAddrPointer_reg[18]/NET0131  & ~n1353 ;
  assign n1356 = ~n1349 & ~n1355 ;
  assign n1357 = ~n1354 & ~n1356 ;
  assign n1358 = ~n1351 & n1357 ;
  assign n1359 = n1346 & n1358 ;
  assign n1360 = n1339 & n1359 ;
  assign n1361 = n1324 & n1360 ;
  assign n1363 = n1332 & n1362 ;
  assign n1364 = ~\InstAddrPointer_reg[23]/NET0131  & ~n1363 ;
  assign n1367 = n1336 & n1366 ;
  assign n1368 = ~n1364 & ~n1367 ;
  assign n1369 = ~\InstAddrPointer_reg[24]/NET0131  & ~n1367 ;
  assign n1371 = n1363 & n1370 ;
  assign n1372 = ~n1369 & ~n1371 ;
  assign n1373 = ~n1368 & ~n1372 ;
  assign n1374 = ~\InstAddrPointer_reg[22]/NET0131  & ~n1334 ;
  assign n1375 = ~n1363 & ~n1374 ;
  assign n1376 = n1373 & ~n1375 ;
  assign n1377 = ~\InstAddrPointer_reg[25]/NET0131  & ~n1371 ;
  assign n1379 = n1363 & n1378 ;
  assign n1380 = ~n1377 & ~n1379 ;
  assign n1381 = n1376 & ~n1380 ;
  assign n1382 = n1361 & n1381 ;
  assign n1384 = n1363 & n1383 ;
  assign n1385 = ~\InstAddrPointer_reg[27]/NET0131  & ~n1384 ;
  assign n1387 = n1379 & n1386 ;
  assign n1388 = ~n1385 & ~n1387 ;
  assign n1389 = ~\InstAddrPointer_reg[28]/NET0131  & ~n1387 ;
  assign n1390 = \InstAddrPointer_reg[28]/NET0131  & n1387 ;
  assign n1391 = ~n1389 & ~n1390 ;
  assign n1392 = ~n1388 & ~n1391 ;
  assign n1393 = ~\InstAddrPointer_reg[29]/NET0131  & ~n1390 ;
  assign n1394 = \InstAddrPointer_reg[29]/NET0131  & n1390 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = n1392 & ~n1395 ;
  assign n1397 = ~\InstAddrPointer_reg[26]/NET0131  & ~n1379 ;
  assign n1398 = ~n1384 & ~n1397 ;
  assign n1399 = n1396 & ~n1398 ;
  assign n1400 = n1382 & n1399 ;
  assign n1401 = ~\InstAddrPointer_reg[30]/NET0131  & ~n1394 ;
  assign n1402 = \InstAddrPointer_reg[30]/NET0131  & n1394 ;
  assign n1403 = ~n1401 & ~n1402 ;
  assign n1404 = ~n1014 & n1403 ;
  assign n1405 = ~n1400 & n1404 ;
  assign n1406 = ~n1014 & ~n1403 ;
  assign n1407 = n1400 & n1406 ;
  assign n1520 = ~n1405 & ~n1407 ;
  assign n1521 = ~n1519 & n1520 ;
  assign n1522 = ~n906 & ~n1521 ;
  assign n1523 = ~n973 & ~n1522 ;
  assign n1524 = n773 & ~n1523 ;
  assign n1525 = \InstAddrPointer_reg[3]/NET0131  & ~n1198 ;
  assign n1526 = \InstAddrPointer_reg[4]/NET0131  & n1525 ;
  assign n1527 = \InstAddrPointer_reg[5]/NET0131  & n1526 ;
  assign n1528 = \InstAddrPointer_reg[6]/NET0131  & n1527 ;
  assign n1529 = \InstAddrPointer_reg[7]/NET0131  & n1528 ;
  assign n1530 = n1294 & n1529 ;
  assign n1531 = n1297 & n1530 ;
  assign n1532 = n1328 & n1531 ;
  assign n1533 = n1326 & n1532 ;
  assign n1534 = \InstAddrPointer_reg[20]/NET0131  & n1533 ;
  assign n1535 = n1365 & n1534 ;
  assign n1536 = \InstAddrPointer_reg[24]/NET0131  & n1535 ;
  assign n1537 = \InstAddrPointer_reg[25]/NET0131  & n1536 ;
  assign n1538 = ~\InstAddrPointer_reg[26]/NET0131  & ~n1537 ;
  assign n1539 = n1362 & n1534 ;
  assign n1540 = n1383 & n1539 ;
  assign n1541 = ~n1538 & ~n1540 ;
  assign n1542 = ~\InstAddrPointer_reg[7]/NET0131  & ~n1528 ;
  assign n1543 = ~n1529 & ~n1542 ;
  assign n1544 = n1014 & ~n1543 ;
  assign n1545 = \InstAddrPointer_reg[8]/NET0131  & n1529 ;
  assign n1546 = ~\InstAddrPointer_reg[8]/NET0131  & ~n1529 ;
  assign n1547 = ~n1545 & ~n1546 ;
  assign n1548 = ~n1544 & n1547 ;
  assign n1549 = ~\InstAddrPointer_reg[6]/NET0131  & ~n1527 ;
  assign n1550 = ~n1528 & ~n1549 ;
  assign n1551 = n1050 & ~n1550 ;
  assign n1552 = ~\InstAddrPointer_reg[5]/NET0131  & ~n1526 ;
  assign n1553 = ~n1527 & ~n1552 ;
  assign n1554 = n1088 & ~n1553 ;
  assign n1555 = ~n1551 & ~n1554 ;
  assign n1556 = ~\InstAddrPointer_reg[4]/NET0131  & ~n1525 ;
  assign n1557 = ~n1526 & ~n1556 ;
  assign n1558 = n1124 & ~n1557 ;
  assign n1559 = ~\InstAddrPointer_reg[3]/NET0131  & n1198 ;
  assign n1560 = ~n1525 & ~n1559 ;
  assign n1561 = n1162 & ~n1560 ;
  assign n1562 = ~n1558 & ~n1561 ;
  assign n1563 = ~n1162 & n1560 ;
  assign n1564 = n1197 & n1199 ;
  assign n1565 = ~n1197 & ~n1199 ;
  assign n1566 = ~n1232 & n1234 ;
  assign n1567 = ~\InstAddrPointer_reg[0]/NET0131  & ~n1267 ;
  assign n1568 = ~n1566 & ~n1567 ;
  assign n1569 = ~n1235 & ~n1568 ;
  assign n1570 = ~n1565 & ~n1569 ;
  assign n1571 = ~n1564 & ~n1570 ;
  assign n1572 = ~n1563 & ~n1571 ;
  assign n1573 = n1562 & ~n1572 ;
  assign n1574 = ~n1124 & n1557 ;
  assign n1575 = ~n1088 & n1553 ;
  assign n1576 = ~n1574 & ~n1575 ;
  assign n1577 = ~n1573 & n1576 ;
  assign n1578 = n1555 & ~n1577 ;
  assign n1579 = ~n1050 & n1550 ;
  assign n1580 = ~n1014 & n1543 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1582 = ~n1578 & n1581 ;
  assign n1583 = n1548 & ~n1582 ;
  assign n1584 = ~\InstAddrPointer_reg[17]/NET0131  & ~n1532 ;
  assign n1585 = \InstAddrPointer_reg[17]/NET0131  & n1532 ;
  assign n1586 = ~n1584 & ~n1585 ;
  assign n1589 = \InstAddrPointer_reg[9]/NET0131  & n1545 ;
  assign n1590 = n1457 & n1589 ;
  assign n1591 = ~\InstAddrPointer_reg[12]/NET0131  & ~n1590 ;
  assign n1592 = \InstAddrPointer_reg[12]/NET0131  & n1590 ;
  assign n1593 = ~n1591 & ~n1592 ;
  assign n1594 = \InstAddrPointer_reg[13]/NET0131  & n1593 ;
  assign n1595 = ~\InstAddrPointer_reg[9]/NET0131  & ~n1545 ;
  assign n1596 = ~n1589 & ~n1595 ;
  assign n1597 = \InstAddrPointer_reg[10]/NET0131  & n1596 ;
  assign n1598 = \InstAddrPointer_reg[14]/NET0131  & n1597 ;
  assign n1599 = n1594 & n1598 ;
  assign n1587 = \InstAddrPointer_reg[14]/NET0131  & n1531 ;
  assign n1588 = ~\InstAddrPointer_reg[15]/NET0131  & ~n1587 ;
  assign n1600 = \InstAddrPointer_reg[11]/NET0131  & ~n1588 ;
  assign n1601 = n1599 & n1600 ;
  assign n1602 = \InstAddrPointer_reg[16]/NET0131  & ~n1530 ;
  assign n1603 = n1601 & n1602 ;
  assign n1604 = n1586 & n1603 ;
  assign n1605 = n1583 & n1604 ;
  assign n1606 = ~\InstAddrPointer_reg[18]/NET0131  & ~n1585 ;
  assign n1607 = \InstAddrPointer_reg[18]/NET0131  & n1585 ;
  assign n1608 = ~n1606 & ~n1607 ;
  assign n1609 = n1605 & n1608 ;
  assign n1610 = \InstAddrPointer_reg[21]/NET0131  & n1534 ;
  assign n1611 = ~\InstAddrPointer_reg[21]/NET0131  & ~n1534 ;
  assign n1612 = ~n1610 & ~n1611 ;
  assign n1613 = \InstAddrPointer_reg[22]/NET0131  & n1612 ;
  assign n1614 = \InstAddrPointer_reg[23]/NET0131  & n1613 ;
  assign n1615 = ~\InstAddrPointer_reg[24]/NET0131  & ~n1535 ;
  assign n1616 = ~n1536 & ~n1615 ;
  assign n1617 = n1614 & n1616 ;
  assign n1618 = ~\InstAddrPointer_reg[19]/NET0131  & ~n1607 ;
  assign n1619 = ~n1533 & ~n1618 ;
  assign n1620 = \InstAddrPointer_reg[20]/NET0131  & n1619 ;
  assign n1621 = \InstAddrPointer_reg[25]/NET0131  & n1620 ;
  assign n1622 = n1617 & n1621 ;
  assign n1623 = n1609 & n1622 ;
  assign n1624 = n1541 & n1623 ;
  assign n1625 = ~\InstAddrPointer_reg[27]/NET0131  & ~n1540 ;
  assign n1626 = \InstAddrPointer_reg[27]/NET0131  & n1540 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = \InstAddrPointer_reg[28]/NET0131  & n1627 ;
  assign n1629 = \InstAddrPointer_reg[29]/NET0131  & n1628 ;
  assign n1630 = n1624 & n1629 ;
  assign n1631 = n1505 & n1537 ;
  assign n1632 = \InstAddrPointer_reg[29]/NET0131  & n1631 ;
  assign n1633 = ~\InstAddrPointer_reg[30]/NET0131  & ~n1632 ;
  assign n1634 = \InstAddrPointer_reg[30]/NET0131  & n1632 ;
  assign n1635 = ~n1633 & ~n1634 ;
  assign n1636 = ~n1630 & ~n1635 ;
  assign n1637 = n1629 & n1635 ;
  assign n1638 = n1624 & n1637 ;
  assign n1639 = n899 & ~n1638 ;
  assign n1640 = ~n1636 & n1639 ;
  assign n1647 = n766 & n1635 ;
  assign n1646 = ~n811 & n1403 ;
  assign n1641 = n828 & ~n836 ;
  assign n1642 = n912 & ~n1641 ;
  assign n1643 = ~n785 & ~n846 ;
  assign n1644 = n1642 & ~n1643 ;
  assign n1645 = \InstAddrPointer_reg[30]/NET0131  & ~n1644 ;
  assign n1648 = ~n873 & n1515 ;
  assign n1649 = ~n1645 & ~n1648 ;
  assign n1650 = ~n1646 & n1649 ;
  assign n1651 = ~n1647 & n1650 ;
  assign n1652 = ~n1640 & n1651 ;
  assign n1653 = ~n1524 & n1652 ;
  assign n1654 = n929 & ~n1653 ;
  assign n1655 = n931 & n935 ;
  assign n1656 = \rEIP_reg[30]/NET0131  & n1655 ;
  assign n1657 = \State2_reg[1]/NET0131  & \State2_reg[3]/NET0131  ;
  assign n1658 = ~\State2_reg[2]/NET0131  & ~n931 ;
  assign n1659 = ~\State2_reg[1]/NET0131  & ~n940 ;
  assign n1660 = ~n1658 & n1659 ;
  assign n1661 = ~n1657 & ~n1660 ;
  assign n1662 = \InstAddrPointer_reg[30]/NET0131  & n1661 ;
  assign n1663 = ~n1656 & ~n1662 ;
  assign n1664 = ~n1654 & n1663 ;
  assign n1665 = \InstAddrPointer_reg[29]/NET0131  & n906 ;
  assign n1674 = ~n1270 & ~n1273 ;
  assign n1675 = ~n1130 & n1201 ;
  assign n1676 = ~n1674 & n1675 ;
  assign n1677 = ~n1130 & n1272 ;
  assign n1678 = ~n1280 & ~n1677 ;
  assign n1679 = ~n1676 & n1678 ;
  assign n1680 = n1054 & ~n1089 ;
  assign n1681 = ~n1679 & n1680 ;
  assign n1671 = ~n1053 & n1279 ;
  assign n1672 = ~n1055 & ~n1671 ;
  assign n1673 = ~n1015 & ~n1672 ;
  assign n1682 = n1290 & ~n1673 ;
  assign n1683 = ~n1681 & n1682 ;
  assign n1684 = n1321 & n1683 ;
  assign n1685 = n1307 & n1346 ;
  assign n1686 = ~n1338 & n1685 ;
  assign n1687 = n1358 & n1686 ;
  assign n1688 = n1684 & n1687 ;
  assign n1689 = ~n1335 & n1688 ;
  assign n1690 = n1376 & n1689 ;
  assign n1691 = ~n1380 & ~n1398 ;
  assign n1692 = n1392 & n1691 ;
  assign n1693 = n1690 & n1692 ;
  assign n1695 = ~n1395 & n1693 ;
  assign n1694 = n1395 & ~n1693 ;
  assign n1696 = ~n1014 & ~n1694 ;
  assign n1697 = ~n1695 & n1696 ;
  assign n1666 = n1487 & n1504 ;
  assign n1668 = n1509 & ~n1666 ;
  assign n1667 = ~n1509 & n1666 ;
  assign n1669 = n1014 & ~n1667 ;
  assign n1670 = ~n1668 & n1669 ;
  assign n1698 = ~n906 & ~n1670 ;
  assign n1699 = ~n1697 & n1698 ;
  assign n1700 = ~n1665 & ~n1699 ;
  assign n1701 = n773 & ~n1700 ;
  assign n1702 = ~\InstAddrPointer_reg[29]/NET0131  & ~n1631 ;
  assign n1703 = ~n1632 & ~n1702 ;
  assign n1704 = n1562 & n1571 ;
  assign n1705 = ~n1558 & n1563 ;
  assign n1706 = ~n1574 & ~n1705 ;
  assign n1707 = ~n1704 & n1706 ;
  assign n1708 = n1555 & ~n1707 ;
  assign n1709 = ~n1551 & n1575 ;
  assign n1710 = ~n1579 & ~n1709 ;
  assign n1711 = ~n1708 & n1710 ;
  assign n1712 = ~n1580 & n1711 ;
  assign n1713 = n1548 & ~n1712 ;
  assign n1714 = n1603 & n1713 ;
  assign n1715 = \InstAddrPointer_reg[18]/NET0131  & n1586 ;
  assign n1716 = n1620 & n1715 ;
  assign n1717 = n1714 & n1716 ;
  assign n1718 = n1617 & n1717 ;
  assign n1719 = ~\InstAddrPointer_reg[25]/NET0131  & ~n1536 ;
  assign n1720 = ~n1537 & ~n1719 ;
  assign n1721 = \InstAddrPointer_reg[26]/NET0131  & n1720 ;
  assign n1722 = n1628 & n1721 ;
  assign n1723 = n1718 & n1722 ;
  assign n1725 = ~n1703 & ~n1723 ;
  assign n1724 = n1703 & n1723 ;
  assign n1726 = n899 & ~n1724 ;
  assign n1727 = ~n1725 & n1726 ;
  assign n1736 = ~\InstAddrPointer_reg[29]/NET0131  & ~n765 ;
  assign n1737 = ~n740 & ~n1736 ;
  assign n1738 = n1703 & n1737 ;
  assign n1732 = ~n785 & n834 ;
  assign n1733 = ~n859 & ~n1732 ;
  assign n1734 = n1642 & n1733 ;
  assign n1735 = \InstAddrPointer_reg[29]/NET0131  & ~n1734 ;
  assign n1728 = ~n811 & n1395 ;
  assign n1729 = ~n858 & ~n1506 ;
  assign n1730 = n873 & ~n1729 ;
  assign n1731 = n1509 & ~n1730 ;
  assign n1739 = ~n1728 & ~n1731 ;
  assign n1740 = ~n1735 & n1739 ;
  assign n1741 = ~n1738 & n1740 ;
  assign n1742 = ~n1727 & n1741 ;
  assign n1743 = ~n1701 & n1742 ;
  assign n1744 = n929 & ~n1743 ;
  assign n1745 = \rEIP_reg[29]/NET0131  & n1655 ;
  assign n1746 = \InstAddrPointer_reg[29]/NET0131  & n1661 ;
  assign n1747 = ~n1745 & ~n1746 ;
  assign n1748 = ~n1744 & n1747 ;
  assign n1749 = \InstAddrPointer_reg[27]/NET0131  & n906 ;
  assign n1766 = ~\InstAddrPointer_reg[11]/NET0131  & ~n1295 ;
  assign n1767 = ~n1458 & ~n1766 ;
  assign n1768 = n1462 & n1767 ;
  assign n1769 = n1429 & n1444 ;
  assign n1770 = n1452 & ~n1769 ;
  assign n1771 = ~\InstAddrPointer_reg[10]/NET0131  & ~n1476 ;
  assign n1772 = ~n1295 & ~n1771 ;
  assign n1773 = \InstAddrPointer_reg[9]/NET0131  & n1436 ;
  assign n1774 = n1772 & n1773 ;
  assign n1775 = ~n1433 & n1774 ;
  assign n1776 = ~n1770 & n1775 ;
  assign n1777 = n1768 & n1776 ;
  assign n1778 = n1474 & n1777 ;
  assign n1779 = ~\InstAddrPointer_reg[26]/NET0131  & ~n1490 ;
  assign n1780 = ~n1493 & ~n1779 ;
  assign n1781 = n1366 & n1465 ;
  assign n1782 = n1498 & n1781 ;
  assign n1783 = n1780 & n1782 ;
  assign n1784 = n1778 & n1783 ;
  assign n1786 = ~n1495 & n1784 ;
  assign n1785 = n1495 & ~n1784 ;
  assign n1787 = n1014 & ~n1785 ;
  assign n1788 = ~n1786 & n1787 ;
  assign n1750 = n1339 & ~n1375 ;
  assign n1751 = ~n1053 & ~n1089 ;
  assign n1752 = n1676 & n1751 ;
  assign n1753 = ~n1678 & n1751 ;
  assign n1754 = n1672 & ~n1753 ;
  assign n1755 = ~n1752 & n1754 ;
  assign n1756 = ~n1015 & ~n1755 ;
  assign n1757 = n1323 & ~n1756 ;
  assign n1758 = n1359 & n1757 ;
  assign n1759 = n1750 & n1758 ;
  assign n1760 = n1373 & n1691 ;
  assign n1761 = n1759 & n1760 ;
  assign n1763 = n1388 & ~n1761 ;
  assign n1762 = ~n1388 & n1761 ;
  assign n1764 = ~n1014 & ~n1762 ;
  assign n1765 = ~n1763 & n1764 ;
  assign n1789 = ~n906 & ~n1765 ;
  assign n1790 = ~n1788 & n1789 ;
  assign n1791 = ~n1749 & ~n1790 ;
  assign n1792 = n773 & ~n1791 ;
  assign n1793 = ~\InstAddrPointer_reg[11]/NET0131  & ~n1530 ;
  assign n1794 = ~n1590 & ~n1793 ;
  assign n1795 = n1599 & n1794 ;
  assign n1796 = n1713 & n1795 ;
  assign n1797 = n1327 & n1531 ;
  assign n1800 = ~n1588 & ~n1797 ;
  assign n1798 = ~\InstAddrPointer_reg[16]/NET0131  & ~n1797 ;
  assign n1799 = ~n1532 & ~n1798 ;
  assign n1801 = n1325 & n1799 ;
  assign n1802 = n1800 & n1801 ;
  assign n1803 = n1796 & n1802 ;
  assign n1804 = n1613 & n1620 ;
  assign n1805 = n1803 & n1804 ;
  assign n1806 = ~\InstAddrPointer_reg[23]/NET0131  & ~n1539 ;
  assign n1807 = ~n1535 & ~n1806 ;
  assign n1808 = \InstAddrPointer_reg[24]/NET0131  & n1807 ;
  assign n1809 = n1721 & n1808 ;
  assign n1810 = n1805 & n1809 ;
  assign n1812 = ~n1627 & ~n1810 ;
  assign n1811 = n1627 & n1810 ;
  assign n1813 = n899 & ~n1811 ;
  assign n1814 = ~n1812 & n1813 ;
  assign n1815 = n863 & ~n911 ;
  assign n1816 = ~n814 & n1815 ;
  assign n1817 = \InstAddrPointer_reg[27]/NET0131  & ~n1816 ;
  assign n1819 = ~n873 & n1495 ;
  assign n1818 = n766 & n1627 ;
  assign n1820 = ~n811 & n1388 ;
  assign n1821 = ~n1818 & ~n1820 ;
  assign n1822 = ~n1819 & n1821 ;
  assign n1823 = ~n1817 & n1822 ;
  assign n1824 = ~n1814 & n1823 ;
  assign n1825 = ~n1792 & n1824 ;
  assign n1826 = n929 & ~n1825 ;
  assign n1827 = \rEIP_reg[27]/NET0131  & n1655 ;
  assign n1828 = \InstAddrPointer_reg[27]/NET0131  & n1661 ;
  assign n1829 = ~n1827 & ~n1828 ;
  assign n1830 = ~n1826 & n1829 ;
  assign n1831 = \PhyAddrPointer_reg[31]/NET0131  & n906 ;
  assign n1839 = n1396 & ~n1403 ;
  assign n1840 = n1761 & n1839 ;
  assign n1841 = ~\InstAddrPointer_reg[31]/NET0131  & ~n1402 ;
  assign n1842 = \InstAddrPointer_reg[31]/NET0131  & n1402 ;
  assign n1843 = ~n1841 & ~n1842 ;
  assign n1845 = ~n1840 & n1843 ;
  assign n1844 = n1840 & ~n1843 ;
  assign n1846 = ~n1014 & ~n1844 ;
  assign n1847 = ~n1845 & n1846 ;
  assign n1832 = ~\InstAddrPointer_reg[31]/NET0131  & ~n1514 ;
  assign n1833 = \InstAddrPointer_reg[31]/NET0131  & n1514 ;
  assign n1834 = ~n1832 & ~n1833 ;
  assign n1836 = ~n1512 & n1834 ;
  assign n1835 = n1512 & ~n1834 ;
  assign n1837 = n1014 & ~n1835 ;
  assign n1838 = ~n1836 & n1837 ;
  assign n1848 = ~n906 & ~n1838 ;
  assign n1849 = ~n1847 & n1848 ;
  assign n1850 = ~n1831 & ~n1849 ;
  assign n1851 = n773 & ~n1850 ;
  assign n1852 = ~n774 & ~n911 ;
  assign n1853 = \PhyAddrPointer_reg[31]/NET0131  & ~n1852 ;
  assign n1854 = n1637 & n1809 ;
  assign n1855 = n1805 & n1854 ;
  assign n1856 = ~\InstAddrPointer_reg[31]/NET0131  & ~n1634 ;
  assign n1857 = \InstAddrPointer_reg[31]/NET0131  & n1634 ;
  assign n1858 = ~n1856 & ~n1857 ;
  assign n1860 = n1855 & n1858 ;
  assign n1859 = ~n1855 & ~n1858 ;
  assign n1861 = n899 & ~n1859 ;
  assign n1862 = ~n1860 & n1861 ;
  assign n1863 = ~n1853 & ~n1862 ;
  assign n1864 = ~n1851 & n1863 ;
  assign n1865 = n929 & ~n1864 ;
  assign n1868 = \PhyAddrPointer_reg[22]/NET0131  & \PhyAddrPointer_reg[23]/NET0131  ;
  assign n1869 = \PhyAddrPointer_reg[24]/NET0131  & n1868 ;
  assign n1870 = \PhyAddrPointer_reg[2]/NET0131  & \PhyAddrPointer_reg[3]/NET0131  ;
  assign n1871 = \PhyAddrPointer_reg[4]/NET0131  & n1870 ;
  assign n1872 = \PhyAddrPointer_reg[5]/NET0131  & n1871 ;
  assign n1873 = \PhyAddrPointer_reg[6]/NET0131  & n1872 ;
  assign n1874 = \PhyAddrPointer_reg[7]/NET0131  & n1873 ;
  assign n1875 = \PhyAddrPointer_reg[8]/NET0131  & n1874 ;
  assign n1876 = \PhyAddrPointer_reg[9]/NET0131  & n1875 ;
  assign n1877 = \PhyAddrPointer_reg[10]/NET0131  & n1876 ;
  assign n1878 = \PhyAddrPointer_reg[11]/NET0131  & \PhyAddrPointer_reg[12]/NET0131  ;
  assign n1879 = \PhyAddrPointer_reg[13]/NET0131  & n1878 ;
  assign n1880 = n1877 & n1879 ;
  assign n1881 = \PhyAddrPointer_reg[14]/NET0131  & n1880 ;
  assign n1882 = \PhyAddrPointer_reg[15]/NET0131  & \PhyAddrPointer_reg[16]/NET0131  ;
  assign n1883 = \PhyAddrPointer_reg[17]/NET0131  & n1882 ;
  assign n1884 = n1881 & n1883 ;
  assign n1885 = \PhyAddrPointer_reg[18]/NET0131  & \PhyAddrPointer_reg[19]/NET0131  ;
  assign n1886 = \PhyAddrPointer_reg[20]/NET0131  & \PhyAddrPointer_reg[21]/NET0131  ;
  assign n1887 = n1885 & n1886 ;
  assign n1888 = n1884 & n1887 ;
  assign n1889 = n1869 & n1888 ;
  assign n1890 = \PhyAddrPointer_reg[25]/NET0131  & n1889 ;
  assign n1891 = \PhyAddrPointer_reg[26]/NET0131  & n1890 ;
  assign n1892 = \PhyAddrPointer_reg[27]/NET0131  & n1891 ;
  assign n1904 = \PhyAddrPointer_reg[28]/NET0131  & n1892 ;
  assign n1905 = \PhyAddrPointer_reg[29]/NET0131  & n1904 ;
  assign n1906 = ~\DataWidth_reg[1]/NET0131  & ~\PhyAddrPointer_reg[1]/NET0131  ;
  assign n1907 = n1905 & ~n1906 ;
  assign n1908 = \PhyAddrPointer_reg[30]/NET0131  & n1907 ;
  assign n1910 = \PhyAddrPointer_reg[31]/NET0131  & n1908 ;
  assign n1909 = ~\PhyAddrPointer_reg[31]/NET0131  & ~n1908 ;
  assign n1911 = n933 & ~n1909 ;
  assign n1912 = ~n1910 & n1911 ;
  assign n1867 = ~\State2_reg[1]/NET0131  & n940 ;
  assign n1893 = \PhyAddrPointer_reg[1]/NET0131  & n1892 ;
  assign n1894 = \PhyAddrPointer_reg[28]/NET0131  & n1893 ;
  assign n1895 = \PhyAddrPointer_reg[29]/NET0131  & n1894 ;
  assign n1896 = \PhyAddrPointer_reg[30]/NET0131  & n1895 ;
  assign n1897 = \PhyAddrPointer_reg[31]/NET0131  & ~n1896 ;
  assign n1898 = ~\PhyAddrPointer_reg[31]/NET0131  & n1896 ;
  assign n1899 = ~n1897 & ~n1898 ;
  assign n1900 = n1867 & ~n1899 ;
  assign n1866 = \rEIP_reg[31]/NET0131  & n1655 ;
  assign n1901 = ~n952 & ~n955 ;
  assign n1902 = ~n939 & n1901 ;
  assign n1903 = \PhyAddrPointer_reg[31]/NET0131  & ~n1902 ;
  assign n1913 = ~n1866 & ~n1903 ;
  assign n1914 = ~n1900 & n1913 ;
  assign n1915 = ~n1912 & n1914 ;
  assign n1916 = ~n1865 & n1915 ;
  assign n1920 = \InstAddrPointer_reg[15]/NET0131  & n906 ;
  assign n1925 = ~n1471 & ~n1777 ;
  assign n1926 = n1471 & n1777 ;
  assign n1927 = ~n1925 & ~n1926 ;
  assign n1928 = n1014 & ~n1927 ;
  assign n1921 = ~n1342 & ~n1757 ;
  assign n1922 = n1342 & n1757 ;
  assign n1923 = ~n1921 & ~n1922 ;
  assign n1924 = ~n1014 & ~n1923 ;
  assign n1929 = ~n906 & ~n1924 ;
  assign n1930 = ~n1928 & n1929 ;
  assign n1931 = ~n1920 & ~n1930 ;
  assign n1932 = n773 & ~n1931 ;
  assign n1934 = ~n1796 & ~n1800 ;
  assign n1933 = n1601 & n1713 ;
  assign n1935 = n899 & ~n1933 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1919 = \InstAddrPointer_reg[15]/NET0131  & ~n1816 ;
  assign n1937 = ~n873 & n1471 ;
  assign n1938 = n766 & n1800 ;
  assign n1939 = ~n811 & n1342 ;
  assign n1940 = ~n1938 & ~n1939 ;
  assign n1941 = ~n1937 & n1940 ;
  assign n1942 = ~n1919 & n1941 ;
  assign n1943 = ~n1936 & n1942 ;
  assign n1944 = ~n1932 & n1943 ;
  assign n1945 = n929 & ~n1944 ;
  assign n1917 = \InstAddrPointer_reg[15]/NET0131  & n1661 ;
  assign n1918 = \rEIP_reg[15]/NET0131  & n1655 ;
  assign n1946 = ~n1917 & ~n1918 ;
  assign n1947 = ~n1945 & n1946 ;
  assign n1965 = \InstAddrPointer_reg[22]/NET0131  & n906 ;
  assign n1950 = ~\InstAddrPointer_reg[22]/NET0131  & ~n1483 ;
  assign n1951 = ~n1492 & ~n1950 ;
  assign n1970 = n1482 & n1485 ;
  assign n1971 = ~n1951 & ~n1970 ;
  assign n1972 = ~n1487 & ~n1971 ;
  assign n1973 = n1014 & ~n1972 ;
  assign n1967 = n1361 & ~n1375 ;
  assign n1966 = ~n1361 & n1375 ;
  assign n1968 = ~n1014 & ~n1966 ;
  assign n1969 = ~n1967 & n1968 ;
  assign n1974 = ~n906 & ~n1969 ;
  assign n1975 = ~n1973 & n1974 ;
  assign n1976 = ~n1965 & ~n1975 ;
  assign n1977 = n773 & ~n1976 ;
  assign n1962 = ~\InstAddrPointer_reg[22]/NET0131  & ~n1610 ;
  assign n1963 = ~n1539 & ~n1962 ;
  assign n1978 = n1609 & n1620 ;
  assign n1980 = n1612 & n1978 ;
  assign n1981 = ~n1963 & ~n1980 ;
  assign n1979 = n1613 & n1978 ;
  assign n1982 = n899 & ~n1979 ;
  assign n1983 = ~n1981 & n1982 ;
  assign n1953 = ~READY_n_pad & ~n1951 ;
  assign n1954 = ~\InstAddrPointer_reg[22]/NET0131  & READY_n_pad ;
  assign n1955 = ~n1953 & ~n1954 ;
  assign n1956 = n840 & n1955 ;
  assign n1957 = ~n862 & n912 ;
  assign n1958 = ~n1956 & n1957 ;
  assign n1959 = \InstAddrPointer_reg[22]/NET0131  & ~n1958 ;
  assign n1952 = n788 & n1951 ;
  assign n1960 = ~n858 & n1955 ;
  assign n1984 = ~n1952 & ~n1960 ;
  assign n1961 = ~n811 & n1375 ;
  assign n1964 = n766 & n1963 ;
  assign n1985 = ~n1961 & ~n1964 ;
  assign n1986 = n1984 & n1985 ;
  assign n1987 = ~n1959 & n1986 ;
  assign n1988 = ~n1983 & n1987 ;
  assign n1989 = ~n1977 & n1988 ;
  assign n1990 = n929 & ~n1989 ;
  assign n1948 = \rEIP_reg[22]/NET0131  & n1655 ;
  assign n1949 = \InstAddrPointer_reg[22]/NET0131  & n1661 ;
  assign n1991 = ~n1948 & ~n1949 ;
  assign n1992 = ~n1990 & n1991 ;
  assign n2035 = n1583 & n1601 ;
  assign n2036 = n1799 & n2035 ;
  assign n2037 = n1716 & n2036 ;
  assign n2038 = n1614 & n2037 ;
  assign n2040 = n1616 & n2038 ;
  assign n2039 = ~n1616 & ~n2038 ;
  assign n2041 = n899 & ~n2039 ;
  assign n2042 = ~n2040 & n2041 ;
  assign n1999 = \InstAddrPointer_reg[24]/NET0131  & n906 ;
  assign n2022 = n1324 & ~n1342 ;
  assign n2023 = ~n1345 & n1358 ;
  assign n2024 = ~n1368 & n2023 ;
  assign n2025 = n1750 & n2024 ;
  assign n2026 = n2022 & n2025 ;
  assign n2028 = ~n1372 & n2026 ;
  assign n2027 = n1372 & ~n2026 ;
  assign n2029 = ~n1014 & ~n2027 ;
  assign n2030 = ~n2028 & n2029 ;
  assign n2000 = n1417 & ~n1422 ;
  assign n2001 = ~n1416 & n1418 ;
  assign n2002 = ~n1426 & ~n2001 ;
  assign n2003 = ~n2000 & n2002 ;
  assign n2004 = ~n1410 & ~n1443 ;
  assign n2005 = ~n2003 & n2004 ;
  assign n2006 = n1425 & ~n1443 ;
  assign n2007 = ~n1449 & ~n2006 ;
  assign n2008 = ~n2005 & n2007 ;
  assign n2009 = ~n1433 & ~n1440 ;
  assign n2010 = ~n2008 & n2009 ;
  assign n2011 = ~n1433 & n1448 ;
  assign n2012 = ~n1447 & ~n2011 ;
  assign n2013 = ~n2010 & n2012 ;
  assign n2014 = n1436 & n1480 ;
  assign n2015 = ~n2013 & n2014 ;
  assign n2016 = n1365 & n1456 ;
  assign n2017 = n2015 & n2016 ;
  assign n2019 = n1497 & ~n2017 ;
  assign n2018 = ~n1497 & n2017 ;
  assign n2020 = n1014 & ~n2018 ;
  assign n2021 = ~n2019 & n2020 ;
  assign n2031 = ~n906 & ~n2021 ;
  assign n2032 = ~n2030 & n2031 ;
  assign n2033 = ~n1999 & ~n2032 ;
  assign n2034 = n773 & ~n2033 ;
  assign n1998 = \InstAddrPointer_reg[24]/NET0131  & ~n1816 ;
  assign n1995 = ~n873 & n1497 ;
  assign n1996 = n766 & n1616 ;
  assign n1997 = ~n811 & n1372 ;
  assign n2043 = ~n1996 & ~n1997 ;
  assign n2044 = ~n1995 & n2043 ;
  assign n2045 = ~n1998 & n2044 ;
  assign n2046 = ~n2034 & n2045 ;
  assign n2047 = ~n2042 & n2046 ;
  assign n2048 = n929 & ~n2047 ;
  assign n1993 = \rEIP_reg[24]/NET0131  & n1655 ;
  assign n1994 = \InstAddrPointer_reg[24]/NET0131  & n1661 ;
  assign n2049 = ~n1993 & ~n1994 ;
  assign n2050 = ~n2048 & n2049 ;
  assign n2051 = \InstAddrPointer_reg[26]/NET0131  & n906 ;
  assign n2056 = n1774 & ~n2013 ;
  assign n2057 = n1768 & n2056 ;
  assign n2058 = n1474 & n2057 ;
  assign n2059 = n1782 & n2058 ;
  assign n2061 = ~n1780 & n2059 ;
  assign n2060 = n1780 & ~n2059 ;
  assign n2062 = n1014 & ~n2060 ;
  assign n2063 = ~n2061 & n2062 ;
  assign n2053 = n1382 & ~n1398 ;
  assign n2052 = ~n1382 & n1398 ;
  assign n2054 = ~n1014 & ~n2052 ;
  assign n2055 = ~n2053 & n2054 ;
  assign n2064 = ~n906 & ~n2055 ;
  assign n2065 = ~n2063 & n2064 ;
  assign n2066 = ~n2051 & ~n2065 ;
  assign n2067 = n773 & ~n2066 ;
  assign n2069 = ~n1541 & ~n1623 ;
  assign n2070 = n899 & ~n1624 ;
  assign n2071 = ~n2069 & n2070 ;
  assign n2077 = n766 & n1541 ;
  assign n2076 = ~n844 & n1780 ;
  assign n2068 = ~n811 & n1398 ;
  assign n2072 = ~n836 & n1780 ;
  assign n2073 = n850 & n912 ;
  assign n2074 = ~n2072 & n2073 ;
  assign n2075 = \InstAddrPointer_reg[26]/NET0131  & ~n2074 ;
  assign n2078 = ~n2068 & ~n2075 ;
  assign n2079 = ~n2076 & n2078 ;
  assign n2080 = ~n2077 & n2079 ;
  assign n2081 = ~n2071 & n2080 ;
  assign n2082 = ~n2067 & n2081 ;
  assign n2083 = n929 & ~n2082 ;
  assign n2084 = \rEIP_reg[26]/NET0131  & n1655 ;
  assign n2085 = \InstAddrPointer_reg[26]/NET0131  & n1661 ;
  assign n2086 = ~n2084 & ~n2085 ;
  assign n2087 = ~n2083 & n2086 ;
  assign n2088 = \PhyAddrPointer_reg[30]/NET0131  & n906 ;
  assign n2089 = ~n1522 & ~n2088 ;
  assign n2090 = n773 & ~n2089 ;
  assign n2091 = \PhyAddrPointer_reg[30]/NET0131  & ~n1852 ;
  assign n2092 = ~n1640 & ~n2091 ;
  assign n2093 = ~n2090 & n2092 ;
  assign n2094 = n929 & ~n2093 ;
  assign n2096 = ~\PhyAddrPointer_reg[30]/NET0131  & ~n1895 ;
  assign n2097 = ~n1896 & ~n2096 ;
  assign n2098 = ~n933 & ~n1867 ;
  assign n2099 = \DataWidth_reg[1]/NET0131  & ~n1867 ;
  assign n2100 = ~n2098 & ~n2099 ;
  assign n2101 = n2097 & n2100 ;
  assign n2103 = ~\PhyAddrPointer_reg[30]/NET0131  & ~n1905 ;
  assign n2102 = \PhyAddrPointer_reg[30]/NET0131  & n1905 ;
  assign n2104 = n969 & ~n2102 ;
  assign n2105 = ~n2103 & n2104 ;
  assign n2095 = \PhyAddrPointer_reg[30]/NET0131  & ~n1902 ;
  assign n2106 = ~n1656 & ~n2095 ;
  assign n2107 = ~n2105 & n2106 ;
  assign n2108 = ~n2101 & n2107 ;
  assign n2109 = ~n2094 & n2108 ;
  assign n2113 = \InstAddrPointer_reg[11]/NET0131  & n906 ;
  assign n2122 = ~n1767 & n1776 ;
  assign n2121 = n1767 & ~n1776 ;
  assign n2123 = n1014 & ~n2121 ;
  assign n2124 = ~n2122 & n2123 ;
  assign n2114 = n1290 & n1317 ;
  assign n2115 = ~n1285 & n2114 ;
  assign n2116 = ~n1319 & n2115 ;
  assign n2117 = n1755 & n2114 ;
  assign n2118 = n1319 & ~n2117 ;
  assign n2119 = ~n1014 & ~n2118 ;
  assign n2120 = ~n2116 & n2119 ;
  assign n2125 = ~n906 & ~n2120 ;
  assign n2126 = ~n2124 & n2125 ;
  assign n2127 = ~n2113 & ~n2126 ;
  assign n2128 = n773 & ~n2127 ;
  assign n2132 = n1597 & n1713 ;
  assign n2134 = ~n1794 & ~n2132 ;
  assign n2133 = \InstAddrPointer_reg[11]/NET0131  & n2132 ;
  assign n2135 = n899 & ~n2133 ;
  assign n2136 = ~n2134 & n2135 ;
  assign n2129 = ~n858 & ~n1295 ;
  assign n2130 = n1816 & ~n2129 ;
  assign n2131 = \InstAddrPointer_reg[11]/NET0131  & ~n2130 ;
  assign n2112 = ~n873 & n1767 ;
  assign n2137 = n766 & n1794 ;
  assign n2138 = ~n811 & n1319 ;
  assign n2139 = ~n2137 & ~n2138 ;
  assign n2140 = ~n2112 & n2139 ;
  assign n2141 = ~n2131 & n2140 ;
  assign n2142 = ~n2136 & n2141 ;
  assign n2143 = ~n2128 & n2142 ;
  assign n2144 = n929 & ~n2143 ;
  assign n2110 = \InstAddrPointer_reg[11]/NET0131  & n1661 ;
  assign n2111 = \rEIP_reg[11]/NET0131  & n1655 ;
  assign n2145 = ~n2110 & ~n2111 ;
  assign n2146 = ~n2144 & n2145 ;
  assign n2147 = \InstAddrPointer_reg[14]/NET0131  & n906 ;
  assign n2148 = ~\InstAddrPointer_reg[14]/NET0131  & ~n1298 ;
  assign n2149 = ~n1468 & ~n2148 ;
  assign n2150 = n1767 & n2056 ;
  assign n2151 = \InstAddrPointer_reg[12]/NET0131  & n2150 ;
  assign n2152 = \InstAddrPointer_reg[13]/NET0131  & n2151 ;
  assign n2153 = ~n2149 & ~n2152 ;
  assign n2154 = ~n2057 & ~n2153 ;
  assign n2155 = n1014 & ~n2154 ;
  assign n2156 = ~n1312 & n2116 ;
  assign n2157 = ~n1306 & n2156 ;
  assign n2158 = n1302 & ~n2157 ;
  assign n2159 = ~n1014 & ~n1324 ;
  assign n2160 = ~n2158 & n2159 ;
  assign n2161 = ~n906 & ~n2160 ;
  assign n2162 = ~n2155 & n2161 ;
  assign n2163 = ~n2147 & ~n2162 ;
  assign n2164 = n773 & ~n2163 ;
  assign n2167 = ~\InstAddrPointer_reg[14]/NET0131  & ~n1531 ;
  assign n2168 = ~n1587 & ~n2167 ;
  assign n2169 = n1583 & n1596 ;
  assign n2170 = \InstAddrPointer_reg[10]/NET0131  & n2169 ;
  assign n2171 = n1594 & n1794 ;
  assign n2172 = n2170 & n2171 ;
  assign n2173 = ~n2168 & ~n2172 ;
  assign n2166 = n1583 & n1795 ;
  assign n2174 = n899 & ~n2166 ;
  assign n2175 = ~n2173 & n2174 ;
  assign n2180 = \InstAddrPointer_reg[14]/NET0131  & ~n1815 ;
  assign n2165 = ~n873 & n2149 ;
  assign n2177 = n765 & ~n2168 ;
  assign n2176 = ~\InstAddrPointer_reg[14]/NET0131  & ~n765 ;
  assign n2178 = ~n740 & ~n2176 ;
  assign n2179 = ~n2177 & n2178 ;
  assign n2181 = ~n811 & n1302 ;
  assign n2182 = ~n2179 & ~n2181 ;
  assign n2183 = ~n2165 & n2182 ;
  assign n2184 = ~n2180 & n2183 ;
  assign n2185 = ~n2175 & n2184 ;
  assign n2186 = ~n2164 & n2185 ;
  assign n2187 = n929 & ~n2186 ;
  assign n2188 = \rEIP_reg[14]/NET0131  & n1655 ;
  assign n2189 = \InstAddrPointer_reg[14]/NET0131  & n1661 ;
  assign n2190 = ~n2188 & ~n2189 ;
  assign n2191 = ~n2187 & n2190 ;
  assign n2192 = \InstAddrPointer_reg[25]/NET0131  & n906 ;
  assign n2202 = ~n1380 & n1690 ;
  assign n2201 = n1380 & ~n1690 ;
  assign n2203 = ~n1014 & ~n2201 ;
  assign n2204 = ~n2202 & n2203 ;
  assign n2193 = \InstAddrPointer_reg[24]/NET0131  & n1502 ;
  assign n2194 = n1487 & n2193 ;
  assign n2196 = ~\InstAddrPointer_reg[25]/NET0131  & ~n1489 ;
  assign n2197 = ~n1490 & ~n2196 ;
  assign n2198 = ~n2194 & n2197 ;
  assign n2195 = ~\InstAddrPointer_reg[25]/NET0131  & n2194 ;
  assign n2199 = n1014 & ~n2195 ;
  assign n2200 = ~n2198 & n2199 ;
  assign n2205 = ~n906 & ~n2200 ;
  assign n2206 = ~n2204 & n2205 ;
  assign n2207 = ~n2192 & ~n2206 ;
  assign n2208 = n773 & ~n2207 ;
  assign n2211 = n1718 & n1720 ;
  assign n2210 = ~n1718 & ~n1720 ;
  assign n2212 = n899 & ~n2210 ;
  assign n2213 = ~n2211 & n2212 ;
  assign n2214 = n836 & ~n842 ;
  assign n2215 = READY_n_pad & ~n2214 ;
  assign n2216 = n1957 & ~n2215 ;
  assign n2217 = ~n836 & ~n1489 ;
  assign n2218 = n2216 & ~n2217 ;
  assign n2219 = \InstAddrPointer_reg[25]/NET0131  & ~n2218 ;
  assign n2221 = ~n873 & n2197 ;
  assign n2209 = n766 & n1720 ;
  assign n2220 = ~n811 & n1380 ;
  assign n2222 = ~n2209 & ~n2220 ;
  assign n2223 = ~n2221 & n2222 ;
  assign n2224 = ~n2219 & n2223 ;
  assign n2225 = ~n2213 & n2224 ;
  assign n2226 = ~n2208 & n2225 ;
  assign n2227 = n929 & ~n2226 ;
  assign n2228 = \rEIP_reg[25]/NET0131  & n1655 ;
  assign n2229 = \InstAddrPointer_reg[25]/NET0131  & n1661 ;
  assign n2230 = ~n2228 & ~n2229 ;
  assign n2231 = ~n2227 & n2230 ;
  assign n2242 = \PhyAddrPointer_reg[15]/NET0131  & n906 ;
  assign n2243 = ~n1930 & ~n2242 ;
  assign n2244 = n773 & ~n2243 ;
  assign n2245 = \PhyAddrPointer_reg[15]/NET0131  & ~n1852 ;
  assign n2246 = ~n1936 & ~n2245 ;
  assign n2247 = ~n2244 & n2246 ;
  assign n2248 = n929 & ~n2247 ;
  assign n2251 = n1881 & ~n1906 ;
  assign n2252 = ~\PhyAddrPointer_reg[15]/NET0131  & ~n2251 ;
  assign n2249 = \PhyAddrPointer_reg[15]/NET0131  & n1881 ;
  assign n2250 = ~n1906 & n2249 ;
  assign n2253 = n933 & ~n2250 ;
  assign n2254 = ~n2252 & n2253 ;
  assign n2232 = \PhyAddrPointer_reg[1]/NET0131  & n1874 ;
  assign n2233 = \PhyAddrPointer_reg[8]/NET0131  & n2232 ;
  assign n2234 = \PhyAddrPointer_reg[9]/NET0131  & n2233 ;
  assign n2235 = \PhyAddrPointer_reg[10]/NET0131  & n2234 ;
  assign n2236 = n1879 & n2235 ;
  assign n2237 = \PhyAddrPointer_reg[14]/NET0131  & n2236 ;
  assign n2238 = ~\PhyAddrPointer_reg[15]/NET0131  & ~n2237 ;
  assign n2239 = \PhyAddrPointer_reg[15]/NET0131  & n2237 ;
  assign n2240 = ~n2238 & ~n2239 ;
  assign n2241 = n1867 & n2240 ;
  assign n2255 = \PhyAddrPointer_reg[15]/NET0131  & ~n1902 ;
  assign n2256 = ~n1918 & ~n2255 ;
  assign n2257 = ~n2241 & n2256 ;
  assign n2258 = ~n2254 & n2257 ;
  assign n2259 = ~n2248 & n2258 ;
  assign n2274 = \PhyAddrPointer_reg[23]/NET0131  & n906 ;
  assign n2279 = ~n1487 & ~n1502 ;
  assign n2280 = ~n2017 & ~n2279 ;
  assign n2281 = n1014 & ~n2280 ;
  assign n2275 = ~n1368 & ~n1759 ;
  assign n2276 = n1368 & n1759 ;
  assign n2277 = ~n2275 & ~n2276 ;
  assign n2278 = ~n1014 & ~n2277 ;
  assign n2282 = ~n906 & ~n2278 ;
  assign n2283 = ~n2281 & n2282 ;
  assign n2284 = ~n2274 & ~n2283 ;
  assign n2285 = n773 & ~n2284 ;
  assign n2286 = \PhyAddrPointer_reg[23]/NET0131  & ~n1852 ;
  assign n2287 = ~n1805 & ~n1807 ;
  assign n2288 = n899 & ~n2038 ;
  assign n2289 = ~n2287 & n2288 ;
  assign n2290 = ~n2286 & ~n2289 ;
  assign n2291 = ~n2285 & n2290 ;
  assign n2292 = n929 & ~n2291 ;
  assign n2265 = \PhyAddrPointer_reg[1]/NET0131  & n1884 ;
  assign n2266 = n1887 & n2265 ;
  assign n2267 = \PhyAddrPointer_reg[22]/NET0131  & n2266 ;
  assign n2268 = ~\PhyAddrPointer_reg[23]/NET0131  & ~n2267 ;
  assign n2269 = n1868 & n2266 ;
  assign n2270 = ~n2268 & ~n2269 ;
  assign n2271 = n2100 & n2270 ;
  assign n2260 = \PhyAddrPointer_reg[22]/NET0131  & n1888 ;
  assign n2262 = \PhyAddrPointer_reg[23]/NET0131  & n2260 ;
  assign n2261 = ~\PhyAddrPointer_reg[23]/NET0131  & ~n2260 ;
  assign n2263 = n969 & ~n2261 ;
  assign n2264 = ~n2262 & n2263 ;
  assign n2272 = \rEIP_reg[23]/NET0131  & n1655 ;
  assign n2273 = \PhyAddrPointer_reg[23]/NET0131  & ~n1902 ;
  assign n2293 = ~n2272 & ~n2273 ;
  assign n2294 = ~n2264 & n2293 ;
  assign n2295 = ~n2271 & n2294 ;
  assign n2296 = ~n2292 & n2295 ;
  assign n2297 = \PhyAddrPointer_reg[27]/NET0131  & n906 ;
  assign n2298 = ~n1790 & ~n2297 ;
  assign n2299 = n773 & ~n2298 ;
  assign n2300 = \PhyAddrPointer_reg[27]/NET0131  & ~n1852 ;
  assign n2301 = ~n1814 & ~n2300 ;
  assign n2302 = ~n2299 & n2301 ;
  assign n2303 = n929 & ~n2302 ;
  assign n2304 = \PhyAddrPointer_reg[1]/NET0131  & n1891 ;
  assign n2305 = ~\PhyAddrPointer_reg[27]/NET0131  & ~n2304 ;
  assign n2306 = ~n1893 & ~n2305 ;
  assign n2311 = ~\DataWidth_reg[1]/NET0131  & ~n2306 ;
  assign n2308 = ~\PhyAddrPointer_reg[27]/NET0131  & ~n1891 ;
  assign n2309 = ~n1892 & ~n2308 ;
  assign n2310 = \DataWidth_reg[1]/NET0131  & ~n2309 ;
  assign n2312 = n933 & ~n2310 ;
  assign n2313 = ~n2311 & n2312 ;
  assign n2307 = n1867 & n2306 ;
  assign n2314 = \PhyAddrPointer_reg[27]/NET0131  & ~n1902 ;
  assign n2315 = ~n1827 & ~n2314 ;
  assign n2316 = ~n2307 & n2315 ;
  assign n2317 = ~n2313 & n2316 ;
  assign n2318 = ~n2303 & n2317 ;
  assign n2319 = \PhyAddrPointer_reg[28]/NET0131  & n906 ;
  assign n2327 = ~n1372 & ~n1388 ;
  assign n2328 = n1691 & n2327 ;
  assign n2329 = n2026 & n2328 ;
  assign n2331 = ~n1391 & n2329 ;
  assign n2330 = n1391 & ~n2329 ;
  assign n2332 = ~n1014 & ~n2330 ;
  assign n2333 = ~n2331 & n2332 ;
  assign n2320 = n1500 & n2017 ;
  assign n2321 = ~\InstAddrPointer_reg[28]/NET0131  & ~n1491 ;
  assign n2322 = ~n1506 & ~n2321 ;
  assign n2324 = n2320 & ~n2322 ;
  assign n2323 = ~n2320 & n2322 ;
  assign n2325 = n1014 & ~n2323 ;
  assign n2326 = ~n2324 & n2325 ;
  assign n2334 = ~n906 & ~n2326 ;
  assign n2335 = ~n2333 & n2334 ;
  assign n2336 = ~n2319 & ~n2335 ;
  assign n2337 = n773 & ~n2336 ;
  assign n2338 = \PhyAddrPointer_reg[28]/NET0131  & ~n1852 ;
  assign n2339 = ~\InstAddrPointer_reg[28]/NET0131  & ~n1626 ;
  assign n2340 = ~n1631 & ~n2339 ;
  assign n2341 = n1326 & n2036 ;
  assign n2342 = ~\InstAddrPointer_reg[20]/NET0131  & ~n1533 ;
  assign n2343 = ~n1534 & ~n2342 ;
  assign n2344 = \InstAddrPointer_reg[25]/NET0131  & n1386 ;
  assign n2345 = n2343 & n2344 ;
  assign n2346 = n1617 & n2345 ;
  assign n2347 = n2341 & n2346 ;
  assign n2349 = n2340 & n2347 ;
  assign n2348 = ~n2340 & ~n2347 ;
  assign n2350 = n899 & ~n2348 ;
  assign n2351 = ~n2349 & n2350 ;
  assign n2352 = ~n2338 & ~n2351 ;
  assign n2353 = ~n2337 & n2352 ;
  assign n2354 = n929 & ~n2353 ;
  assign n2358 = ~\PhyAddrPointer_reg[28]/NET0131  & ~n1893 ;
  assign n2359 = ~n1894 & ~n2358 ;
  assign n2360 = n2100 & n2359 ;
  assign n2355 = ~\PhyAddrPointer_reg[28]/NET0131  & ~n1892 ;
  assign n2356 = n969 & ~n1904 ;
  assign n2357 = ~n2355 & n2356 ;
  assign n2361 = \rEIP_reg[28]/NET0131  & n1655 ;
  assign n2362 = \PhyAddrPointer_reg[28]/NET0131  & ~n1902 ;
  assign n2363 = ~n2361 & ~n2362 ;
  assign n2364 = ~n2357 & n2363 ;
  assign n2365 = ~n2360 & n2364 ;
  assign n2366 = ~n2354 & n2365 ;
  assign n2367 = \PhyAddrPointer_reg[29]/NET0131  & n906 ;
  assign n2368 = ~n1699 & ~n2367 ;
  assign n2369 = n773 & ~n2368 ;
  assign n2370 = \PhyAddrPointer_reg[29]/NET0131  & ~n1852 ;
  assign n2371 = ~n1727 & ~n2370 ;
  assign n2372 = ~n2369 & n2371 ;
  assign n2373 = n929 & ~n2372 ;
  assign n2378 = ~\PhyAddrPointer_reg[29]/NET0131  & ~n1894 ;
  assign n2379 = ~n1895 & ~n2378 ;
  assign n2380 = n1867 & n2379 ;
  assign n2374 = n1904 & ~n1906 ;
  assign n2375 = ~\PhyAddrPointer_reg[29]/NET0131  & ~n2374 ;
  assign n2376 = n933 & ~n1907 ;
  assign n2377 = ~n2375 & n2376 ;
  assign n2381 = \PhyAddrPointer_reg[29]/NET0131  & ~n1902 ;
  assign n2382 = ~n1745 & ~n2381 ;
  assign n2383 = ~n2377 & n2382 ;
  assign n2384 = ~n2380 & n2383 ;
  assign n2385 = ~n2373 & n2384 ;
  assign n2392 = \InstAddrPointer_reg[8]/NET0131  & n906 ;
  assign n2397 = ~n1285 & ~n1289 ;
  assign n2399 = ~n1288 & n2397 ;
  assign n2398 = n1288 & ~n2397 ;
  assign n2400 = ~n1014 & ~n2398 ;
  assign n2401 = ~n2399 & n2400 ;
  assign n2394 = n1436 & n2013 ;
  assign n2393 = ~n1436 & ~n2013 ;
  assign n2395 = n1014 & ~n2393 ;
  assign n2396 = ~n2394 & n2395 ;
  assign n2402 = ~n906 & ~n2396 ;
  assign n2403 = ~n2401 & n2402 ;
  assign n2404 = ~n2392 & ~n2403 ;
  assign n2405 = n773 & ~n2404 ;
  assign n2406 = ~n1544 & ~n1582 ;
  assign n2407 = ~n1547 & ~n2406 ;
  assign n2408 = n899 & ~n1583 ;
  assign n2409 = ~n2407 & n2408 ;
  assign n2388 = \InstAddrPointer_reg[8]/NET0131  & ~n1816 ;
  assign n2390 = ~n873 & n1436 ;
  assign n2389 = ~n811 & n1288 ;
  assign n2391 = n766 & n1547 ;
  assign n2410 = ~n2389 & ~n2391 ;
  assign n2411 = ~n2390 & n2410 ;
  assign n2412 = ~n2388 & n2411 ;
  assign n2413 = ~n2409 & n2412 ;
  assign n2414 = ~n2405 & n2413 ;
  assign n2415 = n929 & ~n2414 ;
  assign n2386 = \rEIP_reg[8]/NET0131  & n1655 ;
  assign n2387 = \InstAddrPointer_reg[8]/NET0131  & n1661 ;
  assign n2416 = ~n2386 & ~n2387 ;
  assign n2417 = ~n2415 & n2416 ;
  assign n2418 = \InstAddrPointer_reg[13]/NET0131  & n906 ;
  assign n2422 = ~\InstAddrPointer_reg[13]/NET0131  & ~n1303 ;
  assign n2423 = ~n1298 & ~n2422 ;
  assign n2424 = ~n1454 & n1477 ;
  assign n2425 = n1296 & n1772 ;
  assign n2426 = n2424 & n2425 ;
  assign n2427 = ~n2423 & ~n2426 ;
  assign n2428 = n2423 & n2426 ;
  assign n2429 = ~n2427 & ~n2428 ;
  assign n2430 = n1014 & ~n2429 ;
  assign n2419 = n1306 & ~n1684 ;
  assign n2420 = ~n1014 & ~n2419 ;
  assign n2421 = ~n2157 & n2420 ;
  assign n2431 = ~n906 & ~n2421 ;
  assign n2432 = ~n2430 & n2431 ;
  assign n2433 = ~n2418 & ~n2432 ;
  assign n2434 = n773 & ~n2433 ;
  assign n2436 = \InstAddrPointer_reg[12]/NET0131  & n2133 ;
  assign n2438 = ~\InstAddrPointer_reg[13]/NET0131  & ~n1592 ;
  assign n2439 = ~n1531 & ~n2438 ;
  assign n2440 = ~n2436 & ~n2439 ;
  assign n2437 = \InstAddrPointer_reg[13]/NET0131  & n2436 ;
  assign n2441 = n899 & ~n2437 ;
  assign n2442 = ~n2440 & n2441 ;
  assign n2444 = \InstAddrPointer_reg[13]/NET0131  & ~n836 ;
  assign n2445 = n873 & ~n2444 ;
  assign n2446 = n2423 & ~n2445 ;
  assign n2443 = \InstAddrPointer_reg[13]/NET0131  & ~n2216 ;
  assign n2435 = ~n811 & n1306 ;
  assign n2447 = n766 & n2439 ;
  assign n2448 = ~n2435 & ~n2447 ;
  assign n2449 = ~n2443 & n2448 ;
  assign n2450 = ~n2446 & n2449 ;
  assign n2451 = ~n2442 & n2450 ;
  assign n2452 = ~n2434 & n2451 ;
  assign n2453 = n929 & ~n2452 ;
  assign n2454 = \rEIP_reg[13]/NET0131  & n1655 ;
  assign n2455 = \InstAddrPointer_reg[13]/NET0131  & n1661 ;
  assign n2456 = ~n2454 & ~n2455 ;
  assign n2457 = ~n2453 & n2456 ;
  assign n2458 = \PhyAddrPointer_reg[11]/NET0131  & n906 ;
  assign n2459 = ~n2126 & ~n2458 ;
  assign n2460 = n773 & ~n2459 ;
  assign n2461 = \PhyAddrPointer_reg[11]/NET0131  & ~n1852 ;
  assign n2462 = ~n2136 & ~n2461 ;
  assign n2463 = ~n2460 & n2462 ;
  assign n2464 = n929 & ~n2463 ;
  assign n2469 = ~\PhyAddrPointer_reg[11]/NET0131  & ~n2235 ;
  assign n2465 = \PhyAddrPointer_reg[11]/NET0131  & n1877 ;
  assign n2470 = \PhyAddrPointer_reg[1]/NET0131  & n2465 ;
  assign n2471 = ~n2469 & ~n2470 ;
  assign n2472 = n2100 & n2471 ;
  assign n2466 = ~\PhyAddrPointer_reg[11]/NET0131  & ~n1877 ;
  assign n2467 = n969 & ~n2465 ;
  assign n2468 = ~n2466 & n2467 ;
  assign n2473 = \PhyAddrPointer_reg[11]/NET0131  & ~n1902 ;
  assign n2474 = ~n2111 & ~n2473 ;
  assign n2475 = ~n2468 & n2474 ;
  assign n2476 = ~n2472 & n2475 ;
  assign n2477 = ~n2464 & n2476 ;
  assign n2478 = \PhyAddrPointer_reg[14]/NET0131  & n906 ;
  assign n2479 = ~n2162 & ~n2478 ;
  assign n2480 = n773 & ~n2479 ;
  assign n2481 = \PhyAddrPointer_reg[14]/NET0131  & ~n1852 ;
  assign n2482 = ~n2175 & ~n2481 ;
  assign n2483 = ~n2480 & n2482 ;
  assign n2484 = n929 & ~n2483 ;
  assign n2485 = ~\PhyAddrPointer_reg[14]/NET0131  & ~n2236 ;
  assign n2486 = ~n2237 & ~n2485 ;
  assign n2491 = ~\DataWidth_reg[1]/NET0131  & ~n2486 ;
  assign n2488 = ~\PhyAddrPointer_reg[14]/NET0131  & ~n1880 ;
  assign n2489 = ~n1881 & ~n2488 ;
  assign n2490 = \DataWidth_reg[1]/NET0131  & ~n2489 ;
  assign n2492 = n933 & ~n2490 ;
  assign n2493 = ~n2491 & n2492 ;
  assign n2487 = n1867 & n2486 ;
  assign n2494 = \PhyAddrPointer_reg[14]/NET0131  & ~n1902 ;
  assign n2495 = ~n2188 & ~n2494 ;
  assign n2496 = ~n2487 & n2495 ;
  assign n2497 = ~n2493 & n2496 ;
  assign n2498 = ~n2484 & n2497 ;
  assign n2512 = \PhyAddrPointer_reg[19]/NET0131  & n906 ;
  assign n2518 = ~n1465 & ~n1778 ;
  assign n2519 = ~n2015 & ~n2518 ;
  assign n2520 = n1014 & ~n2519 ;
  assign n2513 = n1346 & n1357 ;
  assign n2514 = n1757 & n2513 ;
  assign n2515 = n1351 & ~n2514 ;
  assign n2516 = ~n1014 & ~n1758 ;
  assign n2517 = ~n2515 & n2516 ;
  assign n2521 = ~n906 & ~n2517 ;
  assign n2522 = ~n2520 & n2521 ;
  assign n2523 = ~n2512 & ~n2522 ;
  assign n2524 = n773 & ~n2523 ;
  assign n2525 = \PhyAddrPointer_reg[19]/NET0131  & ~n1852 ;
  assign n2527 = n1619 & n1803 ;
  assign n2526 = ~n1619 & ~n1803 ;
  assign n2528 = n899 & ~n2526 ;
  assign n2529 = ~n2527 & n2528 ;
  assign n2530 = ~n2525 & ~n2529 ;
  assign n2531 = ~n2524 & n2530 ;
  assign n2532 = n929 & ~n2531 ;
  assign n2499 = \PhyAddrPointer_reg[18]/NET0131  & n1884 ;
  assign n2506 = \PhyAddrPointer_reg[1]/NET0131  & n2499 ;
  assign n2507 = ~\PhyAddrPointer_reg[19]/NET0131  & ~n2506 ;
  assign n2508 = n1884 & n1885 ;
  assign n2509 = \PhyAddrPointer_reg[1]/NET0131  & n2508 ;
  assign n2510 = ~n2507 & ~n2509 ;
  assign n2511 = n2100 & n2510 ;
  assign n2500 = n969 & ~n2499 ;
  assign n2501 = n1902 & ~n2500 ;
  assign n2502 = \PhyAddrPointer_reg[19]/NET0131  & ~n2501 ;
  assign n2503 = ~\PhyAddrPointer_reg[19]/NET0131  & n969 ;
  assign n2504 = n2499 & n2503 ;
  assign n2505 = \rEIP_reg[19]/NET0131  & n1655 ;
  assign n2533 = ~n2504 & ~n2505 ;
  assign n2534 = ~n2502 & n2533 ;
  assign n2535 = ~n2511 & n2534 ;
  assign n2536 = ~n2532 & n2535 ;
  assign n2537 = \PhyAddrPointer_reg[22]/NET0131  & n906 ;
  assign n2538 = ~n1975 & ~n2537 ;
  assign n2539 = n773 & ~n2538 ;
  assign n2540 = \PhyAddrPointer_reg[22]/NET0131  & ~n1852 ;
  assign n2541 = ~n1983 & ~n2540 ;
  assign n2542 = ~n2539 & n2541 ;
  assign n2543 = n929 & ~n2542 ;
  assign n2544 = ~\PhyAddrPointer_reg[22]/NET0131  & ~n2266 ;
  assign n2545 = ~n2267 & ~n2544 ;
  assign n2550 = ~\DataWidth_reg[1]/NET0131  & ~n2545 ;
  assign n2547 = ~\PhyAddrPointer_reg[22]/NET0131  & ~n1888 ;
  assign n2548 = ~n2260 & ~n2547 ;
  assign n2549 = \DataWidth_reg[1]/NET0131  & ~n2548 ;
  assign n2551 = n933 & ~n2549 ;
  assign n2552 = ~n2550 & n2551 ;
  assign n2546 = n1867 & n2545 ;
  assign n2553 = \PhyAddrPointer_reg[22]/NET0131  & ~n1902 ;
  assign n2554 = ~n1948 & ~n2553 ;
  assign n2555 = ~n2546 & n2554 ;
  assign n2556 = ~n2552 & n2555 ;
  assign n2557 = ~n2543 & n2556 ;
  assign n2558 = \PhyAddrPointer_reg[24]/NET0131  & n906 ;
  assign n2559 = ~n2032 & ~n2558 ;
  assign n2560 = n773 & ~n2559 ;
  assign n2561 = \PhyAddrPointer_reg[24]/NET0131  & ~n1852 ;
  assign n2562 = ~n2042 & ~n2561 ;
  assign n2563 = ~n2560 & n2562 ;
  assign n2564 = n929 & ~n2563 ;
  assign n2568 = ~\PhyAddrPointer_reg[24]/NET0131  & ~n2269 ;
  assign n2569 = n1869 & n2266 ;
  assign n2570 = ~n2568 & ~n2569 ;
  assign n2571 = n2100 & n2570 ;
  assign n2565 = ~\PhyAddrPointer_reg[24]/NET0131  & ~n2262 ;
  assign n2566 = n969 & ~n1889 ;
  assign n2567 = ~n2565 & n2566 ;
  assign n2572 = \PhyAddrPointer_reg[24]/NET0131  & ~n1902 ;
  assign n2573 = ~n1993 & ~n2572 ;
  assign n2574 = ~n2567 & n2573 ;
  assign n2575 = ~n2571 & n2574 ;
  assign n2576 = ~n2564 & n2575 ;
  assign n2577 = \PhyAddrPointer_reg[26]/NET0131  & n906 ;
  assign n2578 = ~n2065 & ~n2577 ;
  assign n2579 = n773 & ~n2578 ;
  assign n2580 = \PhyAddrPointer_reg[26]/NET0131  & ~n1852 ;
  assign n2581 = ~n2071 & ~n2580 ;
  assign n2582 = ~n2579 & n2581 ;
  assign n2583 = n929 & ~n2582 ;
  assign n2587 = \PhyAddrPointer_reg[1]/NET0131  & n1890 ;
  assign n2588 = ~\PhyAddrPointer_reg[26]/NET0131  & ~n2587 ;
  assign n2589 = ~n2304 & ~n2588 ;
  assign n2590 = n2100 & n2589 ;
  assign n2584 = ~\PhyAddrPointer_reg[26]/NET0131  & ~n1890 ;
  assign n2585 = n969 & ~n1891 ;
  assign n2586 = ~n2584 & n2585 ;
  assign n2591 = \PhyAddrPointer_reg[26]/NET0131  & ~n1902 ;
  assign n2592 = ~n2084 & ~n2591 ;
  assign n2593 = ~n2586 & n2592 ;
  assign n2594 = ~n2590 & n2593 ;
  assign n2595 = ~n2583 & n2594 ;
  assign n2618 = \InstAddrPointer_reg[7]/NET0131  & n906 ;
  assign n2619 = n1451 & ~n1769 ;
  assign n2620 = ~n1433 & ~n1447 ;
  assign n2621 = ~n2619 & ~n2620 ;
  assign n2622 = n2619 & n2620 ;
  assign n2623 = ~n2621 & ~n2622 ;
  assign n2624 = ~n906 & ~n2623 ;
  assign n2625 = ~n2618 & ~n2624 ;
  assign n2626 = n773 & ~n2625 ;
  assign n2602 = ~n1544 & ~n1580 ;
  assign n2604 = ~n1711 & n2602 ;
  assign n2603 = n1711 & ~n2602 ;
  assign n2605 = n899 & ~n2603 ;
  assign n2606 = ~n2604 & n2605 ;
  assign n2599 = READY_n_pad & n840 ;
  assign n2600 = n1957 & ~n2599 ;
  assign n2601 = \InstAddrPointer_reg[7]/NET0131  & ~n2600 ;
  assign n2617 = ~n811 & n983 ;
  assign n2611 = ~n828 & ~n836 ;
  assign n2612 = ~n782 & ~n2611 ;
  assign n2610 = ~\InstAddrPointer_reg[7]/NET0131  & READY_n_pad ;
  assign n2613 = ~READY_n_pad & ~n1432 ;
  assign n2614 = ~n2610 & ~n2613 ;
  assign n2615 = ~n834 & n2614 ;
  assign n2616 = ~n2612 & n2615 ;
  assign n2598 = n766 & n1543 ;
  assign n2607 = n840 & n846 ;
  assign n2608 = ~n788 & ~n2607 ;
  assign n2609 = n1432 & ~n2608 ;
  assign n2627 = ~n2598 & ~n2609 ;
  assign n2628 = ~n2616 & n2627 ;
  assign n2629 = ~n2617 & n2628 ;
  assign n2630 = ~n2601 & n2629 ;
  assign n2631 = ~n2606 & n2630 ;
  assign n2632 = ~n2626 & n2631 ;
  assign n2633 = n929 & ~n2632 ;
  assign n2596 = \InstAddrPointer_reg[7]/NET0131  & n1661 ;
  assign n2597 = \rEIP_reg[7]/NET0131  & n1655 ;
  assign n2634 = ~n2596 & ~n2597 ;
  assign n2635 = ~n2633 & n2634 ;
  assign n2639 = \InstAddrPointer_reg[9]/NET0131  & n906 ;
  assign n2644 = n1454 & ~n1477 ;
  assign n2645 = ~n2424 & ~n2644 ;
  assign n2646 = n1014 & ~n2645 ;
  assign n2641 = n1314 & ~n1683 ;
  assign n2640 = ~n1314 & n1683 ;
  assign n2642 = ~n1014 & ~n2640 ;
  assign n2643 = ~n2641 & n2642 ;
  assign n2647 = ~n906 & ~n2643 ;
  assign n2648 = ~n2646 & n2647 ;
  assign n2649 = ~n2639 & ~n2648 ;
  assign n2650 = n773 & ~n2649 ;
  assign n2655 = ~n1596 & ~n1713 ;
  assign n2654 = n1596 & n1713 ;
  assign n2656 = n899 & ~n2654 ;
  assign n2657 = ~n2655 & n2656 ;
  assign n2651 = ~n873 & n1477 ;
  assign n2652 = ~n811 & n1314 ;
  assign n2638 = \InstAddrPointer_reg[9]/NET0131  & ~n2073 ;
  assign n2653 = n766 & n1596 ;
  assign n2658 = ~n2638 & ~n2653 ;
  assign n2659 = ~n2652 & n2658 ;
  assign n2660 = ~n2651 & n2659 ;
  assign n2661 = ~n2657 & n2660 ;
  assign n2662 = ~n2650 & n2661 ;
  assign n2663 = n929 & ~n2662 ;
  assign n2636 = \rEIP_reg[9]/NET0131  & n1655 ;
  assign n2637 = \InstAddrPointer_reg[9]/NET0131  & n1661 ;
  assign n2664 = ~n2636 & ~n2637 ;
  assign n2665 = ~n2663 & n2664 ;
  assign n2666 = \PhyAddrPointer_reg[13]/NET0131  & n906 ;
  assign n2667 = ~n2432 & ~n2666 ;
  assign n2668 = n773 & ~n2667 ;
  assign n2669 = \PhyAddrPointer_reg[13]/NET0131  & ~n1852 ;
  assign n2670 = ~n2442 & ~n2669 ;
  assign n2671 = ~n2668 & n2670 ;
  assign n2672 = n929 & ~n2671 ;
  assign n2678 = \PhyAddrPointer_reg[12]/NET0131  & n2470 ;
  assign n2679 = ~\PhyAddrPointer_reg[13]/NET0131  & ~n2678 ;
  assign n2680 = ~n2236 & ~n2679 ;
  assign n2681 = n2100 & n2680 ;
  assign n2674 = n1877 & n1878 ;
  assign n2675 = ~\PhyAddrPointer_reg[13]/NET0131  & ~n2674 ;
  assign n2676 = n969 & ~n1880 ;
  assign n2677 = ~n2675 & n2676 ;
  assign n2673 = \PhyAddrPointer_reg[13]/NET0131  & ~n1902 ;
  assign n2682 = ~n2454 & ~n2673 ;
  assign n2683 = ~n2677 & n2682 ;
  assign n2684 = ~n2681 & n2683 ;
  assign n2685 = ~n2672 & n2684 ;
  assign n2686 = \PhyAddrPointer_reg[16]/NET0131  & n906 ;
  assign n2687 = n1471 & n2057 ;
  assign n2689 = ~\InstAddrPointer_reg[16]/NET0131  & ~n1470 ;
  assign n2690 = ~n1329 & ~n2689 ;
  assign n2691 = ~n2687 & n2690 ;
  assign n2688 = ~\InstAddrPointer_reg[16]/NET0131  & n2687 ;
  assign n2692 = n1014 & ~n2688 ;
  assign n2693 = ~n2691 & n2692 ;
  assign n2694 = n1345 & ~n2022 ;
  assign n2695 = n1324 & n1346 ;
  assign n2696 = ~n1014 & ~n2695 ;
  assign n2697 = ~n2694 & n2696 ;
  assign n2698 = ~n906 & ~n2697 ;
  assign n2699 = ~n2693 & n2698 ;
  assign n2700 = ~n2686 & ~n2699 ;
  assign n2701 = n773 & ~n2700 ;
  assign n2702 = \PhyAddrPointer_reg[16]/NET0131  & ~n1852 ;
  assign n2703 = ~n1799 & ~n2035 ;
  assign n2704 = n899 & ~n2036 ;
  assign n2705 = ~n2703 & n2704 ;
  assign n2706 = ~n2702 & ~n2705 ;
  assign n2707 = ~n2701 & n2706 ;
  assign n2708 = n929 & ~n2707 ;
  assign n2713 = ~\PhyAddrPointer_reg[16]/NET0131  & ~n2239 ;
  assign n2714 = n1882 & n2237 ;
  assign n2715 = ~n2713 & ~n2714 ;
  assign n2716 = n2100 & n2715 ;
  assign n2710 = \PhyAddrPointer_reg[16]/NET0131  & n2249 ;
  assign n2709 = ~\PhyAddrPointer_reg[16]/NET0131  & ~n2249 ;
  assign n2711 = n969 & ~n2709 ;
  assign n2712 = ~n2710 & n2711 ;
  assign n2717 = \PhyAddrPointer_reg[16]/NET0131  & ~n1902 ;
  assign n2718 = \rEIP_reg[16]/NET0131  & n1655 ;
  assign n2719 = ~n2717 & ~n2718 ;
  assign n2720 = ~n2712 & n2719 ;
  assign n2721 = ~n2716 & n2720 ;
  assign n2722 = ~n2708 & n2721 ;
  assign n2728 = ~\InstAddrPointer_reg[17]/NET0131  & ~n1329 ;
  assign n2729 = ~n1347 & ~n2728 ;
  assign n2730 = n1463 & n1472 ;
  assign n2731 = n2424 & n2730 ;
  assign n2732 = ~n2729 & ~n2731 ;
  assign n2733 = n2729 & n2731 ;
  assign n2734 = ~n2732 & ~n2733 ;
  assign n2735 = n1014 & ~n2734 ;
  assign n2723 = n1684 & n1685 ;
  assign n2725 = ~n1354 & n2723 ;
  assign n2724 = n1354 & ~n2723 ;
  assign n2726 = ~n1014 & ~n2724 ;
  assign n2727 = ~n2725 & n2726 ;
  assign n2736 = ~n906 & ~n2727 ;
  assign n2737 = ~n2735 & n2736 ;
  assign n2738 = n773 & n2737 ;
  assign n2739 = ~n910 & n1852 ;
  assign n2740 = \PhyAddrPointer_reg[17]/NET0131  & ~n2739 ;
  assign n2742 = n1586 & n1714 ;
  assign n2741 = ~n1586 & ~n1714 ;
  assign n2743 = n899 & ~n2741 ;
  assign n2744 = ~n2742 & n2743 ;
  assign n2745 = ~n2740 & ~n2744 ;
  assign n2746 = ~n2738 & n2745 ;
  assign n2747 = n929 & ~n2746 ;
  assign n2751 = ~\PhyAddrPointer_reg[17]/NET0131  & ~n2714 ;
  assign n2752 = ~n2265 & ~n2751 ;
  assign n2753 = n2100 & n2752 ;
  assign n2748 = ~\PhyAddrPointer_reg[17]/NET0131  & ~n2710 ;
  assign n2749 = n969 & ~n1884 ;
  assign n2750 = ~n2748 & n2749 ;
  assign n2754 = \PhyAddrPointer_reg[17]/NET0131  & ~n1902 ;
  assign n2755 = \rEIP_reg[17]/NET0131  & n1655 ;
  assign n2756 = ~n2754 & ~n2755 ;
  assign n2757 = ~n2750 & n2756 ;
  assign n2758 = ~n2753 & n2757 ;
  assign n2759 = ~n2747 & n2758 ;
  assign n2760 = \PhyAddrPointer_reg[18]/NET0131  & n906 ;
  assign n2764 = n1473 & n2057 ;
  assign n2765 = ~n1467 & ~n2764 ;
  assign n2766 = ~n2058 & ~n2765 ;
  assign n2767 = n1014 & ~n2766 ;
  assign n2761 = n1356 & ~n2725 ;
  assign n2762 = ~n1014 & ~n2514 ;
  assign n2763 = ~n2761 & n2762 ;
  assign n2768 = ~n906 & ~n2763 ;
  assign n2769 = ~n2767 & n2768 ;
  assign n2770 = ~n2760 & ~n2769 ;
  assign n2771 = n773 & ~n2770 ;
  assign n2772 = \PhyAddrPointer_reg[18]/NET0131  & ~n1852 ;
  assign n2773 = ~n1605 & ~n1608 ;
  assign n2774 = n899 & ~n1609 ;
  assign n2775 = ~n2773 & n2774 ;
  assign n2776 = ~n2772 & ~n2775 ;
  assign n2777 = ~n2771 & n2776 ;
  assign n2778 = n929 & ~n2777 ;
  assign n2780 = ~\PhyAddrPointer_reg[18]/NET0131  & ~n2265 ;
  assign n2781 = ~n2506 & ~n2780 ;
  assign n2782 = n2100 & n2781 ;
  assign n2783 = ~\PhyAddrPointer_reg[18]/NET0131  & ~n1884 ;
  assign n2784 = n2500 & ~n2783 ;
  assign n2779 = \PhyAddrPointer_reg[18]/NET0131  & ~n1902 ;
  assign n2785 = \rEIP_reg[18]/NET0131  & n1655 ;
  assign n2786 = ~n2779 & ~n2785 ;
  assign n2787 = ~n2784 & n2786 ;
  assign n2788 = ~n2782 & n2787 ;
  assign n2789 = ~n2778 & n2788 ;
  assign n2791 = \PhyAddrPointer_reg[21]/NET0131  & n906 ;
  assign n2795 = ~n1482 & ~n1485 ;
  assign n2796 = ~n1970 & ~n2795 ;
  assign n2797 = n1014 & ~n2796 ;
  assign n2792 = n1335 & ~n1688 ;
  assign n2793 = ~n1014 & ~n1689 ;
  assign n2794 = ~n2792 & n2793 ;
  assign n2798 = ~n906 & ~n2794 ;
  assign n2799 = ~n2797 & n2798 ;
  assign n2800 = ~n2791 & ~n2799 ;
  assign n2801 = n773 & ~n2800 ;
  assign n2802 = \PhyAddrPointer_reg[21]/NET0131  & ~n1852 ;
  assign n2804 = n1612 & n1717 ;
  assign n2803 = ~n1612 & ~n1717 ;
  assign n2805 = n899 & ~n2803 ;
  assign n2806 = ~n2804 & n2805 ;
  assign n2807 = ~n2802 & ~n2806 ;
  assign n2808 = ~n2801 & n2807 ;
  assign n2809 = n929 & ~n2808 ;
  assign n2810 = \PhyAddrPointer_reg[20]/NET0131  & n2509 ;
  assign n2811 = ~\PhyAddrPointer_reg[21]/NET0131  & ~n2810 ;
  assign n2812 = ~n2266 & ~n2811 ;
  assign n2813 = n1867 & n2812 ;
  assign n2816 = \PhyAddrPointer_reg[20]/NET0131  & n2508 ;
  assign n2817 = ~n1906 & n2816 ;
  assign n2818 = ~\PhyAddrPointer_reg[21]/NET0131  & ~n2817 ;
  assign n2815 = n1888 & ~n1906 ;
  assign n2819 = n933 & ~n2815 ;
  assign n2820 = ~n2818 & n2819 ;
  assign n2790 = \PhyAddrPointer_reg[21]/NET0131  & ~n1902 ;
  assign n2814 = \rEIP_reg[21]/NET0131  & n1655 ;
  assign n2821 = ~n2790 & ~n2814 ;
  assign n2822 = ~n2820 & n2821 ;
  assign n2823 = ~n2813 & n2822 ;
  assign n2824 = ~n2809 & n2823 ;
  assign n2825 = \PhyAddrPointer_reg[25]/NET0131  & n906 ;
  assign n2826 = ~n2206 & ~n2825 ;
  assign n2827 = n773 & ~n2826 ;
  assign n2828 = \PhyAddrPointer_reg[25]/NET0131  & ~n1852 ;
  assign n2829 = ~n2213 & ~n2828 ;
  assign n2830 = ~n2827 & n2829 ;
  assign n2831 = n929 & ~n2830 ;
  assign n2832 = ~\PhyAddrPointer_reg[25]/NET0131  & ~n2569 ;
  assign n2833 = ~n2587 & ~n2832 ;
  assign n2838 = ~\DataWidth_reg[1]/NET0131  & ~n2833 ;
  assign n2835 = ~\PhyAddrPointer_reg[25]/NET0131  & ~n1889 ;
  assign n2836 = ~n1890 & ~n2835 ;
  assign n2837 = \DataWidth_reg[1]/NET0131  & ~n2836 ;
  assign n2839 = n933 & ~n2837 ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2834 = n1867 & n2833 ;
  assign n2841 = \PhyAddrPointer_reg[25]/NET0131  & ~n1902 ;
  assign n2842 = ~n2228 & ~n2841 ;
  assign n2843 = ~n2834 & n2842 ;
  assign n2844 = ~n2840 & n2843 ;
  assign n2845 = ~n2831 & n2844 ;
  assign n2846 = \PhyAddrPointer_reg[8]/NET0131  & n906 ;
  assign n2847 = ~n2403 & ~n2846 ;
  assign n2848 = n773 & ~n2847 ;
  assign n2849 = \PhyAddrPointer_reg[8]/NET0131  & ~n1852 ;
  assign n2850 = ~n2409 & ~n2849 ;
  assign n2851 = ~n2848 & n2850 ;
  assign n2852 = n929 & ~n2851 ;
  assign n2856 = ~\PhyAddrPointer_reg[8]/NET0131  & ~n2232 ;
  assign n2857 = ~n2233 & ~n2856 ;
  assign n2858 = n2100 & n2857 ;
  assign n2853 = ~\PhyAddrPointer_reg[8]/NET0131  & ~n1874 ;
  assign n2854 = n969 & ~n1875 ;
  assign n2855 = ~n2853 & n2854 ;
  assign n2859 = \PhyAddrPointer_reg[8]/NET0131  & ~n1902 ;
  assign n2860 = ~n2386 & ~n2859 ;
  assign n2861 = ~n2855 & n2860 ;
  assign n2862 = ~n2858 & n2861 ;
  assign n2863 = ~n2852 & n2862 ;
  assign n2888 = ~READY_n_pad & ~n1409 ;
  assign n2889 = ~n858 & ~n2888 ;
  assign n2886 = ~n849 & ~n911 ;
  assign n2887 = ~n860 & n2886 ;
  assign n2890 = ~n836 & ~n975 ;
  assign n2891 = n2887 & ~n2890 ;
  assign n2892 = ~n2889 & n2891 ;
  assign n2893 = \InstAddrPointer_reg[4]/NET0131  & ~n2892 ;
  assign n2867 = ~n873 & n1409 ;
  assign n2866 = ~n811 & n1129 ;
  assign n2882 = n765 & ~n1557 ;
  assign n2883 = ~\InstAddrPointer_reg[4]/NET0131  & ~n765 ;
  assign n2884 = ~n2882 & ~n2883 ;
  assign n2885 = ~n740 & n2884 ;
  assign n2894 = ~n2866 & ~n2885 ;
  assign n2895 = ~n2867 & n2894 ;
  assign n2868 = \InstAddrPointer_reg[4]/NET0131  & n906 ;
  assign n2869 = ~n1410 & ~n1425 ;
  assign n2870 = ~n2003 & ~n2869 ;
  assign n2871 = n2003 & n2869 ;
  assign n2872 = ~n2870 & ~n2871 ;
  assign n2873 = ~n906 & ~n2872 ;
  assign n2874 = ~n2868 & ~n2873 ;
  assign n2875 = n773 & ~n2874 ;
  assign n2876 = ~n1558 & ~n1574 ;
  assign n2877 = ~n1561 & ~n1572 ;
  assign n2879 = n2876 & n2877 ;
  assign n2878 = ~n2876 & ~n2877 ;
  assign n2880 = n899 & ~n2878 ;
  assign n2881 = ~n2879 & n2880 ;
  assign n2896 = ~n2875 & ~n2881 ;
  assign n2897 = n2895 & n2896 ;
  assign n2898 = ~n2893 & n2897 ;
  assign n2899 = n929 & ~n2898 ;
  assign n2864 = \rEIP_reg[4]/NET0131  & n1655 ;
  assign n2865 = \InstAddrPointer_reg[4]/NET0131  & n1661 ;
  assign n2900 = ~n2864 & ~n2865 ;
  assign n2901 = ~n2899 & n2900 ;
  assign n2903 = \InstAddrPointer_reg[6]/NET0131  & n906 ;
  assign n2909 = ~n1440 & ~n1448 ;
  assign n2910 = ~n2008 & n2909 ;
  assign n2911 = n2008 & ~n2909 ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = n1014 & ~n2912 ;
  assign n2904 = ~n1053 & ~n1055 ;
  assign n2906 = n1283 & n2904 ;
  assign n2905 = ~n1283 & ~n2904 ;
  assign n2907 = ~n1014 & ~n2905 ;
  assign n2908 = ~n2906 & n2907 ;
  assign n2914 = ~n906 & ~n2908 ;
  assign n2915 = ~n2913 & n2914 ;
  assign n2916 = ~n2903 & ~n2915 ;
  assign n2917 = n773 & ~n2916 ;
  assign n2925 = n1578 & ~n1579 ;
  assign n2922 = ~n1551 & ~n1579 ;
  assign n2923 = ~n1554 & ~n1577 ;
  assign n2924 = ~n2922 & ~n2923 ;
  assign n2926 = n899 & ~n2924 ;
  assign n2927 = ~n2925 & n2926 ;
  assign n2919 = \InstAddrPointer_reg[6]/NET0131  & ~n1816 ;
  assign n2920 = ~n873 & n1439 ;
  assign n2918 = n766 & n1550 ;
  assign n2921 = ~n811 & n1052 ;
  assign n2928 = ~n2918 & ~n2921 ;
  assign n2929 = ~n2920 & n2928 ;
  assign n2930 = ~n2919 & n2929 ;
  assign n2931 = ~n2927 & n2930 ;
  assign n2932 = ~n2917 & n2931 ;
  assign n2933 = n929 & ~n2932 ;
  assign n2902 = \rEIP_reg[6]/NET0131  & n1655 ;
  assign n2934 = \InstAddrPointer_reg[6]/NET0131  & n1661 ;
  assign n2935 = ~n2902 & ~n2934 ;
  assign n2936 = ~n2933 & n2935 ;
  assign n2937 = n739 & n765 ;
  assign n3132 = n786 & n792 ;
  assign n3133 = n841 & ~n3132 ;
  assign n3134 = ~n739 & ~n3133 ;
  assign n3135 = ~n2937 & ~n3134 ;
  assign n3136 = \EAX_reg[0]/NET0131  & \EAX_reg[1]/NET0131  ;
  assign n3137 = \EAX_reg[2]/NET0131  & n3136 ;
  assign n3138 = \EAX_reg[3]/NET0131  & n3137 ;
  assign n3139 = \EAX_reg[4]/NET0131  & n3138 ;
  assign n3140 = \EAX_reg[5]/NET0131  & n3139 ;
  assign n3141 = \EAX_reg[6]/NET0131  & n3140 ;
  assign n3142 = \EAX_reg[7]/NET0131  & n3141 ;
  assign n3143 = \EAX_reg[8]/NET0131  & n3142 ;
  assign n3144 = \EAX_reg[9]/NET0131  & n3143 ;
  assign n3145 = \EAX_reg[10]/NET0131  & n3144 ;
  assign n3146 = \EAX_reg[11]/NET0131  & n3145 ;
  assign n3147 = \EAX_reg[12]/NET0131  & n3146 ;
  assign n3148 = \EAX_reg[13]/NET0131  & n3147 ;
  assign n3149 = \EAX_reg[14]/NET0131  & n3148 ;
  assign n3150 = \EAX_reg[15]/NET0131  & n3149 ;
  assign n3151 = \EAX_reg[16]/NET0131  & n3150 ;
  assign n3152 = \EAX_reg[17]/NET0131  & n3151 ;
  assign n3153 = \EAX_reg[18]/NET0131  & n3152 ;
  assign n3154 = \EAX_reg[20]/NET0131  & \EAX_reg[21]/NET0131  ;
  assign n3155 = \EAX_reg[19]/NET0131  & n3154 ;
  assign n3156 = \EAX_reg[22]/NET0131  & n3155 ;
  assign n3157 = n3153 & n3156 ;
  assign n3158 = \EAX_reg[23]/NET0131  & \EAX_reg[24]/NET0131  ;
  assign n3159 = n3157 & n3158 ;
  assign n3160 = \EAX_reg[25]/NET0131  & n3159 ;
  assign n3161 = \EAX_reg[26]/NET0131  & n3160 ;
  assign n3162 = n3132 & ~n3161 ;
  assign n3163 = ~n3135 & ~n3162 ;
  assign n3164 = \EAX_reg[27]/NET0131  & ~n3163 ;
  assign n3172 = ~\EAX_reg[27]/NET0131  & n3132 ;
  assign n3173 = n3161 & n3172 ;
  assign n3165 = \EAX_reg[27]/NET0131  & ~n846 ;
  assign n3169 = \Datai[27]_pad  & n846 ;
  assign n3170 = ~n3165 & ~n3169 ;
  assign n3171 = n840 & ~n3170 ;
  assign n2942 = \InstQueue_reg[13][7]/NET0131  & n461 ;
  assign n2943 = \InstQueue_reg[4][7]/NET0131  & n488 ;
  assign n2956 = ~n2942 & ~n2943 ;
  assign n2944 = \InstQueue_reg[7][7]/NET0131  & n472 ;
  assign n2945 = \InstQueue_reg[11][7]/NET0131  & n486 ;
  assign n2957 = ~n2944 & ~n2945 ;
  assign n2964 = n2956 & n2957 ;
  assign n2938 = \InstQueue_reg[1][7]/NET0131  & n470 ;
  assign n2939 = \InstQueue_reg[9][7]/NET0131  & n482 ;
  assign n2954 = ~n2938 & ~n2939 ;
  assign n2940 = \InstQueue_reg[2][7]/NET0131  & n522 ;
  assign n2941 = \InstQueue_reg[6][7]/NET0131  & n476 ;
  assign n2955 = ~n2940 & ~n2941 ;
  assign n2965 = n2954 & n2955 ;
  assign n2966 = n2964 & n2965 ;
  assign n2950 = \InstQueue_reg[8][7]/NET0131  & n490 ;
  assign n2951 = \InstQueue_reg[5][7]/NET0131  & n458 ;
  assign n2960 = ~n2950 & ~n2951 ;
  assign n2952 = \InstQueue_reg[15][7]/NET0131  & n468 ;
  assign n2953 = \InstQueue_reg[12][7]/NET0131  & n484 ;
  assign n2961 = ~n2952 & ~n2953 ;
  assign n2962 = n2960 & n2961 ;
  assign n2946 = \InstQueue_reg[0][7]/NET0131  & n465 ;
  assign n2947 = \InstQueue_reg[3][7]/NET0131  & n474 ;
  assign n2958 = ~n2946 & ~n2947 ;
  assign n2948 = \InstQueue_reg[14][7]/NET0131  & n492 ;
  assign n2949 = \InstQueue_reg[10][7]/NET0131  & n454 ;
  assign n2959 = ~n2948 & ~n2949 ;
  assign n2963 = n2958 & n2959 ;
  assign n2967 = n2962 & n2963 ;
  assign n2968 = n2966 & n2967 ;
  assign n2973 = \InstQueue_reg[14][0]/NET0131  & n461 ;
  assign n2974 = \InstQueue_reg[6][0]/NET0131  & n458 ;
  assign n2987 = ~n2973 & ~n2974 ;
  assign n2975 = \InstQueue_reg[3][0]/NET0131  & n522 ;
  assign n2976 = \InstQueue_reg[11][0]/NET0131  & n454 ;
  assign n2988 = ~n2975 & ~n2976 ;
  assign n2995 = n2987 & n2988 ;
  assign n2969 = \InstQueue_reg[7][0]/NET0131  & n476 ;
  assign n2970 = \InstQueue_reg[10][0]/NET0131  & n482 ;
  assign n2985 = ~n2969 & ~n2970 ;
  assign n2971 = \InstQueue_reg[1][0]/NET0131  & n465 ;
  assign n2972 = \InstQueue_reg[2][0]/NET0131  & n470 ;
  assign n2986 = ~n2971 & ~n2972 ;
  assign n2996 = n2985 & n2986 ;
  assign n2997 = n2995 & n2996 ;
  assign n2981 = \InstQueue_reg[0][0]/NET0131  & n468 ;
  assign n2982 = \InstQueue_reg[5][0]/NET0131  & n488 ;
  assign n2991 = ~n2981 & ~n2982 ;
  assign n2983 = \InstQueue_reg[9][0]/NET0131  & n490 ;
  assign n2984 = \InstQueue_reg[13][0]/NET0131  & n484 ;
  assign n2992 = ~n2983 & ~n2984 ;
  assign n2993 = n2991 & n2992 ;
  assign n2977 = \InstQueue_reg[8][0]/NET0131  & n472 ;
  assign n2978 = \InstQueue_reg[4][0]/NET0131  & n474 ;
  assign n2989 = ~n2977 & ~n2978 ;
  assign n2979 = \InstQueue_reg[12][0]/NET0131  & n486 ;
  assign n2980 = \InstQueue_reg[15][0]/NET0131  & n492 ;
  assign n2990 = ~n2979 & ~n2980 ;
  assign n2994 = n2989 & n2990 ;
  assign n2998 = n2993 & n2994 ;
  assign n2999 = n2997 & n2998 ;
  assign n3000 = ~n2968 & ~n2999 ;
  assign n3005 = \InstQueue_reg[14][1]/NET0131  & n461 ;
  assign n3006 = \InstQueue_reg[6][1]/NET0131  & n458 ;
  assign n3019 = ~n3005 & ~n3006 ;
  assign n3007 = \InstQueue_reg[3][1]/NET0131  & n522 ;
  assign n3008 = \InstQueue_reg[11][1]/NET0131  & n454 ;
  assign n3020 = ~n3007 & ~n3008 ;
  assign n3027 = n3019 & n3020 ;
  assign n3001 = \InstQueue_reg[7][1]/NET0131  & n476 ;
  assign n3002 = \InstQueue_reg[10][1]/NET0131  & n482 ;
  assign n3017 = ~n3001 & ~n3002 ;
  assign n3003 = \InstQueue_reg[1][1]/NET0131  & n465 ;
  assign n3004 = \InstQueue_reg[2][1]/NET0131  & n470 ;
  assign n3018 = ~n3003 & ~n3004 ;
  assign n3028 = n3017 & n3018 ;
  assign n3029 = n3027 & n3028 ;
  assign n3013 = \InstQueue_reg[0][1]/NET0131  & n468 ;
  assign n3014 = \InstQueue_reg[5][1]/NET0131  & n488 ;
  assign n3023 = ~n3013 & ~n3014 ;
  assign n3015 = \InstQueue_reg[9][1]/NET0131  & n490 ;
  assign n3016 = \InstQueue_reg[13][1]/NET0131  & n484 ;
  assign n3024 = ~n3015 & ~n3016 ;
  assign n3025 = n3023 & n3024 ;
  assign n3009 = \InstQueue_reg[8][1]/NET0131  & n472 ;
  assign n3010 = \InstQueue_reg[4][1]/NET0131  & n474 ;
  assign n3021 = ~n3009 & ~n3010 ;
  assign n3011 = \InstQueue_reg[12][1]/NET0131  & n486 ;
  assign n3012 = \InstQueue_reg[15][1]/NET0131  & n492 ;
  assign n3022 = ~n3011 & ~n3012 ;
  assign n3026 = n3021 & n3022 ;
  assign n3030 = n3025 & n3026 ;
  assign n3031 = n3029 & n3030 ;
  assign n3032 = n3000 & ~n3031 ;
  assign n3037 = \InstQueue_reg[14][2]/NET0131  & n461 ;
  assign n3038 = \InstQueue_reg[5][2]/NET0131  & n488 ;
  assign n3051 = ~n3037 & ~n3038 ;
  assign n3039 = \InstQueue_reg[0][2]/NET0131  & n468 ;
  assign n3040 = \InstQueue_reg[2][2]/NET0131  & n470 ;
  assign n3052 = ~n3039 & ~n3040 ;
  assign n3059 = n3051 & n3052 ;
  assign n3033 = \InstQueue_reg[10][2]/NET0131  & n482 ;
  assign n3034 = \InstQueue_reg[13][2]/NET0131  & n484 ;
  assign n3049 = ~n3033 & ~n3034 ;
  assign n3035 = \InstQueue_reg[9][2]/NET0131  & n490 ;
  assign n3036 = \InstQueue_reg[7][2]/NET0131  & n476 ;
  assign n3050 = ~n3035 & ~n3036 ;
  assign n3060 = n3049 & n3050 ;
  assign n3061 = n3059 & n3060 ;
  assign n3045 = \InstQueue_reg[8][2]/NET0131  & n472 ;
  assign n3046 = \InstQueue_reg[6][2]/NET0131  & n458 ;
  assign n3055 = ~n3045 & ~n3046 ;
  assign n3047 = \InstQueue_reg[3][2]/NET0131  & n522 ;
  assign n3048 = \InstQueue_reg[4][2]/NET0131  & n474 ;
  assign n3056 = ~n3047 & ~n3048 ;
  assign n3057 = n3055 & n3056 ;
  assign n3041 = \InstQueue_reg[12][2]/NET0131  & n486 ;
  assign n3042 = \InstQueue_reg[1][2]/NET0131  & n465 ;
  assign n3053 = ~n3041 & ~n3042 ;
  assign n3043 = \InstQueue_reg[15][2]/NET0131  & n492 ;
  assign n3044 = \InstQueue_reg[11][2]/NET0131  & n454 ;
  assign n3054 = ~n3043 & ~n3044 ;
  assign n3058 = n3053 & n3054 ;
  assign n3062 = n3057 & n3058 ;
  assign n3063 = n3061 & n3062 ;
  assign n3064 = n3032 & ~n3063 ;
  assign n3069 = \InstQueue_reg[14][3]/NET0131  & n461 ;
  assign n3070 = \InstQueue_reg[6][3]/NET0131  & n458 ;
  assign n3083 = ~n3069 & ~n3070 ;
  assign n3071 = \InstQueue_reg[3][3]/NET0131  & n522 ;
  assign n3072 = \InstQueue_reg[11][3]/NET0131  & n454 ;
  assign n3084 = ~n3071 & ~n3072 ;
  assign n3091 = n3083 & n3084 ;
  assign n3065 = \InstQueue_reg[7][3]/NET0131  & n476 ;
  assign n3066 = \InstQueue_reg[10][3]/NET0131  & n482 ;
  assign n3081 = ~n3065 & ~n3066 ;
  assign n3067 = \InstQueue_reg[1][3]/NET0131  & n465 ;
  assign n3068 = \InstQueue_reg[2][3]/NET0131  & n470 ;
  assign n3082 = ~n3067 & ~n3068 ;
  assign n3092 = n3081 & n3082 ;
  assign n3093 = n3091 & n3092 ;
  assign n3077 = \InstQueue_reg[0][3]/NET0131  & n468 ;
  assign n3078 = \InstQueue_reg[5][3]/NET0131  & n488 ;
  assign n3087 = ~n3077 & ~n3078 ;
  assign n3079 = \InstQueue_reg[9][3]/NET0131  & n490 ;
  assign n3080 = \InstQueue_reg[13][3]/NET0131  & n484 ;
  assign n3088 = ~n3079 & ~n3080 ;
  assign n3089 = n3087 & n3088 ;
  assign n3073 = \InstQueue_reg[8][3]/NET0131  & n472 ;
  assign n3074 = \InstQueue_reg[4][3]/NET0131  & n474 ;
  assign n3085 = ~n3073 & ~n3074 ;
  assign n3075 = \InstQueue_reg[12][3]/NET0131  & n486 ;
  assign n3076 = \InstQueue_reg[15][3]/NET0131  & n492 ;
  assign n3086 = ~n3075 & ~n3076 ;
  assign n3090 = n3085 & n3086 ;
  assign n3094 = n3089 & n3090 ;
  assign n3095 = n3093 & n3094 ;
  assign n3096 = n3064 & ~n3095 ;
  assign n3101 = \InstQueue_reg[14][4]/NET0131  & n461 ;
  assign n3102 = \InstQueue_reg[5][4]/NET0131  & n488 ;
  assign n3115 = ~n3101 & ~n3102 ;
  assign n3103 = \InstQueue_reg[0][4]/NET0131  & n468 ;
  assign n3104 = \InstQueue_reg[2][4]/NET0131  & n470 ;
  assign n3116 = ~n3103 & ~n3104 ;
  assign n3123 = n3115 & n3116 ;
  assign n3097 = \InstQueue_reg[10][4]/NET0131  & n482 ;
  assign n3098 = \InstQueue_reg[13][4]/NET0131  & n484 ;
  assign n3113 = ~n3097 & ~n3098 ;
  assign n3099 = \InstQueue_reg[9][4]/NET0131  & n490 ;
  assign n3100 = \InstQueue_reg[7][4]/NET0131  & n476 ;
  assign n3114 = ~n3099 & ~n3100 ;
  assign n3124 = n3113 & n3114 ;
  assign n3125 = n3123 & n3124 ;
  assign n3109 = \InstQueue_reg[8][4]/NET0131  & n472 ;
  assign n3110 = \InstQueue_reg[6][4]/NET0131  & n458 ;
  assign n3119 = ~n3109 & ~n3110 ;
  assign n3111 = \InstQueue_reg[3][4]/NET0131  & n522 ;
  assign n3112 = \InstQueue_reg[4][4]/NET0131  & n474 ;
  assign n3120 = ~n3111 & ~n3112 ;
  assign n3121 = n3119 & n3120 ;
  assign n3105 = \InstQueue_reg[12][4]/NET0131  & n486 ;
  assign n3106 = \InstQueue_reg[1][4]/NET0131  & n465 ;
  assign n3117 = ~n3105 & ~n3106 ;
  assign n3107 = \InstQueue_reg[15][4]/NET0131  & n492 ;
  assign n3108 = \InstQueue_reg[11][4]/NET0131  & n454 ;
  assign n3118 = ~n3107 & ~n3108 ;
  assign n3122 = n3117 & n3118 ;
  assign n3126 = n3121 & n3122 ;
  assign n3127 = n3125 & n3126 ;
  assign n3128 = ~n3096 & n3127 ;
  assign n3129 = n3096 & ~n3127 ;
  assign n3130 = ~n3128 & ~n3129 ;
  assign n3131 = n2937 & n3130 ;
  assign n3166 = \Datai[11]_pad  & n846 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = n782 & ~n3167 ;
  assign n3174 = ~n3131 & ~n3168 ;
  assign n3175 = ~n3171 & n3174 ;
  assign n3176 = ~n3173 & n3175 ;
  assign n3177 = ~n3164 & n3176 ;
  assign n3178 = n929 & ~n3177 ;
  assign n3179 = ~n952 & ~n956 ;
  assign n3180 = ~n931 & ~n939 ;
  assign n3181 = n3179 & n3180 ;
  assign n3182 = \EAX_reg[27]/NET0131  & ~n3181 ;
  assign n3183 = ~n3178 & ~n3182 ;
  assign n3185 = n818 & n929 ;
  assign n3186 = \State2_reg[3]/NET0131  & ~n936 ;
  assign n3187 = ~n928 & ~n3186 ;
  assign n3188 = \InstQueueRd_Addr_reg[0]/NET0131  & n3187 ;
  assign n3184 = ~\InstQueueRd_Addr_reg[0]/NET0131  & n965 ;
  assign n3189 = \Flush_reg/NET0131  & \InstAddrPointer_reg[0]/NET0131  ;
  assign n3190 = ~\Flush_reg/NET0131  & ~\InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n3191 = ~n3189 & ~n3190 ;
  assign n3192 = n956 & n3191 ;
  assign n3193 = ~n3184 & ~n3192 ;
  assign n3194 = ~n3188 & n3193 ;
  assign n3195 = ~n3185 & n3194 ;
  assign n3196 = \PhyAddrPointer_reg[10]/NET0131  & n906 ;
  assign n3200 = n1773 & ~n2013 ;
  assign n3201 = ~n1772 & ~n3200 ;
  assign n3202 = ~n2056 & ~n3201 ;
  assign n3203 = n1014 & ~n3202 ;
  assign n3197 = n1316 & ~n2640 ;
  assign n3198 = ~n1014 & ~n2115 ;
  assign n3199 = ~n3197 & n3198 ;
  assign n3204 = ~n906 & ~n3199 ;
  assign n3205 = ~n3203 & n3204 ;
  assign n3206 = ~n3196 & ~n3205 ;
  assign n3207 = n773 & ~n3206 ;
  assign n3208 = \PhyAddrPointer_reg[10]/NET0131  & ~n1852 ;
  assign n3209 = ~\InstAddrPointer_reg[10]/NET0131  & ~n1589 ;
  assign n3210 = ~n1530 & ~n3209 ;
  assign n3211 = ~n2169 & ~n3210 ;
  assign n3212 = n899 & ~n2170 ;
  assign n3213 = ~n3211 & n3212 ;
  assign n3214 = ~n3208 & ~n3213 ;
  assign n3215 = ~n3207 & n3214 ;
  assign n3216 = n929 & ~n3215 ;
  assign n3220 = ~\PhyAddrPointer_reg[10]/NET0131  & ~n2234 ;
  assign n3221 = ~n2235 & ~n3220 ;
  assign n3222 = n2100 & n3221 ;
  assign n3217 = ~\PhyAddrPointer_reg[10]/NET0131  & ~n1876 ;
  assign n3218 = n969 & ~n1877 ;
  assign n3219 = ~n3217 & n3218 ;
  assign n3223 = \rEIP_reg[10]/NET0131  & n1655 ;
  assign n3224 = \PhyAddrPointer_reg[10]/NET0131  & ~n1902 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = ~n3219 & n3225 ;
  assign n3227 = ~n3222 & n3226 ;
  assign n3228 = ~n3216 & n3227 ;
  assign n3229 = \PhyAddrPointer_reg[7]/NET0131  & n906 ;
  assign n3230 = ~n2624 & ~n3229 ;
  assign n3231 = n773 & ~n3230 ;
  assign n3232 = \PhyAddrPointer_reg[7]/NET0131  & ~n1852 ;
  assign n3233 = ~n2606 & ~n3232 ;
  assign n3234 = ~n3231 & n3233 ;
  assign n3235 = n929 & ~n3234 ;
  assign n3239 = \PhyAddrPointer_reg[1]/NET0131  & n1872 ;
  assign n3240 = \PhyAddrPointer_reg[6]/NET0131  & n3239 ;
  assign n3241 = ~\PhyAddrPointer_reg[7]/NET0131  & ~n3240 ;
  assign n3242 = ~n2232 & ~n3241 ;
  assign n3243 = n2100 & n3242 ;
  assign n3236 = ~\PhyAddrPointer_reg[7]/NET0131  & ~n1873 ;
  assign n3237 = n969 & ~n1874 ;
  assign n3238 = ~n3236 & n3237 ;
  assign n3244 = \PhyAddrPointer_reg[7]/NET0131  & ~n1902 ;
  assign n3245 = ~n2597 & ~n3244 ;
  assign n3246 = ~n3238 & n3245 ;
  assign n3247 = ~n3243 & n3246 ;
  assign n3248 = ~n3235 & n3247 ;
  assign n3249 = \PhyAddrPointer_reg[9]/NET0131  & n906 ;
  assign n3250 = ~n2648 & ~n3249 ;
  assign n3251 = n773 & ~n3250 ;
  assign n3252 = \PhyAddrPointer_reg[9]/NET0131  & ~n1852 ;
  assign n3253 = ~n2657 & ~n3252 ;
  assign n3254 = ~n3251 & n3253 ;
  assign n3255 = n929 & ~n3254 ;
  assign n3259 = ~\PhyAddrPointer_reg[9]/NET0131  & ~n2233 ;
  assign n3260 = ~n2234 & ~n3259 ;
  assign n3261 = n2100 & n3260 ;
  assign n3256 = ~\PhyAddrPointer_reg[9]/NET0131  & ~n1875 ;
  assign n3257 = n969 & ~n1876 ;
  assign n3258 = ~n3256 & n3257 ;
  assign n3262 = \PhyAddrPointer_reg[9]/NET0131  & ~n1902 ;
  assign n3263 = ~n2636 & ~n3262 ;
  assign n3264 = ~n3258 & n3263 ;
  assign n3265 = ~n3261 & n3264 ;
  assign n3266 = ~n3255 & n3265 ;
  assign n3277 = \InstAddrPointer_reg[3]/NET0131  & n906 ;
  assign n3278 = ~n1416 & ~n1426 ;
  assign n3279 = ~n1413 & ~n1423 ;
  assign n3280 = ~n3278 & n3279 ;
  assign n3281 = n3278 & ~n3279 ;
  assign n3282 = ~n3280 & ~n3281 ;
  assign n3283 = ~n906 & ~n3282 ;
  assign n3284 = ~n3277 & ~n3283 ;
  assign n3285 = n773 & ~n3284 ;
  assign n3269 = \InstAddrPointer_reg[3]/NET0131  & ~n2887 ;
  assign n3271 = ~n1561 & ~n1563 ;
  assign n3273 = ~n1571 & ~n3271 ;
  assign n3272 = n1571 & n3271 ;
  assign n3274 = n899 & ~n3272 ;
  assign n3275 = ~n3273 & n3274 ;
  assign n3286 = ~\InstAddrPointer_reg[3]/NET0131  & READY_n_pad ;
  assign n3287 = ~READY_n_pad & ~n1415 ;
  assign n3288 = ~n3286 & ~n3287 ;
  assign n3289 = n842 & n3288 ;
  assign n3290 = ~\InstAddrPointer_reg[3]/NET0131  & ~n765 ;
  assign n3291 = n765 & ~n1560 ;
  assign n3292 = ~n3290 & ~n3291 ;
  assign n3293 = ~n740 & n3292 ;
  assign n3294 = ~n3289 & ~n3293 ;
  assign n3295 = ~n3275 & n3294 ;
  assign n3296 = ~n3269 & n3295 ;
  assign n3270 = ~n839 & n1415 ;
  assign n3276 = ~n811 & n1164 ;
  assign n3297 = ~n3270 & ~n3276 ;
  assign n3298 = n3296 & n3297 ;
  assign n3299 = ~n3285 & n3298 ;
  assign n3300 = n929 & ~n3299 ;
  assign n3267 = \rEIP_reg[3]/NET0131  & n1655 ;
  assign n3268 = \InstAddrPointer_reg[3]/NET0131  & n1661 ;
  assign n3301 = ~n3267 & ~n3268 ;
  assign n3302 = ~n3300 & n3301 ;
  assign n3314 = \InstAddrPointer_reg[5]/NET0131  & n906 ;
  assign n3315 = ~n1443 & ~n1449 ;
  assign n3316 = ~n1429 & n3315 ;
  assign n3317 = n1429 & ~n3315 ;
  assign n3318 = ~n3316 & ~n3317 ;
  assign n3319 = ~n906 & ~n3318 ;
  assign n3320 = ~n3314 & ~n3319 ;
  assign n3321 = n773 & ~n3320 ;
  assign n3307 = \InstAddrPointer_reg[5]/NET0131  & ~n2073 ;
  assign n3306 = ~n811 & n1057 ;
  assign n3308 = n766 & n1553 ;
  assign n3322 = ~n3306 & ~n3308 ;
  assign n3323 = ~n3307 & n3322 ;
  assign n3305 = ~n873 & n1442 ;
  assign n3309 = ~n1554 & ~n1575 ;
  assign n3311 = ~n1707 & n3309 ;
  assign n3310 = n1707 & ~n3309 ;
  assign n3312 = n899 & ~n3310 ;
  assign n3313 = ~n3311 & n3312 ;
  assign n3324 = ~n3305 & ~n3313 ;
  assign n3325 = n3323 & n3324 ;
  assign n3326 = ~n3321 & n3325 ;
  assign n3327 = n929 & ~n3326 ;
  assign n3303 = \rEIP_reg[5]/NET0131  & n1655 ;
  assign n3304 = \InstAddrPointer_reg[5]/NET0131  & n1661 ;
  assign n3328 = ~n3303 & ~n3304 ;
  assign n3329 = ~n3327 & n3328 ;
  assign n3330 = \EAX_reg[30]/NET0131  & ~n3181 ;
  assign n3436 = \EAX_reg[26]/NET0131  & \EAX_reg[27]/NET0131  ;
  assign n3437 = n3160 & n3436 ;
  assign n3438 = \EAX_reg[28]/NET0131  & \EAX_reg[29]/NET0131  ;
  assign n3439 = n3437 & n3438 ;
  assign n3440 = ~\EAX_reg[30]/NET0131  & ~n3439 ;
  assign n3441 = \EAX_reg[30]/NET0131  & n3438 ;
  assign n3442 = n3437 & n3441 ;
  assign n3443 = n3132 & ~n3442 ;
  assign n3444 = ~n3440 & n3443 ;
  assign n3430 = ~n847 & ~n3135 ;
  assign n3431 = \EAX_reg[30]/NET0131  & ~n3430 ;
  assign n3335 = \InstQueue_reg[8][5]/NET0131  & n472 ;
  assign n3336 = \InstQueue_reg[5][5]/NET0131  & n488 ;
  assign n3349 = ~n3335 & ~n3336 ;
  assign n3337 = \InstQueue_reg[0][5]/NET0131  & n468 ;
  assign n3338 = \InstQueue_reg[15][5]/NET0131  & n492 ;
  assign n3350 = ~n3337 & ~n3338 ;
  assign n3357 = n3349 & n3350 ;
  assign n3331 = \InstQueue_reg[2][5]/NET0131  & n470 ;
  assign n3332 = \InstQueue_reg[13][5]/NET0131  & n484 ;
  assign n3347 = ~n3331 & ~n3332 ;
  assign n3333 = \InstQueue_reg[1][5]/NET0131  & n465 ;
  assign n3334 = \InstQueue_reg[7][5]/NET0131  & n476 ;
  assign n3348 = ~n3333 & ~n3334 ;
  assign n3358 = n3347 & n3348 ;
  assign n3359 = n3357 & n3358 ;
  assign n3343 = \InstQueue_reg[14][5]/NET0131  & n461 ;
  assign n3344 = \InstQueue_reg[6][5]/NET0131  & n458 ;
  assign n3353 = ~n3343 & ~n3344 ;
  assign n3345 = \InstQueue_reg[3][5]/NET0131  & n522 ;
  assign n3346 = \InstQueue_reg[10][5]/NET0131  & n482 ;
  assign n3354 = ~n3345 & ~n3346 ;
  assign n3355 = n3353 & n3354 ;
  assign n3339 = \InstQueue_reg[4][5]/NET0131  & n474 ;
  assign n3340 = \InstQueue_reg[9][5]/NET0131  & n490 ;
  assign n3351 = ~n3339 & ~n3340 ;
  assign n3341 = \InstQueue_reg[12][5]/NET0131  & n486 ;
  assign n3342 = \InstQueue_reg[11][5]/NET0131  & n454 ;
  assign n3352 = ~n3341 & ~n3342 ;
  assign n3356 = n3351 & n3352 ;
  assign n3360 = n3355 & n3356 ;
  assign n3361 = n3359 & n3360 ;
  assign n3362 = n3129 & ~n3361 ;
  assign n3367 = \InstQueue_reg[8][6]/NET0131  & n472 ;
  assign n3368 = \InstQueue_reg[5][6]/NET0131  & n488 ;
  assign n3381 = ~n3367 & ~n3368 ;
  assign n3369 = \InstQueue_reg[0][6]/NET0131  & n468 ;
  assign n3370 = \InstQueue_reg[15][6]/NET0131  & n492 ;
  assign n3382 = ~n3369 & ~n3370 ;
  assign n3389 = n3381 & n3382 ;
  assign n3363 = \InstQueue_reg[2][6]/NET0131  & n470 ;
  assign n3364 = \InstQueue_reg[13][6]/NET0131  & n484 ;
  assign n3379 = ~n3363 & ~n3364 ;
  assign n3365 = \InstQueue_reg[1][6]/NET0131  & n465 ;
  assign n3366 = \InstQueue_reg[7][6]/NET0131  & n476 ;
  assign n3380 = ~n3365 & ~n3366 ;
  assign n3390 = n3379 & n3380 ;
  assign n3391 = n3389 & n3390 ;
  assign n3375 = \InstQueue_reg[14][6]/NET0131  & n461 ;
  assign n3376 = \InstQueue_reg[6][6]/NET0131  & n458 ;
  assign n3385 = ~n3375 & ~n3376 ;
  assign n3377 = \InstQueue_reg[3][6]/NET0131  & n522 ;
  assign n3378 = \InstQueue_reg[10][6]/NET0131  & n482 ;
  assign n3386 = ~n3377 & ~n3378 ;
  assign n3387 = n3385 & n3386 ;
  assign n3371 = \InstQueue_reg[4][6]/NET0131  & n474 ;
  assign n3372 = \InstQueue_reg[9][6]/NET0131  & n490 ;
  assign n3383 = ~n3371 & ~n3372 ;
  assign n3373 = \InstQueue_reg[12][6]/NET0131  & n486 ;
  assign n3374 = \InstQueue_reg[11][6]/NET0131  & n454 ;
  assign n3384 = ~n3373 & ~n3374 ;
  assign n3388 = n3383 & n3384 ;
  assign n3392 = n3387 & n3388 ;
  assign n3393 = n3391 & n3392 ;
  assign n3394 = n3362 & ~n3393 ;
  assign n3399 = \InstQueue_reg[14][7]/NET0131  & n461 ;
  assign n3400 = \InstQueue_reg[5][7]/NET0131  & n488 ;
  assign n3413 = ~n3399 & ~n3400 ;
  assign n3401 = \InstQueue_reg[0][7]/NET0131  & n468 ;
  assign n3402 = \InstQueue_reg[2][7]/NET0131  & n470 ;
  assign n3414 = ~n3401 & ~n3402 ;
  assign n3421 = n3413 & n3414 ;
  assign n3395 = \InstQueue_reg[10][7]/NET0131  & n482 ;
  assign n3396 = \InstQueue_reg[13][7]/NET0131  & n484 ;
  assign n3411 = ~n3395 & ~n3396 ;
  assign n3397 = \InstQueue_reg[9][7]/NET0131  & n490 ;
  assign n3398 = \InstQueue_reg[7][7]/NET0131  & n476 ;
  assign n3412 = ~n3397 & ~n3398 ;
  assign n3422 = n3411 & n3412 ;
  assign n3423 = n3421 & n3422 ;
  assign n3407 = \InstQueue_reg[8][7]/NET0131  & n472 ;
  assign n3408 = \InstQueue_reg[6][7]/NET0131  & n458 ;
  assign n3417 = ~n3407 & ~n3408 ;
  assign n3409 = \InstQueue_reg[3][7]/NET0131  & n522 ;
  assign n3410 = \InstQueue_reg[4][7]/NET0131  & n474 ;
  assign n3418 = ~n3409 & ~n3410 ;
  assign n3419 = n3417 & n3418 ;
  assign n3403 = \InstQueue_reg[12][7]/NET0131  & n486 ;
  assign n3404 = \InstQueue_reg[1][7]/NET0131  & n465 ;
  assign n3415 = ~n3403 & ~n3404 ;
  assign n3405 = \InstQueue_reg[15][7]/NET0131  & n492 ;
  assign n3406 = \InstQueue_reg[11][7]/NET0131  & n454 ;
  assign n3416 = ~n3405 & ~n3406 ;
  assign n3420 = n3415 & n3416 ;
  assign n3424 = n3419 & n3420 ;
  assign n3425 = n3423 & n3424 ;
  assign n3426 = n3394 & ~n3425 ;
  assign n3427 = ~n3394 & n3425 ;
  assign n3428 = ~n3426 & ~n3427 ;
  assign n3429 = n2937 & n3428 ;
  assign n3432 = \Datai[14]_pad  & n782 ;
  assign n3433 = \Datai[30]_pad  & n840 ;
  assign n3434 = ~n3432 & ~n3433 ;
  assign n3435 = n846 & ~n3434 ;
  assign n3445 = ~n3429 & ~n3435 ;
  assign n3446 = ~n3431 & n3445 ;
  assign n3447 = ~n3444 & n3446 ;
  assign n3448 = n929 & ~n3447 ;
  assign n3449 = ~n3330 & ~n3448 ;
  assign n3451 = \EAX_reg[31]/NET0131  & n3442 ;
  assign n3450 = ~\EAX_reg[31]/NET0131  & ~n3442 ;
  assign n3452 = n3132 & ~n3450 ;
  assign n3453 = ~n3451 & n3452 ;
  assign n3456 = \EAX_reg[31]/NET0131  & ~n3430 ;
  assign n3454 = n2937 & n3426 ;
  assign n3455 = \Datai[31]_pad  & n2607 ;
  assign n3457 = ~n3454 & ~n3455 ;
  assign n3458 = ~n3456 & n3457 ;
  assign n3459 = ~n3453 & n3458 ;
  assign n3460 = n929 & ~n3459 ;
  assign n3461 = \EAX_reg[31]/NET0131  & ~n3181 ;
  assign n3462 = ~n3460 & ~n3461 ;
  assign n3468 = \EBX_reg[0]/NET0131  & \EBX_reg[1]/NET0131  ;
  assign n3469 = \EBX_reg[2]/NET0131  & n3468 ;
  assign n3470 = \EBX_reg[3]/NET0131  & n3469 ;
  assign n3471 = \EBX_reg[4]/NET0131  & n3470 ;
  assign n3472 = \EBX_reg[5]/NET0131  & n3471 ;
  assign n3473 = \EBX_reg[6]/NET0131  & n3472 ;
  assign n3474 = \EBX_reg[7]/NET0131  & n3473 ;
  assign n3475 = \EBX_reg[8]/NET0131  & n3474 ;
  assign n3476 = \EBX_reg[9]/NET0131  & n3475 ;
  assign n3477 = \EBX_reg[10]/NET0131  & n3476 ;
  assign n3478 = \EBX_reg[11]/NET0131  & n3477 ;
  assign n3479 = \EBX_reg[12]/NET0131  & n3478 ;
  assign n3480 = \EBX_reg[13]/NET0131  & n3479 ;
  assign n3481 = \EBX_reg[14]/NET0131  & n3480 ;
  assign n3482 = \EBX_reg[15]/NET0131  & n3481 ;
  assign n3483 = \EBX_reg[16]/NET0131  & n3482 ;
  assign n3484 = \EBX_reg[17]/NET0131  & n3483 ;
  assign n3485 = \EBX_reg[18]/NET0131  & n3484 ;
  assign n3486 = \EBX_reg[19]/NET0131  & n3485 ;
  assign n3487 = \EBX_reg[20]/NET0131  & \EBX_reg[21]/NET0131  ;
  assign n3488 = \EBX_reg[22]/NET0131  & \EBX_reg[23]/NET0131  ;
  assign n3489 = n3487 & n3488 ;
  assign n3490 = n3486 & n3489 ;
  assign n3491 = \EBX_reg[24]/NET0131  & \EBX_reg[25]/NET0131  ;
  assign n3492 = n3490 & n3491 ;
  assign n3493 = \EBX_reg[26]/NET0131  & \EBX_reg[27]/NET0131  ;
  assign n3494 = n3492 & n3493 ;
  assign n3495 = \EBX_reg[28]/NET0131  & \EBX_reg[29]/NET0131  ;
  assign n3496 = \EBX_reg[30]/NET0131  & n3495 ;
  assign n3497 = n3494 & n3496 ;
  assign n3499 = \EBX_reg[31]/NET0131  & n3497 ;
  assign n3498 = ~\EBX_reg[31]/NET0131  & ~n3497 ;
  assign n3500 = n797 & ~n3498 ;
  assign n3501 = ~n3499 & n3500 ;
  assign n3463 = n735 & n765 ;
  assign n3464 = ~n735 & n797 ;
  assign n3465 = ~n3463 & ~n3464 ;
  assign n3466 = \EBX_reg[31]/NET0131  & n3465 ;
  assign n3467 = n3426 & n3463 ;
  assign n3502 = ~n3466 & ~n3467 ;
  assign n3503 = ~n3501 & n3502 ;
  assign n3504 = n929 & ~n3503 ;
  assign n3505 = \EBX_reg[31]/NET0131  & ~n3181 ;
  assign n3506 = ~n3504 & ~n3505 ;
  assign n3508 = ~n892 & n929 ;
  assign n3509 = \InstAddrPointer_reg[31]/NET0131  & ~n1234 ;
  assign n3510 = ~\InstAddrPointer_reg[1]/NET0131  & ~\InstAddrPointer_reg[31]/NET0131  ;
  assign n3511 = ~n3509 & ~n3510 ;
  assign n3512 = n3189 & n3511 ;
  assign n3513 = ~n957 & ~n3512 ;
  assign n3514 = n956 & ~n3513 ;
  assign n3507 = \InstQueueRd_Addr_reg[2]/NET0131  & n3187 ;
  assign n3515 = n883 & n965 ;
  assign n3516 = ~n3507 & ~n3515 ;
  assign n3517 = ~n3514 & n3516 ;
  assign n3518 = ~n3508 & n3517 ;
  assign n3519 = \PhyAddrPointer_reg[4]/NET0131  & n906 ;
  assign n3520 = ~n2873 & ~n3519 ;
  assign n3521 = n773 & ~n3520 ;
  assign n3522 = \PhyAddrPointer_reg[4]/NET0131  & ~n1852 ;
  assign n3523 = ~n2881 & ~n3522 ;
  assign n3524 = ~n3521 & n3523 ;
  assign n3525 = n929 & ~n3524 ;
  assign n3530 = \PhyAddrPointer_reg[1]/NET0131  & \PhyAddrPointer_reg[2]/NET0131  ;
  assign n3531 = \PhyAddrPointer_reg[3]/NET0131  & n3530 ;
  assign n3532 = ~\PhyAddrPointer_reg[4]/NET0131  & ~n3531 ;
  assign n3533 = \PhyAddrPointer_reg[4]/NET0131  & n3531 ;
  assign n3534 = ~n3532 & ~n3533 ;
  assign n3535 = n2100 & n3534 ;
  assign n3529 = \PhyAddrPointer_reg[4]/NET0131  & ~n1902 ;
  assign n3526 = ~\PhyAddrPointer_reg[4]/NET0131  & ~n1870 ;
  assign n3527 = ~n1871 & ~n3526 ;
  assign n3528 = n969 & n3527 ;
  assign n3536 = ~n2864 & ~n3528 ;
  assign n3537 = ~n3529 & n3536 ;
  assign n3538 = ~n3535 & n3537 ;
  assign n3539 = ~n3525 & n3538 ;
  assign n3549 = ~n873 & n1412 ;
  assign n3542 = ~n900 & n2887 ;
  assign n3543 = \InstAddrPointer_reg[2]/NET0131  & ~n3542 ;
  assign n3548 = ~n811 & n1199 ;
  assign n3550 = \InstAddrPointer_reg[2]/NET0131  & n906 ;
  assign n3551 = ~n1413 & ~n1418 ;
  assign n3552 = ~n1422 & ~n3551 ;
  assign n3553 = n1422 & n3551 ;
  assign n3554 = ~n3552 & ~n3553 ;
  assign n3555 = ~n906 & ~n3554 ;
  assign n3556 = ~n3550 & ~n3555 ;
  assign n3557 = n773 & ~n3556 ;
  assign n3544 = ~\InstAddrPointer_reg[2]/NET0131  & ~n765 ;
  assign n3545 = n765 & n1199 ;
  assign n3546 = ~n3544 & ~n3545 ;
  assign n3547 = ~n740 & n3546 ;
  assign n3558 = ~n1200 & ~n1273 ;
  assign n3560 = n1569 & ~n3558 ;
  assign n3559 = ~n1569 & n3558 ;
  assign n3561 = n899 & ~n3559 ;
  assign n3562 = ~n3560 & n3561 ;
  assign n3563 = ~n3547 & ~n3562 ;
  assign n3564 = ~n3557 & n3563 ;
  assign n3565 = ~n3548 & n3564 ;
  assign n3566 = ~n3543 & n3565 ;
  assign n3567 = ~n3549 & n3566 ;
  assign n3568 = n929 & ~n3567 ;
  assign n3540 = \rEIP_reg[2]/NET0131  & n1655 ;
  assign n3541 = \InstAddrPointer_reg[2]/NET0131  & n1661 ;
  assign n3569 = ~n3540 & ~n3541 ;
  assign n3570 = ~n3568 & n3569 ;
  assign n3578 = ~\InstAddrPointer_reg[0]/NET0131  & n811 ;
  assign n3579 = \InstAddrPointer_reg[0]/NET0131  & ~n911 ;
  assign n3580 = n789 & n3579 ;
  assign n3581 = ~n3578 & ~n3580 ;
  assign n3583 = ~\InstAddrPointer_reg[0]/NET0131  & ~n765 ;
  assign n3584 = \InstAddrPointer_reg[0]/NET0131  & n765 ;
  assign n3585 = ~n3583 & ~n3584 ;
  assign n3586 = ~n740 & n3585 ;
  assign n3573 = \InstAddrPointer_reg[0]/NET0131  & n906 ;
  assign n3574 = ~n1268 & ~n1567 ;
  assign n3575 = ~n906 & ~n3574 ;
  assign n3576 = ~n3573 & ~n3575 ;
  assign n3577 = n773 & ~n3576 ;
  assign n3582 = n899 & n3574 ;
  assign n3587 = ~n3577 & ~n3582 ;
  assign n3588 = ~n3586 & n3587 ;
  assign n3589 = ~n3581 & n3588 ;
  assign n3590 = n929 & ~n3589 ;
  assign n3571 = \rEIP_reg[0]/NET0131  & n1655 ;
  assign n3572 = \InstAddrPointer_reg[0]/NET0131  & n1661 ;
  assign n3591 = ~n3571 & ~n3572 ;
  assign n3592 = ~n3590 & n3591 ;
  assign n3595 = ~n910 & n1816 ;
  assign n3596 = \InstAddrPointer_reg[1]/NET0131  & ~n3595 ;
  assign n3614 = ~n812 & n1234 ;
  assign n3594 = ~\InstAddrPointer_reg[1]/NET0131  & ~n873 ;
  assign n3599 = ~n1235 & ~n1566 ;
  assign n3600 = ~n1268 & n3599 ;
  assign n3597 = ~n1236 & ~n1419 ;
  assign n3598 = n1268 & ~n3597 ;
  assign n3601 = ~n1014 & ~n3598 ;
  assign n3602 = ~n3600 & n3601 ;
  assign n3604 = n1420 & n3597 ;
  assign n3603 = ~n1420 & ~n3597 ;
  assign n3605 = n1014 & ~n3603 ;
  assign n3606 = ~n3604 & n3605 ;
  assign n3607 = ~n3602 & ~n3606 ;
  assign n3608 = n907 & ~n3607 ;
  assign n3609 = ~n1567 & ~n3599 ;
  assign n3610 = n1567 & ~n3597 ;
  assign n3611 = ~n3609 & ~n3610 ;
  assign n3612 = n899 & n3611 ;
  assign n3613 = ~n3608 & ~n3612 ;
  assign n3615 = ~n3594 & n3613 ;
  assign n3616 = ~n3614 & n3615 ;
  assign n3617 = ~n3596 & n3616 ;
  assign n3618 = n929 & ~n3617 ;
  assign n3593 = \rEIP_reg[1]/NET0131  & n1655 ;
  assign n3619 = \InstAddrPointer_reg[1]/NET0131  & n1661 ;
  assign n3620 = ~n3593 & ~n3619 ;
  assign n3621 = ~n3618 & n3620 ;
  assign n3623 = ~n854 & n929 ;
  assign n3624 = ~\Flush_reg/NET0131  & \InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n3625 = n3189 & ~n3511 ;
  assign n3626 = ~n3624 & ~n3625 ;
  assign n3627 = n956 & ~n3626 ;
  assign n3622 = \InstQueueRd_Addr_reg[1]/NET0131  & n3187 ;
  assign n3628 = ~n822 & n965 ;
  assign n3629 = ~n3622 & ~n3628 ;
  assign n3630 = ~n3627 & n3629 ;
  assign n3631 = ~n3623 & n3630 ;
  assign n3632 = \EAX_reg[26]/NET0131  & ~n3181 ;
  assign n3636 = ~\EAX_reg[26]/NET0131  & ~n3160 ;
  assign n3637 = n3162 & ~n3636 ;
  assign n3638 = \EAX_reg[26]/NET0131  & n3135 ;
  assign n3639 = \EAX_reg[26]/NET0131  & ~n846 ;
  assign n3643 = \Datai[10]_pad  & n846 ;
  assign n3644 = ~n3639 & ~n3643 ;
  assign n3645 = n782 & ~n3644 ;
  assign n3633 = ~n3064 & n3095 ;
  assign n3634 = ~n3096 & ~n3633 ;
  assign n3635 = n2937 & n3634 ;
  assign n3640 = \Datai[26]_pad  & n846 ;
  assign n3641 = ~n3639 & ~n3640 ;
  assign n3642 = n840 & ~n3641 ;
  assign n3646 = ~n3635 & ~n3642 ;
  assign n3647 = ~n3645 & n3646 ;
  assign n3648 = ~n3638 & n3647 ;
  assign n3649 = ~n3637 & n3648 ;
  assign n3650 = n929 & ~n3649 ;
  assign n3651 = ~n3632 & ~n3650 ;
  assign n3652 = ~n937 & ~n1655 ;
  assign n3653 = ~n967 & n1901 ;
  assign n3654 = n2098 & n3653 ;
  assign n3655 = n3652 & n3654 ;
  assign n3656 = \uWord_reg[12]/NET0131  & ~n3655 ;
  assign n3666 = ~\EAX_reg[13]/NET0131  & ~\EAX_reg[14]/NET0131  ;
  assign n3667 = ~\EAX_reg[15]/NET0131  & ~\EAX_reg[1]/NET0131  ;
  assign n3674 = n3666 & n3667 ;
  assign n3664 = ~\EAX_reg[0]/NET0131  & ~\EAX_reg[10]/NET0131  ;
  assign n3665 = ~\EAX_reg[11]/NET0131  & ~\EAX_reg[12]/NET0131  ;
  assign n3675 = n3664 & n3665 ;
  assign n3676 = n3674 & n3675 ;
  assign n3670 = ~\EAX_reg[6]/NET0131  & ~\EAX_reg[7]/NET0131  ;
  assign n3671 = ~\EAX_reg[8]/NET0131  & ~\EAX_reg[9]/NET0131  ;
  assign n3672 = n3670 & n3671 ;
  assign n3668 = ~\EAX_reg[2]/NET0131  & ~\EAX_reg[3]/NET0131  ;
  assign n3669 = ~\EAX_reg[4]/NET0131  & ~\EAX_reg[5]/NET0131  ;
  assign n3673 = n3668 & n3669 ;
  assign n3677 = n3672 & n3673 ;
  assign n3678 = n3676 & n3677 ;
  assign n3679 = \EAX_reg[31]/NET0131  & ~n3678 ;
  assign n3680 = \EAX_reg[16]/NET0131  & n3679 ;
  assign n3681 = \EAX_reg[17]/NET0131  & n3680 ;
  assign n3682 = \EAX_reg[18]/NET0131  & n3681 ;
  assign n3683 = n3156 & n3682 ;
  assign n3684 = n3158 & n3683 ;
  assign n3685 = \EAX_reg[25]/NET0131  & n3684 ;
  assign n3686 = n3436 & n3685 ;
  assign n3687 = ~\EAX_reg[28]/NET0131  & ~n3686 ;
  assign n3688 = \EAX_reg[28]/NET0131  & n3686 ;
  assign n3689 = ~n3687 & ~n3688 ;
  assign n3690 = n783 & n3689 ;
  assign n3691 = ~n834 & n3690 ;
  assign n3657 = \Datai[12]_pad  & n846 ;
  assign n3658 = n782 & n3657 ;
  assign n3659 = READY_n_pad & n782 ;
  assign n3660 = n782 & ~n834 ;
  assign n3661 = ~n923 & ~n3660 ;
  assign n3662 = ~n3659 & ~n3661 ;
  assign n3663 = \uWord_reg[12]/NET0131  & ~n3662 ;
  assign n3692 = ~n3658 & ~n3663 ;
  assign n3693 = ~n3691 & n3692 ;
  assign n3694 = n929 & ~n3693 ;
  assign n3695 = ~n3656 & ~n3694 ;
  assign n3696 = \EBX_reg[28]/NET0131  & n3494 ;
  assign n3697 = \EBX_reg[29]/NET0131  & n3696 ;
  assign n3698 = ~\EBX_reg[30]/NET0131  & ~n3697 ;
  assign n3699 = n797 & ~n3497 ;
  assign n3700 = ~n3698 & n3699 ;
  assign n3701 = \EBX_reg[30]/NET0131  & n3465 ;
  assign n3702 = n3428 & n3463 ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = ~n3700 & n3703 ;
  assign n3705 = n929 & ~n3704 ;
  assign n3706 = \EBX_reg[30]/NET0131  & ~n3181 ;
  assign n3707 = ~n3705 & ~n3706 ;
  assign n3711 = \PhyAddrPointer_reg[3]/NET0131  & n906 ;
  assign n3712 = ~n3283 & ~n3711 ;
  assign n3713 = n773 & ~n3712 ;
  assign n3714 = \PhyAddrPointer_reg[3]/NET0131  & ~n1852 ;
  assign n3715 = ~n3275 & ~n3714 ;
  assign n3716 = ~n3713 & n3715 ;
  assign n3717 = n929 & ~n3716 ;
  assign n3718 = \PhyAddrPointer_reg[3]/NET0131  & ~n1902 ;
  assign n3720 = \PhyAddrPointer_reg[2]/NET0131  & ~n1906 ;
  assign n3721 = ~\PhyAddrPointer_reg[3]/NET0131  & ~n3720 ;
  assign n3719 = n1870 & ~n1906 ;
  assign n3722 = n933 & ~n3719 ;
  assign n3723 = ~n3721 & n3722 ;
  assign n3708 = ~\PhyAddrPointer_reg[3]/NET0131  & ~n3530 ;
  assign n3709 = ~n3531 & ~n3708 ;
  assign n3710 = n1867 & n3709 ;
  assign n3724 = ~n3267 & ~n3710 ;
  assign n3725 = ~n3723 & n3724 ;
  assign n3726 = ~n3718 & n3725 ;
  assign n3727 = ~n3717 & n3726 ;
  assign n3728 = \PhyAddrPointer_reg[5]/NET0131  & n906 ;
  assign n3729 = ~n3319 & ~n3728 ;
  assign n3730 = n773 & ~n3729 ;
  assign n3731 = \PhyAddrPointer_reg[5]/NET0131  & ~n1852 ;
  assign n3732 = ~n3313 & ~n3731 ;
  assign n3733 = ~n3730 & n3732 ;
  assign n3734 = n929 & ~n3733 ;
  assign n3738 = ~\PhyAddrPointer_reg[5]/NET0131  & ~n3533 ;
  assign n3739 = ~n3239 & ~n3738 ;
  assign n3740 = n2100 & n3739 ;
  assign n3741 = \PhyAddrPointer_reg[5]/NET0131  & ~n1902 ;
  assign n3735 = ~\PhyAddrPointer_reg[5]/NET0131  & ~n1871 ;
  assign n3736 = n969 & ~n1872 ;
  assign n3737 = ~n3735 & n3736 ;
  assign n3742 = ~n3303 & ~n3737 ;
  assign n3743 = ~n3741 & n3742 ;
  assign n3744 = ~n3740 & n3743 ;
  assign n3745 = ~n3734 & n3744 ;
  assign n3749 = \PhyAddrPointer_reg[6]/NET0131  & n906 ;
  assign n3750 = ~n2915 & ~n3749 ;
  assign n3751 = n773 & ~n3750 ;
  assign n3752 = \PhyAddrPointer_reg[6]/NET0131  & ~n1852 ;
  assign n3753 = ~n2927 & ~n3752 ;
  assign n3754 = ~n3751 & n3753 ;
  assign n3755 = n929 & ~n3754 ;
  assign n3746 = ~\PhyAddrPointer_reg[6]/NET0131  & ~n3239 ;
  assign n3747 = ~n3240 & ~n3746 ;
  assign n3759 = ~\DataWidth_reg[1]/NET0131  & ~n3747 ;
  assign n3756 = ~\PhyAddrPointer_reg[6]/NET0131  & ~n1872 ;
  assign n3757 = ~n1873 & ~n3756 ;
  assign n3758 = \DataWidth_reg[1]/NET0131  & ~n3757 ;
  assign n3760 = n933 & ~n3758 ;
  assign n3761 = ~n3759 & n3760 ;
  assign n3748 = n1867 & n3747 ;
  assign n3762 = \PhyAddrPointer_reg[6]/NET0131  & ~n1902 ;
  assign n3763 = ~n2902 & ~n3762 ;
  assign n3764 = ~n3748 & n3763 ;
  assign n3765 = ~n3761 & n3764 ;
  assign n3766 = ~n3755 & n3765 ;
  assign n3768 = ~n881 & n929 ;
  assign n3769 = ~\Flush_reg/NET0131  & \InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n3770 = ~n3512 & ~n3769 ;
  assign n3771 = n956 & ~n3770 ;
  assign n3767 = \InstQueueRd_Addr_reg[3]/NET0131  & n3187 ;
  assign n3772 = ~n868 & n965 ;
  assign n3773 = ~n3767 & ~n3772 ;
  assign n3774 = ~n3771 & n3773 ;
  assign n3775 = ~n3768 & n3774 ;
  assign n3787 = \EAX_reg[28]/NET0131  & n3437 ;
  assign n3788 = ~\EAX_reg[29]/NET0131  & ~n3787 ;
  assign n3789 = n3132 & ~n3439 ;
  assign n3790 = ~n3788 & n3789 ;
  assign n3777 = n840 & ~n846 ;
  assign n3778 = ~n3135 & ~n3777 ;
  assign n3779 = \EAX_reg[29]/NET0131  & ~n3778 ;
  assign n3780 = ~n3362 & n3393 ;
  assign n3781 = ~n3394 & ~n3780 ;
  assign n3782 = n2937 & n3781 ;
  assign n3776 = \Datai[29]_pad  & n2607 ;
  assign n3783 = \EAX_reg[29]/NET0131  & ~n846 ;
  assign n3784 = \Datai[13]_pad  & n846 ;
  assign n3785 = ~n3783 & ~n3784 ;
  assign n3786 = n782 & ~n3785 ;
  assign n3791 = ~n3776 & ~n3786 ;
  assign n3792 = ~n3782 & n3791 ;
  assign n3793 = ~n3779 & n3792 ;
  assign n3794 = ~n3790 & n3793 ;
  assign n3795 = n929 & ~n3794 ;
  assign n3796 = \EAX_reg[29]/NET0131  & ~n3181 ;
  assign n3797 = ~n3795 & ~n3796 ;
  assign n3799 = ~\EBX_reg[26]/NET0131  & ~n3492 ;
  assign n3800 = \EBX_reg[26]/NET0131  & n3492 ;
  assign n3801 = n797 & ~n3800 ;
  assign n3802 = ~n3799 & n3801 ;
  assign n3798 = n3463 & n3634 ;
  assign n3803 = \EBX_reg[26]/NET0131  & n3465 ;
  assign n3804 = ~n3798 & ~n3803 ;
  assign n3805 = ~n3802 & n3804 ;
  assign n3806 = n929 & ~n3805 ;
  assign n3807 = \EBX_reg[26]/NET0131  & ~n3181 ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3811 = \EAX_reg[23]/NET0131  & n3683 ;
  assign n3812 = ~\EAX_reg[24]/NET0131  & ~n3811 ;
  assign n3813 = n783 & ~n3684 ;
  assign n3814 = ~n3812 & n3813 ;
  assign n3815 = n856 & n3814 ;
  assign n3816 = \Datao[24]_pad  & ~n857 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = n929 & ~n3817 ;
  assign n3809 = ~\State2_reg[0]/NET0131  & n955 ;
  assign n3810 = \uWord_reg[8]/NET0131  & n3809 ;
  assign n3819 = \State2_reg[2]/NET0131  & ~n1867 ;
  assign n3820 = ~n1657 & ~n3819 ;
  assign n3821 = ~n956 & ~n3820 ;
  assign n3822 = \Datao[24]_pad  & ~n3821 ;
  assign n3823 = ~n3810 & ~n3822 ;
  assign n3824 = ~n3818 & n3823 ;
  assign n3826 = n828 & n835 ;
  assign n3827 = n837 & ~n3826 ;
  assign n3828 = ~n828 & ~n3689 ;
  assign n3829 = n923 & ~n3828 ;
  assign n3830 = n3827 & ~n3829 ;
  assign n3831 = \Datao[28]_pad  & ~n3830 ;
  assign n3832 = n856 & n3690 ;
  assign n3833 = ~n3831 & ~n3832 ;
  assign n3834 = n929 & ~n3833 ;
  assign n3825 = \uWord_reg[12]/NET0131  & n3809 ;
  assign n3835 = \Datao[28]_pad  & ~n3821 ;
  assign n3836 = ~n3825 & ~n3835 ;
  assign n3837 = ~n3834 & n3836 ;
  assign n3838 = n929 & ~n3662 ;
  assign n3839 = n3655 & ~n3838 ;
  assign n3840 = \uWord_reg[8]/NET0131  & ~n3839 ;
  assign n3841 = \Datai[8]_pad  & ~READY_n_pad ;
  assign n3842 = n782 & n3841 ;
  assign n3843 = ~n3814 & ~n3842 ;
  assign n3844 = ~n834 & n929 ;
  assign n3845 = ~n3843 & n3844 ;
  assign n3846 = ~n3840 & ~n3845 ;
  assign n3847 = \EBX_reg[29]/NET0131  & ~n3181 ;
  assign n3850 = ~\EBX_reg[29]/NET0131  & ~n3696 ;
  assign n3851 = n797 & ~n3697 ;
  assign n3852 = ~n3850 & n3851 ;
  assign n3848 = \EBX_reg[29]/NET0131  & n3465 ;
  assign n3849 = n3463 & n3781 ;
  assign n3853 = ~n3848 & ~n3849 ;
  assign n3854 = ~n3852 & n3853 ;
  assign n3855 = n929 & ~n3854 ;
  assign n3856 = ~n3847 & ~n3855 ;
  assign n3869 = \InstQueueWr_Addr_reg[0]/NET0131  & ~\InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3870 = \InstQueueWr_Addr_reg[2]/NET0131  & n3869 ;
  assign n3871 = \InstQueueWr_Addr_reg[3]/NET0131  & n3870 ;
  assign n3874 = ~\Datai[13]_pad  & ~\Datai[14]_pad  ;
  assign n3875 = ~\Datai[15]_pad  & ~\Datai[1]_pad  ;
  assign n3882 = n3874 & n3875 ;
  assign n3872 = ~\Datai[0]_pad  & ~\Datai[10]_pad  ;
  assign n3873 = ~\Datai[11]_pad  & ~\Datai[12]_pad  ;
  assign n3883 = n3872 & n3873 ;
  assign n3884 = n3882 & n3883 ;
  assign n3878 = ~\Datai[6]_pad  & ~\Datai[7]_pad  ;
  assign n3879 = ~\Datai[8]_pad  & ~\Datai[9]_pad  ;
  assign n3880 = n3878 & n3879 ;
  assign n3876 = ~\Datai[2]_pad  & ~\Datai[3]_pad  ;
  assign n3877 = ~\Datai[4]_pad  & ~\Datai[5]_pad  ;
  assign n3881 = n3876 & n3877 ;
  assign n3885 = n3880 & n3881 ;
  assign n3886 = n3884 & n3885 ;
  assign n3889 = ~\Datai[20]_pad  & ~\Datai[21]_pad  ;
  assign n3890 = ~\Datai[22]_pad  & ~\Datai[23]_pad  ;
  assign n3891 = n3889 & n3890 ;
  assign n3887 = ~\Datai[16]_pad  & ~\Datai[17]_pad  ;
  assign n3888 = ~\Datai[18]_pad  & ~\Datai[19]_pad  ;
  assign n3892 = n3887 & n3888 ;
  assign n3893 = n3891 & n3892 ;
  assign n3894 = n3886 & n3893 ;
  assign n3895 = \Datai[31]_pad  & ~n3894 ;
  assign n3896 = \Datai[24]_pad  & n3895 ;
  assign n3897 = \Datai[25]_pad  & n3896 ;
  assign n3898 = \Datai[26]_pad  & n3897 ;
  assign n3899 = \Datai[27]_pad  & n3898 ;
  assign n3900 = \Datai[28]_pad  & n3899 ;
  assign n3901 = ~\Datai[28]_pad  & ~n3899 ;
  assign n3902 = ~n3900 & ~n3901 ;
  assign n3903 = n3871 & n3902 ;
  assign n3904 = \Datai[31]_pad  & ~n3886 ;
  assign n3905 = \Datai[16]_pad  & n3904 ;
  assign n3906 = \Datai[17]_pad  & n3905 ;
  assign n3907 = \Datai[18]_pad  & n3906 ;
  assign n3908 = \Datai[19]_pad  & n3907 ;
  assign n3909 = ~\Datai[20]_pad  & ~n3908 ;
  assign n3910 = \Datai[20]_pad  & n3908 ;
  assign n3911 = ~n3909 & ~n3910 ;
  assign n3912 = ~\InstQueueWr_Addr_reg[0]/NET0131  & \InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3913 = \InstQueueWr_Addr_reg[2]/NET0131  & n3912 ;
  assign n3914 = \InstQueueWr_Addr_reg[3]/NET0131  & n3913 ;
  assign n3915 = n3911 & n3914 ;
  assign n3916 = ~n3903 & ~n3915 ;
  assign n3917 = \DataWidth_reg[1]/NET0131  & ~n3916 ;
  assign n3857 = ~\InstQueueWr_Addr_reg[0]/NET0131  & ~\InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3858 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3857 ;
  assign n3859 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3858 ;
  assign n3860 = \InstQueueWr_Addr_reg[0]/NET0131  & \InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3861 = \InstQueueWr_Addr_reg[2]/NET0131  & n3860 ;
  assign n3862 = \InstQueueWr_Addr_reg[3]/NET0131  & n3861 ;
  assign n3863 = ~n3859 & ~n3862 ;
  assign n3864 = \Datai[4]_pad  & ~n3863 ;
  assign n3865 = \InstQueue_reg[0][4]/NET0131  & ~n3859 ;
  assign n3866 = ~n3862 & n3865 ;
  assign n3867 = ~n3864 & ~n3866 ;
  assign n3918 = ~n3871 & ~n3914 ;
  assign n3919 = \DataWidth_reg[1]/NET0131  & ~n3918 ;
  assign n3920 = ~n3867 & ~n3919 ;
  assign n3921 = ~n3917 & ~n3920 ;
  assign n3922 = n933 & ~n3921 ;
  assign n3923 = ~n668 & n3859 ;
  assign n3924 = ~n3865 & ~n3923 ;
  assign n3925 = n965 & ~n3924 ;
  assign n3868 = n1867 & ~n3867 ;
  assign n3926 = ~n936 & ~n967 ;
  assign n3927 = ~n955 & ~n1655 ;
  assign n3928 = ~n929 & n3927 ;
  assign n3929 = n3926 & n3928 ;
  assign n3930 = \InstQueue_reg[0][4]/NET0131  & ~n3929 ;
  assign n3931 = ~n3868 & ~n3930 ;
  assign n3932 = ~n3925 & n3931 ;
  assign n3933 = ~n3922 & n3932 ;
  assign n3944 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3861 ;
  assign n3945 = n3902 & n3944 ;
  assign n3946 = \InstQueueWr_Addr_reg[3]/NET0131  & n3858 ;
  assign n3947 = n3911 & n3946 ;
  assign n3948 = ~n3945 & ~n3947 ;
  assign n3949 = \DataWidth_reg[1]/NET0131  & ~n3948 ;
  assign n3934 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3912 ;
  assign n3935 = \InstQueueWr_Addr_reg[3]/NET0131  & n3934 ;
  assign n3936 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3869 ;
  assign n3937 = \InstQueueWr_Addr_reg[3]/NET0131  & n3936 ;
  assign n3938 = ~n3935 & ~n3937 ;
  assign n3939 = \Datai[4]_pad  & ~n3938 ;
  assign n3940 = \InstQueue_reg[10][4]/NET0131  & ~n3935 ;
  assign n3941 = ~n3937 & n3940 ;
  assign n3942 = ~n3939 & ~n3941 ;
  assign n3950 = ~n3944 & ~n3946 ;
  assign n3951 = \DataWidth_reg[1]/NET0131  & ~n3950 ;
  assign n3952 = ~n3942 & ~n3951 ;
  assign n3953 = ~n3949 & ~n3952 ;
  assign n3954 = n933 & ~n3953 ;
  assign n3955 = ~n668 & n3935 ;
  assign n3956 = ~n3940 & ~n3955 ;
  assign n3957 = n965 & ~n3956 ;
  assign n3943 = n1867 & ~n3942 ;
  assign n3958 = \InstQueue_reg[10][4]/NET0131  & ~n3929 ;
  assign n3959 = ~n3943 & ~n3958 ;
  assign n3960 = ~n3957 & n3959 ;
  assign n3961 = ~n3954 & n3960 ;
  assign n3970 = n3902 & n3946 ;
  assign n3971 = n3911 & n3937 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n3973 = \DataWidth_reg[1]/NET0131  & ~n3972 ;
  assign n3962 = ~\InstQueueWr_Addr_reg[2]/NET0131  & n3860 ;
  assign n3963 = \InstQueueWr_Addr_reg[3]/NET0131  & n3962 ;
  assign n3964 = ~n3935 & ~n3963 ;
  assign n3965 = \Datai[4]_pad  & ~n3964 ;
  assign n3966 = \InstQueue_reg[11][4]/NET0131  & ~n3963 ;
  assign n3967 = ~n3935 & n3966 ;
  assign n3968 = ~n3965 & ~n3967 ;
  assign n3974 = ~n3937 & ~n3946 ;
  assign n3975 = \DataWidth_reg[1]/NET0131  & ~n3974 ;
  assign n3976 = ~n3968 & ~n3975 ;
  assign n3977 = ~n3973 & ~n3976 ;
  assign n3978 = n933 & ~n3977 ;
  assign n3979 = ~n668 & n3963 ;
  assign n3980 = ~n3966 & ~n3979 ;
  assign n3981 = n965 & ~n3980 ;
  assign n3969 = n1867 & ~n3968 ;
  assign n3982 = \InstQueue_reg[11][4]/NET0131  & ~n3929 ;
  assign n3983 = ~n3969 & ~n3982 ;
  assign n3984 = ~n3981 & n3983 ;
  assign n3985 = ~n3978 & n3984 ;
  assign n3994 = n3902 & n3937 ;
  assign n3995 = n3911 & n3935 ;
  assign n3996 = ~n3994 & ~n3995 ;
  assign n3997 = \DataWidth_reg[1]/NET0131  & ~n3996 ;
  assign n3986 = \InstQueueWr_Addr_reg[2]/NET0131  & n3857 ;
  assign n3987 = \InstQueueWr_Addr_reg[3]/NET0131  & n3986 ;
  assign n3988 = ~n3963 & ~n3987 ;
  assign n3989 = \Datai[4]_pad  & ~n3988 ;
  assign n3990 = \InstQueue_reg[12][4]/NET0131  & ~n3987 ;
  assign n3991 = ~n3963 & n3990 ;
  assign n3992 = ~n3989 & ~n3991 ;
  assign n3998 = \DataWidth_reg[1]/NET0131  & ~n3938 ;
  assign n3999 = ~n3992 & ~n3998 ;
  assign n4000 = ~n3997 & ~n3999 ;
  assign n4001 = n933 & ~n4000 ;
  assign n4002 = ~n668 & n3987 ;
  assign n4003 = ~n3990 & ~n4002 ;
  assign n4004 = n965 & ~n4003 ;
  assign n3993 = n1867 & ~n3992 ;
  assign n4005 = \InstQueue_reg[12][4]/NET0131  & ~n3929 ;
  assign n4006 = ~n3993 & ~n4005 ;
  assign n4007 = ~n4004 & n4006 ;
  assign n4008 = ~n4001 & n4007 ;
  assign n4015 = n3902 & n3935 ;
  assign n4016 = n3911 & n3963 ;
  assign n4017 = ~n4015 & ~n4016 ;
  assign n4018 = \DataWidth_reg[1]/NET0131  & ~n4017 ;
  assign n4009 = ~n3871 & ~n3987 ;
  assign n4010 = \Datai[4]_pad  & ~n4009 ;
  assign n4011 = \InstQueue_reg[13][4]/NET0131  & ~n3871 ;
  assign n4012 = ~n3987 & n4011 ;
  assign n4013 = ~n4010 & ~n4012 ;
  assign n4019 = \DataWidth_reg[1]/NET0131  & ~n3964 ;
  assign n4020 = ~n4013 & ~n4019 ;
  assign n4021 = ~n4018 & ~n4020 ;
  assign n4022 = n933 & ~n4021 ;
  assign n4023 = ~n668 & n3871 ;
  assign n4024 = ~n4011 & ~n4023 ;
  assign n4025 = n965 & ~n4024 ;
  assign n4014 = n1867 & ~n4013 ;
  assign n4026 = \InstQueue_reg[13][4]/NET0131  & ~n3929 ;
  assign n4027 = ~n4014 & ~n4026 ;
  assign n4028 = ~n4025 & n4027 ;
  assign n4029 = ~n4022 & n4028 ;
  assign n4035 = n3902 & n3963 ;
  assign n4036 = n3911 & n3987 ;
  assign n4037 = ~n4035 & ~n4036 ;
  assign n4038 = \DataWidth_reg[1]/NET0131  & ~n4037 ;
  assign n4030 = \Datai[4]_pad  & ~n3918 ;
  assign n4031 = \InstQueue_reg[14][4]/NET0131  & ~n3914 ;
  assign n4032 = ~n3871 & n4031 ;
  assign n4033 = ~n4030 & ~n4032 ;
  assign n4039 = \DataWidth_reg[1]/NET0131  & ~n3988 ;
  assign n4040 = ~n4033 & ~n4039 ;
  assign n4041 = ~n4038 & ~n4040 ;
  assign n4042 = n933 & ~n4041 ;
  assign n4043 = ~n668 & n3914 ;
  assign n4044 = ~n4031 & ~n4043 ;
  assign n4045 = n965 & ~n4044 ;
  assign n4034 = n1867 & ~n4033 ;
  assign n4046 = \InstQueue_reg[14][4]/NET0131  & ~n3929 ;
  assign n4047 = ~n4034 & ~n4046 ;
  assign n4048 = ~n4045 & n4047 ;
  assign n4049 = ~n4042 & n4048 ;
  assign n4056 = n3902 & n3987 ;
  assign n4057 = n3871 & n3911 ;
  assign n4058 = ~n4056 & ~n4057 ;
  assign n4059 = \DataWidth_reg[1]/NET0131  & ~n4058 ;
  assign n4050 = ~n3862 & ~n3914 ;
  assign n4051 = \Datai[4]_pad  & ~n4050 ;
  assign n4052 = \InstQueue_reg[15][4]/NET0131  & ~n3862 ;
  assign n4053 = ~n3914 & n4052 ;
  assign n4054 = ~n4051 & ~n4053 ;
  assign n4060 = \DataWidth_reg[1]/NET0131  & ~n4009 ;
  assign n4061 = ~n4054 & ~n4060 ;
  assign n4062 = ~n4059 & ~n4061 ;
  assign n4063 = n933 & ~n4062 ;
  assign n4064 = ~n668 & n3862 ;
  assign n4065 = ~n4052 & ~n4064 ;
  assign n4066 = n965 & ~n4065 ;
  assign n4055 = n1867 & ~n4054 ;
  assign n4067 = \InstQueue_reg[15][4]/NET0131  & ~n3929 ;
  assign n4068 = ~n4055 & ~n4067 ;
  assign n4069 = ~n4066 & n4068 ;
  assign n4070 = ~n4063 & n4069 ;
  assign n4078 = n3902 & n3914 ;
  assign n4079 = n3862 & n3911 ;
  assign n4080 = ~n4078 & ~n4079 ;
  assign n4081 = \DataWidth_reg[1]/NET0131  & ~n4080 ;
  assign n4071 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3936 ;
  assign n4072 = ~n3859 & ~n4071 ;
  assign n4073 = \Datai[4]_pad  & ~n4072 ;
  assign n4074 = \InstQueue_reg[1][4]/NET0131  & ~n4071 ;
  assign n4075 = ~n3859 & n4074 ;
  assign n4076 = ~n4073 & ~n4075 ;
  assign n4082 = \DataWidth_reg[1]/NET0131  & ~n4050 ;
  assign n4083 = ~n4076 & ~n4082 ;
  assign n4084 = ~n4081 & ~n4083 ;
  assign n4085 = n933 & ~n4084 ;
  assign n4086 = ~n668 & n4071 ;
  assign n4087 = ~n4074 & ~n4086 ;
  assign n4088 = n965 & ~n4087 ;
  assign n4077 = n1867 & ~n4076 ;
  assign n4089 = \InstQueue_reg[1][4]/NET0131  & ~n3929 ;
  assign n4090 = ~n4077 & ~n4089 ;
  assign n4091 = ~n4088 & n4090 ;
  assign n4092 = ~n4085 & n4091 ;
  assign n4100 = n3859 & n3911 ;
  assign n4101 = n3862 & n3902 ;
  assign n4102 = ~n4100 & ~n4101 ;
  assign n4103 = \DataWidth_reg[1]/NET0131  & ~n4102 ;
  assign n4093 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3934 ;
  assign n4094 = ~n4071 & ~n4093 ;
  assign n4095 = \Datai[4]_pad  & ~n4094 ;
  assign n4096 = \InstQueue_reg[2][4]/NET0131  & ~n4093 ;
  assign n4097 = ~n4071 & n4096 ;
  assign n4098 = ~n4095 & ~n4097 ;
  assign n4104 = \DataWidth_reg[1]/NET0131  & ~n3863 ;
  assign n4105 = ~n4098 & ~n4104 ;
  assign n4106 = ~n4103 & ~n4105 ;
  assign n4107 = n933 & ~n4106 ;
  assign n4108 = ~n668 & n4093 ;
  assign n4109 = ~n4096 & ~n4108 ;
  assign n4110 = n965 & ~n4109 ;
  assign n4099 = n1867 & ~n4098 ;
  assign n4111 = \InstQueue_reg[2][4]/NET0131  & ~n3929 ;
  assign n4112 = ~n4099 & ~n4111 ;
  assign n4113 = ~n4110 & n4112 ;
  assign n4114 = ~n4107 & n4113 ;
  assign n4122 = n3859 & n3902 ;
  assign n4123 = n3911 & n4071 ;
  assign n4124 = ~n4122 & ~n4123 ;
  assign n4125 = \DataWidth_reg[1]/NET0131  & ~n4124 ;
  assign n4115 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3962 ;
  assign n4116 = ~n4093 & ~n4115 ;
  assign n4117 = \Datai[4]_pad  & ~n4116 ;
  assign n4118 = \InstQueue_reg[3][4]/NET0131  & ~n4115 ;
  assign n4119 = ~n4093 & n4118 ;
  assign n4120 = ~n4117 & ~n4119 ;
  assign n4126 = \DataWidth_reg[1]/NET0131  & ~n4072 ;
  assign n4127 = ~n4120 & ~n4126 ;
  assign n4128 = ~n4125 & ~n4127 ;
  assign n4129 = n933 & ~n4128 ;
  assign n4130 = ~n668 & n4115 ;
  assign n4131 = ~n4118 & ~n4130 ;
  assign n4132 = n965 & ~n4131 ;
  assign n4121 = n1867 & ~n4120 ;
  assign n4133 = \InstQueue_reg[3][4]/NET0131  & ~n3929 ;
  assign n4134 = ~n4121 & ~n4133 ;
  assign n4135 = ~n4132 & n4134 ;
  assign n4136 = ~n4129 & n4135 ;
  assign n4144 = n3902 & n4071 ;
  assign n4145 = n3911 & n4093 ;
  assign n4146 = ~n4144 & ~n4145 ;
  assign n4147 = \DataWidth_reg[1]/NET0131  & ~n4146 ;
  assign n4137 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3986 ;
  assign n4138 = ~n4115 & ~n4137 ;
  assign n4139 = \Datai[4]_pad  & ~n4138 ;
  assign n4140 = \InstQueue_reg[4][4]/NET0131  & ~n4137 ;
  assign n4141 = ~n4115 & n4140 ;
  assign n4142 = ~n4139 & ~n4141 ;
  assign n4148 = \DataWidth_reg[1]/NET0131  & ~n4094 ;
  assign n4149 = ~n4142 & ~n4148 ;
  assign n4150 = ~n4147 & ~n4149 ;
  assign n4151 = n933 & ~n4150 ;
  assign n4152 = ~n668 & n4137 ;
  assign n4153 = ~n4140 & ~n4152 ;
  assign n4154 = n965 & ~n4153 ;
  assign n4143 = n1867 & ~n4142 ;
  assign n4155 = \InstQueue_reg[4][4]/NET0131  & ~n3929 ;
  assign n4156 = ~n4143 & ~n4155 ;
  assign n4157 = ~n4154 & n4156 ;
  assign n4158 = ~n4151 & n4157 ;
  assign n4166 = n3902 & n4093 ;
  assign n4167 = n3911 & n4115 ;
  assign n4168 = ~n4166 & ~n4167 ;
  assign n4169 = \DataWidth_reg[1]/NET0131  & ~n4168 ;
  assign n4159 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3870 ;
  assign n4160 = ~n4137 & ~n4159 ;
  assign n4161 = \Datai[4]_pad  & ~n4160 ;
  assign n4162 = \InstQueue_reg[5][4]/NET0131  & ~n4159 ;
  assign n4163 = ~n4137 & n4162 ;
  assign n4164 = ~n4161 & ~n4163 ;
  assign n4170 = \DataWidth_reg[1]/NET0131  & ~n4116 ;
  assign n4171 = ~n4164 & ~n4170 ;
  assign n4172 = ~n4169 & ~n4171 ;
  assign n4173 = n933 & ~n4172 ;
  assign n4174 = ~n668 & n4159 ;
  assign n4175 = ~n4162 & ~n4174 ;
  assign n4176 = n965 & ~n4175 ;
  assign n4165 = n1867 & ~n4164 ;
  assign n4177 = \InstQueue_reg[5][4]/NET0131  & ~n3929 ;
  assign n4178 = ~n4165 & ~n4177 ;
  assign n4179 = ~n4176 & n4178 ;
  assign n4180 = ~n4173 & n4179 ;
  assign n4188 = n3902 & n4115 ;
  assign n4189 = n3911 & n4137 ;
  assign n4190 = ~n4188 & ~n4189 ;
  assign n4191 = \DataWidth_reg[1]/NET0131  & ~n4190 ;
  assign n4181 = ~\InstQueueWr_Addr_reg[3]/NET0131  & n3913 ;
  assign n4182 = ~n4159 & ~n4181 ;
  assign n4183 = \Datai[4]_pad  & ~n4182 ;
  assign n4184 = \InstQueue_reg[6][4]/NET0131  & ~n4181 ;
  assign n4185 = ~n4159 & n4184 ;
  assign n4186 = ~n4183 & ~n4185 ;
  assign n4192 = \DataWidth_reg[1]/NET0131  & ~n4138 ;
  assign n4193 = ~n4186 & ~n4192 ;
  assign n4194 = ~n4191 & ~n4193 ;
  assign n4195 = n933 & ~n4194 ;
  assign n4196 = ~n668 & n4181 ;
  assign n4197 = ~n4184 & ~n4196 ;
  assign n4198 = n965 & ~n4197 ;
  assign n4187 = n1867 & ~n4186 ;
  assign n4199 = \InstQueue_reg[6][4]/NET0131  & ~n3929 ;
  assign n4200 = ~n4187 & ~n4199 ;
  assign n4201 = ~n4198 & n4200 ;
  assign n4202 = ~n4195 & n4201 ;
  assign n4209 = n3902 & n4137 ;
  assign n4210 = n3911 & n4159 ;
  assign n4211 = ~n4209 & ~n4210 ;
  assign n4212 = \DataWidth_reg[1]/NET0131  & ~n4211 ;
  assign n4203 = ~n3944 & ~n4181 ;
  assign n4204 = \Datai[4]_pad  & ~n4203 ;
  assign n4205 = \InstQueue_reg[7][4]/NET0131  & ~n3944 ;
  assign n4206 = ~n4181 & n4205 ;
  assign n4207 = ~n4204 & ~n4206 ;
  assign n4213 = \DataWidth_reg[1]/NET0131  & ~n4160 ;
  assign n4214 = ~n4207 & ~n4213 ;
  assign n4215 = ~n4212 & ~n4214 ;
  assign n4216 = n933 & ~n4215 ;
  assign n4217 = ~n668 & n3944 ;
  assign n4218 = ~n4205 & ~n4217 ;
  assign n4219 = n965 & ~n4218 ;
  assign n4208 = n1867 & ~n4207 ;
  assign n4220 = \InstQueue_reg[7][4]/NET0131  & ~n3929 ;
  assign n4221 = ~n4208 & ~n4220 ;
  assign n4222 = ~n4219 & n4221 ;
  assign n4223 = ~n4216 & n4222 ;
  assign n4229 = n3902 & n4159 ;
  assign n4230 = n3911 & n4181 ;
  assign n4231 = ~n4229 & ~n4230 ;
  assign n4232 = \DataWidth_reg[1]/NET0131  & ~n4231 ;
  assign n4224 = \Datai[4]_pad  & ~n3950 ;
  assign n4225 = \InstQueue_reg[8][4]/NET0131  & ~n3946 ;
  assign n4226 = ~n3944 & n4225 ;
  assign n4227 = ~n4224 & ~n4226 ;
  assign n4233 = \DataWidth_reg[1]/NET0131  & ~n4182 ;
  assign n4234 = ~n4227 & ~n4233 ;
  assign n4235 = ~n4232 & ~n4234 ;
  assign n4236 = n933 & ~n4235 ;
  assign n4237 = ~n668 & n3946 ;
  assign n4238 = ~n4225 & ~n4237 ;
  assign n4239 = n965 & ~n4238 ;
  assign n4228 = n1867 & ~n4227 ;
  assign n4240 = \InstQueue_reg[8][4]/NET0131  & ~n3929 ;
  assign n4241 = ~n4228 & ~n4240 ;
  assign n4242 = ~n4239 & n4241 ;
  assign n4243 = ~n4236 & n4242 ;
  assign n4249 = n3902 & n4181 ;
  assign n4250 = n3911 & n3944 ;
  assign n4251 = ~n4249 & ~n4250 ;
  assign n4252 = \DataWidth_reg[1]/NET0131  & ~n4251 ;
  assign n4244 = \Datai[4]_pad  & ~n3974 ;
  assign n4245 = \InstQueue_reg[9][4]/NET0131  & ~n3937 ;
  assign n4246 = ~n3946 & n4245 ;
  assign n4247 = ~n4244 & ~n4246 ;
  assign n4253 = \DataWidth_reg[1]/NET0131  & ~n4203 ;
  assign n4254 = ~n4247 & ~n4253 ;
  assign n4255 = ~n4252 & ~n4254 ;
  assign n4256 = n933 & ~n4255 ;
  assign n4257 = ~n668 & n3937 ;
  assign n4258 = ~n4245 & ~n4257 ;
  assign n4259 = n965 & ~n4258 ;
  assign n4248 = n1867 & ~n4247 ;
  assign n4260 = \InstQueue_reg[9][4]/NET0131  & ~n3929 ;
  assign n4261 = ~n4248 & ~n4260 ;
  assign n4262 = ~n4259 & n4261 ;
  assign n4263 = ~n4256 & n4262 ;
  assign n4271 = \PhyAddrPointer_reg[2]/NET0131  & ~n2739 ;
  assign n4272 = n773 & n3555 ;
  assign n4273 = ~n3562 & ~n4272 ;
  assign n4274 = ~n4271 & n4273 ;
  assign n4275 = n929 & ~n4274 ;
  assign n4267 = ~n955 & ~n965 ;
  assign n4268 = n3926 & n4267 ;
  assign n4269 = \PhyAddrPointer_reg[2]/NET0131  & ~n4268 ;
  assign n4264 = ~\PhyAddrPointer_reg[1]/NET0131  & ~\PhyAddrPointer_reg[2]/NET0131  ;
  assign n4265 = ~n3530 & ~n4264 ;
  assign n4266 = n2100 & n4265 ;
  assign n4270 = ~\PhyAddrPointer_reg[2]/NET0131  & n969 ;
  assign n4276 = ~n3540 & ~n4270 ;
  assign n4277 = ~n4266 & n4276 ;
  assign n4278 = ~n4269 & n4277 ;
  assign n4279 = ~n4275 & n4278 ;
  assign n4281 = \EAX_reg[19]/NET0131  & n3682 ;
  assign n4282 = \EAX_reg[20]/NET0131  & n4281 ;
  assign n4283 = ~\EAX_reg[20]/NET0131  & ~n4281 ;
  assign n4284 = ~n4282 & ~n4283 ;
  assign n4285 = ~n828 & ~n4284 ;
  assign n4286 = n923 & ~n4285 ;
  assign n4287 = n3827 & ~n4286 ;
  assign n4288 = \Datao[20]_pad  & ~n4287 ;
  assign n4289 = n923 & n4284 ;
  assign n4290 = ~n828 & n4289 ;
  assign n4291 = ~n4288 & ~n4290 ;
  assign n4292 = n929 & ~n4291 ;
  assign n4280 = \uWord_reg[4]/NET0131  & n3809 ;
  assign n4293 = \Datao[20]_pad  & ~n3821 ;
  assign n4294 = ~n4280 & ~n4293 ;
  assign n4295 = ~n4292 & n4294 ;
  assign n4296 = \uWord_reg[4]/NET0131  & ~n3655 ;
  assign n4297 = READY_n_pad & \uWord_reg[4]/NET0131  ;
  assign n4298 = \Datai[4]_pad  & n846 ;
  assign n4299 = ~n4297 & ~n4298 ;
  assign n4300 = n782 & ~n4299 ;
  assign n4301 = \uWord_reg[4]/NET0131  & n3661 ;
  assign n4302 = ~n4289 & ~n4301 ;
  assign n4303 = ~n4300 & n4302 ;
  assign n4304 = n929 & ~n4303 ;
  assign n4305 = ~n4296 & ~n4304 ;
  assign n4309 = ~\EAX_reg[25]/NET0131  & ~n3159 ;
  assign n4310 = n3132 & ~n3160 ;
  assign n4311 = ~n4309 & n4310 ;
  assign n4312 = \EAX_reg[25]/NET0131  & n3135 ;
  assign n4313 = \EAX_reg[25]/NET0131  & ~n846 ;
  assign n4317 = \Datai[25]_pad  & n846 ;
  assign n4318 = ~n4313 & ~n4317 ;
  assign n4319 = n840 & ~n4318 ;
  assign n4306 = ~n3032 & n3063 ;
  assign n4307 = ~n3064 & ~n4306 ;
  assign n4308 = n2937 & n4307 ;
  assign n4314 = \Datai[9]_pad  & n846 ;
  assign n4315 = ~n4313 & ~n4314 ;
  assign n4316 = n782 & ~n4315 ;
  assign n4320 = ~n4308 & ~n4316 ;
  assign n4321 = ~n4319 & n4320 ;
  assign n4322 = ~n4312 & n4321 ;
  assign n4323 = ~n4311 & n4322 ;
  assign n4324 = n929 & ~n4323 ;
  assign n4325 = \EAX_reg[25]/NET0131  & ~n3181 ;
  assign n4326 = ~n4324 & ~n4325 ;
  assign n4332 = \Datai[29]_pad  & n3900 ;
  assign n4333 = \Datai[30]_pad  & n4332 ;
  assign n4334 = \Datai[31]_pad  & ~n4333 ;
  assign n4335 = n3871 & n4334 ;
  assign n4336 = \Datai[21]_pad  & n3910 ;
  assign n4337 = \Datai[22]_pad  & n4336 ;
  assign n4338 = ~\Datai[23]_pad  & ~n4337 ;
  assign n4339 = \Datai[23]_pad  & n4337 ;
  assign n4340 = ~n4338 & ~n4339 ;
  assign n4341 = n3914 & n4340 ;
  assign n4342 = ~n4335 & ~n4341 ;
  assign n4343 = \DataWidth_reg[1]/NET0131  & ~n4342 ;
  assign n4327 = \Datai[7]_pad  & ~n3863 ;
  assign n4328 = \InstQueue_reg[0][7]/NET0131  & ~n3859 ;
  assign n4329 = ~n3862 & n4328 ;
  assign n4330 = ~n4327 & ~n4329 ;
  assign n4344 = ~n3919 & ~n4330 ;
  assign n4345 = ~n4343 & ~n4344 ;
  assign n4346 = n933 & ~n4345 ;
  assign n4347 = ~n700 & n3859 ;
  assign n4348 = ~n4328 & ~n4347 ;
  assign n4349 = n965 & ~n4348 ;
  assign n4331 = n1867 & ~n4330 ;
  assign n4350 = \InstQueue_reg[0][7]/NET0131  & ~n3929 ;
  assign n4351 = ~n4331 & ~n4350 ;
  assign n4352 = ~n4349 & n4351 ;
  assign n4353 = ~n4346 & n4352 ;
  assign n4359 = n3944 & n4334 ;
  assign n4360 = n3946 & n4340 ;
  assign n4361 = ~n4359 & ~n4360 ;
  assign n4362 = \DataWidth_reg[1]/NET0131  & ~n4361 ;
  assign n4354 = \Datai[7]_pad  & ~n3938 ;
  assign n4355 = \InstQueue_reg[10][7]/NET0131  & ~n3935 ;
  assign n4356 = ~n3937 & n4355 ;
  assign n4357 = ~n4354 & ~n4356 ;
  assign n4363 = ~n3951 & ~n4357 ;
  assign n4364 = ~n4362 & ~n4363 ;
  assign n4365 = n933 & ~n4364 ;
  assign n4366 = ~n700 & n3935 ;
  assign n4367 = ~n4355 & ~n4366 ;
  assign n4368 = n965 & ~n4367 ;
  assign n4358 = n1867 & ~n4357 ;
  assign n4369 = \InstQueue_reg[10][7]/NET0131  & ~n3929 ;
  assign n4370 = ~n4358 & ~n4369 ;
  assign n4371 = ~n4368 & n4370 ;
  assign n4372 = ~n4365 & n4371 ;
  assign n4378 = n3946 & n4334 ;
  assign n4379 = n3937 & n4340 ;
  assign n4380 = ~n4378 & ~n4379 ;
  assign n4381 = \DataWidth_reg[1]/NET0131  & ~n4380 ;
  assign n4373 = \Datai[7]_pad  & ~n3964 ;
  assign n4374 = \InstQueue_reg[11][7]/NET0131  & ~n3963 ;
  assign n4375 = ~n3935 & n4374 ;
  assign n4376 = ~n4373 & ~n4375 ;
  assign n4382 = ~n3975 & ~n4376 ;
  assign n4383 = ~n4381 & ~n4382 ;
  assign n4384 = n933 & ~n4383 ;
  assign n4385 = ~n700 & n3963 ;
  assign n4386 = ~n4374 & ~n4385 ;
  assign n4387 = n965 & ~n4386 ;
  assign n4377 = n1867 & ~n4376 ;
  assign n4388 = \InstQueue_reg[11][7]/NET0131  & ~n3929 ;
  assign n4389 = ~n4377 & ~n4388 ;
  assign n4390 = ~n4387 & n4389 ;
  assign n4391 = ~n4384 & n4390 ;
  assign n4397 = n3937 & n4334 ;
  assign n4398 = n3935 & n4340 ;
  assign n4399 = ~n4397 & ~n4398 ;
  assign n4400 = \DataWidth_reg[1]/NET0131  & ~n4399 ;
  assign n4392 = \Datai[7]_pad  & ~n3988 ;
  assign n4393 = \InstQueue_reg[12][7]/NET0131  & ~n3987 ;
  assign n4394 = ~n3963 & n4393 ;
  assign n4395 = ~n4392 & ~n4394 ;
  assign n4401 = ~n3998 & ~n4395 ;
  assign n4402 = ~n4400 & ~n4401 ;
  assign n4403 = n933 & ~n4402 ;
  assign n4404 = ~n700 & n3987 ;
  assign n4405 = ~n4393 & ~n4404 ;
  assign n4406 = n965 & ~n4405 ;
  assign n4396 = n1867 & ~n4395 ;
  assign n4407 = \InstQueue_reg[12][7]/NET0131  & ~n3929 ;
  assign n4408 = ~n4396 & ~n4407 ;
  assign n4409 = ~n4406 & n4408 ;
  assign n4410 = ~n4403 & n4409 ;
  assign n4416 = n3935 & n4334 ;
  assign n4417 = n3963 & n4340 ;
  assign n4418 = ~n4416 & ~n4417 ;
  assign n4419 = \DataWidth_reg[1]/NET0131  & ~n4418 ;
  assign n4411 = \Datai[7]_pad  & ~n4009 ;
  assign n4412 = \InstQueue_reg[13][7]/NET0131  & ~n3871 ;
  assign n4413 = ~n3987 & n4412 ;
  assign n4414 = ~n4411 & ~n4413 ;
  assign n4420 = ~n4019 & ~n4414 ;
  assign n4421 = ~n4419 & ~n4420 ;
  assign n4422 = n933 & ~n4421 ;
  assign n4423 = ~n700 & n3871 ;
  assign n4424 = ~n4412 & ~n4423 ;
  assign n4425 = n965 & ~n4424 ;
  assign n4415 = n1867 & ~n4414 ;
  assign n4426 = \InstQueue_reg[13][7]/NET0131  & ~n3929 ;
  assign n4427 = ~n4415 & ~n4426 ;
  assign n4428 = ~n4425 & n4427 ;
  assign n4429 = ~n4422 & n4428 ;
  assign n4435 = n3963 & n4334 ;
  assign n4436 = n3987 & n4340 ;
  assign n4437 = ~n4435 & ~n4436 ;
  assign n4438 = \DataWidth_reg[1]/NET0131  & ~n4437 ;
  assign n4430 = \Datai[7]_pad  & ~n3918 ;
  assign n4431 = \InstQueue_reg[14][7]/NET0131  & ~n3914 ;
  assign n4432 = ~n3871 & n4431 ;
  assign n4433 = ~n4430 & ~n4432 ;
  assign n4439 = ~n4039 & ~n4433 ;
  assign n4440 = ~n4438 & ~n4439 ;
  assign n4441 = n933 & ~n4440 ;
  assign n4442 = ~n700 & n3914 ;
  assign n4443 = ~n4431 & ~n4442 ;
  assign n4444 = n965 & ~n4443 ;
  assign n4434 = n1867 & ~n4433 ;
  assign n4445 = \InstQueue_reg[14][7]/NET0131  & ~n3929 ;
  assign n4446 = ~n4434 & ~n4445 ;
  assign n4447 = ~n4444 & n4446 ;
  assign n4448 = ~n4441 & n4447 ;
  assign n4454 = n3987 & n4334 ;
  assign n4455 = n3871 & n4340 ;
  assign n4456 = ~n4454 & ~n4455 ;
  assign n4457 = \DataWidth_reg[1]/NET0131  & ~n4456 ;
  assign n4449 = \Datai[7]_pad  & ~n4050 ;
  assign n4450 = \InstQueue_reg[15][7]/NET0131  & ~n3862 ;
  assign n4451 = ~n3914 & n4450 ;
  assign n4452 = ~n4449 & ~n4451 ;
  assign n4458 = ~n4060 & ~n4452 ;
  assign n4459 = ~n4457 & ~n4458 ;
  assign n4460 = n933 & ~n4459 ;
  assign n4461 = ~n700 & n3862 ;
  assign n4462 = ~n4450 & ~n4461 ;
  assign n4463 = n965 & ~n4462 ;
  assign n4453 = n1867 & ~n4452 ;
  assign n4464 = \InstQueue_reg[15][7]/NET0131  & ~n3929 ;
  assign n4465 = ~n4453 & ~n4464 ;
  assign n4466 = ~n4463 & n4465 ;
  assign n4467 = ~n4460 & n4466 ;
  assign n4473 = n3914 & n4334 ;
  assign n4474 = n3862 & n4340 ;
  assign n4475 = ~n4473 & ~n4474 ;
  assign n4476 = \DataWidth_reg[1]/NET0131  & ~n4475 ;
  assign n4468 = \Datai[7]_pad  & ~n4072 ;
  assign n4469 = \InstQueue_reg[1][7]/NET0131  & ~n4071 ;
  assign n4470 = ~n3859 & n4469 ;
  assign n4471 = ~n4468 & ~n4470 ;
  assign n4477 = ~n4082 & ~n4471 ;
  assign n4478 = ~n4476 & ~n4477 ;
  assign n4479 = n933 & ~n4478 ;
  assign n4480 = ~n700 & n4071 ;
  assign n4481 = ~n4469 & ~n4480 ;
  assign n4482 = n965 & ~n4481 ;
  assign n4472 = n1867 & ~n4471 ;
  assign n4483 = \InstQueue_reg[1][7]/NET0131  & ~n3929 ;
  assign n4484 = ~n4472 & ~n4483 ;
  assign n4485 = ~n4482 & n4484 ;
  assign n4486 = ~n4479 & n4485 ;
  assign n4492 = n3859 & n4340 ;
  assign n4493 = n3862 & n4334 ;
  assign n4494 = ~n4492 & ~n4493 ;
  assign n4495 = \DataWidth_reg[1]/NET0131  & ~n4494 ;
  assign n4487 = \Datai[7]_pad  & ~n4094 ;
  assign n4488 = \InstQueue_reg[2][7]/NET0131  & ~n4093 ;
  assign n4489 = ~n4071 & n4488 ;
  assign n4490 = ~n4487 & ~n4489 ;
  assign n4496 = ~n4104 & ~n4490 ;
  assign n4497 = ~n4495 & ~n4496 ;
  assign n4498 = n933 & ~n4497 ;
  assign n4499 = ~n700 & n4093 ;
  assign n4500 = ~n4488 & ~n4499 ;
  assign n4501 = n965 & ~n4500 ;
  assign n4491 = n1867 & ~n4490 ;
  assign n4502 = \InstQueue_reg[2][7]/NET0131  & ~n3929 ;
  assign n4503 = ~n4491 & ~n4502 ;
  assign n4504 = ~n4501 & n4503 ;
  assign n4505 = ~n4498 & n4504 ;
  assign n4511 = n3859 & n4334 ;
  assign n4512 = n4071 & n4340 ;
  assign n4513 = ~n4511 & ~n4512 ;
  assign n4514 = \DataWidth_reg[1]/NET0131  & ~n4513 ;
  assign n4506 = \Datai[7]_pad  & ~n4116 ;
  assign n4507 = \InstQueue_reg[3][7]/NET0131  & ~n4115 ;
  assign n4508 = ~n4093 & n4507 ;
  assign n4509 = ~n4506 & ~n4508 ;
  assign n4515 = ~n4126 & ~n4509 ;
  assign n4516 = ~n4514 & ~n4515 ;
  assign n4517 = n933 & ~n4516 ;
  assign n4518 = ~n700 & n4115 ;
  assign n4519 = ~n4507 & ~n4518 ;
  assign n4520 = n965 & ~n4519 ;
  assign n4510 = n1867 & ~n4509 ;
  assign n4521 = \InstQueue_reg[3][7]/NET0131  & ~n3929 ;
  assign n4522 = ~n4510 & ~n4521 ;
  assign n4523 = ~n4520 & n4522 ;
  assign n4524 = ~n4517 & n4523 ;
  assign n4530 = n4071 & n4334 ;
  assign n4531 = n4093 & n4340 ;
  assign n4532 = ~n4530 & ~n4531 ;
  assign n4533 = \DataWidth_reg[1]/NET0131  & ~n4532 ;
  assign n4525 = \Datai[7]_pad  & ~n4138 ;
  assign n4526 = \InstQueue_reg[4][7]/NET0131  & ~n4137 ;
  assign n4527 = ~n4115 & n4526 ;
  assign n4528 = ~n4525 & ~n4527 ;
  assign n4534 = ~n4148 & ~n4528 ;
  assign n4535 = ~n4533 & ~n4534 ;
  assign n4536 = n933 & ~n4535 ;
  assign n4537 = ~n700 & n4137 ;
  assign n4538 = ~n4526 & ~n4537 ;
  assign n4539 = n965 & ~n4538 ;
  assign n4529 = n1867 & ~n4528 ;
  assign n4540 = \InstQueue_reg[4][7]/NET0131  & ~n3929 ;
  assign n4541 = ~n4529 & ~n4540 ;
  assign n4542 = ~n4539 & n4541 ;
  assign n4543 = ~n4536 & n4542 ;
  assign n4549 = n4093 & n4334 ;
  assign n4550 = n4115 & n4340 ;
  assign n4551 = ~n4549 & ~n4550 ;
  assign n4552 = \DataWidth_reg[1]/NET0131  & ~n4551 ;
  assign n4544 = \Datai[7]_pad  & ~n4160 ;
  assign n4545 = \InstQueue_reg[5][7]/NET0131  & ~n4159 ;
  assign n4546 = ~n4137 & n4545 ;
  assign n4547 = ~n4544 & ~n4546 ;
  assign n4553 = ~n4170 & ~n4547 ;
  assign n4554 = ~n4552 & ~n4553 ;
  assign n4555 = n933 & ~n4554 ;
  assign n4556 = ~n700 & n4159 ;
  assign n4557 = ~n4545 & ~n4556 ;
  assign n4558 = n965 & ~n4557 ;
  assign n4548 = n1867 & ~n4547 ;
  assign n4559 = \InstQueue_reg[5][7]/NET0131  & ~n3929 ;
  assign n4560 = ~n4548 & ~n4559 ;
  assign n4561 = ~n4558 & n4560 ;
  assign n4562 = ~n4555 & n4561 ;
  assign n4568 = n4115 & n4334 ;
  assign n4569 = n4137 & n4340 ;
  assign n4570 = ~n4568 & ~n4569 ;
  assign n4571 = \DataWidth_reg[1]/NET0131  & ~n4570 ;
  assign n4563 = \Datai[7]_pad  & ~n4182 ;
  assign n4564 = \InstQueue_reg[6][7]/NET0131  & ~n4181 ;
  assign n4565 = ~n4159 & n4564 ;
  assign n4566 = ~n4563 & ~n4565 ;
  assign n4572 = ~n4192 & ~n4566 ;
  assign n4573 = ~n4571 & ~n4572 ;
  assign n4574 = n933 & ~n4573 ;
  assign n4575 = ~n700 & n4181 ;
  assign n4576 = ~n4564 & ~n4575 ;
  assign n4577 = n965 & ~n4576 ;
  assign n4567 = n1867 & ~n4566 ;
  assign n4578 = \InstQueue_reg[6][7]/NET0131  & ~n3929 ;
  assign n4579 = ~n4567 & ~n4578 ;
  assign n4580 = ~n4577 & n4579 ;
  assign n4581 = ~n4574 & n4580 ;
  assign n4587 = n4137 & n4334 ;
  assign n4588 = n4159 & n4340 ;
  assign n4589 = ~n4587 & ~n4588 ;
  assign n4590 = \DataWidth_reg[1]/NET0131  & ~n4589 ;
  assign n4582 = \Datai[7]_pad  & ~n4203 ;
  assign n4583 = \InstQueue_reg[7][7]/NET0131  & ~n3944 ;
  assign n4584 = ~n4181 & n4583 ;
  assign n4585 = ~n4582 & ~n4584 ;
  assign n4591 = ~n4213 & ~n4585 ;
  assign n4592 = ~n4590 & ~n4591 ;
  assign n4593 = n933 & ~n4592 ;
  assign n4594 = ~n700 & n3944 ;
  assign n4595 = ~n4583 & ~n4594 ;
  assign n4596 = n965 & ~n4595 ;
  assign n4586 = n1867 & ~n4585 ;
  assign n4597 = \InstQueue_reg[7][7]/NET0131  & ~n3929 ;
  assign n4598 = ~n4586 & ~n4597 ;
  assign n4599 = ~n4596 & n4598 ;
  assign n4600 = ~n4593 & n4599 ;
  assign n4606 = n4159 & n4334 ;
  assign n4607 = n4181 & n4340 ;
  assign n4608 = ~n4606 & ~n4607 ;
  assign n4609 = \DataWidth_reg[1]/NET0131  & ~n4608 ;
  assign n4601 = \Datai[7]_pad  & ~n3950 ;
  assign n4602 = \InstQueue_reg[8][7]/NET0131  & ~n3946 ;
  assign n4603 = ~n3944 & n4602 ;
  assign n4604 = ~n4601 & ~n4603 ;
  assign n4610 = ~n4233 & ~n4604 ;
  assign n4611 = ~n4609 & ~n4610 ;
  assign n4612 = n933 & ~n4611 ;
  assign n4613 = ~n700 & n3946 ;
  assign n4614 = ~n4602 & ~n4613 ;
  assign n4615 = n965 & ~n4614 ;
  assign n4605 = n1867 & ~n4604 ;
  assign n4616 = \InstQueue_reg[8][7]/NET0131  & ~n3929 ;
  assign n4617 = ~n4605 & ~n4616 ;
  assign n4618 = ~n4615 & n4617 ;
  assign n4619 = ~n4612 & n4618 ;
  assign n4625 = n4181 & n4334 ;
  assign n4626 = n3944 & n4340 ;
  assign n4627 = ~n4625 & ~n4626 ;
  assign n4628 = \DataWidth_reg[1]/NET0131  & ~n4627 ;
  assign n4620 = \Datai[7]_pad  & ~n3974 ;
  assign n4621 = \InstQueue_reg[9][7]/NET0131  & ~n3937 ;
  assign n4622 = ~n3946 & n4621 ;
  assign n4623 = ~n4620 & ~n4622 ;
  assign n4629 = ~n4253 & ~n4623 ;
  assign n4630 = ~n4628 & ~n4629 ;
  assign n4631 = n933 & ~n4630 ;
  assign n4632 = ~n700 & n3937 ;
  assign n4633 = ~n4621 & ~n4632 ;
  assign n4634 = n965 & ~n4633 ;
  assign n4624 = n1867 & ~n4623 ;
  assign n4635 = \InstQueue_reg[9][7]/NET0131  & ~n3929 ;
  assign n4636 = ~n4624 & ~n4635 ;
  assign n4637 = ~n4634 & n4636 ;
  assign n4638 = ~n4631 & n4637 ;
  assign n4640 = \EAX_reg[26]/NET0131  & n3685 ;
  assign n4641 = ~\EAX_reg[27]/NET0131  & ~n4640 ;
  assign n4642 = n923 & ~n3686 ;
  assign n4643 = ~n4641 & n4642 ;
  assign n4644 = ~n828 & n4643 ;
  assign n4645 = \Datao[27]_pad  & ~n857 ;
  assign n4646 = ~n4644 & ~n4645 ;
  assign n4647 = n929 & ~n4646 ;
  assign n4639 = \uWord_reg[11]/NET0131  & n3809 ;
  assign n4648 = \Datao[27]_pad  & ~n3821 ;
  assign n4649 = ~n4639 & ~n4648 ;
  assign n4650 = ~n4647 & n4649 ;
  assign n4651 = \EBX_reg[27]/NET0131  & ~n3181 ;
  assign n4653 = ~n3465 & ~n3801 ;
  assign n4654 = \EBX_reg[27]/NET0131  & ~n4653 ;
  assign n4652 = n3130 & n3463 ;
  assign n4655 = ~\EBX_reg[27]/NET0131  & n797 ;
  assign n4656 = n3800 & n4655 ;
  assign n4657 = ~n4652 & ~n4656 ;
  assign n4658 = ~n4654 & n4657 ;
  assign n4659 = n929 & ~n4658 ;
  assign n4660 = ~n4651 & ~n4659 ;
  assign n4661 = \uWord_reg[11]/NET0131  & ~n3655 ;
  assign n4662 = READY_n_pad & \uWord_reg[11]/NET0131  ;
  assign n4663 = ~n3166 & ~n4662 ;
  assign n4664 = n782 & ~n4663 ;
  assign n4665 = \uWord_reg[11]/NET0131  & n3661 ;
  assign n4666 = ~n4643 & ~n4665 ;
  assign n4667 = ~n4664 & n4666 ;
  assign n4668 = n929 & ~n4667 ;
  assign n4669 = ~n4661 & ~n4668 ;
  assign n4670 = n929 & ~n3430 ;
  assign n4671 = n3181 & ~n4670 ;
  assign n4672 = \EAX_reg[7]/NET0131  & ~n4671 ;
  assign n4674 = \Datai[7]_pad  & n846 ;
  assign n4675 = ~n841 & n4674 ;
  assign n4673 = ~n1014 & n2937 ;
  assign n4676 = ~\EAX_reg[7]/NET0131  & ~n3141 ;
  assign n4677 = ~n3142 & ~n4676 ;
  assign n4678 = n3132 & n4677 ;
  assign n4679 = ~n4673 & ~n4678 ;
  assign n4680 = ~n4675 & n4679 ;
  assign n4681 = n929 & ~n4680 ;
  assign n4682 = ~n4672 & ~n4681 ;
  assign n4683 = \EAX_reg[8]/NET0131  & ~n4671 ;
  assign n4684 = n842 & n3841 ;
  assign n4689 = \InstQueue_reg[9][0]/NET0131  & n454 ;
  assign n4690 = \InstQueue_reg[3][0]/NET0131  & n488 ;
  assign n4703 = ~n4689 & ~n4690 ;
  assign n4691 = \InstQueue_reg[15][0]/NET0131  & n465 ;
  assign n4692 = \InstQueue_reg[10][0]/NET0131  & n486 ;
  assign n4704 = ~n4691 & ~n4692 ;
  assign n4711 = n4703 & n4704 ;
  assign n4685 = \InstQueue_reg[0][0]/NET0131  & n470 ;
  assign n4686 = \InstQueue_reg[11][0]/NET0131  & n484 ;
  assign n4701 = ~n4685 & ~n4686 ;
  assign n4687 = \InstQueue_reg[6][0]/NET0131  & n472 ;
  assign n4688 = \InstQueue_reg[5][0]/NET0131  & n476 ;
  assign n4702 = ~n4687 & ~n4688 ;
  assign n4712 = n4701 & n4702 ;
  assign n4713 = n4711 & n4712 ;
  assign n4697 = \InstQueue_reg[2][0]/NET0131  & n474 ;
  assign n4698 = \InstQueue_reg[4][0]/NET0131  & n458 ;
  assign n4707 = ~n4697 & ~n4698 ;
  assign n4699 = \InstQueue_reg[1][0]/NET0131  & n522 ;
  assign n4700 = \InstQueue_reg[8][0]/NET0131  & n482 ;
  assign n4708 = ~n4699 & ~n4700 ;
  assign n4709 = n4707 & n4708 ;
  assign n4693 = \InstQueue_reg[14][0]/NET0131  & n468 ;
  assign n4694 = \InstQueue_reg[7][0]/NET0131  & n490 ;
  assign n4705 = ~n4693 & ~n4694 ;
  assign n4695 = \InstQueue_reg[13][0]/NET0131  & n492 ;
  assign n4696 = \InstQueue_reg[12][0]/NET0131  & n461 ;
  assign n4706 = ~n4695 & ~n4696 ;
  assign n4710 = n4705 & n4706 ;
  assign n4714 = n4709 & n4710 ;
  assign n4715 = n4713 & n4714 ;
  assign n4716 = n2937 & ~n4715 ;
  assign n4717 = ~\EAX_reg[8]/NET0131  & ~n3142 ;
  assign n4718 = ~n3143 & ~n4717 ;
  assign n4719 = n3132 & n4718 ;
  assign n4720 = ~n4716 & ~n4719 ;
  assign n4721 = ~n4684 & n4720 ;
  assign n4722 = n929 & ~n4721 ;
  assign n4723 = ~n4683 & ~n4722 ;
  assign n4724 = \EAX_reg[9]/NET0131  & ~n4671 ;
  assign n4730 = \InstQueue_reg[9][1]/NET0131  & n454 ;
  assign n4731 = \InstQueue_reg[3][1]/NET0131  & n488 ;
  assign n4744 = ~n4730 & ~n4731 ;
  assign n4732 = \InstQueue_reg[6][1]/NET0131  & n472 ;
  assign n4733 = \InstQueue_reg[5][1]/NET0131  & n476 ;
  assign n4745 = ~n4732 & ~n4733 ;
  assign n4752 = n4744 & n4745 ;
  assign n4726 = \InstQueue_reg[8][1]/NET0131  & n482 ;
  assign n4727 = \InstQueue_reg[11][1]/NET0131  & n484 ;
  assign n4742 = ~n4726 & ~n4727 ;
  assign n4728 = \InstQueue_reg[1][1]/NET0131  & n522 ;
  assign n4729 = \InstQueue_reg[0][1]/NET0131  & n470 ;
  assign n4743 = ~n4728 & ~n4729 ;
  assign n4753 = n4742 & n4743 ;
  assign n4754 = n4752 & n4753 ;
  assign n4738 = \InstQueue_reg[12][1]/NET0131  & n461 ;
  assign n4739 = \InstQueue_reg[4][1]/NET0131  & n458 ;
  assign n4748 = ~n4738 & ~n4739 ;
  assign n4740 = \InstQueue_reg[14][1]/NET0131  & n468 ;
  assign n4741 = \InstQueue_reg[15][1]/NET0131  & n465 ;
  assign n4749 = ~n4740 & ~n4741 ;
  assign n4750 = n4748 & n4749 ;
  assign n4734 = \InstQueue_reg[7][1]/NET0131  & n490 ;
  assign n4735 = \InstQueue_reg[2][1]/NET0131  & n474 ;
  assign n4746 = ~n4734 & ~n4735 ;
  assign n4736 = \InstQueue_reg[13][1]/NET0131  & n492 ;
  assign n4737 = \InstQueue_reg[10][1]/NET0131  & n486 ;
  assign n4747 = ~n4736 & ~n4737 ;
  assign n4751 = n4746 & n4747 ;
  assign n4755 = n4750 & n4751 ;
  assign n4756 = n4754 & n4755 ;
  assign n4757 = n2937 & ~n4756 ;
  assign n4725 = ~n841 & n4314 ;
  assign n4758 = ~\EAX_reg[9]/NET0131  & ~n3143 ;
  assign n4759 = ~n3144 & ~n4758 ;
  assign n4760 = n3132 & n4759 ;
  assign n4761 = ~n4725 & ~n4760 ;
  assign n4762 = ~n4757 & n4761 ;
  assign n4763 = n929 & ~n4762 ;
  assign n4764 = ~n4724 & ~n4763 ;
  assign n4765 = \EAX_reg[10]/NET0131  & ~n3181 ;
  assign n4767 = n3132 & ~n3145 ;
  assign n4768 = n3430 & ~n4767 ;
  assign n4769 = \EAX_reg[10]/NET0131  & ~n4768 ;
  assign n4766 = \Datai[10]_pad  & n843 ;
  assign n4770 = n3144 & n4767 ;
  assign n4775 = \InstQueue_reg[2][2]/NET0131  & n474 ;
  assign n4776 = \InstQueue_reg[3][2]/NET0131  & n488 ;
  assign n4789 = ~n4775 & ~n4776 ;
  assign n4777 = \InstQueue_reg[6][2]/NET0131  & n472 ;
  assign n4778 = \InstQueue_reg[10][2]/NET0131  & n486 ;
  assign n4790 = ~n4777 & ~n4778 ;
  assign n4797 = n4789 & n4790 ;
  assign n4771 = \InstQueue_reg[0][2]/NET0131  & n470 ;
  assign n4772 = \InstQueue_reg[8][2]/NET0131  & n482 ;
  assign n4787 = ~n4771 & ~n4772 ;
  assign n4773 = \InstQueue_reg[12][2]/NET0131  & n461 ;
  assign n4774 = \InstQueue_reg[5][2]/NET0131  & n476 ;
  assign n4788 = ~n4773 & ~n4774 ;
  assign n4798 = n4787 & n4788 ;
  assign n4799 = n4797 & n4798 ;
  assign n4783 = \InstQueue_reg[14][2]/NET0131  & n468 ;
  assign n4784 = \InstQueue_reg[4][2]/NET0131  & n458 ;
  assign n4793 = ~n4783 & ~n4784 ;
  assign n4785 = \InstQueue_reg[15][2]/NET0131  & n465 ;
  assign n4786 = \InstQueue_reg[11][2]/NET0131  & n484 ;
  assign n4794 = ~n4785 & ~n4786 ;
  assign n4795 = n4793 & n4794 ;
  assign n4779 = \InstQueue_reg[7][2]/NET0131  & n490 ;
  assign n4780 = \InstQueue_reg[9][2]/NET0131  & n454 ;
  assign n4791 = ~n4779 & ~n4780 ;
  assign n4781 = \InstQueue_reg[13][2]/NET0131  & n492 ;
  assign n4782 = \InstQueue_reg[1][2]/NET0131  & n522 ;
  assign n4792 = ~n4781 & ~n4782 ;
  assign n4796 = n4791 & n4792 ;
  assign n4800 = n4795 & n4796 ;
  assign n4801 = n4799 & n4800 ;
  assign n4802 = n2937 & ~n4801 ;
  assign n4803 = ~n4770 & ~n4802 ;
  assign n4804 = ~n4766 & n4803 ;
  assign n4805 = ~n4769 & n4804 ;
  assign n4806 = n929 & ~n4805 ;
  assign n4807 = ~n4765 & ~n4806 ;
  assign n4808 = \EAX_reg[11]/NET0131  & ~n3181 ;
  assign n4810 = \EAX_reg[11]/NET0131  & ~n4768 ;
  assign n4809 = \Datai[11]_pad  & n843 ;
  assign n4815 = \InstQueue_reg[12][3]/NET0131  & n461 ;
  assign n4816 = \InstQueue_reg[3][3]/NET0131  & n488 ;
  assign n4829 = ~n4815 & ~n4816 ;
  assign n4817 = \InstQueue_reg[6][3]/NET0131  & n472 ;
  assign n4818 = \InstQueue_reg[10][3]/NET0131  & n486 ;
  assign n4830 = ~n4817 & ~n4818 ;
  assign n4837 = n4829 & n4830 ;
  assign n4811 = \InstQueue_reg[0][3]/NET0131  & n470 ;
  assign n4812 = \InstQueue_reg[8][3]/NET0131  & n482 ;
  assign n4827 = ~n4811 & ~n4812 ;
  assign n4813 = \InstQueue_reg[2][3]/NET0131  & n474 ;
  assign n4814 = \InstQueue_reg[5][3]/NET0131  & n476 ;
  assign n4828 = ~n4813 & ~n4814 ;
  assign n4838 = n4827 & n4828 ;
  assign n4839 = n4837 & n4838 ;
  assign n4823 = \InstQueue_reg[1][3]/NET0131  & n522 ;
  assign n4824 = \InstQueue_reg[4][3]/NET0131  & n458 ;
  assign n4833 = ~n4823 & ~n4824 ;
  assign n4825 = \InstQueue_reg[15][3]/NET0131  & n465 ;
  assign n4826 = \InstQueue_reg[11][3]/NET0131  & n484 ;
  assign n4834 = ~n4825 & ~n4826 ;
  assign n4835 = n4833 & n4834 ;
  assign n4819 = \InstQueue_reg[7][3]/NET0131  & n490 ;
  assign n4820 = \InstQueue_reg[9][3]/NET0131  & n454 ;
  assign n4831 = ~n4819 & ~n4820 ;
  assign n4821 = \InstQueue_reg[13][3]/NET0131  & n492 ;
  assign n4822 = \InstQueue_reg[14][3]/NET0131  & n468 ;
  assign n4832 = ~n4821 & ~n4822 ;
  assign n4836 = n4831 & n4832 ;
  assign n4840 = n4835 & n4836 ;
  assign n4841 = n4839 & n4840 ;
  assign n4842 = n2937 & ~n4841 ;
  assign n4843 = ~\EAX_reg[11]/NET0131  & n3145 ;
  assign n4844 = n3132 & n4843 ;
  assign n4845 = ~n4842 & ~n4844 ;
  assign n4846 = ~n4809 & n4845 ;
  assign n4847 = ~n4810 & n4846 ;
  assign n4848 = n929 & ~n4847 ;
  assign n4849 = ~n4808 & ~n4848 ;
  assign n4850 = \EBX_reg[25]/NET0131  & ~n3181 ;
  assign n4852 = \EBX_reg[24]/NET0131  & n3490 ;
  assign n4853 = n797 & ~n4852 ;
  assign n4854 = ~n3465 & ~n4853 ;
  assign n4855 = \EBX_reg[25]/NET0131  & ~n4854 ;
  assign n4851 = n3463 & n4307 ;
  assign n4856 = ~\EBX_reg[25]/NET0131  & n797 ;
  assign n4857 = n4852 & n4856 ;
  assign n4858 = ~n4851 & ~n4857 ;
  assign n4859 = ~n4855 & n4858 ;
  assign n4860 = n929 & ~n4859 ;
  assign n4861 = ~n4850 & ~n4860 ;
  assign n4862 = \EAX_reg[12]/NET0131  & ~n3181 ;
  assign n4863 = n3132 & ~n3146 ;
  assign n4864 = ~n3135 & ~n4863 ;
  assign n4865 = \EAX_reg[12]/NET0131  & ~n4864 ;
  assign n4900 = \EAX_reg[12]/NET0131  & ~n846 ;
  assign n4901 = ~n3657 & ~n4900 ;
  assign n4902 = ~n841 & ~n4901 ;
  assign n4866 = ~\EAX_reg[12]/NET0131  & n3132 ;
  assign n4867 = n3146 & n4866 ;
  assign n4872 = \InstQueue_reg[14][4]/NET0131  & n468 ;
  assign n4873 = \InstQueue_reg[3][4]/NET0131  & n488 ;
  assign n4886 = ~n4872 & ~n4873 ;
  assign n4874 = \InstQueue_reg[7][4]/NET0131  & n490 ;
  assign n4875 = \InstQueue_reg[10][4]/NET0131  & n486 ;
  assign n4887 = ~n4874 & ~n4875 ;
  assign n4894 = n4886 & n4887 ;
  assign n4868 = \InstQueue_reg[0][4]/NET0131  & n470 ;
  assign n4869 = \InstQueue_reg[8][4]/NET0131  & n482 ;
  assign n4884 = ~n4868 & ~n4869 ;
  assign n4870 = \InstQueue_reg[6][4]/NET0131  & n472 ;
  assign n4871 = \InstQueue_reg[5][4]/NET0131  & n476 ;
  assign n4885 = ~n4870 & ~n4871 ;
  assign n4895 = n4884 & n4885 ;
  assign n4896 = n4894 & n4895 ;
  assign n4880 = \InstQueue_reg[12][4]/NET0131  & n461 ;
  assign n4881 = \InstQueue_reg[4][4]/NET0131  & n458 ;
  assign n4890 = ~n4880 & ~n4881 ;
  assign n4882 = \InstQueue_reg[15][4]/NET0131  & n465 ;
  assign n4883 = \InstQueue_reg[11][4]/NET0131  & n484 ;
  assign n4891 = ~n4882 & ~n4883 ;
  assign n4892 = n4890 & n4891 ;
  assign n4876 = \InstQueue_reg[1][4]/NET0131  & n522 ;
  assign n4877 = \InstQueue_reg[9][4]/NET0131  & n454 ;
  assign n4888 = ~n4876 & ~n4877 ;
  assign n4878 = \InstQueue_reg[13][4]/NET0131  & n492 ;
  assign n4879 = \InstQueue_reg[2][4]/NET0131  & n474 ;
  assign n4889 = ~n4878 & ~n4879 ;
  assign n4893 = n4888 & n4889 ;
  assign n4897 = n4892 & n4893 ;
  assign n4898 = n4896 & n4897 ;
  assign n4899 = n2937 & ~n4898 ;
  assign n4903 = ~n4867 & ~n4899 ;
  assign n4904 = ~n4902 & n4903 ;
  assign n4905 = ~n4865 & n4904 ;
  assign n4906 = n929 & ~n4905 ;
  assign n4907 = ~n4862 & ~n4906 ;
  assign n4908 = \EAX_reg[13]/NET0131  & ~n3181 ;
  assign n4910 = n3132 & ~n3147 ;
  assign n4911 = n3430 & ~n4910 ;
  assign n4912 = \EAX_reg[13]/NET0131  & ~n4911 ;
  assign n4909 = \Datai[13]_pad  & n843 ;
  assign n4917 = \InstQueue_reg[2][5]/NET0131  & n474 ;
  assign n4918 = \InstQueue_reg[4][5]/NET0131  & n458 ;
  assign n4931 = ~n4917 & ~n4918 ;
  assign n4919 = \InstQueue_reg[6][5]/NET0131  & n472 ;
  assign n4920 = \InstQueue_reg[8][5]/NET0131  & n482 ;
  assign n4932 = ~n4919 & ~n4920 ;
  assign n4939 = n4931 & n4932 ;
  assign n4913 = \InstQueue_reg[0][5]/NET0131  & n470 ;
  assign n4914 = \InstQueue_reg[11][5]/NET0131  & n484 ;
  assign n4929 = ~n4913 & ~n4914 ;
  assign n4915 = \InstQueue_reg[15][5]/NET0131  & n465 ;
  assign n4916 = \InstQueue_reg[5][5]/NET0131  & n476 ;
  assign n4930 = ~n4915 & ~n4916 ;
  assign n4940 = n4929 & n4930 ;
  assign n4941 = n4939 & n4940 ;
  assign n4925 = \InstQueue_reg[1][5]/NET0131  & n522 ;
  assign n4926 = \InstQueue_reg[3][5]/NET0131  & n488 ;
  assign n4935 = ~n4925 & ~n4926 ;
  assign n4927 = \InstQueue_reg[12][5]/NET0131  & n461 ;
  assign n4928 = \InstQueue_reg[9][5]/NET0131  & n454 ;
  assign n4936 = ~n4927 & ~n4928 ;
  assign n4937 = n4935 & n4936 ;
  assign n4921 = \InstQueue_reg[7][5]/NET0131  & n490 ;
  assign n4922 = \InstQueue_reg[14][5]/NET0131  & n468 ;
  assign n4933 = ~n4921 & ~n4922 ;
  assign n4923 = \InstQueue_reg[10][5]/NET0131  & n486 ;
  assign n4924 = \InstQueue_reg[13][5]/NET0131  & n492 ;
  assign n4934 = ~n4923 & ~n4924 ;
  assign n4938 = n4933 & n4934 ;
  assign n4942 = n4937 & n4938 ;
  assign n4943 = n4941 & n4942 ;
  assign n4944 = n2937 & ~n4943 ;
  assign n4945 = ~\EAX_reg[13]/NET0131  & n3132 ;
  assign n4946 = n3147 & n4945 ;
  assign n4947 = ~n4944 & ~n4946 ;
  assign n4948 = ~n4909 & n4947 ;
  assign n4949 = ~n4912 & n4948 ;
  assign n4950 = n929 & ~n4949 ;
  assign n4951 = ~n4908 & ~n4950 ;
  assign n4984 = \EAX_reg[14]/NET0131  & ~n3430 ;
  assign n4985 = ~\EAX_reg[14]/NET0131  & ~n3148 ;
  assign n4986 = n3132 & ~n3149 ;
  assign n4987 = ~n4985 & n4986 ;
  assign n4956 = \InstQueue_reg[12][6]/NET0131  & n461 ;
  assign n4957 = \InstQueue_reg[3][6]/NET0131  & n488 ;
  assign n4970 = ~n4956 & ~n4957 ;
  assign n4958 = \InstQueue_reg[6][6]/NET0131  & n472 ;
  assign n4959 = \InstQueue_reg[10][6]/NET0131  & n486 ;
  assign n4971 = ~n4958 & ~n4959 ;
  assign n4978 = n4970 & n4971 ;
  assign n4952 = \InstQueue_reg[0][6]/NET0131  & n470 ;
  assign n4953 = \InstQueue_reg[8][6]/NET0131  & n482 ;
  assign n4968 = ~n4952 & ~n4953 ;
  assign n4954 = \InstQueue_reg[2][6]/NET0131  & n474 ;
  assign n4955 = \InstQueue_reg[5][6]/NET0131  & n476 ;
  assign n4969 = ~n4954 & ~n4955 ;
  assign n4979 = n4968 & n4969 ;
  assign n4980 = n4978 & n4979 ;
  assign n4964 = \InstQueue_reg[1][6]/NET0131  & n522 ;
  assign n4965 = \InstQueue_reg[4][6]/NET0131  & n458 ;
  assign n4974 = ~n4964 & ~n4965 ;
  assign n4966 = \InstQueue_reg[15][6]/NET0131  & n465 ;
  assign n4967 = \InstQueue_reg[11][6]/NET0131  & n484 ;
  assign n4975 = ~n4966 & ~n4967 ;
  assign n4976 = n4974 & n4975 ;
  assign n4960 = \InstQueue_reg[7][6]/NET0131  & n490 ;
  assign n4961 = \InstQueue_reg[9][6]/NET0131  & n454 ;
  assign n4972 = ~n4960 & ~n4961 ;
  assign n4962 = \InstQueue_reg[13][6]/NET0131  & n492 ;
  assign n4963 = \InstQueue_reg[14][6]/NET0131  & n468 ;
  assign n4973 = ~n4962 & ~n4963 ;
  assign n4977 = n4972 & n4973 ;
  assign n4981 = n4976 & n4977 ;
  assign n4982 = n4980 & n4981 ;
  assign n4983 = n2937 & ~n4982 ;
  assign n4988 = \Datai[14]_pad  & n843 ;
  assign n4989 = ~n4983 & ~n4988 ;
  assign n4990 = ~n4987 & n4989 ;
  assign n4991 = ~n4984 & n4990 ;
  assign n4992 = n929 & ~n4991 ;
  assign n4993 = \EAX_reg[14]/NET0131  & ~n3181 ;
  assign n4994 = ~n4992 & ~n4993 ;
  assign n4995 = \EAX_reg[15]/NET0131  & ~n3181 ;
  assign n4998 = n3430 & ~n4986 ;
  assign n4999 = \EAX_reg[15]/NET0131  & ~n4998 ;
  assign n5032 = ~\EAX_reg[15]/NET0131  & n3132 ;
  assign n5033 = n3149 & n5032 ;
  assign n4996 = \Datai[15]_pad  & n846 ;
  assign n4997 = ~n841 & n4996 ;
  assign n5004 = \InstQueue_reg[12][7]/NET0131  & n461 ;
  assign n5005 = \InstQueue_reg[3][7]/NET0131  & n488 ;
  assign n5018 = ~n5004 & ~n5005 ;
  assign n5006 = \InstQueue_reg[6][7]/NET0131  & n472 ;
  assign n5007 = \InstQueue_reg[10][7]/NET0131  & n486 ;
  assign n5019 = ~n5006 & ~n5007 ;
  assign n5026 = n5018 & n5019 ;
  assign n5000 = \InstQueue_reg[0][7]/NET0131  & n470 ;
  assign n5001 = \InstQueue_reg[8][7]/NET0131  & n482 ;
  assign n5016 = ~n5000 & ~n5001 ;
  assign n5002 = \InstQueue_reg[2][7]/NET0131  & n474 ;
  assign n5003 = \InstQueue_reg[5][7]/NET0131  & n476 ;
  assign n5017 = ~n5002 & ~n5003 ;
  assign n5027 = n5016 & n5017 ;
  assign n5028 = n5026 & n5027 ;
  assign n5012 = \InstQueue_reg[1][7]/NET0131  & n522 ;
  assign n5013 = \InstQueue_reg[4][7]/NET0131  & n458 ;
  assign n5022 = ~n5012 & ~n5013 ;
  assign n5014 = \InstQueue_reg[15][7]/NET0131  & n465 ;
  assign n5015 = \InstQueue_reg[11][7]/NET0131  & n484 ;
  assign n5023 = ~n5014 & ~n5015 ;
  assign n5024 = n5022 & n5023 ;
  assign n5008 = \InstQueue_reg[7][7]/NET0131  & n490 ;
  assign n5009 = \InstQueue_reg[9][7]/NET0131  & n454 ;
  assign n5020 = ~n5008 & ~n5009 ;
  assign n5010 = \InstQueue_reg[13][7]/NET0131  & n492 ;
  assign n5011 = \InstQueue_reg[14][7]/NET0131  & n468 ;
  assign n5021 = ~n5010 & ~n5011 ;
  assign n5025 = n5020 & n5021 ;
  assign n5029 = n5024 & n5025 ;
  assign n5030 = n5028 & n5029 ;
  assign n5031 = n2937 & ~n5030 ;
  assign n5034 = ~n4997 & ~n5031 ;
  assign n5035 = ~n5033 & n5034 ;
  assign n5036 = ~n4999 & n5035 ;
  assign n5037 = n929 & ~n5036 ;
  assign n5038 = ~n4995 & ~n5037 ;
  assign n5044 = ~\Datai[27]_pad  & ~n3898 ;
  assign n5045 = ~n3899 & ~n5044 ;
  assign n5046 = n3871 & n5045 ;
  assign n5047 = ~\Datai[19]_pad  & ~n3907 ;
  assign n5048 = ~n3908 & ~n5047 ;
  assign n5049 = n3914 & n5048 ;
  assign n5050 = ~n5046 & ~n5049 ;
  assign n5051 = \DataWidth_reg[1]/NET0131  & ~n5050 ;
  assign n5039 = \Datai[3]_pad  & ~n3863 ;
  assign n5040 = \InstQueue_reg[0][3]/NET0131  & ~n3859 ;
  assign n5041 = ~n3862 & n5040 ;
  assign n5042 = ~n5039 & ~n5041 ;
  assign n5052 = ~n3919 & ~n5042 ;
  assign n5053 = ~n5051 & ~n5052 ;
  assign n5054 = n933 & ~n5053 ;
  assign n5055 = ~n540 & n3859 ;
  assign n5056 = ~n5040 & ~n5055 ;
  assign n5057 = n965 & ~n5056 ;
  assign n5043 = n1867 & ~n5042 ;
  assign n5058 = \InstQueue_reg[0][3]/NET0131  & ~n3929 ;
  assign n5059 = ~n5043 & ~n5058 ;
  assign n5060 = ~n5057 & n5059 ;
  assign n5061 = ~n5054 & n5060 ;
  assign n5067 = ~\Datai[30]_pad  & ~n4332 ;
  assign n5068 = ~n4333 & ~n5067 ;
  assign n5069 = n3871 & n5068 ;
  assign n5070 = ~\Datai[22]_pad  & ~n4336 ;
  assign n5071 = ~n4337 & ~n5070 ;
  assign n5072 = n3914 & n5071 ;
  assign n5073 = ~n5069 & ~n5072 ;
  assign n5074 = \DataWidth_reg[1]/NET0131  & ~n5073 ;
  assign n5062 = \Datai[6]_pad  & ~n3863 ;
  assign n5063 = \InstQueue_reg[0][6]/NET0131  & ~n3859 ;
  assign n5064 = ~n3862 & n5063 ;
  assign n5065 = ~n5062 & ~n5064 ;
  assign n5075 = ~n3919 & ~n5065 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = n933 & ~n5076 ;
  assign n5078 = ~n731 & n3859 ;
  assign n5079 = ~n5063 & ~n5078 ;
  assign n5080 = n965 & ~n5079 ;
  assign n5066 = n1867 & ~n5065 ;
  assign n5081 = \InstQueue_reg[0][6]/NET0131  & ~n3929 ;
  assign n5082 = ~n5066 & ~n5081 ;
  assign n5083 = ~n5080 & n5082 ;
  assign n5084 = ~n5077 & n5083 ;
  assign n5090 = n3944 & n5045 ;
  assign n5091 = n3946 & n5048 ;
  assign n5092 = ~n5090 & ~n5091 ;
  assign n5093 = \DataWidth_reg[1]/NET0131  & ~n5092 ;
  assign n5085 = \Datai[3]_pad  & ~n3938 ;
  assign n5086 = \InstQueue_reg[10][3]/NET0131  & ~n3935 ;
  assign n5087 = ~n3937 & n5086 ;
  assign n5088 = ~n5085 & ~n5087 ;
  assign n5094 = ~n3951 & ~n5088 ;
  assign n5095 = ~n5093 & ~n5094 ;
  assign n5096 = n933 & ~n5095 ;
  assign n5097 = ~n540 & n3935 ;
  assign n5098 = ~n5086 & ~n5097 ;
  assign n5099 = n965 & ~n5098 ;
  assign n5089 = n1867 & ~n5088 ;
  assign n5100 = \InstQueue_reg[10][3]/NET0131  & ~n3929 ;
  assign n5101 = ~n5089 & ~n5100 ;
  assign n5102 = ~n5099 & n5101 ;
  assign n5103 = ~n5096 & n5102 ;
  assign n5109 = n3944 & n5068 ;
  assign n5110 = n3946 & n5071 ;
  assign n5111 = ~n5109 & ~n5110 ;
  assign n5112 = \DataWidth_reg[1]/NET0131  & ~n5111 ;
  assign n5104 = \Datai[6]_pad  & ~n3938 ;
  assign n5105 = \InstQueue_reg[10][6]/NET0131  & ~n3935 ;
  assign n5106 = ~n3937 & n5105 ;
  assign n5107 = ~n5104 & ~n5106 ;
  assign n5113 = ~n3951 & ~n5107 ;
  assign n5114 = ~n5112 & ~n5113 ;
  assign n5115 = n933 & ~n5114 ;
  assign n5116 = ~n731 & n3935 ;
  assign n5117 = ~n5105 & ~n5116 ;
  assign n5118 = n965 & ~n5117 ;
  assign n5108 = n1867 & ~n5107 ;
  assign n5119 = \InstQueue_reg[10][6]/NET0131  & ~n3929 ;
  assign n5120 = ~n5108 & ~n5119 ;
  assign n5121 = ~n5118 & n5120 ;
  assign n5122 = ~n5115 & n5121 ;
  assign n5128 = n3946 & n5045 ;
  assign n5129 = n3937 & n5048 ;
  assign n5130 = ~n5128 & ~n5129 ;
  assign n5131 = \DataWidth_reg[1]/NET0131  & ~n5130 ;
  assign n5123 = \Datai[3]_pad  & ~n3964 ;
  assign n5124 = \InstQueue_reg[11][3]/NET0131  & ~n3963 ;
  assign n5125 = ~n3935 & n5124 ;
  assign n5126 = ~n5123 & ~n5125 ;
  assign n5132 = ~n3975 & ~n5126 ;
  assign n5133 = ~n5131 & ~n5132 ;
  assign n5134 = n933 & ~n5133 ;
  assign n5135 = ~n540 & n3963 ;
  assign n5136 = ~n5124 & ~n5135 ;
  assign n5137 = n965 & ~n5136 ;
  assign n5127 = n1867 & ~n5126 ;
  assign n5138 = \InstQueue_reg[11][3]/NET0131  & ~n3929 ;
  assign n5139 = ~n5127 & ~n5138 ;
  assign n5140 = ~n5137 & n5139 ;
  assign n5141 = ~n5134 & n5140 ;
  assign n5147 = n3946 & n5068 ;
  assign n5148 = n3937 & n5071 ;
  assign n5149 = ~n5147 & ~n5148 ;
  assign n5150 = \DataWidth_reg[1]/NET0131  & ~n5149 ;
  assign n5142 = \Datai[6]_pad  & ~n3964 ;
  assign n5143 = \InstQueue_reg[11][6]/NET0131  & ~n3963 ;
  assign n5144 = ~n3935 & n5143 ;
  assign n5145 = ~n5142 & ~n5144 ;
  assign n5151 = ~n3975 & ~n5145 ;
  assign n5152 = ~n5150 & ~n5151 ;
  assign n5153 = n933 & ~n5152 ;
  assign n5154 = ~n731 & n3963 ;
  assign n5155 = ~n5143 & ~n5154 ;
  assign n5156 = n965 & ~n5155 ;
  assign n5146 = n1867 & ~n5145 ;
  assign n5157 = \InstQueue_reg[11][6]/NET0131  & ~n3929 ;
  assign n5158 = ~n5146 & ~n5157 ;
  assign n5159 = ~n5156 & n5158 ;
  assign n5160 = ~n5153 & n5159 ;
  assign n5166 = n3937 & n5045 ;
  assign n5167 = n3935 & n5048 ;
  assign n5168 = ~n5166 & ~n5167 ;
  assign n5169 = \DataWidth_reg[1]/NET0131  & ~n5168 ;
  assign n5161 = \Datai[3]_pad  & ~n3988 ;
  assign n5162 = \InstQueue_reg[12][3]/NET0131  & ~n3987 ;
  assign n5163 = ~n3963 & n5162 ;
  assign n5164 = ~n5161 & ~n5163 ;
  assign n5170 = ~n3998 & ~n5164 ;
  assign n5171 = ~n5169 & ~n5170 ;
  assign n5172 = n933 & ~n5171 ;
  assign n5173 = ~n540 & n3987 ;
  assign n5174 = ~n5162 & ~n5173 ;
  assign n5175 = n965 & ~n5174 ;
  assign n5165 = n1867 & ~n5164 ;
  assign n5176 = \InstQueue_reg[12][3]/NET0131  & ~n3929 ;
  assign n5177 = ~n5165 & ~n5176 ;
  assign n5178 = ~n5175 & n5177 ;
  assign n5179 = ~n5172 & n5178 ;
  assign n5185 = n3937 & n5068 ;
  assign n5186 = n3935 & n5071 ;
  assign n5187 = ~n5185 & ~n5186 ;
  assign n5188 = \DataWidth_reg[1]/NET0131  & ~n5187 ;
  assign n5180 = \Datai[6]_pad  & ~n3988 ;
  assign n5181 = \InstQueue_reg[12][6]/NET0131  & ~n3987 ;
  assign n5182 = ~n3963 & n5181 ;
  assign n5183 = ~n5180 & ~n5182 ;
  assign n5189 = ~n3998 & ~n5183 ;
  assign n5190 = ~n5188 & ~n5189 ;
  assign n5191 = n933 & ~n5190 ;
  assign n5192 = ~n731 & n3987 ;
  assign n5193 = ~n5181 & ~n5192 ;
  assign n5194 = n965 & ~n5193 ;
  assign n5184 = n1867 & ~n5183 ;
  assign n5195 = \InstQueue_reg[12][6]/NET0131  & ~n3929 ;
  assign n5196 = ~n5184 & ~n5195 ;
  assign n5197 = ~n5194 & n5196 ;
  assign n5198 = ~n5191 & n5197 ;
  assign n5204 = n3935 & n5045 ;
  assign n5205 = n3963 & n5048 ;
  assign n5206 = ~n5204 & ~n5205 ;
  assign n5207 = \DataWidth_reg[1]/NET0131  & ~n5206 ;
  assign n5199 = \Datai[3]_pad  & ~n4009 ;
  assign n5200 = \InstQueue_reg[13][3]/NET0131  & ~n3871 ;
  assign n5201 = ~n3987 & n5200 ;
  assign n5202 = ~n5199 & ~n5201 ;
  assign n5208 = ~n4019 & ~n5202 ;
  assign n5209 = ~n5207 & ~n5208 ;
  assign n5210 = n933 & ~n5209 ;
  assign n5211 = ~n540 & n3871 ;
  assign n5212 = ~n5200 & ~n5211 ;
  assign n5213 = n965 & ~n5212 ;
  assign n5203 = n1867 & ~n5202 ;
  assign n5214 = \InstQueue_reg[13][3]/NET0131  & ~n3929 ;
  assign n5215 = ~n5203 & ~n5214 ;
  assign n5216 = ~n5213 & n5215 ;
  assign n5217 = ~n5210 & n5216 ;
  assign n5223 = n3935 & n5068 ;
  assign n5224 = n3963 & n5071 ;
  assign n5225 = ~n5223 & ~n5224 ;
  assign n5226 = \DataWidth_reg[1]/NET0131  & ~n5225 ;
  assign n5218 = \Datai[6]_pad  & ~n4009 ;
  assign n5219 = \InstQueue_reg[13][6]/NET0131  & ~n3871 ;
  assign n5220 = ~n3987 & n5219 ;
  assign n5221 = ~n5218 & ~n5220 ;
  assign n5227 = ~n4019 & ~n5221 ;
  assign n5228 = ~n5226 & ~n5227 ;
  assign n5229 = n933 & ~n5228 ;
  assign n5230 = ~n731 & n3871 ;
  assign n5231 = ~n5219 & ~n5230 ;
  assign n5232 = n965 & ~n5231 ;
  assign n5222 = n1867 & ~n5221 ;
  assign n5233 = \InstQueue_reg[13][6]/NET0131  & ~n3929 ;
  assign n5234 = ~n5222 & ~n5233 ;
  assign n5235 = ~n5232 & n5234 ;
  assign n5236 = ~n5229 & n5235 ;
  assign n5242 = n3963 & n5045 ;
  assign n5243 = n3987 & n5048 ;
  assign n5244 = ~n5242 & ~n5243 ;
  assign n5245 = \DataWidth_reg[1]/NET0131  & ~n5244 ;
  assign n5237 = \Datai[3]_pad  & ~n3918 ;
  assign n5238 = \InstQueue_reg[14][3]/NET0131  & ~n3914 ;
  assign n5239 = ~n3871 & n5238 ;
  assign n5240 = ~n5237 & ~n5239 ;
  assign n5246 = ~n4039 & ~n5240 ;
  assign n5247 = ~n5245 & ~n5246 ;
  assign n5248 = n933 & ~n5247 ;
  assign n5249 = ~n540 & n3914 ;
  assign n5250 = ~n5238 & ~n5249 ;
  assign n5251 = n965 & ~n5250 ;
  assign n5241 = n1867 & ~n5240 ;
  assign n5252 = \InstQueue_reg[14][3]/NET0131  & ~n3929 ;
  assign n5253 = ~n5241 & ~n5252 ;
  assign n5254 = ~n5251 & n5253 ;
  assign n5255 = ~n5248 & n5254 ;
  assign n5261 = n3963 & n5068 ;
  assign n5262 = n3987 & n5071 ;
  assign n5263 = ~n5261 & ~n5262 ;
  assign n5264 = \DataWidth_reg[1]/NET0131  & ~n5263 ;
  assign n5256 = \Datai[6]_pad  & ~n3918 ;
  assign n5257 = \InstQueue_reg[14][6]/NET0131  & ~n3914 ;
  assign n5258 = ~n3871 & n5257 ;
  assign n5259 = ~n5256 & ~n5258 ;
  assign n5265 = ~n4039 & ~n5259 ;
  assign n5266 = ~n5264 & ~n5265 ;
  assign n5267 = n933 & ~n5266 ;
  assign n5268 = ~n731 & n3914 ;
  assign n5269 = ~n5257 & ~n5268 ;
  assign n5270 = n965 & ~n5269 ;
  assign n5260 = n1867 & ~n5259 ;
  assign n5271 = \InstQueue_reg[14][6]/NET0131  & ~n3929 ;
  assign n5272 = ~n5260 & ~n5271 ;
  assign n5273 = ~n5270 & n5272 ;
  assign n5274 = ~n5267 & n5273 ;
  assign n5280 = n3987 & n5045 ;
  assign n5281 = n3871 & n5048 ;
  assign n5282 = ~n5280 & ~n5281 ;
  assign n5283 = \DataWidth_reg[1]/NET0131  & ~n5282 ;
  assign n5275 = \Datai[3]_pad  & ~n4050 ;
  assign n5276 = \InstQueue_reg[15][3]/NET0131  & ~n3862 ;
  assign n5277 = ~n3914 & n5276 ;
  assign n5278 = ~n5275 & ~n5277 ;
  assign n5284 = ~n4060 & ~n5278 ;
  assign n5285 = ~n5283 & ~n5284 ;
  assign n5286 = n933 & ~n5285 ;
  assign n5287 = ~n540 & n3862 ;
  assign n5288 = ~n5276 & ~n5287 ;
  assign n5289 = n965 & ~n5288 ;
  assign n5279 = n1867 & ~n5278 ;
  assign n5290 = \InstQueue_reg[15][3]/NET0131  & ~n3929 ;
  assign n5291 = ~n5279 & ~n5290 ;
  assign n5292 = ~n5289 & n5291 ;
  assign n5293 = ~n5286 & n5292 ;
  assign n5299 = n3987 & n5068 ;
  assign n5300 = n3871 & n5071 ;
  assign n5301 = ~n5299 & ~n5300 ;
  assign n5302 = \DataWidth_reg[1]/NET0131  & ~n5301 ;
  assign n5294 = \Datai[6]_pad  & ~n4050 ;
  assign n5295 = \InstQueue_reg[15][6]/NET0131  & ~n3862 ;
  assign n5296 = ~n3914 & n5295 ;
  assign n5297 = ~n5294 & ~n5296 ;
  assign n5303 = ~n4060 & ~n5297 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = n933 & ~n5304 ;
  assign n5306 = ~n731 & n3862 ;
  assign n5307 = ~n5295 & ~n5306 ;
  assign n5308 = n965 & ~n5307 ;
  assign n5298 = n1867 & ~n5297 ;
  assign n5309 = \InstQueue_reg[15][6]/NET0131  & ~n3929 ;
  assign n5310 = ~n5298 & ~n5309 ;
  assign n5311 = ~n5308 & n5310 ;
  assign n5312 = ~n5305 & n5311 ;
  assign n5318 = n3914 & n5045 ;
  assign n5319 = n3862 & n5048 ;
  assign n5320 = ~n5318 & ~n5319 ;
  assign n5321 = \DataWidth_reg[1]/NET0131  & ~n5320 ;
  assign n5313 = \Datai[3]_pad  & ~n4072 ;
  assign n5314 = \InstQueue_reg[1][3]/NET0131  & ~n4071 ;
  assign n5315 = ~n3859 & n5314 ;
  assign n5316 = ~n5313 & ~n5315 ;
  assign n5322 = ~n4082 & ~n5316 ;
  assign n5323 = ~n5321 & ~n5322 ;
  assign n5324 = n933 & ~n5323 ;
  assign n5325 = ~n540 & n4071 ;
  assign n5326 = ~n5314 & ~n5325 ;
  assign n5327 = n965 & ~n5326 ;
  assign n5317 = n1867 & ~n5316 ;
  assign n5328 = \InstQueue_reg[1][3]/NET0131  & ~n3929 ;
  assign n5329 = ~n5317 & ~n5328 ;
  assign n5330 = ~n5327 & n5329 ;
  assign n5331 = ~n5324 & n5330 ;
  assign n5337 = n3914 & n5068 ;
  assign n5338 = n3862 & n5071 ;
  assign n5339 = ~n5337 & ~n5338 ;
  assign n5340 = \DataWidth_reg[1]/NET0131  & ~n5339 ;
  assign n5332 = \Datai[6]_pad  & ~n4072 ;
  assign n5333 = \InstQueue_reg[1][6]/NET0131  & ~n4071 ;
  assign n5334 = ~n3859 & n5333 ;
  assign n5335 = ~n5332 & ~n5334 ;
  assign n5341 = ~n4082 & ~n5335 ;
  assign n5342 = ~n5340 & ~n5341 ;
  assign n5343 = n933 & ~n5342 ;
  assign n5344 = ~n731 & n4071 ;
  assign n5345 = ~n5333 & ~n5344 ;
  assign n5346 = n965 & ~n5345 ;
  assign n5336 = n1867 & ~n5335 ;
  assign n5347 = \InstQueue_reg[1][6]/NET0131  & ~n3929 ;
  assign n5348 = ~n5336 & ~n5347 ;
  assign n5349 = ~n5346 & n5348 ;
  assign n5350 = ~n5343 & n5349 ;
  assign n5356 = n3859 & n5048 ;
  assign n5357 = n3862 & n5045 ;
  assign n5358 = ~n5356 & ~n5357 ;
  assign n5359 = \DataWidth_reg[1]/NET0131  & ~n5358 ;
  assign n5351 = \Datai[3]_pad  & ~n4094 ;
  assign n5352 = \InstQueue_reg[2][3]/NET0131  & ~n4093 ;
  assign n5353 = ~n4071 & n5352 ;
  assign n5354 = ~n5351 & ~n5353 ;
  assign n5360 = ~n4104 & ~n5354 ;
  assign n5361 = ~n5359 & ~n5360 ;
  assign n5362 = n933 & ~n5361 ;
  assign n5363 = ~n540 & n4093 ;
  assign n5364 = ~n5352 & ~n5363 ;
  assign n5365 = n965 & ~n5364 ;
  assign n5355 = n1867 & ~n5354 ;
  assign n5366 = \InstQueue_reg[2][3]/NET0131  & ~n3929 ;
  assign n5367 = ~n5355 & ~n5366 ;
  assign n5368 = ~n5365 & n5367 ;
  assign n5369 = ~n5362 & n5368 ;
  assign n5375 = n3859 & n5071 ;
  assign n5376 = n3862 & n5068 ;
  assign n5377 = ~n5375 & ~n5376 ;
  assign n5378 = \DataWidth_reg[1]/NET0131  & ~n5377 ;
  assign n5370 = \Datai[6]_pad  & ~n4094 ;
  assign n5371 = \InstQueue_reg[2][6]/NET0131  & ~n4093 ;
  assign n5372 = ~n4071 & n5371 ;
  assign n5373 = ~n5370 & ~n5372 ;
  assign n5379 = ~n4104 & ~n5373 ;
  assign n5380 = ~n5378 & ~n5379 ;
  assign n5381 = n933 & ~n5380 ;
  assign n5382 = ~n731 & n4093 ;
  assign n5383 = ~n5371 & ~n5382 ;
  assign n5384 = n965 & ~n5383 ;
  assign n5374 = n1867 & ~n5373 ;
  assign n5385 = \InstQueue_reg[2][6]/NET0131  & ~n3929 ;
  assign n5386 = ~n5374 & ~n5385 ;
  assign n5387 = ~n5384 & n5386 ;
  assign n5388 = ~n5381 & n5387 ;
  assign n5394 = n3859 & n5045 ;
  assign n5395 = n4071 & n5048 ;
  assign n5396 = ~n5394 & ~n5395 ;
  assign n5397 = \DataWidth_reg[1]/NET0131  & ~n5396 ;
  assign n5389 = \Datai[3]_pad  & ~n4116 ;
  assign n5390 = \InstQueue_reg[3][3]/NET0131  & ~n4115 ;
  assign n5391 = ~n4093 & n5390 ;
  assign n5392 = ~n5389 & ~n5391 ;
  assign n5398 = ~n4126 & ~n5392 ;
  assign n5399 = ~n5397 & ~n5398 ;
  assign n5400 = n933 & ~n5399 ;
  assign n5401 = ~n540 & n4115 ;
  assign n5402 = ~n5390 & ~n5401 ;
  assign n5403 = n965 & ~n5402 ;
  assign n5393 = n1867 & ~n5392 ;
  assign n5404 = \InstQueue_reg[3][3]/NET0131  & ~n3929 ;
  assign n5405 = ~n5393 & ~n5404 ;
  assign n5406 = ~n5403 & n5405 ;
  assign n5407 = ~n5400 & n5406 ;
  assign n5413 = n3859 & n5068 ;
  assign n5414 = n4071 & n5071 ;
  assign n5415 = ~n5413 & ~n5414 ;
  assign n5416 = \DataWidth_reg[1]/NET0131  & ~n5415 ;
  assign n5408 = \Datai[6]_pad  & ~n4116 ;
  assign n5409 = \InstQueue_reg[3][6]/NET0131  & ~n4115 ;
  assign n5410 = ~n4093 & n5409 ;
  assign n5411 = ~n5408 & ~n5410 ;
  assign n5417 = ~n4126 & ~n5411 ;
  assign n5418 = ~n5416 & ~n5417 ;
  assign n5419 = n933 & ~n5418 ;
  assign n5420 = ~n731 & n4115 ;
  assign n5421 = ~n5409 & ~n5420 ;
  assign n5422 = n965 & ~n5421 ;
  assign n5412 = n1867 & ~n5411 ;
  assign n5423 = \InstQueue_reg[3][6]/NET0131  & ~n3929 ;
  assign n5424 = ~n5412 & ~n5423 ;
  assign n5425 = ~n5422 & n5424 ;
  assign n5426 = ~n5419 & n5425 ;
  assign n5432 = n4071 & n5045 ;
  assign n5433 = n4093 & n5048 ;
  assign n5434 = ~n5432 & ~n5433 ;
  assign n5435 = \DataWidth_reg[1]/NET0131  & ~n5434 ;
  assign n5427 = \Datai[3]_pad  & ~n4138 ;
  assign n5428 = \InstQueue_reg[4][3]/NET0131  & ~n4137 ;
  assign n5429 = ~n4115 & n5428 ;
  assign n5430 = ~n5427 & ~n5429 ;
  assign n5436 = ~n4148 & ~n5430 ;
  assign n5437 = ~n5435 & ~n5436 ;
  assign n5438 = n933 & ~n5437 ;
  assign n5439 = ~n540 & n4137 ;
  assign n5440 = ~n5428 & ~n5439 ;
  assign n5441 = n965 & ~n5440 ;
  assign n5431 = n1867 & ~n5430 ;
  assign n5442 = \InstQueue_reg[4][3]/NET0131  & ~n3929 ;
  assign n5443 = ~n5431 & ~n5442 ;
  assign n5444 = ~n5441 & n5443 ;
  assign n5445 = ~n5438 & n5444 ;
  assign n5451 = n4071 & n5068 ;
  assign n5452 = n4093 & n5071 ;
  assign n5453 = ~n5451 & ~n5452 ;
  assign n5454 = \DataWidth_reg[1]/NET0131  & ~n5453 ;
  assign n5446 = \Datai[6]_pad  & ~n4138 ;
  assign n5447 = \InstQueue_reg[4][6]/NET0131  & ~n4137 ;
  assign n5448 = ~n4115 & n5447 ;
  assign n5449 = ~n5446 & ~n5448 ;
  assign n5455 = ~n4148 & ~n5449 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5457 = n933 & ~n5456 ;
  assign n5458 = ~n731 & n4137 ;
  assign n5459 = ~n5447 & ~n5458 ;
  assign n5460 = n965 & ~n5459 ;
  assign n5450 = n1867 & ~n5449 ;
  assign n5461 = \InstQueue_reg[4][6]/NET0131  & ~n3929 ;
  assign n5462 = ~n5450 & ~n5461 ;
  assign n5463 = ~n5460 & n5462 ;
  assign n5464 = ~n5457 & n5463 ;
  assign n5470 = n4093 & n5045 ;
  assign n5471 = n4115 & n5048 ;
  assign n5472 = ~n5470 & ~n5471 ;
  assign n5473 = \DataWidth_reg[1]/NET0131  & ~n5472 ;
  assign n5465 = \Datai[3]_pad  & ~n4160 ;
  assign n5466 = \InstQueue_reg[5][3]/NET0131  & ~n4159 ;
  assign n5467 = ~n4137 & n5466 ;
  assign n5468 = ~n5465 & ~n5467 ;
  assign n5474 = ~n4170 & ~n5468 ;
  assign n5475 = ~n5473 & ~n5474 ;
  assign n5476 = n933 & ~n5475 ;
  assign n5477 = ~n540 & n4159 ;
  assign n5478 = ~n5466 & ~n5477 ;
  assign n5479 = n965 & ~n5478 ;
  assign n5469 = n1867 & ~n5468 ;
  assign n5480 = \InstQueue_reg[5][3]/NET0131  & ~n3929 ;
  assign n5481 = ~n5469 & ~n5480 ;
  assign n5482 = ~n5479 & n5481 ;
  assign n5483 = ~n5476 & n5482 ;
  assign n5489 = n4093 & n5068 ;
  assign n5490 = n4115 & n5071 ;
  assign n5491 = ~n5489 & ~n5490 ;
  assign n5492 = \DataWidth_reg[1]/NET0131  & ~n5491 ;
  assign n5484 = \Datai[6]_pad  & ~n4160 ;
  assign n5485 = \InstQueue_reg[5][6]/NET0131  & ~n4159 ;
  assign n5486 = ~n4137 & n5485 ;
  assign n5487 = ~n5484 & ~n5486 ;
  assign n5493 = ~n4170 & ~n5487 ;
  assign n5494 = ~n5492 & ~n5493 ;
  assign n5495 = n933 & ~n5494 ;
  assign n5496 = ~n731 & n4159 ;
  assign n5497 = ~n5485 & ~n5496 ;
  assign n5498 = n965 & ~n5497 ;
  assign n5488 = n1867 & ~n5487 ;
  assign n5499 = \InstQueue_reg[5][6]/NET0131  & ~n3929 ;
  assign n5500 = ~n5488 & ~n5499 ;
  assign n5501 = ~n5498 & n5500 ;
  assign n5502 = ~n5495 & n5501 ;
  assign n5508 = n4115 & n5045 ;
  assign n5509 = n4137 & n5048 ;
  assign n5510 = ~n5508 & ~n5509 ;
  assign n5511 = \DataWidth_reg[1]/NET0131  & ~n5510 ;
  assign n5503 = \Datai[3]_pad  & ~n4182 ;
  assign n5504 = \InstQueue_reg[6][3]/NET0131  & ~n4181 ;
  assign n5505 = ~n4159 & n5504 ;
  assign n5506 = ~n5503 & ~n5505 ;
  assign n5512 = ~n4192 & ~n5506 ;
  assign n5513 = ~n5511 & ~n5512 ;
  assign n5514 = n933 & ~n5513 ;
  assign n5515 = ~n540 & n4181 ;
  assign n5516 = ~n5504 & ~n5515 ;
  assign n5517 = n965 & ~n5516 ;
  assign n5507 = n1867 & ~n5506 ;
  assign n5518 = \InstQueue_reg[6][3]/NET0131  & ~n3929 ;
  assign n5519 = ~n5507 & ~n5518 ;
  assign n5520 = ~n5517 & n5519 ;
  assign n5521 = ~n5514 & n5520 ;
  assign n5527 = n4115 & n5068 ;
  assign n5528 = n4137 & n5071 ;
  assign n5529 = ~n5527 & ~n5528 ;
  assign n5530 = \DataWidth_reg[1]/NET0131  & ~n5529 ;
  assign n5522 = \Datai[6]_pad  & ~n4182 ;
  assign n5523 = \InstQueue_reg[6][6]/NET0131  & ~n4181 ;
  assign n5524 = ~n4159 & n5523 ;
  assign n5525 = ~n5522 & ~n5524 ;
  assign n5531 = ~n4192 & ~n5525 ;
  assign n5532 = ~n5530 & ~n5531 ;
  assign n5533 = n933 & ~n5532 ;
  assign n5534 = ~n731 & n4181 ;
  assign n5535 = ~n5523 & ~n5534 ;
  assign n5536 = n965 & ~n5535 ;
  assign n5526 = n1867 & ~n5525 ;
  assign n5537 = \InstQueue_reg[6][6]/NET0131  & ~n3929 ;
  assign n5538 = ~n5526 & ~n5537 ;
  assign n5539 = ~n5536 & n5538 ;
  assign n5540 = ~n5533 & n5539 ;
  assign n5546 = n4137 & n5045 ;
  assign n5547 = n4159 & n5048 ;
  assign n5548 = ~n5546 & ~n5547 ;
  assign n5549 = \DataWidth_reg[1]/NET0131  & ~n5548 ;
  assign n5541 = \Datai[3]_pad  & ~n4203 ;
  assign n5542 = \InstQueue_reg[7][3]/NET0131  & ~n3944 ;
  assign n5543 = ~n4181 & n5542 ;
  assign n5544 = ~n5541 & ~n5543 ;
  assign n5550 = ~n4213 & ~n5544 ;
  assign n5551 = ~n5549 & ~n5550 ;
  assign n5552 = n933 & ~n5551 ;
  assign n5553 = ~n540 & n3944 ;
  assign n5554 = ~n5542 & ~n5553 ;
  assign n5555 = n965 & ~n5554 ;
  assign n5545 = n1867 & ~n5544 ;
  assign n5556 = \InstQueue_reg[7][3]/NET0131  & ~n3929 ;
  assign n5557 = ~n5545 & ~n5556 ;
  assign n5558 = ~n5555 & n5557 ;
  assign n5559 = ~n5552 & n5558 ;
  assign n5565 = n4137 & n5068 ;
  assign n5566 = n4159 & n5071 ;
  assign n5567 = ~n5565 & ~n5566 ;
  assign n5568 = \DataWidth_reg[1]/NET0131  & ~n5567 ;
  assign n5560 = \Datai[6]_pad  & ~n4203 ;
  assign n5561 = \InstQueue_reg[7][6]/NET0131  & ~n3944 ;
  assign n5562 = ~n4181 & n5561 ;
  assign n5563 = ~n5560 & ~n5562 ;
  assign n5569 = ~n4213 & ~n5563 ;
  assign n5570 = ~n5568 & ~n5569 ;
  assign n5571 = n933 & ~n5570 ;
  assign n5572 = ~n731 & n3944 ;
  assign n5573 = ~n5561 & ~n5572 ;
  assign n5574 = n965 & ~n5573 ;
  assign n5564 = n1867 & ~n5563 ;
  assign n5575 = \InstQueue_reg[7][6]/NET0131  & ~n3929 ;
  assign n5576 = ~n5564 & ~n5575 ;
  assign n5577 = ~n5574 & n5576 ;
  assign n5578 = ~n5571 & n5577 ;
  assign n5584 = n4159 & n5045 ;
  assign n5585 = n4181 & n5048 ;
  assign n5586 = ~n5584 & ~n5585 ;
  assign n5587 = \DataWidth_reg[1]/NET0131  & ~n5586 ;
  assign n5579 = \Datai[3]_pad  & ~n3950 ;
  assign n5580 = \InstQueue_reg[8][3]/NET0131  & ~n3946 ;
  assign n5581 = ~n3944 & n5580 ;
  assign n5582 = ~n5579 & ~n5581 ;
  assign n5588 = ~n4233 & ~n5582 ;
  assign n5589 = ~n5587 & ~n5588 ;
  assign n5590 = n933 & ~n5589 ;
  assign n5591 = ~n540 & n3946 ;
  assign n5592 = ~n5580 & ~n5591 ;
  assign n5593 = n965 & ~n5592 ;
  assign n5583 = n1867 & ~n5582 ;
  assign n5594 = \InstQueue_reg[8][3]/NET0131  & ~n3929 ;
  assign n5595 = ~n5583 & ~n5594 ;
  assign n5596 = ~n5593 & n5595 ;
  assign n5597 = ~n5590 & n5596 ;
  assign n5603 = n4159 & n5068 ;
  assign n5604 = n4181 & n5071 ;
  assign n5605 = ~n5603 & ~n5604 ;
  assign n5606 = \DataWidth_reg[1]/NET0131  & ~n5605 ;
  assign n5598 = \Datai[6]_pad  & ~n3950 ;
  assign n5599 = \InstQueue_reg[8][6]/NET0131  & ~n3946 ;
  assign n5600 = ~n3944 & n5599 ;
  assign n5601 = ~n5598 & ~n5600 ;
  assign n5607 = ~n4233 & ~n5601 ;
  assign n5608 = ~n5606 & ~n5607 ;
  assign n5609 = n933 & ~n5608 ;
  assign n5610 = ~n731 & n3946 ;
  assign n5611 = ~n5599 & ~n5610 ;
  assign n5612 = n965 & ~n5611 ;
  assign n5602 = n1867 & ~n5601 ;
  assign n5613 = \InstQueue_reg[8][6]/NET0131  & ~n3929 ;
  assign n5614 = ~n5602 & ~n5613 ;
  assign n5615 = ~n5612 & n5614 ;
  assign n5616 = ~n5609 & n5615 ;
  assign n5622 = n4181 & n5045 ;
  assign n5623 = n3944 & n5048 ;
  assign n5624 = ~n5622 & ~n5623 ;
  assign n5625 = \DataWidth_reg[1]/NET0131  & ~n5624 ;
  assign n5617 = \Datai[3]_pad  & ~n3974 ;
  assign n5618 = \InstQueue_reg[9][3]/NET0131  & ~n3937 ;
  assign n5619 = ~n3946 & n5618 ;
  assign n5620 = ~n5617 & ~n5619 ;
  assign n5626 = ~n4253 & ~n5620 ;
  assign n5627 = ~n5625 & ~n5626 ;
  assign n5628 = n933 & ~n5627 ;
  assign n5629 = ~n540 & n3937 ;
  assign n5630 = ~n5618 & ~n5629 ;
  assign n5631 = n965 & ~n5630 ;
  assign n5621 = n1867 & ~n5620 ;
  assign n5632 = \InstQueue_reg[9][3]/NET0131  & ~n3929 ;
  assign n5633 = ~n5621 & ~n5632 ;
  assign n5634 = ~n5631 & n5633 ;
  assign n5635 = ~n5628 & n5634 ;
  assign n5641 = n4181 & n5068 ;
  assign n5642 = n3944 & n5071 ;
  assign n5643 = ~n5641 & ~n5642 ;
  assign n5644 = \DataWidth_reg[1]/NET0131  & ~n5643 ;
  assign n5636 = \Datai[6]_pad  & ~n3974 ;
  assign n5637 = \InstQueue_reg[9][6]/NET0131  & ~n3937 ;
  assign n5638 = ~n3946 & n5637 ;
  assign n5639 = ~n5636 & ~n5638 ;
  assign n5645 = ~n4253 & ~n5639 ;
  assign n5646 = ~n5644 & ~n5645 ;
  assign n5647 = n933 & ~n5646 ;
  assign n5648 = ~n731 & n3937 ;
  assign n5649 = ~n5637 & ~n5648 ;
  assign n5650 = n965 & ~n5649 ;
  assign n5640 = n1867 & ~n5639 ;
  assign n5651 = \InstQueue_reg[9][6]/NET0131  & ~n3929 ;
  assign n5652 = ~n5640 & ~n5651 ;
  assign n5653 = ~n5650 & n5652 ;
  assign n5654 = ~n5647 & n5653 ;
  assign n5659 = n929 & ~n2739 ;
  assign n5658 = n941 & n966 ;
  assign n5660 = ~n933 & ~n953 ;
  assign n5661 = n5658 & n5660 ;
  assign n5662 = ~n5659 & n5661 ;
  assign n5663 = \PhyAddrPointer_reg[0]/NET0131  & ~n5662 ;
  assign n5655 = n773 & n3575 ;
  assign n5656 = ~n3582 & ~n5655 ;
  assign n5657 = n929 & ~n5656 ;
  assign n5664 = ~n3571 & ~n5657 ;
  assign n5665 = ~n5663 & n5664 ;
  assign n5693 = \PhyAddrPointer_reg[0]/NET0131  & ~n1899 ;
  assign n5695 = \PhyAddrPointer_reg[1]/NET0131  & n5693 ;
  assign n5694 = ~\PhyAddrPointer_reg[1]/NET0131  & ~n5693 ;
  assign n5696 = ~\DataWidth_reg[1]/NET0131  & ~n5694 ;
  assign n5697 = ~n5695 & n5696 ;
  assign n5692 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[1]/NET0131  ;
  assign n5698 = n933 & ~n5692 ;
  assign n5699 = ~n5697 & n5698 ;
  assign n5684 = ~n785 & ~n834 ;
  assign n5685 = \rEIP_reg[1]/NET0131  & ~n5684 ;
  assign n5671 = ~\EBX_reg[1]/NET0131  & ~n924 ;
  assign n5672 = n923 & ~n5671 ;
  assign n5673 = ~\EBX_reg[0]/NET0131  & ~\EBX_reg[1]/NET0131  ;
  assign n5674 = ~n3468 & ~n5673 ;
  assign n5675 = \EBX_reg[31]/NET0131  & n5674 ;
  assign n5676 = ~\DataWidth_reg[1]/NET0131  & ~READY_n_pad ;
  assign n5677 = \EBX_reg[1]/NET0131  & ~\EBX_reg[31]/NET0131  ;
  assign n5678 = ~n5676 & ~n5677 ;
  assign n5679 = ~n5675 & n5678 ;
  assign n5680 = n3660 & ~n5679 ;
  assign n5681 = ~n5672 & ~n5680 ;
  assign n5682 = \rEIP_reg[1]/NET0131  & n5676 ;
  assign n5683 = ~n5681 & ~n5682 ;
  assign n5669 = n778 & ~n834 ;
  assign n5670 = ~n822 & n5669 ;
  assign n5686 = n828 & n5672 ;
  assign n5687 = ~n5670 & ~n5686 ;
  assign n5688 = ~n5683 & n5687 ;
  assign n5689 = ~n5685 & n5688 ;
  assign n5690 = n929 & ~n5689 ;
  assign n5666 = ~n939 & ~n1867 ;
  assign n5667 = n4267 & n5666 ;
  assign n5668 = \rEIP_reg[1]/NET0131  & ~n5667 ;
  assign n5691 = \PhyAddrPointer_reg[1]/NET0131  & n953 ;
  assign n5700 = ~n5668 & ~n5691 ;
  assign n5701 = ~n5690 & n5700 ;
  assign n5702 = ~n5699 & n5701 ;
  assign n5704 = ~\PhyAddrPointer_reg[20]/NET0131  & ~n2509 ;
  assign n5705 = ~n2810 & ~n5704 ;
  assign n5706 = ~\PhyAddrPointer_reg[0]/NET0131  & n2232 ;
  assign n5707 = n1880 & n5706 ;
  assign n5708 = ~n2486 & n5707 ;
  assign n5709 = ~n2240 & n5708 ;
  assign n5710 = ~n2715 & n5709 ;
  assign n5711 = ~n2752 & n5710 ;
  assign n5712 = ~n2510 & ~n2781 ;
  assign n5713 = n5711 & n5712 ;
  assign n5714 = n3531 & n5713 ;
  assign n5715 = ~n1899 & ~n5714 ;
  assign n5717 = ~n5705 & n5715 ;
  assign n5716 = n5705 & ~n5715 ;
  assign n5718 = ~\DataWidth_reg[1]/NET0131  & ~n5716 ;
  assign n5719 = ~n5717 & n5718 ;
  assign n5703 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[20]/NET0131  ;
  assign n5720 = n933 & ~n5703 ;
  assign n5721 = ~n5719 & n5720 ;
  assign n5747 = ~\EBX_reg[2]/NET0131  & n5673 ;
  assign n5748 = ~\EBX_reg[3]/NET0131  & n5747 ;
  assign n5749 = ~\EBX_reg[4]/NET0131  & n5748 ;
  assign n5750 = ~\EBX_reg[5]/NET0131  & n5749 ;
  assign n5751 = ~\EBX_reg[6]/NET0131  & n5750 ;
  assign n5752 = ~\EBX_reg[7]/NET0131  & n5751 ;
  assign n5753 = ~\EBX_reg[8]/NET0131  & n5752 ;
  assign n5754 = ~\EBX_reg[10]/NET0131  & ~\EBX_reg[9]/NET0131  ;
  assign n5755 = n5753 & n5754 ;
  assign n5756 = ~\EBX_reg[11]/NET0131  & ~\EBX_reg[12]/NET0131  ;
  assign n5757 = n5755 & n5756 ;
  assign n5758 = ~\EBX_reg[13]/NET0131  & n5757 ;
  assign n5759 = ~\EBX_reg[14]/NET0131  & n5758 ;
  assign n5760 = ~\EBX_reg[15]/NET0131  & ~\EBX_reg[16]/NET0131  ;
  assign n5761 = n5759 & n5760 ;
  assign n5762 = ~\EBX_reg[17]/NET0131  & n5761 ;
  assign n5763 = ~\EBX_reg[18]/NET0131  & n5762 ;
  assign n5764 = ~\EBX_reg[19]/NET0131  & n5763 ;
  assign n5765 = \EBX_reg[31]/NET0131  & ~n5764 ;
  assign n5767 = ~\EBX_reg[20]/NET0131  & n5765 ;
  assign n5766 = \EBX_reg[20]/NET0131  & ~n5765 ;
  assign n5768 = ~n5676 & ~n5766 ;
  assign n5769 = ~n5767 & n5768 ;
  assign n5724 = \rEIP_reg[1]/NET0131  & \rEIP_reg[2]/NET0131  ;
  assign n5725 = \rEIP_reg[3]/NET0131  & n5724 ;
  assign n5726 = \rEIP_reg[4]/NET0131  & n5725 ;
  assign n5727 = \rEIP_reg[5]/NET0131  & n5726 ;
  assign n5728 = \rEIP_reg[6]/NET0131  & n5727 ;
  assign n5729 = \rEIP_reg[7]/NET0131  & n5728 ;
  assign n5730 = \rEIP_reg[8]/NET0131  & n5729 ;
  assign n5731 = \rEIP_reg[9]/NET0131  & n5730 ;
  assign n5732 = \rEIP_reg[10]/NET0131  & n5731 ;
  assign n5733 = \rEIP_reg[11]/NET0131  & n5732 ;
  assign n5734 = \rEIP_reg[12]/NET0131  & \rEIP_reg[13]/NET0131  ;
  assign n5735 = \rEIP_reg[14]/NET0131  & n5734 ;
  assign n5736 = \rEIP_reg[15]/NET0131  & n5735 ;
  assign n5737 = n5733 & n5736 ;
  assign n5738 = \rEIP_reg[16]/NET0131  & n5737 ;
  assign n5739 = \rEIP_reg[17]/NET0131  & \rEIP_reg[18]/NET0131  ;
  assign n5740 = n5738 & n5739 ;
  assign n5741 = \rEIP_reg[19]/NET0131  & n5740 ;
  assign n5742 = ~\rEIP_reg[20]/NET0131  & ~n5741 ;
  assign n5743 = \rEIP_reg[19]/NET0131  & \rEIP_reg[20]/NET0131  ;
  assign n5744 = n5740 & n5743 ;
  assign n5745 = ~n5742 & ~n5744 ;
  assign n5746 = n5676 & ~n5745 ;
  assign n5770 = n3660 & ~n5746 ;
  assign n5771 = ~n5769 & n5770 ;
  assign n5772 = \rEIP_reg[20]/NET0131  & ~n5684 ;
  assign n5774 = ~n828 & n5746 ;
  assign n5773 = ~\EBX_reg[20]/NET0131  & ~n924 ;
  assign n5775 = n923 & ~n5773 ;
  assign n5776 = ~n5774 & n5775 ;
  assign n5777 = ~n5772 & ~n5776 ;
  assign n5778 = ~n5771 & n5777 ;
  assign n5779 = n929 & ~n5778 ;
  assign n5722 = \PhyAddrPointer_reg[20]/NET0131  & n953 ;
  assign n5723 = \rEIP_reg[20]/NET0131  & ~n5667 ;
  assign n5780 = ~n5722 & ~n5723 ;
  assign n5781 = ~n5779 & n5780 ;
  assign n5782 = ~n5721 & n5781 ;
  assign n5784 = ~n5705 & n5713 ;
  assign n5785 = ~n1899 & ~n5784 ;
  assign n5787 = ~n2812 & n5785 ;
  assign n5786 = n2812 & ~n5785 ;
  assign n5788 = ~\DataWidth_reg[1]/NET0131  & ~n5786 ;
  assign n5789 = ~n5787 & n5788 ;
  assign n5783 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[21]/NET0131  ;
  assign n5790 = n933 & ~n5783 ;
  assign n5791 = ~n5789 & n5790 ;
  assign n5799 = ~\EBX_reg[20]/NET0131  & n5764 ;
  assign n5800 = \EBX_reg[31]/NET0131  & ~n5799 ;
  assign n5802 = ~\EBX_reg[21]/NET0131  & n5800 ;
  assign n5801 = \EBX_reg[21]/NET0131  & ~n5800 ;
  assign n5803 = ~n5676 & ~n5801 ;
  assign n5804 = ~n5802 & n5803 ;
  assign n5794 = ~\rEIP_reg[21]/NET0131  & ~n5744 ;
  assign n5795 = \rEIP_reg[21]/NET0131  & n5743 ;
  assign n5796 = n5740 & n5795 ;
  assign n5797 = ~n5794 & ~n5796 ;
  assign n5798 = n5676 & ~n5797 ;
  assign n5805 = n3660 & ~n5798 ;
  assign n5806 = ~n5804 & n5805 ;
  assign n5807 = \rEIP_reg[21]/NET0131  & ~n5684 ;
  assign n5809 = ~n828 & n5798 ;
  assign n5808 = ~\EBX_reg[21]/NET0131  & ~n924 ;
  assign n5810 = n923 & ~n5808 ;
  assign n5811 = ~n5809 & n5810 ;
  assign n5812 = ~n5807 & ~n5811 ;
  assign n5813 = ~n5806 & n5812 ;
  assign n5814 = n929 & ~n5813 ;
  assign n5792 = \rEIP_reg[21]/NET0131  & ~n5667 ;
  assign n5793 = \PhyAddrPointer_reg[21]/NET0131  & n953 ;
  assign n5815 = ~n5792 & ~n5793 ;
  assign n5816 = ~n5814 & n5815 ;
  assign n5817 = ~n5791 & n5816 ;
  assign n5841 = ~n2812 & ~n5705 ;
  assign n5842 = n5714 & n5841 ;
  assign n5843 = ~n1899 & ~n5842 ;
  assign n5845 = ~n2545 & n5843 ;
  assign n5844 = n2545 & ~n5843 ;
  assign n5846 = ~\DataWidth_reg[1]/NET0131  & ~n5844 ;
  assign n5847 = ~n5845 & n5846 ;
  assign n5840 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[22]/NET0131  ;
  assign n5848 = n933 & ~n5840 ;
  assign n5849 = ~n5847 & n5848 ;
  assign n5818 = \rEIP_reg[22]/NET0131  & ~n5684 ;
  assign n5819 = ~\EBX_reg[22]/NET0131  & ~n924 ;
  assign n5820 = n923 & ~n5819 ;
  assign n5821 = ~\EBX_reg[21]/NET0131  & n5799 ;
  assign n5822 = \EBX_reg[31]/NET0131  & ~n5821 ;
  assign n5824 = ~\EBX_reg[22]/NET0131  & n5822 ;
  assign n5823 = \EBX_reg[22]/NET0131  & ~n5822 ;
  assign n5825 = ~n5676 & ~n5823 ;
  assign n5826 = ~n5824 & n5825 ;
  assign n5827 = n3660 & ~n5826 ;
  assign n5828 = ~n5820 & ~n5827 ;
  assign n5829 = ~\rEIP_reg[22]/NET0131  & ~n5796 ;
  assign n5830 = \rEIP_reg[22]/NET0131  & n5739 ;
  assign n5831 = n5795 & n5830 ;
  assign n5832 = n5738 & n5831 ;
  assign n5833 = ~n5829 & ~n5832 ;
  assign n5834 = n828 & n5820 ;
  assign n5835 = n5676 & ~n5834 ;
  assign n5836 = ~n5833 & n5835 ;
  assign n5837 = ~n5828 & ~n5836 ;
  assign n5838 = ~n5818 & ~n5837 ;
  assign n5839 = n929 & ~n5838 ;
  assign n5850 = \rEIP_reg[22]/NET0131  & ~n5667 ;
  assign n5851 = \PhyAddrPointer_reg[22]/NET0131  & n953 ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = ~n5839 & n5852 ;
  assign n5854 = ~n5849 & n5853 ;
  assign n5878 = ~n2545 & n5841 ;
  assign n5879 = n5714 & n5878 ;
  assign n5880 = ~n1899 & ~n5879 ;
  assign n5882 = n2270 & ~n5880 ;
  assign n5881 = ~n2270 & n5880 ;
  assign n5883 = ~\DataWidth_reg[1]/NET0131  & ~n5881 ;
  assign n5884 = ~n5882 & n5883 ;
  assign n5877 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[23]/NET0131  ;
  assign n5885 = n933 & ~n5877 ;
  assign n5886 = ~n5884 & n5885 ;
  assign n5864 = ~\EBX_reg[22]/NET0131  & n5821 ;
  assign n5865 = \EBX_reg[31]/NET0131  & ~n5864 ;
  assign n5867 = ~\EBX_reg[23]/NET0131  & n5865 ;
  assign n5866 = \EBX_reg[23]/NET0131  & ~n5865 ;
  assign n5868 = ~n5676 & ~n5866 ;
  assign n5869 = ~n5867 & n5868 ;
  assign n5857 = ~\rEIP_reg[23]/NET0131  & ~n5832 ;
  assign n5858 = \rEIP_reg[23]/NET0131  & n5832 ;
  assign n5859 = ~n5857 & ~n5858 ;
  assign n5863 = n5676 & ~n5859 ;
  assign n5870 = n3660 & ~n5863 ;
  assign n5871 = ~n5869 & n5870 ;
  assign n5855 = \rEIP_reg[23]/NET0131  & ~n5684 ;
  assign n5860 = n924 & ~n5859 ;
  assign n5856 = ~\EBX_reg[23]/NET0131  & ~n924 ;
  assign n5861 = n923 & ~n5856 ;
  assign n5862 = ~n5860 & n5861 ;
  assign n5872 = ~n5855 & ~n5862 ;
  assign n5873 = ~n5871 & n5872 ;
  assign n5874 = n929 & ~n5873 ;
  assign n5875 = \PhyAddrPointer_reg[23]/NET0131  & n953 ;
  assign n5876 = \rEIP_reg[23]/NET0131  & ~n5667 ;
  assign n5887 = ~n5875 & ~n5876 ;
  assign n5888 = ~n5874 & n5887 ;
  assign n5889 = ~n5886 & n5888 ;
  assign n5894 = ~\EBX_reg[23]/NET0131  & n5864 ;
  assign n5895 = \EBX_reg[31]/NET0131  & ~n5894 ;
  assign n5897 = ~\EBX_reg[24]/NET0131  & ~n5895 ;
  assign n5896 = \EBX_reg[24]/NET0131  & n5895 ;
  assign n5898 = ~n5676 & ~n5896 ;
  assign n5899 = ~n5897 & n5898 ;
  assign n5890 = ~\rEIP_reg[24]/NET0131  & ~n5858 ;
  assign n5891 = \rEIP_reg[24]/NET0131  & n5858 ;
  assign n5892 = ~n5890 & ~n5891 ;
  assign n5893 = n5676 & n5892 ;
  assign n5900 = ~n834 & ~n5893 ;
  assign n5901 = ~n5899 & n5900 ;
  assign n5902 = ~\rEIP_reg[24]/NET0131  & n834 ;
  assign n5903 = n782 & ~n5902 ;
  assign n5904 = ~n5901 & n5903 ;
  assign n5906 = n924 & ~n5892 ;
  assign n5905 = ~\EBX_reg[24]/NET0131  & ~n924 ;
  assign n5907 = n923 & ~n5905 ;
  assign n5908 = ~n5906 & n5907 ;
  assign n5909 = ~n778 & n782 ;
  assign n5910 = \rEIP_reg[24]/NET0131  & ~n5909 ;
  assign n5911 = ~n5684 & n5910 ;
  assign n5912 = ~n5908 & ~n5911 ;
  assign n5913 = ~n5904 & n5912 ;
  assign n5914 = n929 & ~n5913 ;
  assign n5916 = ~n2270 & n5879 ;
  assign n5917 = ~n1899 & ~n5916 ;
  assign n5919 = ~n2570 & n5917 ;
  assign n5918 = n2570 & ~n5917 ;
  assign n5920 = ~\DataWidth_reg[1]/NET0131  & ~n5918 ;
  assign n5921 = ~n5919 & n5920 ;
  assign n5915 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[24]/NET0131  ;
  assign n5922 = n933 & ~n5915 ;
  assign n5923 = ~n5921 & n5922 ;
  assign n5924 = \rEIP_reg[24]/NET0131  & ~n5667 ;
  assign n5925 = \PhyAddrPointer_reg[24]/NET0131  & n953 ;
  assign n5926 = ~n5924 & ~n5925 ;
  assign n5927 = ~n5923 & n5926 ;
  assign n5928 = ~n5914 & n5927 ;
  assign n5952 = ~n2270 & ~n2570 ;
  assign n5953 = n5713 & n5952 ;
  assign n5954 = n5878 & n5953 ;
  assign n5955 = ~n1899 & ~n5954 ;
  assign n5957 = ~n2833 & n5955 ;
  assign n5956 = n2833 & ~n5955 ;
  assign n5958 = ~\DataWidth_reg[1]/NET0131  & ~n5956 ;
  assign n5959 = ~n5957 & n5958 ;
  assign n5951 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[25]/NET0131  ;
  assign n5960 = n933 & ~n5951 ;
  assign n5961 = ~n5959 & n5960 ;
  assign n5939 = ~\EBX_reg[23]/NET0131  & ~\EBX_reg[24]/NET0131  ;
  assign n5940 = n5864 & n5939 ;
  assign n5941 = \EBX_reg[31]/NET0131  & ~n5940 ;
  assign n5943 = \EBX_reg[25]/NET0131  & ~n5941 ;
  assign n5942 = ~\EBX_reg[25]/NET0131  & n5941 ;
  assign n5944 = ~n5676 & ~n5942 ;
  assign n5945 = ~n5943 & n5944 ;
  assign n5931 = ~\rEIP_reg[25]/NET0131  & ~n5891 ;
  assign n5932 = \rEIP_reg[24]/NET0131  & \rEIP_reg[25]/NET0131  ;
  assign n5933 = n5858 & n5932 ;
  assign n5934 = ~n5931 & ~n5933 ;
  assign n5938 = n5676 & ~n5934 ;
  assign n5946 = n3660 & ~n5938 ;
  assign n5947 = ~n5945 & n5946 ;
  assign n5929 = \rEIP_reg[25]/NET0131  & ~n5684 ;
  assign n5935 = n924 & ~n5934 ;
  assign n5930 = ~\EBX_reg[25]/NET0131  & ~n924 ;
  assign n5936 = n923 & ~n5930 ;
  assign n5937 = ~n5935 & n5936 ;
  assign n5948 = ~n5929 & ~n5937 ;
  assign n5949 = ~n5947 & n5948 ;
  assign n5950 = n929 & ~n5949 ;
  assign n5962 = \rEIP_reg[25]/NET0131  & ~n5667 ;
  assign n5963 = \PhyAddrPointer_reg[25]/NET0131  & n953 ;
  assign n5964 = ~n5962 & ~n5963 ;
  assign n5965 = ~n5950 & n5964 ;
  assign n5966 = ~n5961 & n5965 ;
  assign n5993 = ~n2833 & n5952 ;
  assign n5994 = n5879 & n5993 ;
  assign n5995 = ~n1899 & ~n5994 ;
  assign n5997 = ~n2589 & n5995 ;
  assign n5996 = n2589 & ~n5995 ;
  assign n5998 = ~\DataWidth_reg[1]/NET0131  & ~n5996 ;
  assign n5999 = ~n5997 & n5998 ;
  assign n5992 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[26]/NET0131  ;
  assign n6000 = n933 & ~n5992 ;
  assign n6001 = ~n5999 & n6000 ;
  assign n5977 = ~\EBX_reg[22]/NET0131  & ~\EBX_reg[25]/NET0131  ;
  assign n5978 = n5939 & n5977 ;
  assign n5979 = n5821 & n5978 ;
  assign n5980 = \EBX_reg[31]/NET0131  & ~n5979 ;
  assign n5982 = \EBX_reg[26]/NET0131  & ~n5980 ;
  assign n5981 = ~\EBX_reg[26]/NET0131  & n5980 ;
  assign n5983 = ~n5676 & ~n5981 ;
  assign n5984 = ~n5982 & n5983 ;
  assign n5969 = ~\rEIP_reg[26]/NET0131  & ~n5933 ;
  assign n5970 = \rEIP_reg[26]/NET0131  & n5932 ;
  assign n5971 = n5858 & n5970 ;
  assign n5972 = ~n5969 & ~n5971 ;
  assign n5976 = n5676 & ~n5972 ;
  assign n5985 = n3660 & ~n5976 ;
  assign n5986 = ~n5984 & n5985 ;
  assign n5967 = \rEIP_reg[26]/NET0131  & ~n5684 ;
  assign n5973 = n924 & ~n5972 ;
  assign n5968 = ~\EBX_reg[26]/NET0131  & ~n924 ;
  assign n5974 = n923 & ~n5968 ;
  assign n5975 = ~n5973 & n5974 ;
  assign n5987 = ~n5967 & ~n5975 ;
  assign n5988 = ~n5986 & n5987 ;
  assign n5989 = n929 & ~n5988 ;
  assign n5990 = \rEIP_reg[26]/NET0131  & ~n5667 ;
  assign n5991 = \PhyAddrPointer_reg[26]/NET0131  & n953 ;
  assign n6002 = ~n5990 & ~n5991 ;
  assign n6003 = ~n5989 & n6002 ;
  assign n6004 = ~n6001 & n6003 ;
  assign n6026 = ~n2589 & n5994 ;
  assign n6027 = ~n1899 & ~n6026 ;
  assign n6029 = ~n2306 & n6027 ;
  assign n6028 = n2306 & ~n6027 ;
  assign n6030 = ~\DataWidth_reg[1]/NET0131  & ~n6028 ;
  assign n6031 = ~n6029 & n6030 ;
  assign n6025 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[27]/NET0131  ;
  assign n6032 = n933 & ~n6025 ;
  assign n6033 = ~n6031 & n6032 ;
  assign n6014 = ~\EBX_reg[26]/NET0131  & n5979 ;
  assign n6015 = \EBX_reg[31]/NET0131  & ~n6014 ;
  assign n6017 = ~\EBX_reg[27]/NET0131  & n6015 ;
  assign n6016 = \EBX_reg[27]/NET0131  & ~n6015 ;
  assign n6018 = ~n5676 & ~n6016 ;
  assign n6019 = ~n6017 & n6018 ;
  assign n6007 = ~\rEIP_reg[27]/NET0131  & ~n5971 ;
  assign n6008 = \rEIP_reg[27]/NET0131  & n5971 ;
  assign n6009 = ~n6007 & ~n6008 ;
  assign n6010 = n5676 & ~n6009 ;
  assign n6020 = n3660 & ~n6010 ;
  assign n6021 = ~n6019 & n6020 ;
  assign n6005 = \rEIP_reg[27]/NET0131  & ~n5684 ;
  assign n6011 = ~n828 & n6010 ;
  assign n6006 = ~\EBX_reg[27]/NET0131  & ~n924 ;
  assign n6012 = n923 & ~n6006 ;
  assign n6013 = ~n6011 & n6012 ;
  assign n6022 = ~n6005 & ~n6013 ;
  assign n6023 = ~n6021 & n6022 ;
  assign n6024 = n929 & ~n6023 ;
  assign n6034 = \PhyAddrPointer_reg[27]/NET0131  & n953 ;
  assign n6035 = \rEIP_reg[27]/NET0131  & ~n5667 ;
  assign n6036 = ~n6034 & ~n6035 ;
  assign n6037 = ~n6024 & n6036 ;
  assign n6038 = ~n6033 & n6037 ;
  assign n6043 = ~\EBX_reg[27]/NET0131  & n6014 ;
  assign n6044 = \EBX_reg[31]/NET0131  & ~n6043 ;
  assign n6046 = ~\EBX_reg[28]/NET0131  & n6044 ;
  assign n6045 = \EBX_reg[28]/NET0131  & ~n6044 ;
  assign n6047 = ~n5676 & ~n6045 ;
  assign n6048 = ~n6046 & n6047 ;
  assign n6039 = \rEIP_reg[28]/NET0131  & n6008 ;
  assign n6040 = ~\rEIP_reg[28]/NET0131  & ~n6008 ;
  assign n6041 = ~n6039 & ~n6040 ;
  assign n6042 = n5676 & ~n6041 ;
  assign n6049 = n3660 & ~n6042 ;
  assign n6050 = ~n6048 & n6049 ;
  assign n6051 = \rEIP_reg[28]/NET0131  & ~n5684 ;
  assign n6053 = n924 & ~n6041 ;
  assign n6052 = ~\EBX_reg[28]/NET0131  & ~n924 ;
  assign n6054 = n923 & ~n6052 ;
  assign n6055 = ~n6053 & n6054 ;
  assign n6056 = ~n6051 & ~n6055 ;
  assign n6057 = ~n6050 & n6056 ;
  assign n6058 = n929 & ~n6057 ;
  assign n6060 = ~n2306 & n6026 ;
  assign n6061 = ~n1899 & ~n6060 ;
  assign n6063 = ~n2359 & n6061 ;
  assign n6062 = n2359 & ~n6061 ;
  assign n6064 = ~\DataWidth_reg[1]/NET0131  & ~n6062 ;
  assign n6065 = ~n6063 & n6064 ;
  assign n6059 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[28]/NET0131  ;
  assign n6066 = n933 & ~n6059 ;
  assign n6067 = ~n6065 & n6066 ;
  assign n6068 = \rEIP_reg[28]/NET0131  & ~n5667 ;
  assign n6069 = \PhyAddrPointer_reg[28]/NET0131  & n953 ;
  assign n6070 = ~n6068 & ~n6069 ;
  assign n6071 = ~n6067 & n6070 ;
  assign n6072 = ~n6058 & n6071 ;
  assign n6077 = ~\EBX_reg[27]/NET0131  & ~\EBX_reg[28]/NET0131  ;
  assign n6078 = n6014 & n6077 ;
  assign n6079 = \EBX_reg[31]/NET0131  & ~n6078 ;
  assign n6081 = \EBX_reg[29]/NET0131  & ~n6079 ;
  assign n6080 = ~\EBX_reg[29]/NET0131  & n6079 ;
  assign n6082 = ~n5676 & ~n6080 ;
  assign n6083 = ~n6081 & n6082 ;
  assign n6073 = ~\rEIP_reg[29]/NET0131  & ~n6039 ;
  assign n6074 = \rEIP_reg[29]/NET0131  & n6039 ;
  assign n6075 = ~n6073 & ~n6074 ;
  assign n6076 = n5676 & ~n6075 ;
  assign n6084 = n3660 & ~n6076 ;
  assign n6085 = ~n6083 & n6084 ;
  assign n6086 = \rEIP_reg[29]/NET0131  & ~n5684 ;
  assign n6088 = n924 & ~n6075 ;
  assign n6087 = ~\EBX_reg[29]/NET0131  & ~n924 ;
  assign n6089 = n923 & ~n6087 ;
  assign n6090 = ~n6088 & n6089 ;
  assign n6091 = ~n6086 & ~n6090 ;
  assign n6092 = ~n6085 & n6091 ;
  assign n6093 = n929 & ~n6092 ;
  assign n6095 = ~n2589 & ~n2833 ;
  assign n6096 = ~n2306 & n6095 ;
  assign n6097 = ~n2359 & n6096 ;
  assign n6098 = n5954 & n6097 ;
  assign n6099 = ~n1899 & ~n6098 ;
  assign n6101 = n2379 & ~n6099 ;
  assign n6100 = ~n2379 & n6099 ;
  assign n6102 = ~\DataWidth_reg[1]/NET0131  & ~n6100 ;
  assign n6103 = ~n6101 & n6102 ;
  assign n6094 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[29]/NET0131  ;
  assign n6104 = n933 & ~n6094 ;
  assign n6105 = ~n6103 & n6104 ;
  assign n6106 = \PhyAddrPointer_reg[29]/NET0131  & n953 ;
  assign n6107 = \rEIP_reg[29]/NET0131  & ~n5667 ;
  assign n6108 = ~n6106 & ~n6107 ;
  assign n6109 = ~n6105 & n6108 ;
  assign n6110 = ~n6093 & n6109 ;
  assign n6112 = ~\PhyAddrPointer_reg[0]/NET0131  & \PhyAddrPointer_reg[1]/NET0131  ;
  assign n6113 = ~n1899 & ~n6112 ;
  assign n6115 = ~n4265 & n6113 ;
  assign n6114 = n4265 & ~n6113 ;
  assign n6116 = ~\DataWidth_reg[1]/NET0131  & ~n6114 ;
  assign n6117 = ~n6115 & n6116 ;
  assign n6111 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[2]/NET0131  ;
  assign n6118 = n933 & ~n6111 ;
  assign n6119 = ~n6117 & n6118 ;
  assign n6123 = \rEIP_reg[2]/NET0131  & ~n5684 ;
  assign n6135 = \EBX_reg[2]/NET0131  & ~n924 ;
  assign n6124 = ~\rEIP_reg[1]/NET0131  & ~\rEIP_reg[2]/NET0131  ;
  assign n6125 = ~\DataWidth_reg[1]/NET0131  & ~n5724 ;
  assign n6126 = ~n6124 & n6125 ;
  assign n6136 = n829 & n6126 ;
  assign n6137 = ~n6135 & ~n6136 ;
  assign n6138 = n923 & ~n6137 ;
  assign n6122 = n883 & n5669 ;
  assign n6127 = ~READY_n_pad & n6126 ;
  assign n6128 = \EBX_reg[31]/NET0131  & ~n5673 ;
  assign n6130 = \EBX_reg[2]/NET0131  & n6128 ;
  assign n6129 = ~\EBX_reg[2]/NET0131  & ~n6128 ;
  assign n6131 = ~n5676 & ~n6129 ;
  assign n6132 = ~n6130 & n6131 ;
  assign n6133 = ~n6127 & ~n6132 ;
  assign n6134 = n3660 & ~n6133 ;
  assign n6139 = ~n6122 & ~n6134 ;
  assign n6140 = ~n6138 & n6139 ;
  assign n6141 = ~n6123 & n6140 ;
  assign n6142 = n929 & ~n6141 ;
  assign n6120 = \PhyAddrPointer_reg[2]/NET0131  & n953 ;
  assign n6121 = \rEIP_reg[2]/NET0131  & ~n5667 ;
  assign n6143 = ~n6120 & ~n6121 ;
  assign n6144 = ~n6142 & n6143 ;
  assign n6145 = ~n6119 & n6144 ;
  assign n6146 = \rEIP_reg[31]/NET0131  & ~n5684 ;
  assign n6147 = ~\EBX_reg[29]/NET0131  & n6077 ;
  assign n6148 = n6014 & n6147 ;
  assign n6149 = ~\EBX_reg[30]/NET0131  & \EBX_reg[31]/NET0131  ;
  assign n6150 = ~n5676 & n6149 ;
  assign n6151 = n6148 & n6150 ;
  assign n6152 = \rEIP_reg[30]/NET0131  & n6074 ;
  assign n6153 = \rEIP_reg[31]/NET0131  & ~n6152 ;
  assign n6154 = ~\rEIP_reg[31]/NET0131  & n6152 ;
  assign n6155 = ~n6153 & ~n6154 ;
  assign n6156 = n5676 & ~n6155 ;
  assign n6157 = ~n6151 & ~n6156 ;
  assign n6158 = n782 & ~n6157 ;
  assign n6160 = n924 & n6155 ;
  assign n6159 = ~\EBX_reg[31]/NET0131  & ~n924 ;
  assign n6161 = n783 & ~n6159 ;
  assign n6162 = ~n6160 & n6161 ;
  assign n6163 = ~n6158 & ~n6162 ;
  assign n6164 = ~n834 & ~n6163 ;
  assign n6165 = ~n6146 & ~n6164 ;
  assign n6166 = n929 & ~n6165 ;
  assign n6167 = \DataWidth_reg[1]/NET0131  & \rEIP_reg[31]/NET0131  ;
  assign n6168 = ~n2379 & n3531 ;
  assign n6169 = n6098 & n6168 ;
  assign n6170 = ~\DataWidth_reg[1]/NET0131  & ~n2097 ;
  assign n6171 = ~n1899 & n6170 ;
  assign n6172 = n6169 & n6171 ;
  assign n6173 = ~n6167 & ~n6172 ;
  assign n6174 = n933 & ~n6173 ;
  assign n6175 = \PhyAddrPointer_reg[31]/NET0131  & n953 ;
  assign n6176 = \rEIP_reg[31]/NET0131  & ~n5667 ;
  assign n6177 = ~n6175 & ~n6176 ;
  assign n6178 = ~n6174 & n6177 ;
  assign n6179 = ~n6166 & n6178 ;
  assign n6181 = \PhyAddrPointer_reg[2]/NET0131  & n6112 ;
  assign n6182 = ~n1899 & ~n6181 ;
  assign n6184 = n3709 & ~n6182 ;
  assign n6183 = ~n3709 & n6182 ;
  assign n6185 = ~\DataWidth_reg[1]/NET0131  & ~n6183 ;
  assign n6186 = ~n6184 & n6185 ;
  assign n6180 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[3]/NET0131  ;
  assign n6187 = n933 & ~n6180 ;
  assign n6188 = ~n6186 & n6187 ;
  assign n6192 = \rEIP_reg[3]/NET0131  & ~n5684 ;
  assign n6200 = \EBX_reg[31]/NET0131  & ~n5747 ;
  assign n6202 = \EBX_reg[3]/NET0131  & n6200 ;
  assign n6201 = ~\EBX_reg[3]/NET0131  & ~n6200 ;
  assign n6203 = ~n5676 & ~n6201 ;
  assign n6204 = ~n6202 & n6203 ;
  assign n6194 = ~\rEIP_reg[3]/NET0131  & ~n5724 ;
  assign n6195 = ~\DataWidth_reg[1]/NET0131  & ~n5725 ;
  assign n6196 = ~n6194 & n6195 ;
  assign n6205 = ~READY_n_pad & n6196 ;
  assign n6206 = ~n6204 & ~n6205 ;
  assign n6207 = n3660 & ~n6206 ;
  assign n6191 = ~n868 & n5669 ;
  assign n6193 = \EBX_reg[3]/NET0131  & ~n924 ;
  assign n6197 = n829 & n6196 ;
  assign n6198 = ~n6193 & ~n6197 ;
  assign n6199 = n923 & ~n6198 ;
  assign n6208 = ~n6191 & ~n6199 ;
  assign n6209 = ~n6207 & n6208 ;
  assign n6210 = ~n6192 & n6209 ;
  assign n6211 = n929 & ~n6210 ;
  assign n6189 = \PhyAddrPointer_reg[3]/NET0131  & n953 ;
  assign n6190 = \rEIP_reg[3]/NET0131  & ~n5667 ;
  assign n6212 = ~n6189 & ~n6190 ;
  assign n6213 = ~n6211 & n6212 ;
  assign n6214 = ~n6188 & n6213 ;
  assign n6216 = ~\PhyAddrPointer_reg[0]/NET0131  & n3531 ;
  assign n6217 = ~n1899 & ~n6216 ;
  assign n6219 = ~n3534 & n6217 ;
  assign n6218 = n3534 & ~n6217 ;
  assign n6220 = ~\DataWidth_reg[1]/NET0131  & ~n6218 ;
  assign n6221 = ~n6219 & n6220 ;
  assign n6215 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[4]/NET0131  ;
  assign n6222 = n933 & ~n6215 ;
  assign n6223 = ~n6221 & n6222 ;
  assign n6225 = \rEIP_reg[4]/NET0131  & ~n5684 ;
  assign n6226 = \EBX_reg[31]/NET0131  & ~n5748 ;
  assign n6228 = ~\EBX_reg[4]/NET0131  & n6226 ;
  assign n6227 = \EBX_reg[4]/NET0131  & ~n6226 ;
  assign n6229 = ~n5676 & ~n6227 ;
  assign n6230 = ~n6228 & n6229 ;
  assign n6231 = ~\rEIP_reg[4]/NET0131  & ~n5725 ;
  assign n6232 = ~n5726 & ~n6231 ;
  assign n6233 = n5676 & ~n6232 ;
  assign n6234 = ~n6230 & ~n6233 ;
  assign n6235 = n3660 & n6234 ;
  assign n6236 = ~\EBX_reg[4]/NET0131  & ~n924 ;
  assign n6237 = n924 & ~n6232 ;
  assign n6238 = ~n6236 & ~n6237 ;
  assign n6239 = n923 & n6238 ;
  assign n6240 = ~n6235 & ~n6239 ;
  assign n6241 = ~n6225 & n6240 ;
  assign n6242 = n929 & ~n6241 ;
  assign n6224 = \rEIP_reg[4]/NET0131  & ~n5658 ;
  assign n6243 = \PhyAddrPointer_reg[4]/NET0131  & n953 ;
  assign n6244 = ~n1655 & ~n6243 ;
  assign n6245 = ~n6224 & n6244 ;
  assign n6246 = ~n6242 & n6245 ;
  assign n6247 = ~n6223 & n6246 ;
  assign n6249 = ~n1871 & ~n1899 ;
  assign n6250 = ~n6113 & ~n6249 ;
  assign n6252 = n3739 & n6250 ;
  assign n6251 = ~n3739 & ~n6250 ;
  assign n6253 = ~\DataWidth_reg[1]/NET0131  & ~n6251 ;
  assign n6254 = ~n6252 & n6253 ;
  assign n6248 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[5]/NET0131  ;
  assign n6255 = n933 & ~n6248 ;
  assign n6256 = ~n6254 & n6255 ;
  assign n6258 = \rEIP_reg[5]/NET0131  & ~n5684 ;
  assign n6259 = \EBX_reg[31]/NET0131  & ~n5749 ;
  assign n6261 = \EBX_reg[5]/NET0131  & n6259 ;
  assign n6260 = ~\EBX_reg[5]/NET0131  & ~n6259 ;
  assign n6262 = ~n5676 & ~n6260 ;
  assign n6263 = ~n6261 & n6262 ;
  assign n6264 = ~\rEIP_reg[5]/NET0131  & ~n5726 ;
  assign n6265 = ~n5727 & ~n6264 ;
  assign n6266 = ~\DataWidth_reg[1]/NET0131  & n6265 ;
  assign n6267 = ~READY_n_pad & n6266 ;
  assign n6268 = ~n6263 & ~n6267 ;
  assign n6269 = n3660 & ~n6268 ;
  assign n6270 = \EBX_reg[5]/NET0131  & ~n924 ;
  assign n6271 = n829 & n6266 ;
  assign n6272 = ~n6270 & ~n6271 ;
  assign n6273 = n923 & ~n6272 ;
  assign n6274 = ~n6269 & ~n6273 ;
  assign n6275 = ~n6258 & n6274 ;
  assign n6276 = n929 & ~n6275 ;
  assign n6257 = \rEIP_reg[5]/NET0131  & ~n5658 ;
  assign n6277 = \PhyAddrPointer_reg[5]/NET0131  & n953 ;
  assign n6278 = ~n1655 & ~n6277 ;
  assign n6279 = ~n6257 & n6278 ;
  assign n6280 = ~n6276 & n6279 ;
  assign n6281 = ~n6256 & n6280 ;
  assign n6283 = ~\PhyAddrPointer_reg[0]/NET0131  & n3239 ;
  assign n6284 = ~n1899 & ~n6283 ;
  assign n6286 = n3747 & ~n6284 ;
  assign n6285 = ~n3747 & n6284 ;
  assign n6287 = ~\DataWidth_reg[1]/NET0131  & ~n6285 ;
  assign n6288 = ~n6286 & n6287 ;
  assign n6282 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[6]/NET0131  ;
  assign n6289 = n933 & ~n6282 ;
  assign n6290 = ~n6288 & n6289 ;
  assign n6292 = \rEIP_reg[6]/NET0131  & ~n5684 ;
  assign n6293 = ~\EBX_reg[6]/NET0131  & ~n924 ;
  assign n6294 = ~\rEIP_reg[6]/NET0131  & ~n5727 ;
  assign n6295 = ~n5728 & ~n6294 ;
  assign n6296 = n924 & ~n6295 ;
  assign n6297 = ~n6293 & ~n6296 ;
  assign n6298 = n923 & n6297 ;
  assign n6299 = n5676 & ~n6295 ;
  assign n6300 = \EBX_reg[31]/NET0131  & ~n5750 ;
  assign n6302 = ~\EBX_reg[6]/NET0131  & n6300 ;
  assign n6301 = \EBX_reg[6]/NET0131  & ~n6300 ;
  assign n6303 = ~n5676 & ~n6301 ;
  assign n6304 = ~n6302 & n6303 ;
  assign n6305 = ~n6299 & ~n6304 ;
  assign n6306 = n3660 & n6305 ;
  assign n6307 = ~n6298 & ~n6306 ;
  assign n6308 = ~n6292 & n6307 ;
  assign n6309 = n929 & ~n6308 ;
  assign n6291 = \rEIP_reg[6]/NET0131  & ~n5658 ;
  assign n6310 = \PhyAddrPointer_reg[6]/NET0131  & n953 ;
  assign n6311 = ~n1655 & ~n6310 ;
  assign n6312 = ~n6291 & n6311 ;
  assign n6313 = ~n6309 & n6312 ;
  assign n6314 = ~n6290 & n6313 ;
  assign n6316 = ~n1873 & ~n1899 ;
  assign n6317 = ~n6113 & ~n6316 ;
  assign n6319 = ~n3242 & ~n6317 ;
  assign n6318 = n3242 & n6317 ;
  assign n6320 = ~\DataWidth_reg[1]/NET0131  & ~n6318 ;
  assign n6321 = ~n6319 & n6320 ;
  assign n6315 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[7]/NET0131  ;
  assign n6322 = n933 & ~n6315 ;
  assign n6323 = ~n6321 & n6322 ;
  assign n6325 = \rEIP_reg[7]/NET0131  & ~n5684 ;
  assign n6326 = ~\EBX_reg[7]/NET0131  & ~n924 ;
  assign n6327 = ~\rEIP_reg[7]/NET0131  & ~n5728 ;
  assign n6328 = ~n5729 & ~n6327 ;
  assign n6329 = n924 & ~n6328 ;
  assign n6330 = ~n6326 & ~n6329 ;
  assign n6331 = n783 & n6330 ;
  assign n6333 = \EBX_reg[31]/NET0131  & ~n5751 ;
  assign n6335 = ~\EBX_reg[7]/NET0131  & n6333 ;
  assign n6334 = \EBX_reg[7]/NET0131  & ~n6333 ;
  assign n6336 = ~n5676 & ~n6334 ;
  assign n6337 = ~n6335 & n6336 ;
  assign n6332 = n5676 & ~n6328 ;
  assign n6338 = n782 & ~n6332 ;
  assign n6339 = ~n6337 & n6338 ;
  assign n6340 = ~n6331 & ~n6339 ;
  assign n6341 = ~n834 & ~n6340 ;
  assign n6342 = ~n6325 & ~n6341 ;
  assign n6343 = n929 & ~n6342 ;
  assign n6324 = \rEIP_reg[7]/NET0131  & ~n5658 ;
  assign n6344 = \PhyAddrPointer_reg[7]/NET0131  & n953 ;
  assign n6345 = ~n1655 & ~n6344 ;
  assign n6346 = ~n6324 & n6345 ;
  assign n6347 = ~n6343 & n6346 ;
  assign n6348 = ~n6323 & n6347 ;
  assign n6350 = ~n1899 & ~n5706 ;
  assign n6352 = n2857 & ~n6350 ;
  assign n6351 = ~n2857 & n6350 ;
  assign n6353 = ~\DataWidth_reg[1]/NET0131  & ~n6351 ;
  assign n6354 = ~n6352 & n6353 ;
  assign n6349 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[8]/NET0131  ;
  assign n6355 = n933 & ~n6349 ;
  assign n6356 = ~n6354 & n6355 ;
  assign n6358 = \rEIP_reg[8]/NET0131  & ~n5684 ;
  assign n6359 = ~\EBX_reg[8]/NET0131  & ~n924 ;
  assign n6360 = ~\rEIP_reg[8]/NET0131  & ~n5729 ;
  assign n6361 = ~n5730 & ~n6360 ;
  assign n6362 = n924 & ~n6361 ;
  assign n6363 = ~n6359 & ~n6362 ;
  assign n6364 = n923 & n6363 ;
  assign n6366 = \EBX_reg[31]/NET0131  & ~n5752 ;
  assign n6368 = ~\EBX_reg[8]/NET0131  & n6366 ;
  assign n6367 = \EBX_reg[8]/NET0131  & ~n6366 ;
  assign n6369 = ~n5676 & ~n6367 ;
  assign n6370 = ~n6368 & n6369 ;
  assign n6365 = n5676 & ~n6361 ;
  assign n6371 = n3660 & ~n6365 ;
  assign n6372 = ~n6370 & n6371 ;
  assign n6373 = ~n6364 & ~n6372 ;
  assign n6374 = ~n6358 & n6373 ;
  assign n6375 = n929 & ~n6374 ;
  assign n6357 = \rEIP_reg[8]/NET0131  & ~n5658 ;
  assign n6376 = \PhyAddrPointer_reg[8]/NET0131  & n953 ;
  assign n6377 = ~n1655 & ~n6376 ;
  assign n6378 = ~n6357 & n6377 ;
  assign n6379 = ~n6375 & n6378 ;
  assign n6380 = ~n6356 & n6379 ;
  assign n6382 = ~\PhyAddrPointer_reg[0]/NET0131  & n2233 ;
  assign n6383 = ~n1899 & ~n6382 ;
  assign n6385 = ~n3260 & n6383 ;
  assign n6384 = n3260 & ~n6383 ;
  assign n6386 = ~\DataWidth_reg[1]/NET0131  & ~n6384 ;
  assign n6387 = ~n6385 & n6386 ;
  assign n6381 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[9]/NET0131  ;
  assign n6388 = n933 & ~n6381 ;
  assign n6389 = ~n6387 & n6388 ;
  assign n6392 = \EBX_reg[31]/NET0131  & ~n5753 ;
  assign n6394 = \EBX_reg[9]/NET0131  & n6392 ;
  assign n6393 = ~\EBX_reg[9]/NET0131  & ~n6392 ;
  assign n6395 = ~n5676 & ~n6393 ;
  assign n6396 = ~n6394 & n6395 ;
  assign n6397 = ~\rEIP_reg[9]/NET0131  & ~n5730 ;
  assign n6398 = ~n5731 & ~n6397 ;
  assign n6399 = ~\DataWidth_reg[1]/NET0131  & n6398 ;
  assign n6400 = ~READY_n_pad & n6399 ;
  assign n6401 = ~n6396 & ~n6400 ;
  assign n6402 = n3660 & ~n6401 ;
  assign n6391 = \rEIP_reg[9]/NET0131  & ~n5684 ;
  assign n6403 = \EBX_reg[9]/NET0131  & ~n924 ;
  assign n6404 = n829 & n6399 ;
  assign n6405 = ~n6403 & ~n6404 ;
  assign n6406 = n923 & ~n6405 ;
  assign n6407 = ~n6391 & ~n6406 ;
  assign n6408 = ~n6402 & n6407 ;
  assign n6409 = n929 & ~n6408 ;
  assign n6390 = \rEIP_reg[9]/NET0131  & ~n5658 ;
  assign n6410 = \PhyAddrPointer_reg[9]/NET0131  & n953 ;
  assign n6411 = ~n1655 & ~n6410 ;
  assign n6412 = ~n6390 & n6411 ;
  assign n6413 = ~n6409 & n6412 ;
  assign n6414 = ~n6389 & n6413 ;
  assign n6416 = \PhyAddrPointer_reg[1]/NET0131  & ~n2739 ;
  assign n6417 = n3613 & ~n6416 ;
  assign n6418 = n929 & ~n6417 ;
  assign n6419 = ~n969 & n1902 ;
  assign n6420 = \PhyAddrPointer_reg[1]/NET0131  & ~n6419 ;
  assign n6415 = ~\PhyAddrPointer_reg[1]/NET0131  & n2100 ;
  assign n6421 = ~n3593 & ~n6415 ;
  assign n6422 = ~n6420 & n6421 ;
  assign n6423 = ~n6418 & n6422 ;
  assign n6425 = \PhyAddrPointer_reg[9]/NET0131  & n6382 ;
  assign n6426 = ~n1899 & ~n6425 ;
  assign n6428 = n3221 & ~n6426 ;
  assign n6427 = ~n3221 & n6426 ;
  assign n6429 = ~\DataWidth_reg[1]/NET0131  & ~n6427 ;
  assign n6430 = ~n6428 & n6429 ;
  assign n6424 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[10]/NET0131  ;
  assign n6431 = n933 & ~n6424 ;
  assign n6432 = ~n6430 & n6431 ;
  assign n6442 = ~\EBX_reg[9]/NET0131  & n5753 ;
  assign n6443 = \EBX_reg[31]/NET0131  & ~n6442 ;
  assign n6445 = \EBX_reg[10]/NET0131  & ~n6443 ;
  assign n6444 = ~\EBX_reg[10]/NET0131  & n6443 ;
  assign n6446 = ~n5676 & ~n6444 ;
  assign n6447 = ~n6445 & n6446 ;
  assign n6436 = ~\rEIP_reg[10]/NET0131  & ~n5731 ;
  assign n6437 = ~n5732 & ~n6436 ;
  assign n6441 = n5676 & ~n6437 ;
  assign n6448 = n3660 & ~n6441 ;
  assign n6449 = ~n6447 & n6448 ;
  assign n6434 = \rEIP_reg[10]/NET0131  & ~n5684 ;
  assign n6438 = n924 & ~n6437 ;
  assign n6435 = ~\EBX_reg[10]/NET0131  & ~n924 ;
  assign n6439 = n923 & ~n6435 ;
  assign n6440 = ~n6438 & n6439 ;
  assign n6450 = ~n6434 & ~n6440 ;
  assign n6451 = ~n6449 & n6450 ;
  assign n6452 = n929 & ~n6451 ;
  assign n6433 = \rEIP_reg[10]/NET0131  & ~n5658 ;
  assign n6453 = \PhyAddrPointer_reg[10]/NET0131  & n953 ;
  assign n6454 = ~n1655 & ~n6453 ;
  assign n6455 = ~n6433 & n6454 ;
  assign n6456 = ~n6452 & n6455 ;
  assign n6457 = ~n6432 & n6456 ;
  assign n6459 = n3531 & n5706 ;
  assign n6460 = n1877 & n6459 ;
  assign n6461 = ~n1899 & ~n6460 ;
  assign n6463 = ~n2471 & n6461 ;
  assign n6462 = n2471 & ~n6461 ;
  assign n6464 = ~\DataWidth_reg[1]/NET0131  & ~n6462 ;
  assign n6465 = ~n6463 & n6464 ;
  assign n6458 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[11]/NET0131  ;
  assign n6466 = n933 & ~n6458 ;
  assign n6467 = ~n6465 & n6466 ;
  assign n6477 = \EBX_reg[31]/NET0131  & ~n5755 ;
  assign n6479 = ~\EBX_reg[11]/NET0131  & n6477 ;
  assign n6478 = \EBX_reg[11]/NET0131  & ~n6477 ;
  assign n6480 = ~n5676 & ~n6478 ;
  assign n6481 = ~n6479 & n6480 ;
  assign n6471 = ~\rEIP_reg[11]/NET0131  & ~n5732 ;
  assign n6472 = ~n5733 & ~n6471 ;
  assign n6476 = n5676 & ~n6472 ;
  assign n6482 = n3660 & ~n6476 ;
  assign n6483 = ~n6481 & n6482 ;
  assign n6469 = \rEIP_reg[11]/NET0131  & ~n5684 ;
  assign n6473 = n924 & ~n6472 ;
  assign n6470 = ~\EBX_reg[11]/NET0131  & ~n924 ;
  assign n6474 = n923 & ~n6470 ;
  assign n6475 = ~n6473 & n6474 ;
  assign n6484 = ~n6469 & ~n6475 ;
  assign n6485 = ~n6483 & n6484 ;
  assign n6486 = n929 & ~n6485 ;
  assign n6468 = \rEIP_reg[11]/NET0131  & ~n5658 ;
  assign n6487 = \PhyAddrPointer_reg[11]/NET0131  & n953 ;
  assign n6488 = ~n1655 & ~n6487 ;
  assign n6489 = ~n6468 & n6488 ;
  assign n6490 = ~n6486 & n6489 ;
  assign n6491 = ~n6467 & n6490 ;
  assign n6493 = ~\PhyAddrPointer_reg[12]/NET0131  & ~n2470 ;
  assign n6494 = ~n2678 & ~n6493 ;
  assign n6495 = n2465 & n6459 ;
  assign n6496 = ~n1899 & ~n6495 ;
  assign n6498 = n6494 & ~n6496 ;
  assign n6497 = ~n6494 & n6496 ;
  assign n6499 = ~\DataWidth_reg[1]/NET0131  & ~n6497 ;
  assign n6500 = ~n6498 & n6499 ;
  assign n6492 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[12]/NET0131  ;
  assign n6501 = n933 & ~n6492 ;
  assign n6502 = ~n6500 & n6501 ;
  assign n6504 = \rEIP_reg[12]/NET0131  & ~n5684 ;
  assign n6506 = \rEIP_reg[12]/NET0131  & n5733 ;
  assign n6507 = ~\rEIP_reg[12]/NET0131  & ~n5733 ;
  assign n6508 = ~n6506 & ~n6507 ;
  assign n6509 = n924 & ~n6508 ;
  assign n6505 = ~\EBX_reg[12]/NET0131  & ~n924 ;
  assign n6510 = n783 & ~n6505 ;
  assign n6511 = ~n6509 & n6510 ;
  assign n6513 = ~\EBX_reg[11]/NET0131  & n5755 ;
  assign n6514 = \EBX_reg[31]/NET0131  & ~n6513 ;
  assign n6516 = ~\EBX_reg[12]/NET0131  & n6514 ;
  assign n6515 = \EBX_reg[12]/NET0131  & ~n6514 ;
  assign n6517 = ~n5676 & ~n6515 ;
  assign n6518 = ~n6516 & n6517 ;
  assign n6512 = n5676 & ~n6508 ;
  assign n6519 = n782 & ~n6512 ;
  assign n6520 = ~n6518 & n6519 ;
  assign n6521 = ~n6511 & ~n6520 ;
  assign n6522 = ~n834 & ~n6521 ;
  assign n6523 = ~n6504 & ~n6522 ;
  assign n6524 = n929 & ~n6523 ;
  assign n6503 = \rEIP_reg[12]/NET0131  & ~n5658 ;
  assign n6525 = \PhyAddrPointer_reg[12]/NET0131  & n953 ;
  assign n6526 = ~n1655 & ~n6525 ;
  assign n6527 = ~n6503 & n6526 ;
  assign n6528 = ~n6524 & n6527 ;
  assign n6529 = ~n6502 & n6528 ;
  assign n6531 = ~n1899 & ~n2674 ;
  assign n6532 = ~n6350 & ~n6531 ;
  assign n6534 = ~n2680 & ~n6532 ;
  assign n6533 = n2680 & n6532 ;
  assign n6535 = ~\DataWidth_reg[1]/NET0131  & ~n6533 ;
  assign n6536 = ~n6534 & n6535 ;
  assign n6530 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[13]/NET0131  ;
  assign n6537 = n933 & ~n6530 ;
  assign n6538 = ~n6536 & n6537 ;
  assign n6540 = \rEIP_reg[13]/NET0131  & ~n5684 ;
  assign n6542 = ~\rEIP_reg[13]/NET0131  & ~n6506 ;
  assign n6543 = n5733 & n5734 ;
  assign n6544 = ~n6542 & ~n6543 ;
  assign n6545 = n924 & ~n6544 ;
  assign n6541 = ~\EBX_reg[13]/NET0131  & ~n924 ;
  assign n6546 = n783 & ~n6541 ;
  assign n6547 = ~n6545 & n6546 ;
  assign n6549 = \EBX_reg[31]/NET0131  & ~n5757 ;
  assign n6551 = ~\EBX_reg[13]/NET0131  & n6549 ;
  assign n6550 = \EBX_reg[13]/NET0131  & ~n6549 ;
  assign n6552 = ~n5676 & ~n6550 ;
  assign n6553 = ~n6551 & n6552 ;
  assign n6548 = n5676 & ~n6544 ;
  assign n6554 = n782 & ~n6548 ;
  assign n6555 = ~n6553 & n6554 ;
  assign n6556 = ~n6547 & ~n6555 ;
  assign n6557 = ~n834 & ~n6556 ;
  assign n6558 = ~n6540 & ~n6557 ;
  assign n6559 = n929 & ~n6558 ;
  assign n6539 = \rEIP_reg[13]/NET0131  & ~n5658 ;
  assign n6560 = \PhyAddrPointer_reg[13]/NET0131  & n953 ;
  assign n6561 = ~n1655 & ~n6560 ;
  assign n6562 = ~n6539 & n6561 ;
  assign n6563 = ~n6559 & n6562 ;
  assign n6564 = ~n6538 & n6563 ;
  assign n6566 = n1880 & n6459 ;
  assign n6567 = ~n1899 & ~n6566 ;
  assign n6569 = ~n2486 & n6567 ;
  assign n6568 = n2486 & ~n6567 ;
  assign n6570 = ~\DataWidth_reg[1]/NET0131  & ~n6568 ;
  assign n6571 = ~n6569 & n6570 ;
  assign n6565 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[14]/NET0131  ;
  assign n6572 = n933 & ~n6565 ;
  assign n6573 = ~n6571 & n6572 ;
  assign n6575 = \rEIP_reg[14]/NET0131  & ~n5684 ;
  assign n6577 = ~\rEIP_reg[14]/NET0131  & ~n6543 ;
  assign n6578 = n5733 & n5735 ;
  assign n6579 = ~n6577 & ~n6578 ;
  assign n6580 = n924 & ~n6579 ;
  assign n6576 = ~\EBX_reg[14]/NET0131  & ~n924 ;
  assign n6581 = n783 & ~n6576 ;
  assign n6582 = ~n6580 & n6581 ;
  assign n6584 = \EBX_reg[31]/NET0131  & ~n5758 ;
  assign n6586 = \EBX_reg[14]/NET0131  & ~n6584 ;
  assign n6585 = ~\EBX_reg[14]/NET0131  & n6584 ;
  assign n6587 = ~n5676 & ~n6585 ;
  assign n6588 = ~n6586 & n6587 ;
  assign n6583 = n5676 & ~n6579 ;
  assign n6589 = n782 & ~n6583 ;
  assign n6590 = ~n6588 & n6589 ;
  assign n6591 = ~n6582 & ~n6590 ;
  assign n6592 = ~n834 & ~n6591 ;
  assign n6593 = ~n6575 & ~n6592 ;
  assign n6594 = n929 & ~n6593 ;
  assign n6574 = \rEIP_reg[14]/NET0131  & ~n5658 ;
  assign n6595 = \PhyAddrPointer_reg[14]/NET0131  & n953 ;
  assign n6596 = ~n1655 & ~n6595 ;
  assign n6597 = ~n6574 & n6596 ;
  assign n6598 = ~n6594 & n6597 ;
  assign n6599 = ~n6573 & n6598 ;
  assign n6601 = ~n2486 & n6566 ;
  assign n6602 = ~n1899 & ~n6601 ;
  assign n6604 = ~n2240 & n6602 ;
  assign n6603 = n2240 & ~n6602 ;
  assign n6605 = ~\DataWidth_reg[1]/NET0131  & ~n6603 ;
  assign n6606 = ~n6604 & n6605 ;
  assign n6600 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[15]/NET0131  ;
  assign n6607 = n933 & ~n6600 ;
  assign n6608 = ~n6606 & n6607 ;
  assign n6610 = \rEIP_reg[15]/NET0131  & ~n5684 ;
  assign n6611 = ~\EBX_reg[15]/NET0131  & ~n924 ;
  assign n6612 = n783 & ~n6611 ;
  assign n6613 = \EBX_reg[31]/NET0131  & ~n5759 ;
  assign n6615 = ~\EBX_reg[15]/NET0131  & n6613 ;
  assign n6614 = \EBX_reg[15]/NET0131  & ~n6613 ;
  assign n6616 = ~n5676 & ~n6614 ;
  assign n6617 = ~n6615 & n6616 ;
  assign n6618 = n782 & ~n6617 ;
  assign n6619 = ~n6612 & ~n6618 ;
  assign n6621 = ~\rEIP_reg[15]/NET0131  & ~n6578 ;
  assign n6622 = ~n5737 & ~n6621 ;
  assign n6620 = n828 & n6612 ;
  assign n6623 = n5676 & ~n6620 ;
  assign n6624 = ~n6622 & n6623 ;
  assign n6625 = ~n834 & ~n6624 ;
  assign n6626 = ~n6619 & n6625 ;
  assign n6627 = ~n6610 & ~n6626 ;
  assign n6628 = n929 & ~n6627 ;
  assign n6609 = \rEIP_reg[15]/NET0131  & ~n5658 ;
  assign n6629 = \PhyAddrPointer_reg[15]/NET0131  & n953 ;
  assign n6630 = ~n1655 & ~n6629 ;
  assign n6631 = ~n6609 & n6630 ;
  assign n6632 = ~n6628 & n6631 ;
  assign n6633 = ~n6608 & n6632 ;
  assign n6635 = ~n1899 & n2240 ;
  assign n6636 = ~n6602 & ~n6635 ;
  assign n6638 = ~n2715 & ~n6636 ;
  assign n6637 = n2715 & n6636 ;
  assign n6639 = ~\DataWidth_reg[1]/NET0131  & ~n6637 ;
  assign n6640 = ~n6638 & n6639 ;
  assign n6634 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[16]/NET0131  ;
  assign n6641 = n933 & ~n6634 ;
  assign n6642 = ~n6640 & n6641 ;
  assign n6644 = \rEIP_reg[16]/NET0131  & ~n5684 ;
  assign n6646 = ~\rEIP_reg[16]/NET0131  & ~n5737 ;
  assign n6647 = ~n5738 & ~n6646 ;
  assign n6648 = n924 & ~n6647 ;
  assign n6645 = ~\EBX_reg[16]/NET0131  & ~n924 ;
  assign n6649 = n783 & ~n6645 ;
  assign n6650 = ~n6648 & n6649 ;
  assign n6652 = ~\EBX_reg[15]/NET0131  & n5759 ;
  assign n6653 = \EBX_reg[31]/NET0131  & ~n6652 ;
  assign n6655 = \EBX_reg[16]/NET0131  & ~n6653 ;
  assign n6654 = ~\EBX_reg[16]/NET0131  & n6653 ;
  assign n6656 = ~n5676 & ~n6654 ;
  assign n6657 = ~n6655 & n6656 ;
  assign n6651 = n5676 & ~n6647 ;
  assign n6658 = n782 & ~n6651 ;
  assign n6659 = ~n6657 & n6658 ;
  assign n6660 = ~n6650 & ~n6659 ;
  assign n6661 = ~n834 & ~n6660 ;
  assign n6662 = ~n6644 & ~n6661 ;
  assign n6663 = n929 & ~n6662 ;
  assign n6643 = \rEIP_reg[16]/NET0131  & ~n5658 ;
  assign n6664 = \PhyAddrPointer_reg[16]/NET0131  & n953 ;
  assign n6665 = ~n1655 & ~n6664 ;
  assign n6666 = ~n6643 & n6665 ;
  assign n6667 = ~n6663 & n6666 ;
  assign n6668 = ~n6642 & n6667 ;
  assign n6670 = ~n1899 & ~n5710 ;
  assign n6672 = ~n2752 & n6670 ;
  assign n6671 = n2752 & ~n6670 ;
  assign n6673 = ~\DataWidth_reg[1]/NET0131  & ~n6671 ;
  assign n6674 = ~n6672 & n6673 ;
  assign n6669 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[17]/NET0131  ;
  assign n6675 = n933 & ~n6669 ;
  assign n6676 = ~n6674 & n6675 ;
  assign n6681 = n783 & ~n828 ;
  assign n6688 = \EBX_reg[31]/NET0131  & ~n5761 ;
  assign n6689 = ~n6681 & n6688 ;
  assign n6682 = ~n782 & ~n6681 ;
  assign n6690 = \EBX_reg[17]/NET0131  & ~n6682 ;
  assign n6691 = ~n6689 & n6690 ;
  assign n6692 = ~\EBX_reg[17]/NET0131  & n782 ;
  assign n6693 = n6688 & n6692 ;
  assign n6694 = ~n5676 & ~n6693 ;
  assign n6695 = ~n6691 & n6694 ;
  assign n6684 = ~\rEIP_reg[17]/NET0131  & ~n5738 ;
  assign n6683 = \rEIP_reg[17]/NET0131  & n5738 ;
  assign n6685 = ~n6682 & ~n6683 ;
  assign n6686 = ~n6684 & n6685 ;
  assign n6687 = n5676 & ~n6686 ;
  assign n6696 = ~n834 & ~n6687 ;
  assign n6697 = ~n6695 & n6696 ;
  assign n6678 = \EBX_reg[17]/NET0131  & n828 ;
  assign n6679 = n923 & n6678 ;
  assign n6680 = \rEIP_reg[17]/NET0131  & ~n5684 ;
  assign n6698 = ~n6679 & ~n6680 ;
  assign n6699 = ~n6697 & n6698 ;
  assign n6700 = n929 & ~n6699 ;
  assign n6677 = \rEIP_reg[17]/NET0131  & ~n5658 ;
  assign n6701 = \PhyAddrPointer_reg[17]/NET0131  & n953 ;
  assign n6702 = ~n1655 & ~n6701 ;
  assign n6703 = ~n6677 & n6702 ;
  assign n6704 = ~n6700 & n6703 ;
  assign n6705 = ~n6676 & n6704 ;
  assign n6707 = n3531 & n5711 ;
  assign n6708 = ~n1899 & ~n6707 ;
  assign n6710 = ~n2781 & n6708 ;
  assign n6709 = n2781 & ~n6708 ;
  assign n6711 = ~\DataWidth_reg[1]/NET0131  & ~n6709 ;
  assign n6712 = ~n6710 & n6711 ;
  assign n6706 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[18]/NET0131  ;
  assign n6713 = n933 & ~n6706 ;
  assign n6714 = ~n6712 & n6713 ;
  assign n6716 = \rEIP_reg[18]/NET0131  & ~n5684 ;
  assign n6717 = ~\EBX_reg[18]/NET0131  & ~n924 ;
  assign n6718 = n783 & ~n6717 ;
  assign n6719 = \EBX_reg[31]/NET0131  & ~n5762 ;
  assign n6721 = ~\EBX_reg[18]/NET0131  & n6719 ;
  assign n6720 = \EBX_reg[18]/NET0131  & ~n6719 ;
  assign n6722 = ~n5676 & ~n6720 ;
  assign n6723 = ~n6721 & n6722 ;
  assign n6724 = n782 & ~n6723 ;
  assign n6725 = ~n6718 & ~n6724 ;
  assign n6727 = ~\rEIP_reg[18]/NET0131  & ~n6683 ;
  assign n6728 = ~n5740 & ~n6727 ;
  assign n6726 = n828 & n6718 ;
  assign n6729 = n5676 & ~n6726 ;
  assign n6730 = ~n6728 & n6729 ;
  assign n6731 = ~n834 & ~n6730 ;
  assign n6732 = ~n6725 & n6731 ;
  assign n6733 = ~n6716 & ~n6732 ;
  assign n6734 = n929 & ~n6733 ;
  assign n6715 = \rEIP_reg[18]/NET0131  & ~n5658 ;
  assign n6735 = \PhyAddrPointer_reg[18]/NET0131  & n953 ;
  assign n6736 = ~n1655 & ~n6735 ;
  assign n6737 = ~n6715 & n6736 ;
  assign n6738 = ~n6734 & n6737 ;
  assign n6739 = ~n6714 & n6738 ;
  assign n6741 = ~n1899 & n2781 ;
  assign n6742 = ~n6708 & ~n6741 ;
  assign n6744 = ~n2510 & ~n6742 ;
  assign n6743 = n2510 & n6742 ;
  assign n6745 = ~\DataWidth_reg[1]/NET0131  & ~n6743 ;
  assign n6746 = ~n6744 & n6745 ;
  assign n6740 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[19]/NET0131  ;
  assign n6747 = n933 & ~n6740 ;
  assign n6748 = ~n6746 & n6747 ;
  assign n6753 = \EBX_reg[31]/NET0131  & ~n5763 ;
  assign n6755 = ~\EBX_reg[19]/NET0131  & n6753 ;
  assign n6754 = \EBX_reg[19]/NET0131  & ~n6753 ;
  assign n6756 = ~n5676 & ~n6754 ;
  assign n6757 = ~n6755 & n6756 ;
  assign n6750 = ~\rEIP_reg[19]/NET0131  & ~n5740 ;
  assign n6751 = ~n5741 & ~n6750 ;
  assign n6752 = n5676 & ~n6751 ;
  assign n6758 = n3660 & ~n6752 ;
  assign n6759 = ~n6757 & n6758 ;
  assign n6760 = \rEIP_reg[19]/NET0131  & ~n5684 ;
  assign n6762 = ~n828 & n6752 ;
  assign n6761 = ~\EBX_reg[19]/NET0131  & ~n924 ;
  assign n6763 = n923 & ~n6761 ;
  assign n6764 = ~n6762 & n6763 ;
  assign n6765 = ~n6760 & ~n6764 ;
  assign n6766 = ~n6759 & n6765 ;
  assign n6767 = n929 & ~n6766 ;
  assign n6749 = \rEIP_reg[19]/NET0131  & ~n5658 ;
  assign n6768 = \PhyAddrPointer_reg[19]/NET0131  & n953 ;
  assign n6769 = ~n1655 & ~n6768 ;
  assign n6770 = ~n6749 & n6769 ;
  assign n6771 = ~n6767 & n6770 ;
  assign n6772 = ~n6748 & n6771 ;
  assign n6776 = ~\RequestPending_reg/NET0131  & n834 ;
  assign n6777 = ~n850 & ~n6776 ;
  assign n6774 = \RequestPending_reg/NET0131  & n785 ;
  assign n6775 = ~\DataWidth_reg[1]/NET0131  & n923 ;
  assign n6778 = ~n6774 & ~n6775 ;
  assign n6779 = ~n6777 & n6778 ;
  assign n6780 = n929 & ~n6779 ;
  assign n6773 = ~n939 & ~n1655 ;
  assign n6781 = n931 & n950 ;
  assign n6782 = n3179 & ~n6781 ;
  assign n6783 = \RequestPending_reg/NET0131  & ~n6782 ;
  assign n6784 = n6773 & ~n6783 ;
  assign n6785 = ~n6780 & n6784 ;
  assign n6787 = ~\EAX_reg[23]/NET0131  & ~n3683 ;
  assign n6788 = ~n3811 & ~n6787 ;
  assign n6789 = ~n828 & ~n6788 ;
  assign n6790 = n923 & ~n6789 ;
  assign n6791 = n3827 & ~n6790 ;
  assign n6792 = \Datao[23]_pad  & ~n6791 ;
  assign n6793 = n923 & n6788 ;
  assign n6794 = ~n828 & n6793 ;
  assign n6795 = ~n6792 & ~n6794 ;
  assign n6796 = n929 & ~n6795 ;
  assign n6786 = \uWord_reg[7]/NET0131  & n3809 ;
  assign n6797 = \Datao[23]_pad  & ~n3821 ;
  assign n6798 = ~n6786 & ~n6797 ;
  assign n6799 = ~n6796 & n6798 ;
  assign n6801 = ~\EAX_reg[19]/NET0131  & ~n3682 ;
  assign n6802 = ~n4281 & ~n6801 ;
  assign n6803 = ~n828 & ~n6802 ;
  assign n6804 = n923 & ~n6803 ;
  assign n6805 = n3827 & ~n6804 ;
  assign n6806 = \Datao[19]_pad  & ~n6805 ;
  assign n6807 = n923 & n6802 ;
  assign n6808 = ~n828 & n6807 ;
  assign n6809 = ~n6806 & ~n6808 ;
  assign n6810 = n929 & ~n6809 ;
  assign n6800 = \uWord_reg[3]/NET0131  & n3809 ;
  assign n6811 = \Datao[19]_pad  & ~n3821 ;
  assign n6812 = ~n6800 & ~n6811 ;
  assign n6813 = ~n6810 & n6812 ;
  assign n6814 = \EAX_reg[2]/NET0131  & ~n4671 ;
  assign n6816 = \Datai[2]_pad  & n846 ;
  assign n6817 = ~n841 & n6816 ;
  assign n6815 = ~n1197 & n2937 ;
  assign n6818 = ~\EAX_reg[2]/NET0131  & ~n3136 ;
  assign n6819 = ~n3137 & ~n6818 ;
  assign n6820 = n3132 & n6819 ;
  assign n6821 = ~n6815 & ~n6820 ;
  assign n6822 = ~n6817 & n6821 ;
  assign n6823 = n929 & ~n6822 ;
  assign n6824 = ~n6814 & ~n6823 ;
  assign n6825 = \uWord_reg[3]/NET0131  & ~n3655 ;
  assign n6826 = \Datai[3]_pad  & n846 ;
  assign n6827 = READY_n_pad & \uWord_reg[3]/NET0131  ;
  assign n6828 = ~n6826 & ~n6827 ;
  assign n6829 = n782 & ~n6828 ;
  assign n6830 = \uWord_reg[3]/NET0131  & n3661 ;
  assign n6831 = ~n6807 & ~n6830 ;
  assign n6832 = ~n6829 & n6831 ;
  assign n6833 = n929 & ~n6832 ;
  assign n6834 = ~n6825 & ~n6833 ;
  assign n6835 = \uWord_reg[7]/NET0131  & ~n3655 ;
  assign n6836 = READY_n_pad & \uWord_reg[7]/NET0131  ;
  assign n6837 = ~n4674 & ~n6836 ;
  assign n6838 = n782 & ~n6837 ;
  assign n6839 = \uWord_reg[7]/NET0131  & n3661 ;
  assign n6840 = ~n6793 & ~n6839 ;
  assign n6841 = ~n6838 & n6840 ;
  assign n6842 = n929 & ~n6841 ;
  assign n6843 = ~n6835 & ~n6842 ;
  assign n6844 = \EAX_reg[3]/NET0131  & ~n4671 ;
  assign n6846 = ~n841 & n6826 ;
  assign n6845 = ~n1162 & n2937 ;
  assign n6847 = ~\EAX_reg[3]/NET0131  & ~n3137 ;
  assign n6848 = ~n3138 & ~n6847 ;
  assign n6849 = n3132 & n6848 ;
  assign n6850 = ~n6845 & ~n6849 ;
  assign n6851 = ~n6846 & n6850 ;
  assign n6852 = n929 & ~n6851 ;
  assign n6853 = ~n6844 & ~n6852 ;
  assign n6854 = \EAX_reg[4]/NET0131  & ~n4671 ;
  assign n6856 = ~n841 & n4298 ;
  assign n6855 = ~n1124 & n2937 ;
  assign n6857 = ~\EAX_reg[4]/NET0131  & ~n3138 ;
  assign n6858 = ~n3139 & ~n6857 ;
  assign n6859 = n3132 & n6858 ;
  assign n6860 = ~n6855 & ~n6859 ;
  assign n6861 = ~n6856 & n6860 ;
  assign n6862 = n929 & ~n6861 ;
  assign n6863 = ~n6854 & ~n6862 ;
  assign n6864 = \EAX_reg[5]/NET0131  & ~n4671 ;
  assign n6866 = \Datai[5]_pad  & n846 ;
  assign n6867 = ~n841 & n6866 ;
  assign n6865 = ~n1088 & n2937 ;
  assign n6868 = ~\EAX_reg[5]/NET0131  & ~n3139 ;
  assign n6869 = ~n3140 & ~n6868 ;
  assign n6870 = n3132 & n6869 ;
  assign n6871 = ~n6865 & ~n6870 ;
  assign n6872 = ~n6867 & n6871 ;
  assign n6873 = n929 & ~n6872 ;
  assign n6874 = ~n6864 & ~n6873 ;
  assign n6875 = \EAX_reg[6]/NET0131  & ~n4671 ;
  assign n6877 = \Datai[6]_pad  & n843 ;
  assign n6876 = ~n1050 & n2937 ;
  assign n6878 = ~\EAX_reg[6]/NET0131  & ~n3140 ;
  assign n6879 = ~n3141 & ~n6878 ;
  assign n6880 = n3132 & n6879 ;
  assign n6881 = ~n6876 & ~n6880 ;
  assign n6882 = ~n6877 & n6881 ;
  assign n6883 = n929 & ~n6882 ;
  assign n6884 = ~n6875 & ~n6883 ;
  assign n6885 = \EAX_reg[1]/NET0131  & ~n3181 ;
  assign n6888 = ~\EAX_reg[0]/NET0131  & n3132 ;
  assign n6889 = n3430 & ~n6888 ;
  assign n6890 = \EAX_reg[1]/NET0131  & ~n6889 ;
  assign n6891 = ~n1232 & n2937 ;
  assign n6886 = \Datai[1]_pad  & n846 ;
  assign n6887 = ~n841 & n6886 ;
  assign n6892 = \EAX_reg[0]/NET0131  & ~\EAX_reg[1]/NET0131  ;
  assign n6893 = n3132 & n6892 ;
  assign n6894 = ~n6887 & ~n6893 ;
  assign n6895 = ~n6891 & n6894 ;
  assign n6896 = ~n6890 & n6895 ;
  assign n6897 = n929 & ~n6896 ;
  assign n6898 = ~n6885 & ~n6897 ;
  assign n6900 = \MemoryFetch_reg/NET0131  & ~n5669 ;
  assign n6901 = n3661 & ~n6900 ;
  assign n6902 = n929 & ~n6901 ;
  assign n6899 = \MemoryFetch_reg/NET0131  & ~n3654 ;
  assign n6903 = n3652 & ~n6899 ;
  assign n6904 = ~n6902 & n6903 ;
  assign n6906 = \ReadRequest_reg/NET0131  & ~n837 ;
  assign n6907 = ~n842 & ~n6906 ;
  assign n6908 = n929 & ~n6907 ;
  assign n6905 = \ReadRequest_reg/NET0131  & ~n3654 ;
  assign n6909 = n3652 & ~n6905 ;
  assign n6910 = ~n6908 & n6909 ;
  assign n6911 = \rEIP_reg[0]/NET0131  & ~n5684 ;
  assign n6915 = ~\EBX_reg[0]/NET0131  & ~n5676 ;
  assign n6916 = ~\rEIP_reg[0]/NET0131  & n5676 ;
  assign n6917 = ~n6915 & ~n6916 ;
  assign n6918 = ~n6682 & n6917 ;
  assign n6912 = ~\InstQueueRd_Addr_reg[0]/NET0131  & n778 ;
  assign n6913 = \EBX_reg[0]/NET0131  & n828 ;
  assign n6914 = n783 & n6913 ;
  assign n6919 = ~n6912 & ~n6914 ;
  assign n6920 = ~n6918 & n6919 ;
  assign n6921 = ~n834 & ~n6920 ;
  assign n6922 = ~n6911 & ~n6921 ;
  assign n6923 = n929 & ~n6922 ;
  assign n6924 = ~n934 & ~n953 ;
  assign n6925 = \PhyAddrPointer_reg[0]/NET0131  & ~n6924 ;
  assign n6926 = ~n969 & n5667 ;
  assign n6927 = \rEIP_reg[0]/NET0131  & ~n6926 ;
  assign n6928 = ~n6925 & ~n6927 ;
  assign n6929 = ~n6923 & n6928 ;
  assign n6931 = n3438 & n3686 ;
  assign n6932 = ~\EAX_reg[30]/NET0131  & ~n6931 ;
  assign n6933 = \EAX_reg[30]/NET0131  & n6931 ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6935 = ~n828 & ~n6934 ;
  assign n6936 = n923 & ~n6935 ;
  assign n6937 = n3827 & ~n6936 ;
  assign n6938 = \Datao[30]_pad  & ~n6937 ;
  assign n6939 = n783 & n6934 ;
  assign n6940 = n856 & n6939 ;
  assign n6941 = ~n6938 & ~n6940 ;
  assign n6942 = n929 & ~n6941 ;
  assign n6930 = \uWord_reg[14]/NET0131  & n3809 ;
  assign n6943 = \Datao[30]_pad  & ~n3821 ;
  assign n6944 = ~n6930 & ~n6943 ;
  assign n6945 = ~n6942 & n6944 ;
  assign n6946 = \EAX_reg[28]/NET0131  & ~n3181 ;
  assign n6957 = ~\EAX_reg[28]/NET0131  & ~n3437 ;
  assign n6958 = n3132 & ~n3787 ;
  assign n6959 = ~n6957 & n6958 ;
  assign n6951 = \EAX_reg[28]/NET0131  & n3135 ;
  assign n6952 = ~n3129 & n3361 ;
  assign n6953 = ~n3362 & ~n6952 ;
  assign n6954 = n2937 & n6953 ;
  assign n6947 = \EAX_reg[28]/NET0131  & ~n846 ;
  assign n6948 = \Datai[28]_pad  & n846 ;
  assign n6949 = ~n6947 & ~n6948 ;
  assign n6950 = n840 & ~n6949 ;
  assign n6955 = ~n3657 & ~n6947 ;
  assign n6956 = n782 & ~n6955 ;
  assign n6960 = ~n6950 & ~n6956 ;
  assign n6961 = ~n6954 & n6960 ;
  assign n6962 = ~n6951 & n6961 ;
  assign n6963 = ~n6959 & n6962 ;
  assign n6964 = n929 & ~n6963 ;
  assign n6965 = ~n6946 & ~n6964 ;
  assign n6966 = \uWord_reg[14]/NET0131  & ~n3655 ;
  assign n6969 = ~n834 & n6939 ;
  assign n6967 = \uWord_reg[14]/NET0131  & ~n3662 ;
  assign n6968 = n846 & n3432 ;
  assign n6970 = ~n6967 & ~n6968 ;
  assign n6971 = ~n6969 & n6970 ;
  assign n6972 = n929 & ~n6971 ;
  assign n6973 = ~n6966 & ~n6972 ;
  assign n6974 = \EAX_reg[0]/NET0131  & ~n4671 ;
  assign n6976 = \Datai[0]_pad  & n843 ;
  assign n6975 = ~n1267 & n2937 ;
  assign n6977 = ~n6888 & ~n6975 ;
  assign n6978 = ~n6976 & n6977 ;
  assign n6979 = n929 & ~n6978 ;
  assign n6980 = ~n6974 & ~n6979 ;
  assign n6983 = ~\EBX_reg[28]/NET0131  & ~n3494 ;
  assign n6984 = n797 & ~n3696 ;
  assign n6985 = ~n6983 & n6984 ;
  assign n6981 = n3463 & n6953 ;
  assign n6982 = \EBX_reg[28]/NET0131  & n3465 ;
  assign n6986 = ~n6981 & ~n6982 ;
  assign n6987 = ~n6985 & n6986 ;
  assign n6988 = n929 & ~n6987 ;
  assign n6989 = \EBX_reg[28]/NET0131  & ~n3181 ;
  assign n6990 = ~n6988 & ~n6989 ;
  assign n7023 = ~\EAX_reg[16]/NET0131  & ~n3150 ;
  assign n7024 = n3132 & ~n3151 ;
  assign n7025 = ~n7023 & n7024 ;
  assign n7026 = \EAX_reg[16]/NET0131  & n3135 ;
  assign n7028 = \EAX_reg[16]/NET0131  & ~n846 ;
  assign n7031 = \Datai[16]_pad  & n846 ;
  assign n7032 = ~n7028 & ~n7031 ;
  assign n7033 = n840 & ~n7032 ;
  assign n6995 = \InstQueue_reg[0][0]/NET0131  & n465 ;
  assign n6996 = \InstQueue_reg[4][0]/NET0131  & n488 ;
  assign n7009 = ~n6995 & ~n6996 ;
  assign n6997 = \InstQueue_reg[8][0]/NET0131  & n490 ;
  assign n6998 = \InstQueue_reg[14][0]/NET0131  & n492 ;
  assign n7010 = ~n6997 & ~n6998 ;
  assign n7017 = n7009 & n7010 ;
  assign n6991 = \InstQueue_reg[1][0]/NET0131  & n470 ;
  assign n6992 = \InstQueue_reg[9][0]/NET0131  & n482 ;
  assign n7007 = ~n6991 & ~n6992 ;
  assign n6993 = \InstQueue_reg[2][0]/NET0131  & n522 ;
  assign n6994 = \InstQueue_reg[6][0]/NET0131  & n476 ;
  assign n7008 = ~n6993 & ~n6994 ;
  assign n7018 = n7007 & n7008 ;
  assign n7019 = n7017 & n7018 ;
  assign n7003 = \InstQueue_reg[15][0]/NET0131  & n468 ;
  assign n7004 = \InstQueue_reg[5][0]/NET0131  & n458 ;
  assign n7013 = ~n7003 & ~n7004 ;
  assign n7005 = \InstQueue_reg[13][0]/NET0131  & n461 ;
  assign n7006 = \InstQueue_reg[12][0]/NET0131  & n484 ;
  assign n7014 = ~n7005 & ~n7006 ;
  assign n7015 = n7013 & n7014 ;
  assign n6999 = \InstQueue_reg[7][0]/NET0131  & n472 ;
  assign n7000 = \InstQueue_reg[3][0]/NET0131  & n474 ;
  assign n7011 = ~n6999 & ~n7000 ;
  assign n7001 = \InstQueue_reg[11][0]/NET0131  & n486 ;
  assign n7002 = \InstQueue_reg[10][0]/NET0131  & n454 ;
  assign n7012 = ~n7001 & ~n7002 ;
  assign n7016 = n7011 & n7012 ;
  assign n7020 = n7015 & n7016 ;
  assign n7021 = n7019 & n7020 ;
  assign n7022 = n2937 & ~n7021 ;
  assign n7027 = \Datai[0]_pad  & n846 ;
  assign n7029 = ~n7027 & ~n7028 ;
  assign n7030 = n782 & ~n7029 ;
  assign n7034 = ~n7022 & ~n7030 ;
  assign n7035 = ~n7033 & n7034 ;
  assign n7036 = ~n7026 & n7035 ;
  assign n7037 = ~n7025 & n7036 ;
  assign n7038 = n929 & ~n7037 ;
  assign n7039 = \EAX_reg[16]/NET0131  & ~n3181 ;
  assign n7040 = ~n7038 & ~n7039 ;
  assign n7041 = \EAX_reg[17]/NET0131  & ~n3181 ;
  assign n7074 = ~\EAX_reg[17]/NET0131  & ~n3151 ;
  assign n7075 = n3132 & ~n3152 ;
  assign n7076 = ~n7074 & n7075 ;
  assign n7077 = \EAX_reg[17]/NET0131  & n3135 ;
  assign n7078 = \EAX_reg[17]/NET0131  & ~n846 ;
  assign n7081 = \Datai[17]_pad  & n846 ;
  assign n7082 = ~n7078 & ~n7081 ;
  assign n7083 = n840 & ~n7082 ;
  assign n7046 = \InstQueue_reg[3][1]/NET0131  & n474 ;
  assign n7047 = \InstQueue_reg[5][1]/NET0131  & n458 ;
  assign n7060 = ~n7046 & ~n7047 ;
  assign n7048 = \InstQueue_reg[15][1]/NET0131  & n468 ;
  assign n7049 = \InstQueue_reg[7][1]/NET0131  & n472 ;
  assign n7061 = ~n7048 & ~n7049 ;
  assign n7068 = n7060 & n7061 ;
  assign n7042 = \InstQueue_reg[1][1]/NET0131  & n470 ;
  assign n7043 = \InstQueue_reg[9][1]/NET0131  & n482 ;
  assign n7058 = ~n7042 & ~n7043 ;
  assign n7044 = \InstQueue_reg[13][1]/NET0131  & n461 ;
  assign n7045 = \InstQueue_reg[6][1]/NET0131  & n476 ;
  assign n7059 = ~n7044 & ~n7045 ;
  assign n7069 = n7058 & n7059 ;
  assign n7070 = n7068 & n7069 ;
  assign n7054 = \InstQueue_reg[2][1]/NET0131  & n522 ;
  assign n7055 = \InstQueue_reg[4][1]/NET0131  & n488 ;
  assign n7064 = ~n7054 & ~n7055 ;
  assign n7056 = \InstQueue_reg[8][1]/NET0131  & n490 ;
  assign n7057 = \InstQueue_reg[12][1]/NET0131  & n484 ;
  assign n7065 = ~n7056 & ~n7057 ;
  assign n7066 = n7064 & n7065 ;
  assign n7050 = \InstQueue_reg[10][1]/NET0131  & n454 ;
  assign n7051 = \InstQueue_reg[0][1]/NET0131  & n465 ;
  assign n7062 = ~n7050 & ~n7051 ;
  assign n7052 = \InstQueue_reg[11][1]/NET0131  & n486 ;
  assign n7053 = \InstQueue_reg[14][1]/NET0131  & n492 ;
  assign n7063 = ~n7052 & ~n7053 ;
  assign n7067 = n7062 & n7063 ;
  assign n7071 = n7066 & n7067 ;
  assign n7072 = n7070 & n7071 ;
  assign n7073 = n2937 & ~n7072 ;
  assign n7079 = ~n6886 & ~n7078 ;
  assign n7080 = n782 & ~n7079 ;
  assign n7084 = ~n7073 & ~n7080 ;
  assign n7085 = ~n7083 & n7084 ;
  assign n7086 = ~n7077 & n7085 ;
  assign n7087 = ~n7076 & n7086 ;
  assign n7088 = n929 & ~n7087 ;
  assign n7089 = ~n7041 & ~n7088 ;
  assign n7090 = \EAX_reg[18]/NET0131  & ~n3181 ;
  assign n7123 = ~\EAX_reg[18]/NET0131  & ~n3152 ;
  assign n7124 = n3132 & ~n3153 ;
  assign n7125 = ~n7123 & n7124 ;
  assign n7126 = \EAX_reg[18]/NET0131  & n3135 ;
  assign n7127 = \EAX_reg[18]/NET0131  & ~n846 ;
  assign n7131 = ~n6816 & ~n7127 ;
  assign n7132 = n782 & ~n7131 ;
  assign n7095 = \InstQueue_reg[5][2]/NET0131  & n458 ;
  assign n7096 = \InstQueue_reg[0][2]/NET0131  & n465 ;
  assign n7109 = ~n7095 & ~n7096 ;
  assign n7097 = \InstQueue_reg[12][2]/NET0131  & n484 ;
  assign n7098 = \InstQueue_reg[7][2]/NET0131  & n472 ;
  assign n7110 = ~n7097 & ~n7098 ;
  assign n7117 = n7109 & n7110 ;
  assign n7091 = \InstQueue_reg[11][2]/NET0131  & n486 ;
  assign n7092 = \InstQueue_reg[2][2]/NET0131  & n522 ;
  assign n7107 = ~n7091 & ~n7092 ;
  assign n7093 = \InstQueue_reg[1][2]/NET0131  & n470 ;
  assign n7094 = \InstQueue_reg[8][2]/NET0131  & n490 ;
  assign n7108 = ~n7093 & ~n7094 ;
  assign n7118 = n7107 & n7108 ;
  assign n7119 = n7117 & n7118 ;
  assign n7103 = \InstQueue_reg[9][2]/NET0131  & n482 ;
  assign n7104 = \InstQueue_reg[10][2]/NET0131  & n454 ;
  assign n7113 = ~n7103 & ~n7104 ;
  assign n7105 = \InstQueue_reg[14][2]/NET0131  & n492 ;
  assign n7106 = \InstQueue_reg[15][2]/NET0131  & n468 ;
  assign n7114 = ~n7105 & ~n7106 ;
  assign n7115 = n7113 & n7114 ;
  assign n7099 = \InstQueue_reg[13][2]/NET0131  & n461 ;
  assign n7100 = \InstQueue_reg[6][2]/NET0131  & n476 ;
  assign n7111 = ~n7099 & ~n7100 ;
  assign n7101 = \InstQueue_reg[4][2]/NET0131  & n488 ;
  assign n7102 = \InstQueue_reg[3][2]/NET0131  & n474 ;
  assign n7112 = ~n7101 & ~n7102 ;
  assign n7116 = n7111 & n7112 ;
  assign n7120 = n7115 & n7116 ;
  assign n7121 = n7119 & n7120 ;
  assign n7122 = n2937 & ~n7121 ;
  assign n7128 = \Datai[18]_pad  & n846 ;
  assign n7129 = ~n7127 & ~n7128 ;
  assign n7130 = n840 & ~n7129 ;
  assign n7133 = ~n7122 & ~n7130 ;
  assign n7134 = ~n7132 & n7133 ;
  assign n7135 = ~n7126 & n7134 ;
  assign n7136 = ~n7125 & n7135 ;
  assign n7137 = n929 & ~n7136 ;
  assign n7138 = ~n7090 & ~n7137 ;
  assign n7172 = \EAX_reg[19]/NET0131  & n3153 ;
  assign n7171 = ~\EAX_reg[19]/NET0131  & ~n3153 ;
  assign n7173 = n3132 & ~n7171 ;
  assign n7174 = ~n7172 & n7173 ;
  assign n7175 = \EAX_reg[19]/NET0131  & n3135 ;
  assign n7176 = \EAX_reg[19]/NET0131  & ~n846 ;
  assign n7180 = ~n6826 & ~n7176 ;
  assign n7181 = n782 & ~n7180 ;
  assign n7143 = \InstQueue_reg[3][3]/NET0131  & n474 ;
  assign n7144 = \InstQueue_reg[4][3]/NET0131  & n488 ;
  assign n7157 = ~n7143 & ~n7144 ;
  assign n7145 = \InstQueue_reg[13][3]/NET0131  & n461 ;
  assign n7146 = \InstQueue_reg[14][3]/NET0131  & n492 ;
  assign n7158 = ~n7145 & ~n7146 ;
  assign n7165 = n7157 & n7158 ;
  assign n7139 = \InstQueue_reg[1][3]/NET0131  & n470 ;
  assign n7140 = \InstQueue_reg[12][3]/NET0131  & n484 ;
  assign n7155 = ~n7139 & ~n7140 ;
  assign n7141 = \InstQueue_reg[8][3]/NET0131  & n490 ;
  assign n7142 = \InstQueue_reg[6][3]/NET0131  & n476 ;
  assign n7156 = ~n7141 & ~n7142 ;
  assign n7166 = n7155 & n7156 ;
  assign n7167 = n7165 & n7166 ;
  assign n7151 = \InstQueue_reg[2][3]/NET0131  & n522 ;
  assign n7152 = \InstQueue_reg[5][3]/NET0131  & n458 ;
  assign n7161 = ~n7151 & ~n7152 ;
  assign n7153 = \InstQueue_reg[0][3]/NET0131  & n465 ;
  assign n7154 = \InstQueue_reg[9][3]/NET0131  & n482 ;
  assign n7162 = ~n7153 & ~n7154 ;
  assign n7163 = n7161 & n7162 ;
  assign n7147 = \InstQueue_reg[15][3]/NET0131  & n468 ;
  assign n7148 = \InstQueue_reg[7][3]/NET0131  & n472 ;
  assign n7159 = ~n7147 & ~n7148 ;
  assign n7149 = \InstQueue_reg[11][3]/NET0131  & n486 ;
  assign n7150 = \InstQueue_reg[10][3]/NET0131  & n454 ;
  assign n7160 = ~n7149 & ~n7150 ;
  assign n7164 = n7159 & n7160 ;
  assign n7168 = n7163 & n7164 ;
  assign n7169 = n7167 & n7168 ;
  assign n7170 = n2937 & ~n7169 ;
  assign n7177 = \Datai[19]_pad  & n846 ;
  assign n7178 = ~n7176 & ~n7177 ;
  assign n7179 = n840 & ~n7178 ;
  assign n7182 = ~n7170 & ~n7179 ;
  assign n7183 = ~n7181 & n7182 ;
  assign n7184 = ~n7175 & n7183 ;
  assign n7185 = ~n7174 & n7184 ;
  assign n7186 = n929 & ~n7185 ;
  assign n7187 = \EAX_reg[19]/NET0131  & ~n3181 ;
  assign n7188 = ~n7186 & ~n7187 ;
  assign n7189 = ~n916 & n929 ;
  assign n7190 = \More_reg/NET0131  & ~n3181 ;
  assign n7191 = ~n7189 & ~n7190 ;
  assign n7224 = ~\EAX_reg[20]/NET0131  & ~n7172 ;
  assign n7225 = \EAX_reg[20]/NET0131  & n7172 ;
  assign n7226 = n3132 & ~n7225 ;
  assign n7227 = ~n7224 & n7226 ;
  assign n7228 = \EAX_reg[20]/NET0131  & n3135 ;
  assign n7229 = \EAX_reg[20]/NET0131  & ~n846 ;
  assign n7233 = ~n4298 & ~n7229 ;
  assign n7234 = n782 & ~n7233 ;
  assign n7196 = \InstQueue_reg[5][4]/NET0131  & n458 ;
  assign n7197 = \InstQueue_reg[7][4]/NET0131  & n472 ;
  assign n7210 = ~n7196 & ~n7197 ;
  assign n7198 = \InstQueue_reg[9][4]/NET0131  & n482 ;
  assign n7199 = \InstQueue_reg[2][4]/NET0131  & n522 ;
  assign n7211 = ~n7198 & ~n7199 ;
  assign n7218 = n7210 & n7211 ;
  assign n7192 = \InstQueue_reg[10][4]/NET0131  & n454 ;
  assign n7193 = \InstQueue_reg[8][4]/NET0131  & n490 ;
  assign n7208 = ~n7192 & ~n7193 ;
  assign n7194 = \InstQueue_reg[6][4]/NET0131  & n476 ;
  assign n7195 = \InstQueue_reg[12][4]/NET0131  & n484 ;
  assign n7209 = ~n7194 & ~n7195 ;
  assign n7219 = n7208 & n7209 ;
  assign n7220 = n7218 & n7219 ;
  assign n7204 = \InstQueue_reg[1][4]/NET0131  & n470 ;
  assign n7205 = \InstQueue_reg[15][4]/NET0131  & n468 ;
  assign n7214 = ~n7204 & ~n7205 ;
  assign n7206 = \InstQueue_reg[11][4]/NET0131  & n486 ;
  assign n7207 = \InstQueue_reg[0][4]/NET0131  & n465 ;
  assign n7215 = ~n7206 & ~n7207 ;
  assign n7216 = n7214 & n7215 ;
  assign n7200 = \InstQueue_reg[3][4]/NET0131  & n474 ;
  assign n7201 = \InstQueue_reg[14][4]/NET0131  & n492 ;
  assign n7212 = ~n7200 & ~n7201 ;
  assign n7202 = \InstQueue_reg[4][4]/NET0131  & n488 ;
  assign n7203 = \InstQueue_reg[13][4]/NET0131  & n461 ;
  assign n7213 = ~n7202 & ~n7203 ;
  assign n7217 = n7212 & n7213 ;
  assign n7221 = n7216 & n7217 ;
  assign n7222 = n7220 & n7221 ;
  assign n7223 = n2937 & ~n7222 ;
  assign n7230 = \Datai[20]_pad  & n846 ;
  assign n7231 = ~n7229 & ~n7230 ;
  assign n7232 = n840 & ~n7231 ;
  assign n7235 = ~n7223 & ~n7232 ;
  assign n7236 = ~n7234 & n7235 ;
  assign n7237 = ~n7228 & n7236 ;
  assign n7238 = ~n7227 & n7237 ;
  assign n7239 = n929 & ~n7238 ;
  assign n7240 = \EAX_reg[20]/NET0131  & ~n3181 ;
  assign n7241 = ~n7239 & ~n7240 ;
  assign n7242 = \EAX_reg[21]/NET0131  & ~n3181 ;
  assign n7275 = ~n3135 & ~n7226 ;
  assign n7276 = \EAX_reg[21]/NET0131  & ~n7275 ;
  assign n7283 = ~\EAX_reg[21]/NET0131  & n3132 ;
  assign n7284 = n7225 & n7283 ;
  assign n7277 = \EAX_reg[21]/NET0131  & ~n846 ;
  assign n7280 = \Datai[21]_pad  & n846 ;
  assign n7281 = ~n7277 & ~n7280 ;
  assign n7282 = n840 & ~n7281 ;
  assign n7247 = \InstQueue_reg[15][5]/NET0131  & n468 ;
  assign n7248 = \InstQueue_reg[4][5]/NET0131  & n488 ;
  assign n7261 = ~n7247 & ~n7248 ;
  assign n7249 = \InstQueue_reg[0][5]/NET0131  & n465 ;
  assign n7250 = \InstQueue_reg[11][5]/NET0131  & n486 ;
  assign n7262 = ~n7249 & ~n7250 ;
  assign n7269 = n7261 & n7262 ;
  assign n7243 = \InstQueue_reg[1][5]/NET0131  & n470 ;
  assign n7244 = \InstQueue_reg[9][5]/NET0131  & n482 ;
  assign n7259 = ~n7243 & ~n7244 ;
  assign n7245 = \InstQueue_reg[7][5]/NET0131  & n472 ;
  assign n7246 = \InstQueue_reg[6][5]/NET0131  & n476 ;
  assign n7260 = ~n7245 & ~n7246 ;
  assign n7270 = n7259 & n7260 ;
  assign n7271 = n7269 & n7270 ;
  assign n7255 = \InstQueue_reg[3][5]/NET0131  & n474 ;
  assign n7256 = \InstQueue_reg[5][5]/NET0131  & n458 ;
  assign n7265 = ~n7255 & ~n7256 ;
  assign n7257 = \InstQueue_reg[2][5]/NET0131  & n522 ;
  assign n7258 = \InstQueue_reg[12][5]/NET0131  & n484 ;
  assign n7266 = ~n7257 & ~n7258 ;
  assign n7267 = n7265 & n7266 ;
  assign n7251 = \InstQueue_reg[13][5]/NET0131  & n461 ;
  assign n7252 = \InstQueue_reg[8][5]/NET0131  & n490 ;
  assign n7263 = ~n7251 & ~n7252 ;
  assign n7253 = \InstQueue_reg[14][5]/NET0131  & n492 ;
  assign n7254 = \InstQueue_reg[10][5]/NET0131  & n454 ;
  assign n7264 = ~n7253 & ~n7254 ;
  assign n7268 = n7263 & n7264 ;
  assign n7272 = n7267 & n7268 ;
  assign n7273 = n7271 & n7272 ;
  assign n7274 = n2937 & ~n7273 ;
  assign n7278 = ~n6866 & ~n7277 ;
  assign n7279 = n782 & ~n7278 ;
  assign n7285 = ~n7274 & ~n7279 ;
  assign n7286 = ~n7282 & n7285 ;
  assign n7287 = ~n7284 & n7286 ;
  assign n7288 = ~n7276 & n7287 ;
  assign n7289 = n929 & ~n7288 ;
  assign n7290 = ~n7242 & ~n7289 ;
  assign n7291 = \EAX_reg[22]/NET0131  & ~n3181 ;
  assign n7324 = n3154 & n7172 ;
  assign n7325 = ~\EAX_reg[22]/NET0131  & ~n7324 ;
  assign n7326 = n3132 & ~n3157 ;
  assign n7327 = ~n7325 & n7326 ;
  assign n7328 = \EAX_reg[22]/NET0131  & ~n3430 ;
  assign n7296 = \InstQueue_reg[5][6]/NET0131  & n458 ;
  assign n7297 = \InstQueue_reg[3][6]/NET0131  & n474 ;
  assign n7310 = ~n7296 & ~n7297 ;
  assign n7298 = \InstQueue_reg[12][6]/NET0131  & n484 ;
  assign n7299 = \InstQueue_reg[2][6]/NET0131  & n522 ;
  assign n7311 = ~n7298 & ~n7299 ;
  assign n7318 = n7310 & n7311 ;
  assign n7292 = \InstQueue_reg[10][6]/NET0131  & n454 ;
  assign n7293 = \InstQueue_reg[8][6]/NET0131  & n490 ;
  assign n7308 = ~n7292 & ~n7293 ;
  assign n7294 = \InstQueue_reg[6][6]/NET0131  & n476 ;
  assign n7295 = \InstQueue_reg[9][6]/NET0131  & n482 ;
  assign n7309 = ~n7294 & ~n7295 ;
  assign n7319 = n7308 & n7309 ;
  assign n7320 = n7318 & n7319 ;
  assign n7304 = \InstQueue_reg[1][6]/NET0131  & n470 ;
  assign n7305 = \InstQueue_reg[15][6]/NET0131  & n468 ;
  assign n7314 = ~n7304 & ~n7305 ;
  assign n7306 = \InstQueue_reg[11][6]/NET0131  & n486 ;
  assign n7307 = \InstQueue_reg[0][6]/NET0131  & n465 ;
  assign n7315 = ~n7306 & ~n7307 ;
  assign n7316 = n7314 & n7315 ;
  assign n7300 = \InstQueue_reg[7][6]/NET0131  & n472 ;
  assign n7301 = \InstQueue_reg[14][6]/NET0131  & n492 ;
  assign n7312 = ~n7300 & ~n7301 ;
  assign n7302 = \InstQueue_reg[4][6]/NET0131  & n488 ;
  assign n7303 = \InstQueue_reg[13][6]/NET0131  & n461 ;
  assign n7313 = ~n7302 & ~n7303 ;
  assign n7317 = n7312 & n7313 ;
  assign n7321 = n7316 & n7317 ;
  assign n7322 = n7320 & n7321 ;
  assign n7323 = n2937 & ~n7322 ;
  assign n7329 = \Datai[6]_pad  & n782 ;
  assign n7330 = \Datai[22]_pad  & n840 ;
  assign n7331 = ~n7329 & ~n7330 ;
  assign n7332 = n846 & ~n7331 ;
  assign n7333 = ~n7323 & ~n7332 ;
  assign n7334 = ~n7328 & n7333 ;
  assign n7335 = ~n7327 & n7334 ;
  assign n7336 = n929 & ~n7335 ;
  assign n7337 = ~n7291 & ~n7336 ;
  assign n7338 = \EAX_reg[23]/NET0131  & ~n3181 ;
  assign n7343 = ~\EAX_reg[23]/NET0131  & ~n3157 ;
  assign n7342 = \EAX_reg[23]/NET0131  & n3157 ;
  assign n7344 = n3132 & ~n7342 ;
  assign n7345 = ~n7343 & n7344 ;
  assign n7346 = \EAX_reg[23]/NET0131  & n3135 ;
  assign n7347 = \EAX_reg[23]/NET0131  & ~n846 ;
  assign n7351 = ~n4674 & ~n7347 ;
  assign n7352 = n782 & ~n7351 ;
  assign n7339 = n2968 & n2999 ;
  assign n7340 = ~n3000 & ~n7339 ;
  assign n7341 = n2937 & n7340 ;
  assign n7348 = \Datai[23]_pad  & n846 ;
  assign n7349 = ~n7347 & ~n7348 ;
  assign n7350 = n840 & ~n7349 ;
  assign n7353 = ~n7341 & ~n7350 ;
  assign n7354 = ~n7352 & n7353 ;
  assign n7355 = ~n7346 & n7354 ;
  assign n7356 = ~n7345 & n7355 ;
  assign n7357 = n929 & ~n7356 ;
  assign n7358 = ~n7338 & ~n7357 ;
  assign n7362 = ~\EAX_reg[24]/NET0131  & ~n7342 ;
  assign n7363 = n3132 & ~n3159 ;
  assign n7364 = ~n7362 & n7363 ;
  assign n7365 = \EAX_reg[24]/NET0131  & n3135 ;
  assign n7366 = \EAX_reg[24]/NET0131  & ~n846 ;
  assign n7370 = \Datai[8]_pad  & n846 ;
  assign n7371 = ~n7366 & ~n7370 ;
  assign n7372 = n782 & ~n7371 ;
  assign n7359 = ~n3000 & n3031 ;
  assign n7360 = ~n3032 & ~n7359 ;
  assign n7361 = n2937 & n7360 ;
  assign n7367 = \Datai[24]_pad  & n846 ;
  assign n7368 = ~n7366 & ~n7367 ;
  assign n7369 = n840 & ~n7368 ;
  assign n7373 = ~n7361 & ~n7369 ;
  assign n7374 = ~n7372 & n7373 ;
  assign n7375 = ~n7365 & n7374 ;
  assign n7376 = ~n7364 & n7375 ;
  assign n7377 = n929 & ~n7376 ;
  assign n7378 = \EAX_reg[24]/NET0131  & ~n3181 ;
  assign n7379 = ~n7377 & ~n7378 ;
  assign n7381 = ~\EAX_reg[26]/NET0131  & ~n3685 ;
  assign n7382 = n783 & ~n4640 ;
  assign n7383 = ~n7381 & n7382 ;
  assign n7384 = n856 & n7383 ;
  assign n7385 = \Datao[26]_pad  & ~n857 ;
  assign n7386 = ~n7384 & ~n7385 ;
  assign n7387 = n929 & ~n7386 ;
  assign n7380 = \uWord_reg[10]/NET0131  & n3809 ;
  assign n7388 = \Datao[26]_pad  & ~n3821 ;
  assign n7389 = ~n7380 & ~n7388 ;
  assign n7390 = ~n7387 & n7389 ;
  assign n7391 = \uWord_reg[0]/NET0131  & ~n3655 ;
  assign n7393 = READY_n_pad & \uWord_reg[0]/NET0131  ;
  assign n7394 = ~n7027 & ~n7393 ;
  assign n7395 = n782 & ~n7394 ;
  assign n7392 = \uWord_reg[0]/NET0131  & n3661 ;
  assign n7396 = ~\EAX_reg[16]/NET0131  & ~n3679 ;
  assign n7397 = ~n3680 & ~n7396 ;
  assign n7398 = n923 & n7397 ;
  assign n7399 = ~n7392 & ~n7398 ;
  assign n7400 = ~n7395 & n7399 ;
  assign n7401 = n929 & ~n7400 ;
  assign n7402 = ~n7391 & ~n7401 ;
  assign n7403 = \uWord_reg[10]/NET0131  & ~n3839 ;
  assign n7404 = \Datai[10]_pad  & ~READY_n_pad ;
  assign n7405 = n782 & n7404 ;
  assign n7406 = ~n7383 & ~n7405 ;
  assign n7407 = n3844 & ~n7406 ;
  assign n7408 = ~n7403 & ~n7407 ;
  assign n7409 = \uWord_reg[13]/NET0131  & ~n3655 ;
  assign n7414 = ~\EAX_reg[29]/NET0131  & ~n3688 ;
  assign n7415 = n923 & ~n6931 ;
  assign n7416 = ~n7414 & n7415 ;
  assign n7410 = READY_n_pad & \uWord_reg[13]/NET0131  ;
  assign n7411 = ~n3784 & ~n7410 ;
  assign n7412 = n782 & ~n7411 ;
  assign n7413 = \uWord_reg[13]/NET0131  & n3661 ;
  assign n7417 = ~n7412 & ~n7413 ;
  assign n7418 = ~n7416 & n7417 ;
  assign n7419 = n929 & ~n7418 ;
  assign n7420 = ~n7409 & ~n7419 ;
  assign n7421 = \uWord_reg[1]/NET0131  & ~n3655 ;
  assign n7422 = READY_n_pad & \uWord_reg[1]/NET0131  ;
  assign n7423 = ~n6886 & ~n7422 ;
  assign n7424 = n782 & ~n7423 ;
  assign n7425 = \uWord_reg[1]/NET0131  & n3661 ;
  assign n7426 = ~\EAX_reg[17]/NET0131  & ~n3680 ;
  assign n7427 = ~n3681 & ~n7426 ;
  assign n7428 = n923 & n7427 ;
  assign n7429 = ~n7425 & ~n7428 ;
  assign n7430 = ~n7424 & n7429 ;
  assign n7431 = n929 & ~n7430 ;
  assign n7432 = ~n7421 & ~n7431 ;
  assign n7433 = \uWord_reg[2]/NET0131  & ~n3655 ;
  assign n7434 = READY_n_pad & \uWord_reg[2]/NET0131  ;
  assign n7435 = ~n6816 & ~n7434 ;
  assign n7436 = n782 & ~n7435 ;
  assign n7437 = \uWord_reg[2]/NET0131  & n3661 ;
  assign n7438 = ~\EAX_reg[18]/NET0131  & ~n3681 ;
  assign n7439 = ~n3682 & ~n7438 ;
  assign n7440 = n923 & n7439 ;
  assign n7441 = ~n7437 & ~n7440 ;
  assign n7442 = ~n7436 & n7441 ;
  assign n7443 = n929 & ~n7442 ;
  assign n7444 = ~n7433 & ~n7443 ;
  assign n7445 = \uWord_reg[5]/NET0131  & ~n3655 ;
  assign n7446 = READY_n_pad & \uWord_reg[5]/NET0131  ;
  assign n7447 = ~n6866 & ~n7446 ;
  assign n7448 = n782 & ~n7447 ;
  assign n7449 = \uWord_reg[5]/NET0131  & n3661 ;
  assign n7451 = ~\EAX_reg[21]/NET0131  & ~n4282 ;
  assign n7450 = n3155 & n3682 ;
  assign n7452 = n923 & ~n7450 ;
  assign n7453 = ~n7451 & n7452 ;
  assign n7454 = ~n7449 & ~n7453 ;
  assign n7455 = ~n7448 & n7454 ;
  assign n7456 = n929 & ~n7455 ;
  assign n7457 = ~n7445 & ~n7456 ;
  assign n7458 = \uWord_reg[6]/NET0131  & ~n3839 ;
  assign n7459 = ~\EAX_reg[22]/NET0131  & ~n7450 ;
  assign n7460 = ~n3683 & ~n7459 ;
  assign n7461 = n783 & n7460 ;
  assign n7462 = ~READY_n_pad & n7329 ;
  assign n7463 = ~n7461 & ~n7462 ;
  assign n7464 = n3844 & ~n7463 ;
  assign n7465 = ~n7458 & ~n7464 ;
  assign n7466 = \uWord_reg[9]/NET0131  & ~n3655 ;
  assign n7467 = \uWord_reg[9]/NET0131  & ~n3662 ;
  assign n7468 = ~\EAX_reg[25]/NET0131  & ~n3684 ;
  assign n7469 = ~n3685 & ~n7468 ;
  assign n7470 = n923 & n7469 ;
  assign n7471 = n782 & n4314 ;
  assign n7472 = ~n7470 & ~n7471 ;
  assign n7473 = ~n7467 & n7472 ;
  assign n7474 = n929 & ~n7473 ;
  assign n7475 = ~n7466 & ~n7474 ;
  assign n7477 = \EBX_reg[10]/NET0131  & n3465 ;
  assign n7476 = n3463 & ~n4801 ;
  assign n7478 = ~\EBX_reg[10]/NET0131  & ~n3476 ;
  assign n7479 = ~n3477 & ~n7478 ;
  assign n7480 = n797 & n7479 ;
  assign n7481 = ~n7476 & ~n7480 ;
  assign n7482 = ~n7477 & n7481 ;
  assign n7483 = n929 & ~n7482 ;
  assign n7484 = \EBX_reg[10]/NET0131  & ~n3181 ;
  assign n7485 = ~n7483 & ~n7484 ;
  assign n7487 = \EBX_reg[11]/NET0131  & n3465 ;
  assign n7486 = n3463 & ~n4841 ;
  assign n7488 = ~\EBX_reg[11]/NET0131  & ~n3477 ;
  assign n7489 = n797 & ~n3478 ;
  assign n7490 = ~n7488 & n7489 ;
  assign n7491 = ~n7486 & ~n7490 ;
  assign n7492 = ~n7487 & n7491 ;
  assign n7493 = n929 & ~n7492 ;
  assign n7494 = \EBX_reg[11]/NET0131  & ~n3181 ;
  assign n7495 = ~n7493 & ~n7494 ;
  assign n7498 = ~\EBX_reg[12]/NET0131  & ~n3478 ;
  assign n7499 = n797 & ~n3479 ;
  assign n7500 = ~n7498 & n7499 ;
  assign n7496 = \EBX_reg[12]/NET0131  & n3465 ;
  assign n7497 = n3463 & ~n4898 ;
  assign n7501 = ~n7496 & ~n7497 ;
  assign n7502 = ~n7500 & n7501 ;
  assign n7503 = n929 & ~n7502 ;
  assign n7504 = \EBX_reg[12]/NET0131  & ~n3181 ;
  assign n7505 = ~n7503 & ~n7504 ;
  assign n7508 = ~\EBX_reg[14]/NET0131  & ~n3480 ;
  assign n7509 = n797 & ~n3481 ;
  assign n7510 = ~n7508 & n7509 ;
  assign n7506 = n3463 & ~n4982 ;
  assign n7507 = \EBX_reg[14]/NET0131  & n3465 ;
  assign n7511 = ~n7506 & ~n7507 ;
  assign n7512 = ~n7510 & n7511 ;
  assign n7513 = n929 & ~n7512 ;
  assign n7514 = \EBX_reg[14]/NET0131  & ~n3181 ;
  assign n7515 = ~n7513 & ~n7514 ;
  assign n7518 = ~\EBX_reg[13]/NET0131  & ~n3479 ;
  assign n7519 = n797 & ~n3480 ;
  assign n7520 = ~n7518 & n7519 ;
  assign n7516 = n3463 & ~n4943 ;
  assign n7517 = \EBX_reg[13]/NET0131  & n3465 ;
  assign n7521 = ~n7516 & ~n7517 ;
  assign n7522 = ~n7520 & n7521 ;
  assign n7523 = n929 & ~n7522 ;
  assign n7524 = \EBX_reg[13]/NET0131  & ~n3181 ;
  assign n7525 = ~n7523 & ~n7524 ;
  assign n7528 = ~\EBX_reg[15]/NET0131  & ~n3481 ;
  assign n7529 = n797 & ~n3482 ;
  assign n7530 = ~n7528 & n7529 ;
  assign n7526 = \EBX_reg[15]/NET0131  & n3465 ;
  assign n7527 = n3463 & ~n5030 ;
  assign n7531 = ~n7526 & ~n7527 ;
  assign n7532 = ~n7530 & n7531 ;
  assign n7533 = n929 & ~n7532 ;
  assign n7534 = \EBX_reg[15]/NET0131  & ~n3181 ;
  assign n7535 = ~n7533 & ~n7534 ;
  assign n7538 = ~\EBX_reg[16]/NET0131  & ~n3482 ;
  assign n7539 = n797 & ~n3483 ;
  assign n7540 = ~n7538 & n7539 ;
  assign n7536 = \EBX_reg[16]/NET0131  & n3465 ;
  assign n7537 = n3463 & ~n7021 ;
  assign n7541 = ~n7536 & ~n7537 ;
  assign n7542 = ~n7540 & n7541 ;
  assign n7543 = n929 & ~n7542 ;
  assign n7544 = \EBX_reg[16]/NET0131  & ~n3181 ;
  assign n7545 = ~n7543 & ~n7544 ;
  assign n7548 = ~\EBX_reg[17]/NET0131  & ~n3483 ;
  assign n7549 = n797 & ~n3484 ;
  assign n7550 = ~n7548 & n7549 ;
  assign n7546 = \EBX_reg[17]/NET0131  & n3465 ;
  assign n7547 = n3463 & ~n7072 ;
  assign n7551 = ~n7546 & ~n7547 ;
  assign n7552 = ~n7550 & n7551 ;
  assign n7553 = n929 & ~n7552 ;
  assign n7554 = \EBX_reg[17]/NET0131  & ~n3181 ;
  assign n7555 = ~n7553 & ~n7554 ;
  assign n7558 = ~\EBX_reg[18]/NET0131  & ~n3484 ;
  assign n7559 = n797 & ~n3485 ;
  assign n7560 = ~n7558 & n7559 ;
  assign n7556 = \EBX_reg[18]/NET0131  & n3465 ;
  assign n7557 = n3463 & ~n7121 ;
  assign n7561 = ~n7556 & ~n7557 ;
  assign n7562 = ~n7560 & n7561 ;
  assign n7563 = n929 & ~n7562 ;
  assign n7564 = \EBX_reg[18]/NET0131  & ~n3181 ;
  assign n7565 = ~n7563 & ~n7564 ;
  assign n7568 = ~\EBX_reg[19]/NET0131  & ~n3485 ;
  assign n7569 = n797 & ~n3486 ;
  assign n7570 = ~n7568 & n7569 ;
  assign n7566 = n3463 & ~n7169 ;
  assign n7567 = \EBX_reg[19]/NET0131  & n3465 ;
  assign n7571 = ~n7566 & ~n7567 ;
  assign n7572 = ~n7570 & n7571 ;
  assign n7573 = n929 & ~n7572 ;
  assign n7574 = \EBX_reg[19]/NET0131  & ~n3181 ;
  assign n7575 = ~n7573 & ~n7574 ;
  assign n7579 = ~\EBX_reg[20]/NET0131  & ~n3486 ;
  assign n7578 = \EBX_reg[20]/NET0131  & n3486 ;
  assign n7580 = n797 & ~n7578 ;
  assign n7581 = ~n7579 & n7580 ;
  assign n7576 = \EBX_reg[20]/NET0131  & n3465 ;
  assign n7577 = n3463 & ~n7222 ;
  assign n7582 = ~n7576 & ~n7577 ;
  assign n7583 = ~n7581 & n7582 ;
  assign n7584 = n929 & ~n7583 ;
  assign n7585 = \EBX_reg[20]/NET0131  & ~n3181 ;
  assign n7586 = ~n7584 & ~n7585 ;
  assign n7590 = ~\EBX_reg[21]/NET0131  & ~n7578 ;
  assign n7589 = \EBX_reg[21]/NET0131  & n7578 ;
  assign n7591 = n797 & ~n7589 ;
  assign n7592 = ~n7590 & n7591 ;
  assign n7587 = n3463 & ~n7273 ;
  assign n7588 = \EBX_reg[21]/NET0131  & n3465 ;
  assign n7593 = ~n7587 & ~n7588 ;
  assign n7594 = ~n7592 & n7593 ;
  assign n7595 = n929 & ~n7594 ;
  assign n7596 = \EBX_reg[21]/NET0131  & ~n3181 ;
  assign n7597 = ~n7595 & ~n7596 ;
  assign n7601 = \EBX_reg[22]/NET0131  & n7589 ;
  assign n7600 = ~\EBX_reg[22]/NET0131  & ~n7589 ;
  assign n7602 = n797 & ~n7600 ;
  assign n7603 = ~n7601 & n7602 ;
  assign n7598 = n3463 & ~n7322 ;
  assign n7599 = \EBX_reg[22]/NET0131  & n3465 ;
  assign n7604 = ~n7598 & ~n7599 ;
  assign n7605 = ~n7603 & n7604 ;
  assign n7606 = n929 & ~n7605 ;
  assign n7607 = \EBX_reg[22]/NET0131  & ~n3181 ;
  assign n7608 = ~n7606 & ~n7607 ;
  assign n7611 = ~\EBX_reg[23]/NET0131  & ~n7601 ;
  assign n7612 = n797 & ~n3490 ;
  assign n7613 = ~n7611 & n7612 ;
  assign n7609 = \EBX_reg[23]/NET0131  & n3465 ;
  assign n7610 = n3463 & n7340 ;
  assign n7614 = ~n7609 & ~n7610 ;
  assign n7615 = ~n7613 & n7614 ;
  assign n7616 = n929 & ~n7615 ;
  assign n7617 = \EBX_reg[23]/NET0131  & ~n3181 ;
  assign n7618 = ~n7616 & ~n7617 ;
  assign n7620 = ~\EBX_reg[24]/NET0131  & ~n3490 ;
  assign n7621 = n4853 & ~n7620 ;
  assign n7619 = n3463 & n7360 ;
  assign n7622 = \EBX_reg[24]/NET0131  & n3465 ;
  assign n7623 = ~n7619 & ~n7622 ;
  assign n7624 = ~n7621 & n7623 ;
  assign n7625 = n929 & ~n7624 ;
  assign n7626 = \EBX_reg[24]/NET0131  & ~n3181 ;
  assign n7627 = ~n7625 & ~n7626 ;
  assign n7629 = \EBX_reg[8]/NET0131  & n3465 ;
  assign n7628 = n3463 & ~n4715 ;
  assign n7630 = ~\EBX_reg[8]/NET0131  & ~n3474 ;
  assign n7631 = ~n3475 & ~n7630 ;
  assign n7632 = n797 & n7631 ;
  assign n7633 = ~n7628 & ~n7632 ;
  assign n7634 = ~n7629 & n7633 ;
  assign n7635 = n929 & ~n7634 ;
  assign n7636 = \EBX_reg[8]/NET0131  & ~n3181 ;
  assign n7637 = ~n7635 & ~n7636 ;
  assign n7639 = \EBX_reg[9]/NET0131  & n3465 ;
  assign n7638 = n3463 & ~n4756 ;
  assign n7640 = ~\EBX_reg[9]/NET0131  & ~n3475 ;
  assign n7641 = ~n3476 & ~n7640 ;
  assign n7642 = n797 & n7641 ;
  assign n7643 = ~n7638 & ~n7642 ;
  assign n7644 = ~n7639 & n7643 ;
  assign n7645 = n929 & ~n7644 ;
  assign n7646 = \EBX_reg[9]/NET0131  & ~n3181 ;
  assign n7647 = ~n7645 & ~n7646 ;
  assign n7648 = ~n909 & n929 ;
  assign n7649 = \Flush_reg/NET0131  & ~n3181 ;
  assign n7650 = ~n7648 & ~n7649 ;
  assign n7656 = ~\Datai[26]_pad  & ~n3897 ;
  assign n7657 = ~n3898 & ~n7656 ;
  assign n7658 = n3871 & n7657 ;
  assign n7659 = ~\Datai[18]_pad  & ~n3906 ;
  assign n7660 = ~n3907 & ~n7659 ;
  assign n7661 = n3914 & n7660 ;
  assign n7662 = ~n7658 & ~n7661 ;
  assign n7663 = \DataWidth_reg[1]/NET0131  & ~n7662 ;
  assign n7651 = \Datai[2]_pad  & ~n3863 ;
  assign n7652 = \InstQueue_reg[0][2]/NET0131  & ~n3859 ;
  assign n7653 = ~n3862 & n7652 ;
  assign n7654 = ~n7651 & ~n7653 ;
  assign n7664 = ~n3919 & ~n7654 ;
  assign n7665 = ~n7663 & ~n7664 ;
  assign n7666 = n933 & ~n7665 ;
  assign n7667 = ~n572 & n3859 ;
  assign n7668 = ~n7652 & ~n7667 ;
  assign n7669 = n965 & ~n7668 ;
  assign n7655 = n1867 & ~n7654 ;
  assign n7670 = \InstQueue_reg[0][2]/NET0131  & ~n3929 ;
  assign n7671 = ~n7655 & ~n7670 ;
  assign n7672 = ~n7669 & n7671 ;
  assign n7673 = ~n7666 & n7672 ;
  assign n7679 = n3944 & n7657 ;
  assign n7680 = n3946 & n7660 ;
  assign n7681 = ~n7679 & ~n7680 ;
  assign n7682 = \DataWidth_reg[1]/NET0131  & ~n7681 ;
  assign n7674 = \Datai[2]_pad  & ~n3938 ;
  assign n7675 = \InstQueue_reg[10][2]/NET0131  & ~n3935 ;
  assign n7676 = ~n3937 & n7675 ;
  assign n7677 = ~n7674 & ~n7676 ;
  assign n7683 = ~n3951 & ~n7677 ;
  assign n7684 = ~n7682 & ~n7683 ;
  assign n7685 = n933 & ~n7684 ;
  assign n7686 = ~n572 & n3935 ;
  assign n7687 = ~n7675 & ~n7686 ;
  assign n7688 = n965 & ~n7687 ;
  assign n7678 = n1867 & ~n7677 ;
  assign n7689 = \InstQueue_reg[10][2]/NET0131  & ~n3929 ;
  assign n7690 = ~n7678 & ~n7689 ;
  assign n7691 = ~n7688 & n7690 ;
  assign n7692 = ~n7685 & n7691 ;
  assign n7698 = n3946 & n7657 ;
  assign n7699 = n3937 & n7660 ;
  assign n7700 = ~n7698 & ~n7699 ;
  assign n7701 = \DataWidth_reg[1]/NET0131  & ~n7700 ;
  assign n7693 = \Datai[2]_pad  & ~n3964 ;
  assign n7694 = \InstQueue_reg[11][2]/NET0131  & ~n3963 ;
  assign n7695 = ~n3935 & n7694 ;
  assign n7696 = ~n7693 & ~n7695 ;
  assign n7702 = ~n3975 & ~n7696 ;
  assign n7703 = ~n7701 & ~n7702 ;
  assign n7704 = n933 & ~n7703 ;
  assign n7705 = ~n572 & n3963 ;
  assign n7706 = ~n7694 & ~n7705 ;
  assign n7707 = n965 & ~n7706 ;
  assign n7697 = n1867 & ~n7696 ;
  assign n7708 = \InstQueue_reg[11][2]/NET0131  & ~n3929 ;
  assign n7709 = ~n7697 & ~n7708 ;
  assign n7710 = ~n7707 & n7709 ;
  assign n7711 = ~n7704 & n7710 ;
  assign n7717 = n3937 & n7657 ;
  assign n7718 = n3935 & n7660 ;
  assign n7719 = ~n7717 & ~n7718 ;
  assign n7720 = \DataWidth_reg[1]/NET0131  & ~n7719 ;
  assign n7712 = \Datai[2]_pad  & ~n3988 ;
  assign n7713 = \InstQueue_reg[12][2]/NET0131  & ~n3987 ;
  assign n7714 = ~n3963 & n7713 ;
  assign n7715 = ~n7712 & ~n7714 ;
  assign n7721 = ~n3998 & ~n7715 ;
  assign n7722 = ~n7720 & ~n7721 ;
  assign n7723 = n933 & ~n7722 ;
  assign n7724 = ~n572 & n3987 ;
  assign n7725 = ~n7713 & ~n7724 ;
  assign n7726 = n965 & ~n7725 ;
  assign n7716 = n1867 & ~n7715 ;
  assign n7727 = \InstQueue_reg[12][2]/NET0131  & ~n3929 ;
  assign n7728 = ~n7716 & ~n7727 ;
  assign n7729 = ~n7726 & n7728 ;
  assign n7730 = ~n7723 & n7729 ;
  assign n7736 = n3935 & n7657 ;
  assign n7737 = n3963 & n7660 ;
  assign n7738 = ~n7736 & ~n7737 ;
  assign n7739 = \DataWidth_reg[1]/NET0131  & ~n7738 ;
  assign n7731 = \Datai[2]_pad  & ~n4009 ;
  assign n7732 = \InstQueue_reg[13][2]/NET0131  & ~n3871 ;
  assign n7733 = ~n3987 & n7732 ;
  assign n7734 = ~n7731 & ~n7733 ;
  assign n7740 = ~n4019 & ~n7734 ;
  assign n7741 = ~n7739 & ~n7740 ;
  assign n7742 = n933 & ~n7741 ;
  assign n7743 = ~n572 & n3871 ;
  assign n7744 = ~n7732 & ~n7743 ;
  assign n7745 = n965 & ~n7744 ;
  assign n7735 = n1867 & ~n7734 ;
  assign n7746 = \InstQueue_reg[13][2]/NET0131  & ~n3929 ;
  assign n7747 = ~n7735 & ~n7746 ;
  assign n7748 = ~n7745 & n7747 ;
  assign n7749 = ~n7742 & n7748 ;
  assign n7755 = n3963 & n7657 ;
  assign n7756 = n3987 & n7660 ;
  assign n7757 = ~n7755 & ~n7756 ;
  assign n7758 = \DataWidth_reg[1]/NET0131  & ~n7757 ;
  assign n7750 = \Datai[2]_pad  & ~n3918 ;
  assign n7751 = \InstQueue_reg[14][2]/NET0131  & ~n3914 ;
  assign n7752 = ~n3871 & n7751 ;
  assign n7753 = ~n7750 & ~n7752 ;
  assign n7759 = ~n4039 & ~n7753 ;
  assign n7760 = ~n7758 & ~n7759 ;
  assign n7761 = n933 & ~n7760 ;
  assign n7762 = ~n572 & n3914 ;
  assign n7763 = ~n7751 & ~n7762 ;
  assign n7764 = n965 & ~n7763 ;
  assign n7754 = n1867 & ~n7753 ;
  assign n7765 = \InstQueue_reg[14][2]/NET0131  & ~n3929 ;
  assign n7766 = ~n7754 & ~n7765 ;
  assign n7767 = ~n7764 & n7766 ;
  assign n7768 = ~n7761 & n7767 ;
  assign n7774 = n3987 & n7657 ;
  assign n7775 = n3871 & n7660 ;
  assign n7776 = ~n7774 & ~n7775 ;
  assign n7777 = \DataWidth_reg[1]/NET0131  & ~n7776 ;
  assign n7769 = \Datai[2]_pad  & ~n4050 ;
  assign n7770 = \InstQueue_reg[15][2]/NET0131  & ~n3862 ;
  assign n7771 = ~n3914 & n7770 ;
  assign n7772 = ~n7769 & ~n7771 ;
  assign n7778 = ~n4060 & ~n7772 ;
  assign n7779 = ~n7777 & ~n7778 ;
  assign n7780 = n933 & ~n7779 ;
  assign n7781 = ~n572 & n3862 ;
  assign n7782 = ~n7770 & ~n7781 ;
  assign n7783 = n965 & ~n7782 ;
  assign n7773 = n1867 & ~n7772 ;
  assign n7784 = \InstQueue_reg[15][2]/NET0131  & ~n3929 ;
  assign n7785 = ~n7773 & ~n7784 ;
  assign n7786 = ~n7783 & n7785 ;
  assign n7787 = ~n7780 & n7786 ;
  assign n7793 = n3914 & n7657 ;
  assign n7794 = n3862 & n7660 ;
  assign n7795 = ~n7793 & ~n7794 ;
  assign n7796 = \DataWidth_reg[1]/NET0131  & ~n7795 ;
  assign n7788 = \Datai[2]_pad  & ~n4072 ;
  assign n7789 = \InstQueue_reg[1][2]/NET0131  & ~n4071 ;
  assign n7790 = ~n3859 & n7789 ;
  assign n7791 = ~n7788 & ~n7790 ;
  assign n7797 = ~n4082 & ~n7791 ;
  assign n7798 = ~n7796 & ~n7797 ;
  assign n7799 = n933 & ~n7798 ;
  assign n7800 = ~n572 & n4071 ;
  assign n7801 = ~n7789 & ~n7800 ;
  assign n7802 = n965 & ~n7801 ;
  assign n7792 = n1867 & ~n7791 ;
  assign n7803 = \InstQueue_reg[1][2]/NET0131  & ~n3929 ;
  assign n7804 = ~n7792 & ~n7803 ;
  assign n7805 = ~n7802 & n7804 ;
  assign n7806 = ~n7799 & n7805 ;
  assign n7812 = n3859 & n7660 ;
  assign n7813 = n3862 & n7657 ;
  assign n7814 = ~n7812 & ~n7813 ;
  assign n7815 = \DataWidth_reg[1]/NET0131  & ~n7814 ;
  assign n7807 = \Datai[2]_pad  & ~n4094 ;
  assign n7808 = \InstQueue_reg[2][2]/NET0131  & ~n4093 ;
  assign n7809 = ~n4071 & n7808 ;
  assign n7810 = ~n7807 & ~n7809 ;
  assign n7816 = ~n4104 & ~n7810 ;
  assign n7817 = ~n7815 & ~n7816 ;
  assign n7818 = n933 & ~n7817 ;
  assign n7819 = ~n572 & n4093 ;
  assign n7820 = ~n7808 & ~n7819 ;
  assign n7821 = n965 & ~n7820 ;
  assign n7811 = n1867 & ~n7810 ;
  assign n7822 = \InstQueue_reg[2][2]/NET0131  & ~n3929 ;
  assign n7823 = ~n7811 & ~n7822 ;
  assign n7824 = ~n7821 & n7823 ;
  assign n7825 = ~n7818 & n7824 ;
  assign n7831 = n3859 & n7657 ;
  assign n7832 = n4071 & n7660 ;
  assign n7833 = ~n7831 & ~n7832 ;
  assign n7834 = \DataWidth_reg[1]/NET0131  & ~n7833 ;
  assign n7826 = \Datai[2]_pad  & ~n4116 ;
  assign n7827 = \InstQueue_reg[3][2]/NET0131  & ~n4115 ;
  assign n7828 = ~n4093 & n7827 ;
  assign n7829 = ~n7826 & ~n7828 ;
  assign n7835 = ~n4126 & ~n7829 ;
  assign n7836 = ~n7834 & ~n7835 ;
  assign n7837 = n933 & ~n7836 ;
  assign n7838 = ~n572 & n4115 ;
  assign n7839 = ~n7827 & ~n7838 ;
  assign n7840 = n965 & ~n7839 ;
  assign n7830 = n1867 & ~n7829 ;
  assign n7841 = \InstQueue_reg[3][2]/NET0131  & ~n3929 ;
  assign n7842 = ~n7830 & ~n7841 ;
  assign n7843 = ~n7840 & n7842 ;
  assign n7844 = ~n7837 & n7843 ;
  assign n7850 = n4071 & n7657 ;
  assign n7851 = n4093 & n7660 ;
  assign n7852 = ~n7850 & ~n7851 ;
  assign n7853 = \DataWidth_reg[1]/NET0131  & ~n7852 ;
  assign n7845 = \Datai[2]_pad  & ~n4138 ;
  assign n7846 = \InstQueue_reg[4][2]/NET0131  & ~n4137 ;
  assign n7847 = ~n4115 & n7846 ;
  assign n7848 = ~n7845 & ~n7847 ;
  assign n7854 = ~n4148 & ~n7848 ;
  assign n7855 = ~n7853 & ~n7854 ;
  assign n7856 = n933 & ~n7855 ;
  assign n7857 = ~n572 & n4137 ;
  assign n7858 = ~n7846 & ~n7857 ;
  assign n7859 = n965 & ~n7858 ;
  assign n7849 = n1867 & ~n7848 ;
  assign n7860 = \InstQueue_reg[4][2]/NET0131  & ~n3929 ;
  assign n7861 = ~n7849 & ~n7860 ;
  assign n7862 = ~n7859 & n7861 ;
  assign n7863 = ~n7856 & n7862 ;
  assign n7869 = n4093 & n7657 ;
  assign n7870 = n4115 & n7660 ;
  assign n7871 = ~n7869 & ~n7870 ;
  assign n7872 = \DataWidth_reg[1]/NET0131  & ~n7871 ;
  assign n7864 = \Datai[2]_pad  & ~n4160 ;
  assign n7865 = \InstQueue_reg[5][2]/NET0131  & ~n4159 ;
  assign n7866 = ~n4137 & n7865 ;
  assign n7867 = ~n7864 & ~n7866 ;
  assign n7873 = ~n4170 & ~n7867 ;
  assign n7874 = ~n7872 & ~n7873 ;
  assign n7875 = n933 & ~n7874 ;
  assign n7876 = ~n572 & n4159 ;
  assign n7877 = ~n7865 & ~n7876 ;
  assign n7878 = n965 & ~n7877 ;
  assign n7868 = n1867 & ~n7867 ;
  assign n7879 = \InstQueue_reg[5][2]/NET0131  & ~n3929 ;
  assign n7880 = ~n7868 & ~n7879 ;
  assign n7881 = ~n7878 & n7880 ;
  assign n7882 = ~n7875 & n7881 ;
  assign n7888 = n4115 & n7657 ;
  assign n7889 = n4137 & n7660 ;
  assign n7890 = ~n7888 & ~n7889 ;
  assign n7891 = \DataWidth_reg[1]/NET0131  & ~n7890 ;
  assign n7883 = \Datai[2]_pad  & ~n4182 ;
  assign n7884 = \InstQueue_reg[6][2]/NET0131  & ~n4181 ;
  assign n7885 = ~n4159 & n7884 ;
  assign n7886 = ~n7883 & ~n7885 ;
  assign n7892 = ~n4192 & ~n7886 ;
  assign n7893 = ~n7891 & ~n7892 ;
  assign n7894 = n933 & ~n7893 ;
  assign n7895 = ~n572 & n4181 ;
  assign n7896 = ~n7884 & ~n7895 ;
  assign n7897 = n965 & ~n7896 ;
  assign n7887 = n1867 & ~n7886 ;
  assign n7898 = \InstQueue_reg[6][2]/NET0131  & ~n3929 ;
  assign n7899 = ~n7887 & ~n7898 ;
  assign n7900 = ~n7897 & n7899 ;
  assign n7901 = ~n7894 & n7900 ;
  assign n7907 = n4137 & n7657 ;
  assign n7908 = n4159 & n7660 ;
  assign n7909 = ~n7907 & ~n7908 ;
  assign n7910 = \DataWidth_reg[1]/NET0131  & ~n7909 ;
  assign n7902 = \Datai[2]_pad  & ~n4203 ;
  assign n7903 = \InstQueue_reg[7][2]/NET0131  & ~n3944 ;
  assign n7904 = ~n4181 & n7903 ;
  assign n7905 = ~n7902 & ~n7904 ;
  assign n7911 = ~n4213 & ~n7905 ;
  assign n7912 = ~n7910 & ~n7911 ;
  assign n7913 = n933 & ~n7912 ;
  assign n7914 = ~n572 & n3944 ;
  assign n7915 = ~n7903 & ~n7914 ;
  assign n7916 = n965 & ~n7915 ;
  assign n7906 = n1867 & ~n7905 ;
  assign n7917 = \InstQueue_reg[7][2]/NET0131  & ~n3929 ;
  assign n7918 = ~n7906 & ~n7917 ;
  assign n7919 = ~n7916 & n7918 ;
  assign n7920 = ~n7913 & n7919 ;
  assign n7926 = n4159 & n7657 ;
  assign n7927 = n4181 & n7660 ;
  assign n7928 = ~n7926 & ~n7927 ;
  assign n7929 = \DataWidth_reg[1]/NET0131  & ~n7928 ;
  assign n7921 = \Datai[2]_pad  & ~n3950 ;
  assign n7922 = \InstQueue_reg[8][2]/NET0131  & ~n3946 ;
  assign n7923 = ~n3944 & n7922 ;
  assign n7924 = ~n7921 & ~n7923 ;
  assign n7930 = ~n4233 & ~n7924 ;
  assign n7931 = ~n7929 & ~n7930 ;
  assign n7932 = n933 & ~n7931 ;
  assign n7933 = ~n572 & n3946 ;
  assign n7934 = ~n7922 & ~n7933 ;
  assign n7935 = n965 & ~n7934 ;
  assign n7925 = n1867 & ~n7924 ;
  assign n7936 = \InstQueue_reg[8][2]/NET0131  & ~n3929 ;
  assign n7937 = ~n7925 & ~n7936 ;
  assign n7938 = ~n7935 & n7937 ;
  assign n7939 = ~n7932 & n7938 ;
  assign n7945 = n4181 & n7657 ;
  assign n7946 = n3944 & n7660 ;
  assign n7947 = ~n7945 & ~n7946 ;
  assign n7948 = \DataWidth_reg[1]/NET0131  & ~n7947 ;
  assign n7940 = \Datai[2]_pad  & ~n3974 ;
  assign n7941 = \InstQueue_reg[9][2]/NET0131  & ~n3937 ;
  assign n7942 = ~n3946 & n7941 ;
  assign n7943 = ~n7940 & ~n7942 ;
  assign n7949 = ~n4253 & ~n7943 ;
  assign n7950 = ~n7948 & ~n7949 ;
  assign n7951 = n933 & ~n7950 ;
  assign n7952 = ~n572 & n3937 ;
  assign n7953 = ~n7941 & ~n7952 ;
  assign n7954 = n965 & ~n7953 ;
  assign n7944 = n1867 & ~n7943 ;
  assign n7955 = \InstQueue_reg[9][2]/NET0131  & ~n3929 ;
  assign n7956 = ~n7944 & ~n7955 ;
  assign n7957 = ~n7954 & n7956 ;
  assign n7958 = ~n7951 & n7957 ;
  assign n7960 = ~n828 & n7416 ;
  assign n7961 = \Datao[29]_pad  & ~n857 ;
  assign n7962 = ~n7960 & ~n7961 ;
  assign n7963 = n929 & ~n7962 ;
  assign n7959 = \uWord_reg[13]/NET0131  & n3809 ;
  assign n7964 = \Datao[29]_pad  & ~n3821 ;
  assign n7965 = ~n7959 & ~n7964 ;
  assign n7966 = ~n7963 & n7965 ;
  assign n7969 = \CodeFetch_reg/NET0131  & n929 ;
  assign n7970 = ~n5684 & n7969 ;
  assign n7967 = ~n955 & ~n3820 ;
  assign n7968 = \CodeFetch_reg/NET0131  & ~n7967 ;
  assign n7971 = ~n937 & ~n7968 ;
  assign n7972 = ~n7970 & n7971 ;
  assign n7974 = ~n828 & n7440 ;
  assign n7975 = \Datao[18]_pad  & ~n857 ;
  assign n7976 = ~n7974 & ~n7975 ;
  assign n7977 = n929 & ~n7976 ;
  assign n7973 = \uWord_reg[2]/NET0131  & n3809 ;
  assign n7978 = \Datao[18]_pad  & ~n3821 ;
  assign n7979 = ~n7973 & ~n7978 ;
  assign n7980 = ~n7977 & n7979 ;
  assign n7982 = ~n828 & ~n7460 ;
  assign n7983 = n923 & ~n7982 ;
  assign n7984 = n3827 & ~n7983 ;
  assign n7985 = \Datao[22]_pad  & ~n7984 ;
  assign n7986 = n856 & n7461 ;
  assign n7987 = ~n7985 & ~n7986 ;
  assign n7988 = n929 & ~n7987 ;
  assign n7981 = \uWord_reg[6]/NET0131  & n3809 ;
  assign n7989 = \Datao[22]_pad  & ~n3821 ;
  assign n7990 = ~n7981 & ~n7989 ;
  assign n7991 = ~n7988 & n7990 ;
  assign n7992 = n929 & n3465 ;
  assign n7993 = n3181 & ~n7992 ;
  assign n7994 = \EBX_reg[0]/NET0131  & ~n7993 ;
  assign n7995 = \InstQueue_reg[0][0]/NET0131  & n3463 ;
  assign n7996 = ~\EBX_reg[0]/NET0131  & n797 ;
  assign n7997 = ~n7995 & ~n7996 ;
  assign n7998 = n929 & ~n7997 ;
  assign n7999 = ~n7994 & ~n7998 ;
  assign n8004 = ~\InstQueue_reg[0][1]/NET0131  & n765 ;
  assign n8003 = ~\EBX_reg[1]/NET0131  & ~n765 ;
  assign n8005 = n735 & ~n8003 ;
  assign n8006 = ~n8004 & n8005 ;
  assign n8000 = n797 & n5674 ;
  assign n8001 = \EBX_reg[1]/NET0131  & ~n735 ;
  assign n8002 = ~n797 & n8001 ;
  assign n8007 = ~n8000 & ~n8002 ;
  assign n8008 = ~n8006 & n8007 ;
  assign n8009 = n929 & ~n8008 ;
  assign n8010 = \EBX_reg[1]/NET0131  & ~n3181 ;
  assign n8011 = ~n8009 & ~n8010 ;
  assign n8013 = \EBX_reg[2]/NET0131  & n3465 ;
  assign n8012 = \InstQueue_reg[0][2]/NET0131  & n3463 ;
  assign n8014 = ~\EBX_reg[2]/NET0131  & ~n3468 ;
  assign n8015 = ~n3469 & ~n8014 ;
  assign n8016 = n797 & n8015 ;
  assign n8017 = ~n8012 & ~n8016 ;
  assign n8018 = ~n8013 & n8017 ;
  assign n8019 = n929 & ~n8018 ;
  assign n8020 = \EBX_reg[2]/NET0131  & ~n3181 ;
  assign n8021 = ~n8019 & ~n8020 ;
  assign n8023 = \EBX_reg[3]/NET0131  & n3465 ;
  assign n8022 = \InstQueue_reg[0][3]/NET0131  & n3463 ;
  assign n8024 = ~\EBX_reg[3]/NET0131  & ~n3469 ;
  assign n8025 = ~n3470 & ~n8024 ;
  assign n8026 = n797 & n8025 ;
  assign n8027 = ~n8022 & ~n8026 ;
  assign n8028 = ~n8023 & n8027 ;
  assign n8029 = n929 & ~n8028 ;
  assign n8030 = \EBX_reg[3]/NET0131  & ~n3181 ;
  assign n8031 = ~n8029 & ~n8030 ;
  assign n8033 = \EBX_reg[4]/NET0131  & n3465 ;
  assign n8032 = \InstQueue_reg[0][4]/NET0131  & n3463 ;
  assign n8034 = ~\EBX_reg[4]/NET0131  & ~n3470 ;
  assign n8035 = ~n3471 & ~n8034 ;
  assign n8036 = n797 & n8035 ;
  assign n8037 = ~n8032 & ~n8036 ;
  assign n8038 = ~n8033 & n8037 ;
  assign n8039 = n929 & ~n8038 ;
  assign n8040 = \EBX_reg[4]/NET0131  & ~n3181 ;
  assign n8041 = ~n8039 & ~n8040 ;
  assign n8043 = \EBX_reg[5]/NET0131  & n3465 ;
  assign n8042 = \InstQueue_reg[0][5]/NET0131  & n3463 ;
  assign n8044 = ~\EBX_reg[5]/NET0131  & ~n3471 ;
  assign n8045 = ~n3472 & ~n8044 ;
  assign n8046 = n797 & n8045 ;
  assign n8047 = ~n8042 & ~n8046 ;
  assign n8048 = ~n8043 & n8047 ;
  assign n8049 = n929 & ~n8048 ;
  assign n8050 = \EBX_reg[5]/NET0131  & ~n3181 ;
  assign n8051 = ~n8049 & ~n8050 ;
  assign n8053 = \EBX_reg[6]/NET0131  & n3465 ;
  assign n8052 = \InstQueue_reg[0][6]/NET0131  & n3463 ;
  assign n8054 = ~\EBX_reg[6]/NET0131  & ~n3472 ;
  assign n8055 = ~n3473 & ~n8054 ;
  assign n8056 = n797 & n8055 ;
  assign n8057 = ~n8052 & ~n8056 ;
  assign n8058 = ~n8053 & n8057 ;
  assign n8059 = n929 & ~n8058 ;
  assign n8060 = \EBX_reg[6]/NET0131  & ~n3181 ;
  assign n8061 = ~n8059 & ~n8060 ;
  assign n8063 = \EBX_reg[7]/NET0131  & n3465 ;
  assign n8062 = \InstQueue_reg[0][7]/NET0131  & n3463 ;
  assign n8064 = ~\EBX_reg[7]/NET0131  & ~n3473 ;
  assign n8065 = ~n3474 & ~n8064 ;
  assign n8066 = n797 & n8065 ;
  assign n8067 = ~n8062 & ~n8066 ;
  assign n8068 = ~n8063 & n8067 ;
  assign n8069 = n929 & ~n8068 ;
  assign n8070 = \EBX_reg[7]/NET0131  & ~n3181 ;
  assign n8071 = ~n8069 & ~n8070 ;
  assign n8073 = READY_n_pad & \lWord_reg[0]/NET0131  ;
  assign n8074 = ~n7027 & ~n8073 ;
  assign n8075 = n782 & ~n8074 ;
  assign n8072 = \lWord_reg[0]/NET0131  & n3661 ;
  assign n8076 = \EAX_reg[0]/NET0131  & n923 ;
  assign n8077 = ~n8072 & ~n8076 ;
  assign n8078 = ~n8075 & n8077 ;
  assign n8079 = n929 & ~n8078 ;
  assign n8080 = \lWord_reg[0]/NET0131  & ~n3655 ;
  assign n8081 = ~n8079 & ~n8080 ;
  assign n8082 = \lWord_reg[10]/NET0131  & ~n3839 ;
  assign n8083 = \EAX_reg[10]/NET0131  & n923 ;
  assign n8084 = ~n834 & n7405 ;
  assign n8085 = ~n8083 & ~n8084 ;
  assign n8086 = n929 & ~n8085 ;
  assign n8087 = ~n8082 & ~n8086 ;
  assign n8089 = READY_n_pad & \lWord_reg[11]/NET0131  ;
  assign n8090 = ~n3166 & ~n8089 ;
  assign n8091 = n782 & ~n8090 ;
  assign n8088 = \lWord_reg[11]/NET0131  & n3661 ;
  assign n8092 = \EAX_reg[11]/NET0131  & n923 ;
  assign n8093 = ~n8088 & ~n8092 ;
  assign n8094 = ~n8091 & n8093 ;
  assign n8095 = n929 & ~n8094 ;
  assign n8096 = \lWord_reg[11]/NET0131  & ~n3655 ;
  assign n8097 = ~n8095 & ~n8096 ;
  assign n8098 = \lWord_reg[12]/NET0131  & ~n3839 ;
  assign n8099 = \EAX_reg[12]/NET0131  & n923 ;
  assign n8100 = ~n3658 & ~n8099 ;
  assign n8101 = n929 & ~n8100 ;
  assign n8102 = ~n8098 & ~n8101 ;
  assign n8104 = READY_n_pad & \lWord_reg[13]/NET0131  ;
  assign n8105 = ~n3784 & ~n8104 ;
  assign n8106 = n782 & ~n8105 ;
  assign n8103 = \lWord_reg[13]/NET0131  & n3661 ;
  assign n8107 = \EAX_reg[13]/NET0131  & n923 ;
  assign n8108 = ~n8103 & ~n8107 ;
  assign n8109 = ~n8106 & n8108 ;
  assign n8110 = n929 & ~n8109 ;
  assign n8111 = \lWord_reg[13]/NET0131  & ~n3655 ;
  assign n8112 = ~n8110 & ~n8111 ;
  assign n8113 = \lWord_reg[14]/NET0131  & ~n3839 ;
  assign n8114 = \EAX_reg[14]/NET0131  & n923 ;
  assign n8115 = ~n6968 & ~n8114 ;
  assign n8116 = n929 & ~n8115 ;
  assign n8117 = ~n8113 & ~n8116 ;
  assign n8119 = READY_n_pad & \lWord_reg[15]/NET0131  ;
  assign n8120 = ~n4996 & ~n8119 ;
  assign n8121 = n782 & ~n8120 ;
  assign n8118 = \lWord_reg[15]/NET0131  & n3661 ;
  assign n8122 = \EAX_reg[15]/NET0131  & n923 ;
  assign n8123 = ~n8118 & ~n8122 ;
  assign n8124 = ~n8121 & n8123 ;
  assign n8125 = n929 & ~n8124 ;
  assign n8126 = \lWord_reg[15]/NET0131  & ~n3655 ;
  assign n8127 = ~n8125 & ~n8126 ;
  assign n8129 = READY_n_pad & \lWord_reg[1]/NET0131  ;
  assign n8130 = ~n6886 & ~n8129 ;
  assign n8131 = n782 & ~n8130 ;
  assign n8128 = \lWord_reg[1]/NET0131  & n3661 ;
  assign n8132 = \EAX_reg[1]/NET0131  & n923 ;
  assign n8133 = ~n8128 & ~n8132 ;
  assign n8134 = ~n8131 & n8133 ;
  assign n8135 = n929 & ~n8134 ;
  assign n8136 = \lWord_reg[1]/NET0131  & ~n3655 ;
  assign n8137 = ~n8135 & ~n8136 ;
  assign n8139 = READY_n_pad & \lWord_reg[2]/NET0131  ;
  assign n8140 = ~n6816 & ~n8139 ;
  assign n8141 = n782 & ~n8140 ;
  assign n8138 = \lWord_reg[2]/NET0131  & n3661 ;
  assign n8142 = \EAX_reg[2]/NET0131  & n923 ;
  assign n8143 = ~n8138 & ~n8142 ;
  assign n8144 = ~n8141 & n8143 ;
  assign n8145 = n929 & ~n8144 ;
  assign n8146 = \lWord_reg[2]/NET0131  & ~n3655 ;
  assign n8147 = ~n8145 & ~n8146 ;
  assign n8149 = READY_n_pad & \lWord_reg[3]/NET0131  ;
  assign n8150 = ~n6826 & ~n8149 ;
  assign n8151 = n782 & ~n8150 ;
  assign n8148 = \lWord_reg[3]/NET0131  & n3661 ;
  assign n8152 = \EAX_reg[3]/NET0131  & n923 ;
  assign n8153 = ~n8148 & ~n8152 ;
  assign n8154 = ~n8151 & n8153 ;
  assign n8155 = n929 & ~n8154 ;
  assign n8156 = \lWord_reg[3]/NET0131  & ~n3655 ;
  assign n8157 = ~n8155 & ~n8156 ;
  assign n8159 = READY_n_pad & \lWord_reg[4]/NET0131  ;
  assign n8160 = ~n4298 & ~n8159 ;
  assign n8161 = n782 & ~n8160 ;
  assign n8158 = \lWord_reg[4]/NET0131  & n3661 ;
  assign n8162 = \EAX_reg[4]/NET0131  & n923 ;
  assign n8163 = ~n8158 & ~n8162 ;
  assign n8164 = ~n8161 & n8163 ;
  assign n8165 = n929 & ~n8164 ;
  assign n8166 = \lWord_reg[4]/NET0131  & ~n3655 ;
  assign n8167 = ~n8165 & ~n8166 ;
  assign n8169 = READY_n_pad & \lWord_reg[5]/NET0131  ;
  assign n8170 = ~n6866 & ~n8169 ;
  assign n8171 = n782 & ~n8170 ;
  assign n8168 = \lWord_reg[5]/NET0131  & n3661 ;
  assign n8172 = \EAX_reg[5]/NET0131  & n923 ;
  assign n8173 = ~n8168 & ~n8172 ;
  assign n8174 = ~n8171 & n8173 ;
  assign n8175 = n929 & ~n8174 ;
  assign n8176 = \lWord_reg[5]/NET0131  & ~n3655 ;
  assign n8177 = ~n8175 & ~n8176 ;
  assign n8179 = \Datai[6]_pad  & n846 ;
  assign n8180 = READY_n_pad & \lWord_reg[6]/NET0131  ;
  assign n8181 = ~n8179 & ~n8180 ;
  assign n8182 = n782 & ~n8181 ;
  assign n8178 = \lWord_reg[6]/NET0131  & n3661 ;
  assign n8183 = \EAX_reg[6]/NET0131  & n923 ;
  assign n8184 = ~n8178 & ~n8183 ;
  assign n8185 = ~n8182 & n8184 ;
  assign n8186 = n929 & ~n8185 ;
  assign n8187 = \lWord_reg[6]/NET0131  & ~n3655 ;
  assign n8188 = ~n8186 & ~n8187 ;
  assign n8190 = READY_n_pad & \lWord_reg[7]/NET0131  ;
  assign n8191 = ~n4674 & ~n8190 ;
  assign n8192 = n782 & ~n8191 ;
  assign n8189 = \lWord_reg[7]/NET0131  & n3661 ;
  assign n8193 = \EAX_reg[7]/NET0131  & n923 ;
  assign n8194 = ~n8189 & ~n8193 ;
  assign n8195 = ~n8192 & n8194 ;
  assign n8196 = n929 & ~n8195 ;
  assign n8197 = \lWord_reg[7]/NET0131  & ~n3655 ;
  assign n8198 = ~n8196 & ~n8197 ;
  assign n8199 = \lWord_reg[8]/NET0131  & ~n3839 ;
  assign n8200 = \EAX_reg[8]/NET0131  & n923 ;
  assign n8201 = ~n834 & n3842 ;
  assign n8202 = ~n8200 & ~n8201 ;
  assign n8203 = n929 & ~n8202 ;
  assign n8204 = ~n8199 & ~n8203 ;
  assign n8206 = READY_n_pad & \lWord_reg[9]/NET0131  ;
  assign n8207 = ~n4314 & ~n8206 ;
  assign n8208 = n782 & ~n8207 ;
  assign n8205 = \lWord_reg[9]/NET0131  & n3661 ;
  assign n8209 = \EAX_reg[9]/NET0131  & n923 ;
  assign n8210 = ~n8205 & ~n8209 ;
  assign n8211 = ~n8208 & n8210 ;
  assign n8212 = n929 & ~n8211 ;
  assign n8213 = \lWord_reg[9]/NET0131  & ~n3655 ;
  assign n8214 = ~n8212 & ~n8213 ;
  assign n8220 = ~\Datai[29]_pad  & ~n3900 ;
  assign n8221 = ~n4332 & ~n8220 ;
  assign n8222 = n3871 & n8221 ;
  assign n8223 = ~\Datai[21]_pad  & ~n3910 ;
  assign n8224 = ~n4336 & ~n8223 ;
  assign n8225 = n3914 & n8224 ;
  assign n8226 = ~n8222 & ~n8225 ;
  assign n8227 = \DataWidth_reg[1]/NET0131  & ~n8226 ;
  assign n8215 = \Datai[5]_pad  & ~n3863 ;
  assign n8216 = \InstQueue_reg[0][5]/NET0131  & ~n3859 ;
  assign n8217 = ~n3862 & n8216 ;
  assign n8218 = ~n8215 & ~n8217 ;
  assign n8228 = ~n3919 & ~n8218 ;
  assign n8229 = ~n8227 & ~n8228 ;
  assign n8230 = n933 & ~n8229 ;
  assign n8231 = ~n637 & n3859 ;
  assign n8232 = ~n8216 & ~n8231 ;
  assign n8233 = n965 & ~n8232 ;
  assign n8219 = n1867 & ~n8218 ;
  assign n8234 = \InstQueue_reg[0][5]/NET0131  & ~n3929 ;
  assign n8235 = ~n8219 & ~n8234 ;
  assign n8236 = ~n8233 & n8235 ;
  assign n8237 = ~n8230 & n8236 ;
  assign n8243 = n3944 & n8221 ;
  assign n8244 = n3946 & n8224 ;
  assign n8245 = ~n8243 & ~n8244 ;
  assign n8246 = \DataWidth_reg[1]/NET0131  & ~n8245 ;
  assign n8238 = \Datai[5]_pad  & ~n3938 ;
  assign n8239 = \InstQueue_reg[10][5]/NET0131  & ~n3935 ;
  assign n8240 = ~n3937 & n8239 ;
  assign n8241 = ~n8238 & ~n8240 ;
  assign n8247 = ~n3951 & ~n8241 ;
  assign n8248 = ~n8246 & ~n8247 ;
  assign n8249 = n933 & ~n8248 ;
  assign n8250 = ~n637 & n3935 ;
  assign n8251 = ~n8239 & ~n8250 ;
  assign n8252 = n965 & ~n8251 ;
  assign n8242 = n1867 & ~n8241 ;
  assign n8253 = \InstQueue_reg[10][5]/NET0131  & ~n3929 ;
  assign n8254 = ~n8242 & ~n8253 ;
  assign n8255 = ~n8252 & n8254 ;
  assign n8256 = ~n8249 & n8255 ;
  assign n8262 = n3946 & n8221 ;
  assign n8263 = n3937 & n8224 ;
  assign n8264 = ~n8262 & ~n8263 ;
  assign n8265 = \DataWidth_reg[1]/NET0131  & ~n8264 ;
  assign n8257 = \Datai[5]_pad  & ~n3964 ;
  assign n8258 = \InstQueue_reg[11][5]/NET0131  & ~n3963 ;
  assign n8259 = ~n3935 & n8258 ;
  assign n8260 = ~n8257 & ~n8259 ;
  assign n8266 = ~n3975 & ~n8260 ;
  assign n8267 = ~n8265 & ~n8266 ;
  assign n8268 = n933 & ~n8267 ;
  assign n8269 = ~n637 & n3963 ;
  assign n8270 = ~n8258 & ~n8269 ;
  assign n8271 = n965 & ~n8270 ;
  assign n8261 = n1867 & ~n8260 ;
  assign n8272 = \InstQueue_reg[11][5]/NET0131  & ~n3929 ;
  assign n8273 = ~n8261 & ~n8272 ;
  assign n8274 = ~n8271 & n8273 ;
  assign n8275 = ~n8268 & n8274 ;
  assign n8281 = n3937 & n8221 ;
  assign n8282 = n3935 & n8224 ;
  assign n8283 = ~n8281 & ~n8282 ;
  assign n8284 = \DataWidth_reg[1]/NET0131  & ~n8283 ;
  assign n8276 = \Datai[5]_pad  & ~n3988 ;
  assign n8277 = \InstQueue_reg[12][5]/NET0131  & ~n3987 ;
  assign n8278 = ~n3963 & n8277 ;
  assign n8279 = ~n8276 & ~n8278 ;
  assign n8285 = ~n3998 & ~n8279 ;
  assign n8286 = ~n8284 & ~n8285 ;
  assign n8287 = n933 & ~n8286 ;
  assign n8288 = ~n637 & n3987 ;
  assign n8289 = ~n8277 & ~n8288 ;
  assign n8290 = n965 & ~n8289 ;
  assign n8280 = n1867 & ~n8279 ;
  assign n8291 = \InstQueue_reg[12][5]/NET0131  & ~n3929 ;
  assign n8292 = ~n8280 & ~n8291 ;
  assign n8293 = ~n8290 & n8292 ;
  assign n8294 = ~n8287 & n8293 ;
  assign n8300 = n3935 & n8221 ;
  assign n8301 = n3963 & n8224 ;
  assign n8302 = ~n8300 & ~n8301 ;
  assign n8303 = \DataWidth_reg[1]/NET0131  & ~n8302 ;
  assign n8295 = \Datai[5]_pad  & ~n4009 ;
  assign n8296 = \InstQueue_reg[13][5]/NET0131  & ~n3871 ;
  assign n8297 = ~n3987 & n8296 ;
  assign n8298 = ~n8295 & ~n8297 ;
  assign n8304 = ~n4019 & ~n8298 ;
  assign n8305 = ~n8303 & ~n8304 ;
  assign n8306 = n933 & ~n8305 ;
  assign n8307 = ~n637 & n3871 ;
  assign n8308 = ~n8296 & ~n8307 ;
  assign n8309 = n965 & ~n8308 ;
  assign n8299 = n1867 & ~n8298 ;
  assign n8310 = \InstQueue_reg[13][5]/NET0131  & ~n3929 ;
  assign n8311 = ~n8299 & ~n8310 ;
  assign n8312 = ~n8309 & n8311 ;
  assign n8313 = ~n8306 & n8312 ;
  assign n8319 = n3963 & n8221 ;
  assign n8320 = n3987 & n8224 ;
  assign n8321 = ~n8319 & ~n8320 ;
  assign n8322 = \DataWidth_reg[1]/NET0131  & ~n8321 ;
  assign n8314 = \Datai[5]_pad  & ~n3918 ;
  assign n8315 = \InstQueue_reg[14][5]/NET0131  & ~n3914 ;
  assign n8316 = ~n3871 & n8315 ;
  assign n8317 = ~n8314 & ~n8316 ;
  assign n8323 = ~n4039 & ~n8317 ;
  assign n8324 = ~n8322 & ~n8323 ;
  assign n8325 = n933 & ~n8324 ;
  assign n8326 = ~n637 & n3914 ;
  assign n8327 = ~n8315 & ~n8326 ;
  assign n8328 = n965 & ~n8327 ;
  assign n8318 = n1867 & ~n8317 ;
  assign n8329 = \InstQueue_reg[14][5]/NET0131  & ~n3929 ;
  assign n8330 = ~n8318 & ~n8329 ;
  assign n8331 = ~n8328 & n8330 ;
  assign n8332 = ~n8325 & n8331 ;
  assign n8338 = n3987 & n8221 ;
  assign n8339 = n3871 & n8224 ;
  assign n8340 = ~n8338 & ~n8339 ;
  assign n8341 = \DataWidth_reg[1]/NET0131  & ~n8340 ;
  assign n8333 = \Datai[5]_pad  & ~n4050 ;
  assign n8334 = \InstQueue_reg[15][5]/NET0131  & ~n3862 ;
  assign n8335 = ~n3914 & n8334 ;
  assign n8336 = ~n8333 & ~n8335 ;
  assign n8342 = ~n4060 & ~n8336 ;
  assign n8343 = ~n8341 & ~n8342 ;
  assign n8344 = n933 & ~n8343 ;
  assign n8345 = ~n637 & n3862 ;
  assign n8346 = ~n8334 & ~n8345 ;
  assign n8347 = n965 & ~n8346 ;
  assign n8337 = n1867 & ~n8336 ;
  assign n8348 = \InstQueue_reg[15][5]/NET0131  & ~n3929 ;
  assign n8349 = ~n8337 & ~n8348 ;
  assign n8350 = ~n8347 & n8349 ;
  assign n8351 = ~n8344 & n8350 ;
  assign n8357 = n3914 & n8221 ;
  assign n8358 = n3862 & n8224 ;
  assign n8359 = ~n8357 & ~n8358 ;
  assign n8360 = \DataWidth_reg[1]/NET0131  & ~n8359 ;
  assign n8352 = \Datai[5]_pad  & ~n4072 ;
  assign n8353 = \InstQueue_reg[1][5]/NET0131  & ~n4071 ;
  assign n8354 = ~n3859 & n8353 ;
  assign n8355 = ~n8352 & ~n8354 ;
  assign n8361 = ~n4082 & ~n8355 ;
  assign n8362 = ~n8360 & ~n8361 ;
  assign n8363 = n933 & ~n8362 ;
  assign n8364 = ~n637 & n4071 ;
  assign n8365 = ~n8353 & ~n8364 ;
  assign n8366 = n965 & ~n8365 ;
  assign n8356 = n1867 & ~n8355 ;
  assign n8367 = \InstQueue_reg[1][5]/NET0131  & ~n3929 ;
  assign n8368 = ~n8356 & ~n8367 ;
  assign n8369 = ~n8366 & n8368 ;
  assign n8370 = ~n8363 & n8369 ;
  assign n8376 = n3859 & n8224 ;
  assign n8377 = n3862 & n8221 ;
  assign n8378 = ~n8376 & ~n8377 ;
  assign n8379 = \DataWidth_reg[1]/NET0131  & ~n8378 ;
  assign n8371 = \Datai[5]_pad  & ~n4094 ;
  assign n8372 = \InstQueue_reg[2][5]/NET0131  & ~n4093 ;
  assign n8373 = ~n4071 & n8372 ;
  assign n8374 = ~n8371 & ~n8373 ;
  assign n8380 = ~n4104 & ~n8374 ;
  assign n8381 = ~n8379 & ~n8380 ;
  assign n8382 = n933 & ~n8381 ;
  assign n8383 = ~n637 & n4093 ;
  assign n8384 = ~n8372 & ~n8383 ;
  assign n8385 = n965 & ~n8384 ;
  assign n8375 = n1867 & ~n8374 ;
  assign n8386 = \InstQueue_reg[2][5]/NET0131  & ~n3929 ;
  assign n8387 = ~n8375 & ~n8386 ;
  assign n8388 = ~n8385 & n8387 ;
  assign n8389 = ~n8382 & n8388 ;
  assign n8395 = n3859 & n8221 ;
  assign n8396 = n4071 & n8224 ;
  assign n8397 = ~n8395 & ~n8396 ;
  assign n8398 = \DataWidth_reg[1]/NET0131  & ~n8397 ;
  assign n8390 = \Datai[5]_pad  & ~n4116 ;
  assign n8391 = \InstQueue_reg[3][5]/NET0131  & ~n4115 ;
  assign n8392 = ~n4093 & n8391 ;
  assign n8393 = ~n8390 & ~n8392 ;
  assign n8399 = ~n4126 & ~n8393 ;
  assign n8400 = ~n8398 & ~n8399 ;
  assign n8401 = n933 & ~n8400 ;
  assign n8402 = ~n637 & n4115 ;
  assign n8403 = ~n8391 & ~n8402 ;
  assign n8404 = n965 & ~n8403 ;
  assign n8394 = n1867 & ~n8393 ;
  assign n8405 = \InstQueue_reg[3][5]/NET0131  & ~n3929 ;
  assign n8406 = ~n8394 & ~n8405 ;
  assign n8407 = ~n8404 & n8406 ;
  assign n8408 = ~n8401 & n8407 ;
  assign n8414 = n4071 & n8221 ;
  assign n8415 = n4093 & n8224 ;
  assign n8416 = ~n8414 & ~n8415 ;
  assign n8417 = \DataWidth_reg[1]/NET0131  & ~n8416 ;
  assign n8409 = \Datai[5]_pad  & ~n4138 ;
  assign n8410 = \InstQueue_reg[4][5]/NET0131  & ~n4137 ;
  assign n8411 = ~n4115 & n8410 ;
  assign n8412 = ~n8409 & ~n8411 ;
  assign n8418 = ~n4148 & ~n8412 ;
  assign n8419 = ~n8417 & ~n8418 ;
  assign n8420 = n933 & ~n8419 ;
  assign n8421 = ~n637 & n4137 ;
  assign n8422 = ~n8410 & ~n8421 ;
  assign n8423 = n965 & ~n8422 ;
  assign n8413 = n1867 & ~n8412 ;
  assign n8424 = \InstQueue_reg[4][5]/NET0131  & ~n3929 ;
  assign n8425 = ~n8413 & ~n8424 ;
  assign n8426 = ~n8423 & n8425 ;
  assign n8427 = ~n8420 & n8426 ;
  assign n8433 = n4093 & n8221 ;
  assign n8434 = n4115 & n8224 ;
  assign n8435 = ~n8433 & ~n8434 ;
  assign n8436 = \DataWidth_reg[1]/NET0131  & ~n8435 ;
  assign n8428 = \Datai[5]_pad  & ~n4160 ;
  assign n8429 = \InstQueue_reg[5][5]/NET0131  & ~n4159 ;
  assign n8430 = ~n4137 & n8429 ;
  assign n8431 = ~n8428 & ~n8430 ;
  assign n8437 = ~n4170 & ~n8431 ;
  assign n8438 = ~n8436 & ~n8437 ;
  assign n8439 = n933 & ~n8438 ;
  assign n8440 = ~n637 & n4159 ;
  assign n8441 = ~n8429 & ~n8440 ;
  assign n8442 = n965 & ~n8441 ;
  assign n8432 = n1867 & ~n8431 ;
  assign n8443 = \InstQueue_reg[5][5]/NET0131  & ~n3929 ;
  assign n8444 = ~n8432 & ~n8443 ;
  assign n8445 = ~n8442 & n8444 ;
  assign n8446 = ~n8439 & n8445 ;
  assign n8452 = n4115 & n8221 ;
  assign n8453 = n4137 & n8224 ;
  assign n8454 = ~n8452 & ~n8453 ;
  assign n8455 = \DataWidth_reg[1]/NET0131  & ~n8454 ;
  assign n8447 = \Datai[5]_pad  & ~n4182 ;
  assign n8448 = \InstQueue_reg[6][5]/NET0131  & ~n4181 ;
  assign n8449 = ~n4159 & n8448 ;
  assign n8450 = ~n8447 & ~n8449 ;
  assign n8456 = ~n4192 & ~n8450 ;
  assign n8457 = ~n8455 & ~n8456 ;
  assign n8458 = n933 & ~n8457 ;
  assign n8459 = ~n637 & n4181 ;
  assign n8460 = ~n8448 & ~n8459 ;
  assign n8461 = n965 & ~n8460 ;
  assign n8451 = n1867 & ~n8450 ;
  assign n8462 = \InstQueue_reg[6][5]/NET0131  & ~n3929 ;
  assign n8463 = ~n8451 & ~n8462 ;
  assign n8464 = ~n8461 & n8463 ;
  assign n8465 = ~n8458 & n8464 ;
  assign n8471 = n4137 & n8221 ;
  assign n8472 = n4159 & n8224 ;
  assign n8473 = ~n8471 & ~n8472 ;
  assign n8474 = \DataWidth_reg[1]/NET0131  & ~n8473 ;
  assign n8466 = \Datai[5]_pad  & ~n4203 ;
  assign n8467 = \InstQueue_reg[7][5]/NET0131  & ~n3944 ;
  assign n8468 = ~n4181 & n8467 ;
  assign n8469 = ~n8466 & ~n8468 ;
  assign n8475 = ~n4213 & ~n8469 ;
  assign n8476 = ~n8474 & ~n8475 ;
  assign n8477 = n933 & ~n8476 ;
  assign n8478 = ~n637 & n3944 ;
  assign n8479 = ~n8467 & ~n8478 ;
  assign n8480 = n965 & ~n8479 ;
  assign n8470 = n1867 & ~n8469 ;
  assign n8481 = \InstQueue_reg[7][5]/NET0131  & ~n3929 ;
  assign n8482 = ~n8470 & ~n8481 ;
  assign n8483 = ~n8480 & n8482 ;
  assign n8484 = ~n8477 & n8483 ;
  assign n8490 = n4159 & n8221 ;
  assign n8491 = n4181 & n8224 ;
  assign n8492 = ~n8490 & ~n8491 ;
  assign n8493 = \DataWidth_reg[1]/NET0131  & ~n8492 ;
  assign n8485 = \Datai[5]_pad  & ~n3950 ;
  assign n8486 = \InstQueue_reg[8][5]/NET0131  & ~n3946 ;
  assign n8487 = ~n3944 & n8486 ;
  assign n8488 = ~n8485 & ~n8487 ;
  assign n8494 = ~n4233 & ~n8488 ;
  assign n8495 = ~n8493 & ~n8494 ;
  assign n8496 = n933 & ~n8495 ;
  assign n8497 = ~n637 & n3946 ;
  assign n8498 = ~n8486 & ~n8497 ;
  assign n8499 = n965 & ~n8498 ;
  assign n8489 = n1867 & ~n8488 ;
  assign n8500 = \InstQueue_reg[8][5]/NET0131  & ~n3929 ;
  assign n8501 = ~n8489 & ~n8500 ;
  assign n8502 = ~n8499 & n8501 ;
  assign n8503 = ~n8496 & n8502 ;
  assign n8509 = n4181 & n8221 ;
  assign n8510 = n3944 & n8224 ;
  assign n8511 = ~n8509 & ~n8510 ;
  assign n8512 = \DataWidth_reg[1]/NET0131  & ~n8511 ;
  assign n8504 = \Datai[5]_pad  & ~n3974 ;
  assign n8505 = \InstQueue_reg[9][5]/NET0131  & ~n3937 ;
  assign n8506 = ~n3946 & n8505 ;
  assign n8507 = ~n8504 & ~n8506 ;
  assign n8513 = ~n4253 & ~n8507 ;
  assign n8514 = ~n8512 & ~n8513 ;
  assign n8515 = n933 & ~n8514 ;
  assign n8516 = ~n637 & n3937 ;
  assign n8517 = ~n8505 & ~n8516 ;
  assign n8518 = n965 & ~n8517 ;
  assign n8508 = n1867 & ~n8507 ;
  assign n8519 = \InstQueue_reg[9][5]/NET0131  & ~n3929 ;
  assign n8520 = ~n8508 & ~n8519 ;
  assign n8521 = ~n8518 & n8520 ;
  assign n8522 = ~n8515 & n8521 ;
  assign n8534 = ~\rEIP_reg[0]/NET0131  & ~\rEIP_reg[1]/NET0131  ;
  assign n8535 = \rEIP_reg[31]/NET0131  & ~n8534 ;
  assign n8536 = \rEIP_reg[2]/NET0131  & n8535 ;
  assign n8537 = \rEIP_reg[3]/NET0131  & n8536 ;
  assign n8538 = \rEIP_reg[4]/NET0131  & n8537 ;
  assign n8539 = \rEIP_reg[5]/NET0131  & n8538 ;
  assign n8540 = \rEIP_reg[6]/NET0131  & n8539 ;
  assign n8541 = \rEIP_reg[7]/NET0131  & n8540 ;
  assign n8542 = \rEIP_reg[8]/NET0131  & n8541 ;
  assign n8543 = \rEIP_reg[9]/NET0131  & n8542 ;
  assign n8544 = \rEIP_reg[10]/NET0131  & n8543 ;
  assign n8545 = \rEIP_reg[11]/NET0131  & n8544 ;
  assign n8546 = n5734 & n8545 ;
  assign n8547 = \rEIP_reg[14]/NET0131  & n8546 ;
  assign n8548 = \rEIP_reg[15]/NET0131  & n8547 ;
  assign n8549 = \rEIP_reg[16]/NET0131  & n8548 ;
  assign n8550 = n5831 & n8549 ;
  assign n8551 = \rEIP_reg[23]/NET0131  & n8550 ;
  assign n8552 = n5932 & n8551 ;
  assign n8553 = \rEIP_reg[26]/NET0131  & n8552 ;
  assign n8554 = \rEIP_reg[27]/NET0131  & n8553 ;
  assign n8555 = \rEIP_reg[28]/NET0131  & n8554 ;
  assign n8556 = \rEIP_reg[29]/NET0131  & n8555 ;
  assign n8558 = \rEIP_reg[30]/NET0131  & n8556 ;
  assign n8557 = ~\rEIP_reg[30]/NET0131  & ~n8556 ;
  assign n8559 = n825 & ~n8557 ;
  assign n8560 = ~n8558 & n8559 ;
  assign n8523 = \Address[28]_pad  & ~n824 ;
  assign n8525 = \rEIP_reg[0]/NET0131  & \rEIP_reg[31]/NET0131  ;
  assign n8526 = n5858 & n8525 ;
  assign n8527 = n5970 & n8526 ;
  assign n8528 = \rEIP_reg[27]/NET0131  & n8527 ;
  assign n8529 = \rEIP_reg[28]/NET0131  & n8528 ;
  assign n8531 = \rEIP_reg[29]/NET0131  & n8529 ;
  assign n8524 = \State_reg[2]/NET0131  & n824 ;
  assign n8530 = ~\rEIP_reg[29]/NET0131  & ~n8529 ;
  assign n8532 = n8524 & ~n8530 ;
  assign n8533 = ~n8531 & n8532 ;
  assign n8561 = ~n8523 & ~n8533 ;
  assign n8562 = ~n8560 & n8561 ;
  assign n8564 = ~n828 & ~n7469 ;
  assign n8565 = n923 & ~n8564 ;
  assign n8566 = n3827 & ~n8565 ;
  assign n8567 = \Datao[25]_pad  & ~n8566 ;
  assign n8568 = ~n828 & n7470 ;
  assign n8569 = ~n8567 & ~n8568 ;
  assign n8570 = n929 & ~n8569 ;
  assign n8563 = \uWord_reg[9]/NET0131  & n3809 ;
  assign n8571 = \Datao[25]_pad  & ~n3821 ;
  assign n8572 = ~n8563 & ~n8571 ;
  assign n8573 = ~n8570 & n8572 ;
  assign n8575 = ~n857 & n929 ;
  assign n8576 = n3821 & ~n8575 ;
  assign n8577 = \Datao[17]_pad  & ~n8576 ;
  assign n8574 = \uWord_reg[1]/NET0131  & n3809 ;
  assign n8578 = ~n828 & n929 ;
  assign n8579 = n7428 & n8578 ;
  assign n8580 = ~n8574 & ~n8579 ;
  assign n8581 = ~n8577 & n8580 ;
  assign n8583 = ~n828 & ~n7397 ;
  assign n8584 = n923 & ~n8583 ;
  assign n8585 = n3827 & ~n8584 ;
  assign n8586 = \Datao[16]_pad  & ~n8585 ;
  assign n8587 = ~n828 & n7398 ;
  assign n8588 = ~n8586 & ~n8587 ;
  assign n8589 = n929 & ~n8588 ;
  assign n8582 = \uWord_reg[0]/NET0131  & n3809 ;
  assign n8590 = \Datao[16]_pad  & ~n3821 ;
  assign n8591 = ~n8582 & ~n8590 ;
  assign n8592 = ~n8589 & n8591 ;
  assign n8594 = ~n828 & n7453 ;
  assign n8595 = \Datao[21]_pad  & ~n857 ;
  assign n8596 = ~n8594 & ~n8595 ;
  assign n8597 = n929 & ~n8596 ;
  assign n8593 = \uWord_reg[5]/NET0131  & n3809 ;
  assign n8598 = \Datao[21]_pad  & ~n3821 ;
  assign n8599 = ~n8593 & ~n8598 ;
  assign n8600 = ~n8597 & n8599 ;
  assign n8601 = ~\Flush_reg/NET0131  & n960 ;
  assign n8602 = ~n929 & ~n953 ;
  assign n8603 = ~n3809 & n8602 ;
  assign n8604 = ~n8601 & n8603 ;
  assign n8605 = n6773 & n8604 ;
  assign n8606 = \InstQueueWr_Addr_reg[2]/NET0131  & ~n8605 ;
  assign n8607 = ~n2099 & ~n3912 ;
  assign n8608 = \InstQueueWr_Addr_reg[2]/NET0131  & ~n8607 ;
  assign n8609 = ~n2098 & ~n8608 ;
  assign n8610 = ~n965 & ~n8609 ;
  assign n8611 = ~n2098 & n3912 ;
  assign n8612 = ~\InstQueueWr_Addr_reg[2]/NET0131  & ~n3860 ;
  assign n8613 = ~n969 & n8612 ;
  assign n8614 = ~n8611 & n8613 ;
  assign n8615 = ~n3861 & ~n8614 ;
  assign n8616 = ~n8610 & n8615 ;
  assign n8617 = ~n8606 & ~n8616 ;
  assign n8625 = \rEIP_reg[17]/NET0131  & n8549 ;
  assign n8626 = ~\rEIP_reg[18]/NET0131  & ~n8625 ;
  assign n8624 = n5739 & n8549 ;
  assign n8627 = n825 & ~n8624 ;
  assign n8628 = ~n8626 & n8627 ;
  assign n8618 = \Address[16]_pad  & ~n824 ;
  assign n8621 = n6683 & n8525 ;
  assign n8619 = n5738 & n8525 ;
  assign n8620 = ~\rEIP_reg[17]/NET0131  & ~n8619 ;
  assign n8622 = n8524 & ~n8620 ;
  assign n8623 = ~n8621 & n8622 ;
  assign n8629 = ~n8618 & ~n8623 ;
  assign n8630 = ~n8628 & n8629 ;
  assign n8634 = ~\EAX_reg[2]/NET0131  & n857 ;
  assign n8633 = ~\Datao[2]_pad  & ~n857 ;
  assign n8635 = n929 & ~n8633 ;
  assign n8636 = ~n8634 & n8635 ;
  assign n8631 = \lWord_reg[2]/NET0131  & n3809 ;
  assign n8632 = \Datao[2]_pad  & ~n3821 ;
  assign n8637 = ~n8631 & ~n8632 ;
  assign n8638 = ~n8636 & n8637 ;
  assign n8642 = ~\EAX_reg[4]/NET0131  & n857 ;
  assign n8641 = ~\Datao[4]_pad  & ~n857 ;
  assign n8643 = n929 & ~n8641 ;
  assign n8644 = ~n8642 & n8643 ;
  assign n8639 = \lWord_reg[4]/NET0131  & n3809 ;
  assign n8640 = \Datao[4]_pad  & ~n3821 ;
  assign n8645 = ~n8639 & ~n8640 ;
  assign n8646 = ~n8644 & n8645 ;
  assign n8650 = ~\EAX_reg[3]/NET0131  & n857 ;
  assign n8649 = ~\Datao[3]_pad  & ~n857 ;
  assign n8651 = n929 & ~n8649 ;
  assign n8652 = ~n8650 & n8651 ;
  assign n8647 = \lWord_reg[3]/NET0131  & n3809 ;
  assign n8648 = \Datao[3]_pad  & ~n3821 ;
  assign n8653 = ~n8647 & ~n8648 ;
  assign n8654 = ~n8652 & n8653 ;
  assign n8658 = ~\EAX_reg[5]/NET0131  & n857 ;
  assign n8657 = ~\Datao[5]_pad  & ~n857 ;
  assign n8659 = n929 & ~n8657 ;
  assign n8660 = ~n8658 & n8659 ;
  assign n8655 = \lWord_reg[5]/NET0131  & n3809 ;
  assign n8656 = \Datao[5]_pad  & ~n3821 ;
  assign n8661 = ~n8655 & ~n8656 ;
  assign n8662 = ~n8660 & n8661 ;
  assign n8666 = ~\EAX_reg[6]/NET0131  & n857 ;
  assign n8665 = ~\Datao[6]_pad  & ~n857 ;
  assign n8667 = n929 & ~n8665 ;
  assign n8668 = ~n8666 & n8667 ;
  assign n8663 = \lWord_reg[6]/NET0131  & n3809 ;
  assign n8664 = \Datao[6]_pad  & ~n3821 ;
  assign n8669 = ~n8663 & ~n8664 ;
  assign n8670 = ~n8668 & n8669 ;
  assign n8674 = ~\EAX_reg[7]/NET0131  & n857 ;
  assign n8673 = ~\Datao[7]_pad  & ~n857 ;
  assign n8675 = n929 & ~n8673 ;
  assign n8676 = ~n8674 & n8675 ;
  assign n8671 = \lWord_reg[7]/NET0131  & n3809 ;
  assign n8672 = \Datao[7]_pad  & ~n3821 ;
  assign n8677 = ~n8671 & ~n8672 ;
  assign n8678 = ~n8676 & n8677 ;
  assign n8682 = ~\EAX_reg[8]/NET0131  & n857 ;
  assign n8681 = ~\Datao[8]_pad  & ~n857 ;
  assign n8683 = n929 & ~n8681 ;
  assign n8684 = ~n8682 & n8683 ;
  assign n8679 = \lWord_reg[8]/NET0131  & n3809 ;
  assign n8680 = \Datao[8]_pad  & ~n3821 ;
  assign n8685 = ~n8679 & ~n8680 ;
  assign n8686 = ~n8684 & n8685 ;
  assign n8690 = ~\EAX_reg[9]/NET0131  & n857 ;
  assign n8689 = ~\Datao[9]_pad  & ~n857 ;
  assign n8691 = n929 & ~n8689 ;
  assign n8692 = ~n8690 & n8691 ;
  assign n8687 = \lWord_reg[9]/NET0131  & n3809 ;
  assign n8688 = \Datao[9]_pad  & ~n3821 ;
  assign n8693 = ~n8687 & ~n8688 ;
  assign n8694 = ~n8692 & n8693 ;
  assign n8698 = ~\EAX_reg[0]/NET0131  & n857 ;
  assign n8697 = ~\Datao[0]_pad  & ~n857 ;
  assign n8699 = n929 & ~n8697 ;
  assign n8700 = ~n8698 & n8699 ;
  assign n8695 = \lWord_reg[0]/NET0131  & n3809 ;
  assign n8696 = \Datao[0]_pad  & ~n3821 ;
  assign n8701 = ~n8695 & ~n8696 ;
  assign n8702 = ~n8700 & n8701 ;
  assign n8706 = ~\EAX_reg[10]/NET0131  & n857 ;
  assign n8705 = ~\Datao[10]_pad  & ~n857 ;
  assign n8707 = n929 & ~n8705 ;
  assign n8708 = ~n8706 & n8707 ;
  assign n8703 = \lWord_reg[10]/NET0131  & n3809 ;
  assign n8704 = \Datao[10]_pad  & ~n3821 ;
  assign n8709 = ~n8703 & ~n8704 ;
  assign n8710 = ~n8708 & n8709 ;
  assign n8714 = ~\EAX_reg[12]/NET0131  & n857 ;
  assign n8713 = ~\Datao[12]_pad  & ~n857 ;
  assign n8715 = n929 & ~n8713 ;
  assign n8716 = ~n8714 & n8715 ;
  assign n8711 = \lWord_reg[12]/NET0131  & n3809 ;
  assign n8712 = \Datao[12]_pad  & ~n3821 ;
  assign n8717 = ~n8711 & ~n8712 ;
  assign n8718 = ~n8716 & n8717 ;
  assign n8722 = ~\EAX_reg[11]/NET0131  & n857 ;
  assign n8721 = ~\Datao[11]_pad  & ~n857 ;
  assign n8723 = n929 & ~n8721 ;
  assign n8724 = ~n8722 & n8723 ;
  assign n8719 = \lWord_reg[11]/NET0131  & n3809 ;
  assign n8720 = \Datao[11]_pad  & ~n3821 ;
  assign n8725 = ~n8719 & ~n8720 ;
  assign n8726 = ~n8724 & n8725 ;
  assign n8730 = ~\EAX_reg[13]/NET0131  & n857 ;
  assign n8729 = ~\Datao[13]_pad  & ~n857 ;
  assign n8731 = n929 & ~n8729 ;
  assign n8732 = ~n8730 & n8731 ;
  assign n8727 = \lWord_reg[13]/NET0131  & n3809 ;
  assign n8728 = \Datao[13]_pad  & ~n3821 ;
  assign n8733 = ~n8727 & ~n8728 ;
  assign n8734 = ~n8732 & n8733 ;
  assign n8738 = ~\EAX_reg[14]/NET0131  & n857 ;
  assign n8737 = ~\Datao[14]_pad  & ~n857 ;
  assign n8739 = n929 & ~n8737 ;
  assign n8740 = ~n8738 & n8739 ;
  assign n8735 = \lWord_reg[14]/NET0131  & n3809 ;
  assign n8736 = \Datao[14]_pad  & ~n3821 ;
  assign n8741 = ~n8735 & ~n8736 ;
  assign n8742 = ~n8740 & n8741 ;
  assign n8746 = ~\EAX_reg[15]/NET0131  & n857 ;
  assign n8745 = ~\Datao[15]_pad  & ~n857 ;
  assign n8747 = n929 & ~n8745 ;
  assign n8748 = ~n8746 & n8747 ;
  assign n8743 = \lWord_reg[15]/NET0131  & n3809 ;
  assign n8744 = \Datao[15]_pad  & ~n3821 ;
  assign n8749 = ~n8743 & ~n8744 ;
  assign n8750 = ~n8748 & n8749 ;
  assign n8754 = ~\EAX_reg[1]/NET0131  & n857 ;
  assign n8753 = ~\Datao[1]_pad  & ~n857 ;
  assign n8755 = n929 & ~n8753 ;
  assign n8756 = ~n8754 & n8755 ;
  assign n8751 = \lWord_reg[1]/NET0131  & n3809 ;
  assign n8752 = \Datao[1]_pad  & ~n3821 ;
  assign n8757 = ~n8751 & ~n8752 ;
  assign n8758 = ~n8756 & n8757 ;
  assign n8759 = \InstQueueWr_Addr_reg[3]/NET0131  & ~n3861 ;
  assign n8760 = ~n3944 & ~n8759 ;
  assign n8762 = ~n3913 & ~n8760 ;
  assign n8763 = ~n4181 & ~n8762 ;
  assign n8764 = ~n3870 & ~n8763 ;
  assign n8765 = ~n3986 & ~n4159 ;
  assign n8766 = ~n8764 & n8765 ;
  assign n8767 = n969 & ~n3987 ;
  assign n8768 = ~n8766 & n8767 ;
  assign n8769 = \InstQueueWr_Addr_reg[3]/NET0131  & ~n8605 ;
  assign n8761 = n965 & ~n8760 ;
  assign n8770 = n2100 & ~n8763 ;
  assign n8771 = ~n8761 & ~n8770 ;
  assign n8772 = ~n8769 & n8771 ;
  assign n8773 = ~n8768 & n8772 ;
  assign n8774 = \InstQueueWr_Addr_reg[1]/NET0131  & ~n8604 ;
  assign n8775 = ~\InstQueueWr_Addr_reg[0]/NET0131  & n965 ;
  assign n8776 = \InstQueueWr_Addr_reg[1]/NET0131  & ~n969 ;
  assign n8777 = n6773 & n8776 ;
  assign n8778 = ~n8775 & n8777 ;
  assign n8779 = \InstQueueWr_Addr_reg[0]/NET0131  & n965 ;
  assign n8780 = ~\InstQueueWr_Addr_reg[1]/NET0131  & ~n8779 ;
  assign n8781 = ~n2100 & n8780 ;
  assign n8782 = ~n8778 & ~n8781 ;
  assign n8783 = ~n8774 & ~n8782 ;
  assign n8786 = ~n929 & ~n3187 ;
  assign n8787 = \InstQueueWr_Addr_reg[0]/NET0131  & ~n8786 ;
  assign n8784 = ~\Flush_reg/NET0131  & ~\InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n8785 = n960 & ~n8784 ;
  assign n8788 = ~n8775 & ~n8785 ;
  assign n8789 = ~n8787 & n8788 ;
  assign n8795 = ~\Datai[25]_pad  & ~n3896 ;
  assign n8796 = ~n3897 & ~n8795 ;
  assign n8797 = n3871 & n8796 ;
  assign n8798 = ~\Datai[17]_pad  & ~n3905 ;
  assign n8799 = ~n3906 & ~n8798 ;
  assign n8800 = n3914 & n8799 ;
  assign n8801 = ~n8797 & ~n8800 ;
  assign n8802 = \DataWidth_reg[1]/NET0131  & ~n8801 ;
  assign n8790 = \Datai[1]_pad  & ~n3863 ;
  assign n8791 = \InstQueue_reg[0][1]/NET0131  & ~n3859 ;
  assign n8792 = ~n3862 & n8791 ;
  assign n8793 = ~n8790 & ~n8792 ;
  assign n8803 = ~n3919 & ~n8793 ;
  assign n8804 = ~n8802 & ~n8803 ;
  assign n8805 = n933 & ~n8804 ;
  assign n8806 = ~n604 & n3859 ;
  assign n8807 = ~n8791 & ~n8806 ;
  assign n8808 = n965 & ~n8807 ;
  assign n8794 = n1867 & ~n8793 ;
  assign n8809 = \InstQueue_reg[0][1]/NET0131  & ~n3929 ;
  assign n8810 = ~n8794 & ~n8809 ;
  assign n8811 = ~n8808 & n8810 ;
  assign n8812 = ~n8805 & n8811 ;
  assign n8818 = n3944 & n8796 ;
  assign n8819 = n3946 & n8799 ;
  assign n8820 = ~n8818 & ~n8819 ;
  assign n8821 = \DataWidth_reg[1]/NET0131  & ~n8820 ;
  assign n8813 = \Datai[1]_pad  & ~n3938 ;
  assign n8814 = \InstQueue_reg[10][1]/NET0131  & ~n3935 ;
  assign n8815 = ~n3937 & n8814 ;
  assign n8816 = ~n8813 & ~n8815 ;
  assign n8822 = ~n3951 & ~n8816 ;
  assign n8823 = ~n8821 & ~n8822 ;
  assign n8824 = n933 & ~n8823 ;
  assign n8825 = ~n604 & n3935 ;
  assign n8826 = ~n8814 & ~n8825 ;
  assign n8827 = n965 & ~n8826 ;
  assign n8817 = n1867 & ~n8816 ;
  assign n8828 = \InstQueue_reg[10][1]/NET0131  & ~n3929 ;
  assign n8829 = ~n8817 & ~n8828 ;
  assign n8830 = ~n8827 & n8829 ;
  assign n8831 = ~n8824 & n8830 ;
  assign n8837 = ~\Datai[24]_pad  & ~n3895 ;
  assign n8838 = ~n3896 & ~n8837 ;
  assign n8839 = n3946 & n8838 ;
  assign n8840 = ~\Datai[16]_pad  & ~n3904 ;
  assign n8841 = ~n3905 & ~n8840 ;
  assign n8842 = n3937 & n8841 ;
  assign n8843 = ~n8839 & ~n8842 ;
  assign n8844 = \DataWidth_reg[1]/NET0131  & ~n8843 ;
  assign n8832 = \Datai[0]_pad  & ~n3964 ;
  assign n8833 = \InstQueue_reg[11][0]/NET0131  & ~n3963 ;
  assign n8834 = ~n3935 & n8833 ;
  assign n8835 = ~n8832 & ~n8834 ;
  assign n8845 = ~n3975 & ~n8835 ;
  assign n8846 = ~n8844 & ~n8845 ;
  assign n8847 = n933 & ~n8846 ;
  assign n8848 = ~n508 & n3963 ;
  assign n8849 = ~n8833 & ~n8848 ;
  assign n8850 = n965 & ~n8849 ;
  assign n8836 = n1867 & ~n8835 ;
  assign n8851 = \InstQueue_reg[11][0]/NET0131  & ~n3929 ;
  assign n8852 = ~n8836 & ~n8851 ;
  assign n8853 = ~n8850 & n8852 ;
  assign n8854 = ~n8847 & n8853 ;
  assign n8860 = n3946 & n8796 ;
  assign n8861 = n3937 & n8799 ;
  assign n8862 = ~n8860 & ~n8861 ;
  assign n8863 = \DataWidth_reg[1]/NET0131  & ~n8862 ;
  assign n8855 = \Datai[1]_pad  & ~n3964 ;
  assign n8856 = \InstQueue_reg[11][1]/NET0131  & ~n3963 ;
  assign n8857 = ~n3935 & n8856 ;
  assign n8858 = ~n8855 & ~n8857 ;
  assign n8864 = ~n3975 & ~n8858 ;
  assign n8865 = ~n8863 & ~n8864 ;
  assign n8866 = n933 & ~n8865 ;
  assign n8867 = ~n604 & n3963 ;
  assign n8868 = ~n8856 & ~n8867 ;
  assign n8869 = n965 & ~n8868 ;
  assign n8859 = n1867 & ~n8858 ;
  assign n8870 = \InstQueue_reg[11][1]/NET0131  & ~n3929 ;
  assign n8871 = ~n8859 & ~n8870 ;
  assign n8872 = ~n8869 & n8871 ;
  assign n8873 = ~n8866 & n8872 ;
  assign n8879 = n3937 & n8796 ;
  assign n8880 = n3935 & n8799 ;
  assign n8881 = ~n8879 & ~n8880 ;
  assign n8882 = \DataWidth_reg[1]/NET0131  & ~n8881 ;
  assign n8874 = \Datai[1]_pad  & ~n3988 ;
  assign n8875 = \InstQueue_reg[12][1]/NET0131  & ~n3987 ;
  assign n8876 = ~n3963 & n8875 ;
  assign n8877 = ~n8874 & ~n8876 ;
  assign n8883 = ~n3998 & ~n8877 ;
  assign n8884 = ~n8882 & ~n8883 ;
  assign n8885 = n933 & ~n8884 ;
  assign n8886 = ~n604 & n3987 ;
  assign n8887 = ~n8875 & ~n8886 ;
  assign n8888 = n965 & ~n8887 ;
  assign n8878 = n1867 & ~n8877 ;
  assign n8889 = \InstQueue_reg[12][1]/NET0131  & ~n3929 ;
  assign n8890 = ~n8878 & ~n8889 ;
  assign n8891 = ~n8888 & n8890 ;
  assign n8892 = ~n8885 & n8891 ;
  assign n8898 = n3935 & n8796 ;
  assign n8899 = n3963 & n8799 ;
  assign n8900 = ~n8898 & ~n8899 ;
  assign n8901 = \DataWidth_reg[1]/NET0131  & ~n8900 ;
  assign n8893 = \Datai[1]_pad  & ~n4009 ;
  assign n8894 = \InstQueue_reg[13][1]/NET0131  & ~n3871 ;
  assign n8895 = ~n3987 & n8894 ;
  assign n8896 = ~n8893 & ~n8895 ;
  assign n8902 = ~n4019 & ~n8896 ;
  assign n8903 = ~n8901 & ~n8902 ;
  assign n8904 = n933 & ~n8903 ;
  assign n8905 = ~n604 & n3871 ;
  assign n8906 = ~n8894 & ~n8905 ;
  assign n8907 = n965 & ~n8906 ;
  assign n8897 = n1867 & ~n8896 ;
  assign n8908 = \InstQueue_reg[13][1]/NET0131  & ~n3929 ;
  assign n8909 = ~n8897 & ~n8908 ;
  assign n8910 = ~n8907 & n8909 ;
  assign n8911 = ~n8904 & n8910 ;
  assign n8917 = n3963 & n8796 ;
  assign n8918 = n3987 & n8799 ;
  assign n8919 = ~n8917 & ~n8918 ;
  assign n8920 = \DataWidth_reg[1]/NET0131  & ~n8919 ;
  assign n8912 = \Datai[1]_pad  & ~n3918 ;
  assign n8913 = \InstQueue_reg[14][1]/NET0131  & ~n3914 ;
  assign n8914 = ~n3871 & n8913 ;
  assign n8915 = ~n8912 & ~n8914 ;
  assign n8921 = ~n4039 & ~n8915 ;
  assign n8922 = ~n8920 & ~n8921 ;
  assign n8923 = n933 & ~n8922 ;
  assign n8924 = ~n604 & n3914 ;
  assign n8925 = ~n8913 & ~n8924 ;
  assign n8926 = n965 & ~n8925 ;
  assign n8916 = n1867 & ~n8915 ;
  assign n8927 = \InstQueue_reg[14][1]/NET0131  & ~n3929 ;
  assign n8928 = ~n8916 & ~n8927 ;
  assign n8929 = ~n8926 & n8928 ;
  assign n8930 = ~n8923 & n8929 ;
  assign n8936 = n3987 & n8796 ;
  assign n8937 = n3871 & n8799 ;
  assign n8938 = ~n8936 & ~n8937 ;
  assign n8939 = \DataWidth_reg[1]/NET0131  & ~n8938 ;
  assign n8931 = \Datai[1]_pad  & ~n4050 ;
  assign n8932 = \InstQueue_reg[15][1]/NET0131  & ~n3862 ;
  assign n8933 = ~n3914 & n8932 ;
  assign n8934 = ~n8931 & ~n8933 ;
  assign n8940 = ~n4060 & ~n8934 ;
  assign n8941 = ~n8939 & ~n8940 ;
  assign n8942 = n933 & ~n8941 ;
  assign n8943 = ~n604 & n3862 ;
  assign n8944 = ~n8932 & ~n8943 ;
  assign n8945 = n965 & ~n8944 ;
  assign n8935 = n1867 & ~n8934 ;
  assign n8946 = \InstQueue_reg[15][1]/NET0131  & ~n3929 ;
  assign n8947 = ~n8935 & ~n8946 ;
  assign n8948 = ~n8945 & n8947 ;
  assign n8949 = ~n8942 & n8948 ;
  assign n8955 = n3914 & n8796 ;
  assign n8956 = n3862 & n8799 ;
  assign n8957 = ~n8955 & ~n8956 ;
  assign n8958 = \DataWidth_reg[1]/NET0131  & ~n8957 ;
  assign n8950 = \Datai[1]_pad  & ~n4072 ;
  assign n8951 = \InstQueue_reg[1][1]/NET0131  & ~n4071 ;
  assign n8952 = ~n3859 & n8951 ;
  assign n8953 = ~n8950 & ~n8952 ;
  assign n8959 = ~n4082 & ~n8953 ;
  assign n8960 = ~n8958 & ~n8959 ;
  assign n8961 = n933 & ~n8960 ;
  assign n8962 = ~n604 & n4071 ;
  assign n8963 = ~n8951 & ~n8962 ;
  assign n8964 = n965 & ~n8963 ;
  assign n8954 = n1867 & ~n8953 ;
  assign n8965 = \InstQueue_reg[1][1]/NET0131  & ~n3929 ;
  assign n8966 = ~n8954 & ~n8965 ;
  assign n8967 = ~n8964 & n8966 ;
  assign n8968 = ~n8961 & n8967 ;
  assign n8974 = n3859 & n8799 ;
  assign n8975 = n3862 & n8796 ;
  assign n8976 = ~n8974 & ~n8975 ;
  assign n8977 = \DataWidth_reg[1]/NET0131  & ~n8976 ;
  assign n8969 = \Datai[1]_pad  & ~n4094 ;
  assign n8970 = \InstQueue_reg[2][1]/NET0131  & ~n4093 ;
  assign n8971 = ~n4071 & n8970 ;
  assign n8972 = ~n8969 & ~n8971 ;
  assign n8978 = ~n4104 & ~n8972 ;
  assign n8979 = ~n8977 & ~n8978 ;
  assign n8980 = n933 & ~n8979 ;
  assign n8981 = ~n604 & n4093 ;
  assign n8982 = ~n8970 & ~n8981 ;
  assign n8983 = n965 & ~n8982 ;
  assign n8973 = n1867 & ~n8972 ;
  assign n8984 = \InstQueue_reg[2][1]/NET0131  & ~n3929 ;
  assign n8985 = ~n8973 & ~n8984 ;
  assign n8986 = ~n8983 & n8985 ;
  assign n8987 = ~n8980 & n8986 ;
  assign n8993 = n3859 & n8838 ;
  assign n8994 = n4071 & n8841 ;
  assign n8995 = ~n8993 & ~n8994 ;
  assign n8996 = \DataWidth_reg[1]/NET0131  & ~n8995 ;
  assign n8988 = \Datai[0]_pad  & ~n4116 ;
  assign n8989 = \InstQueue_reg[3][0]/NET0131  & ~n4115 ;
  assign n8990 = ~n4093 & n8989 ;
  assign n8991 = ~n8988 & ~n8990 ;
  assign n8997 = ~n4126 & ~n8991 ;
  assign n8998 = ~n8996 & ~n8997 ;
  assign n8999 = n933 & ~n8998 ;
  assign n9000 = ~n508 & n4115 ;
  assign n9001 = ~n8989 & ~n9000 ;
  assign n9002 = n965 & ~n9001 ;
  assign n8992 = n1867 & ~n8991 ;
  assign n9003 = \InstQueue_reg[3][0]/NET0131  & ~n3929 ;
  assign n9004 = ~n8992 & ~n9003 ;
  assign n9005 = ~n9002 & n9004 ;
  assign n9006 = ~n8999 & n9005 ;
  assign n9012 = n3859 & n8796 ;
  assign n9013 = n4071 & n8799 ;
  assign n9014 = ~n9012 & ~n9013 ;
  assign n9015 = \DataWidth_reg[1]/NET0131  & ~n9014 ;
  assign n9007 = \Datai[1]_pad  & ~n4116 ;
  assign n9008 = \InstQueue_reg[3][1]/NET0131  & ~n4115 ;
  assign n9009 = ~n4093 & n9008 ;
  assign n9010 = ~n9007 & ~n9009 ;
  assign n9016 = ~n4126 & ~n9010 ;
  assign n9017 = ~n9015 & ~n9016 ;
  assign n9018 = n933 & ~n9017 ;
  assign n9019 = ~n604 & n4115 ;
  assign n9020 = ~n9008 & ~n9019 ;
  assign n9021 = n965 & ~n9020 ;
  assign n9011 = n1867 & ~n9010 ;
  assign n9022 = \InstQueue_reg[3][1]/NET0131  & ~n3929 ;
  assign n9023 = ~n9011 & ~n9022 ;
  assign n9024 = ~n9021 & n9023 ;
  assign n9025 = ~n9018 & n9024 ;
  assign n9031 = n4071 & n8796 ;
  assign n9032 = n4093 & n8799 ;
  assign n9033 = ~n9031 & ~n9032 ;
  assign n9034 = \DataWidth_reg[1]/NET0131  & ~n9033 ;
  assign n9026 = \Datai[1]_pad  & ~n4138 ;
  assign n9027 = \InstQueue_reg[4][1]/NET0131  & ~n4137 ;
  assign n9028 = ~n4115 & n9027 ;
  assign n9029 = ~n9026 & ~n9028 ;
  assign n9035 = ~n4148 & ~n9029 ;
  assign n9036 = ~n9034 & ~n9035 ;
  assign n9037 = n933 & ~n9036 ;
  assign n9038 = ~n604 & n4137 ;
  assign n9039 = ~n9027 & ~n9038 ;
  assign n9040 = n965 & ~n9039 ;
  assign n9030 = n1867 & ~n9029 ;
  assign n9041 = \InstQueue_reg[4][1]/NET0131  & ~n3929 ;
  assign n9042 = ~n9030 & ~n9041 ;
  assign n9043 = ~n9040 & n9042 ;
  assign n9044 = ~n9037 & n9043 ;
  assign n9050 = n4093 & n8796 ;
  assign n9051 = n4115 & n8799 ;
  assign n9052 = ~n9050 & ~n9051 ;
  assign n9053 = \DataWidth_reg[1]/NET0131  & ~n9052 ;
  assign n9045 = \Datai[1]_pad  & ~n4160 ;
  assign n9046 = \InstQueue_reg[5][1]/NET0131  & ~n4159 ;
  assign n9047 = ~n4137 & n9046 ;
  assign n9048 = ~n9045 & ~n9047 ;
  assign n9054 = ~n4170 & ~n9048 ;
  assign n9055 = ~n9053 & ~n9054 ;
  assign n9056 = n933 & ~n9055 ;
  assign n9057 = ~n604 & n4159 ;
  assign n9058 = ~n9046 & ~n9057 ;
  assign n9059 = n965 & ~n9058 ;
  assign n9049 = n1867 & ~n9048 ;
  assign n9060 = \InstQueue_reg[5][1]/NET0131  & ~n3929 ;
  assign n9061 = ~n9049 & ~n9060 ;
  assign n9062 = ~n9059 & n9061 ;
  assign n9063 = ~n9056 & n9062 ;
  assign n9069 = n4115 & n8796 ;
  assign n9070 = n4137 & n8799 ;
  assign n9071 = ~n9069 & ~n9070 ;
  assign n9072 = \DataWidth_reg[1]/NET0131  & ~n9071 ;
  assign n9064 = \Datai[1]_pad  & ~n4182 ;
  assign n9065 = \InstQueue_reg[6][1]/NET0131  & ~n4181 ;
  assign n9066 = ~n4159 & n9065 ;
  assign n9067 = ~n9064 & ~n9066 ;
  assign n9073 = ~n4192 & ~n9067 ;
  assign n9074 = ~n9072 & ~n9073 ;
  assign n9075 = n933 & ~n9074 ;
  assign n9076 = ~n604 & n4181 ;
  assign n9077 = ~n9065 & ~n9076 ;
  assign n9078 = n965 & ~n9077 ;
  assign n9068 = n1867 & ~n9067 ;
  assign n9079 = \InstQueue_reg[6][1]/NET0131  & ~n3929 ;
  assign n9080 = ~n9068 & ~n9079 ;
  assign n9081 = ~n9078 & n9080 ;
  assign n9082 = ~n9075 & n9081 ;
  assign n9088 = n4137 & n8838 ;
  assign n9089 = n4159 & n8841 ;
  assign n9090 = ~n9088 & ~n9089 ;
  assign n9091 = \DataWidth_reg[1]/NET0131  & ~n9090 ;
  assign n9083 = \Datai[0]_pad  & ~n4203 ;
  assign n9084 = \InstQueue_reg[7][0]/NET0131  & ~n3944 ;
  assign n9085 = ~n4181 & n9084 ;
  assign n9086 = ~n9083 & ~n9085 ;
  assign n9092 = ~n4213 & ~n9086 ;
  assign n9093 = ~n9091 & ~n9092 ;
  assign n9094 = n933 & ~n9093 ;
  assign n9095 = ~n508 & n3944 ;
  assign n9096 = ~n9084 & ~n9095 ;
  assign n9097 = n965 & ~n9096 ;
  assign n9087 = n1867 & ~n9086 ;
  assign n9098 = \InstQueue_reg[7][0]/NET0131  & ~n3929 ;
  assign n9099 = ~n9087 & ~n9098 ;
  assign n9100 = ~n9097 & n9099 ;
  assign n9101 = ~n9094 & n9100 ;
  assign n9107 = n4137 & n8796 ;
  assign n9108 = n4159 & n8799 ;
  assign n9109 = ~n9107 & ~n9108 ;
  assign n9110 = \DataWidth_reg[1]/NET0131  & ~n9109 ;
  assign n9102 = \Datai[1]_pad  & ~n4203 ;
  assign n9103 = \InstQueue_reg[7][1]/NET0131  & ~n3944 ;
  assign n9104 = ~n4181 & n9103 ;
  assign n9105 = ~n9102 & ~n9104 ;
  assign n9111 = ~n4213 & ~n9105 ;
  assign n9112 = ~n9110 & ~n9111 ;
  assign n9113 = n933 & ~n9112 ;
  assign n9114 = ~n604 & n3944 ;
  assign n9115 = ~n9103 & ~n9114 ;
  assign n9116 = n965 & ~n9115 ;
  assign n9106 = n1867 & ~n9105 ;
  assign n9117 = \InstQueue_reg[7][1]/NET0131  & ~n3929 ;
  assign n9118 = ~n9106 & ~n9117 ;
  assign n9119 = ~n9116 & n9118 ;
  assign n9120 = ~n9113 & n9119 ;
  assign n9126 = n4159 & n8796 ;
  assign n9127 = n4181 & n8799 ;
  assign n9128 = ~n9126 & ~n9127 ;
  assign n9129 = \DataWidth_reg[1]/NET0131  & ~n9128 ;
  assign n9121 = \Datai[1]_pad  & ~n3950 ;
  assign n9122 = \InstQueue_reg[8][1]/NET0131  & ~n3946 ;
  assign n9123 = ~n3944 & n9122 ;
  assign n9124 = ~n9121 & ~n9123 ;
  assign n9130 = ~n4233 & ~n9124 ;
  assign n9131 = ~n9129 & ~n9130 ;
  assign n9132 = n933 & ~n9131 ;
  assign n9133 = ~n604 & n3946 ;
  assign n9134 = ~n9122 & ~n9133 ;
  assign n9135 = n965 & ~n9134 ;
  assign n9125 = n1867 & ~n9124 ;
  assign n9136 = \InstQueue_reg[8][1]/NET0131  & ~n3929 ;
  assign n9137 = ~n9125 & ~n9136 ;
  assign n9138 = ~n9135 & n9137 ;
  assign n9139 = ~n9132 & n9138 ;
  assign n9145 = n4181 & n8796 ;
  assign n9146 = n3944 & n8799 ;
  assign n9147 = ~n9145 & ~n9146 ;
  assign n9148 = \DataWidth_reg[1]/NET0131  & ~n9147 ;
  assign n9140 = \Datai[1]_pad  & ~n3974 ;
  assign n9141 = \InstQueue_reg[9][1]/NET0131  & ~n3937 ;
  assign n9142 = ~n3946 & n9141 ;
  assign n9143 = ~n9140 & ~n9142 ;
  assign n9149 = ~n4253 & ~n9143 ;
  assign n9150 = ~n9148 & ~n9149 ;
  assign n9151 = n933 & ~n9150 ;
  assign n9152 = ~n604 & n3937 ;
  assign n9153 = ~n9141 & ~n9152 ;
  assign n9154 = n965 & ~n9153 ;
  assign n9144 = n1867 & ~n9143 ;
  assign n9155 = \InstQueue_reg[9][1]/NET0131  & ~n3929 ;
  assign n9156 = ~n9144 & ~n9155 ;
  assign n9157 = ~n9154 & n9156 ;
  assign n9158 = ~n9151 & n9157 ;
  assign n9165 = ~\rEIP_reg[26]/NET0131  & ~n8552 ;
  assign n9166 = n825 & ~n8553 ;
  assign n9167 = ~n9165 & n9166 ;
  assign n9159 = \Address[24]_pad  & ~n824 ;
  assign n9160 = \rEIP_reg[24]/NET0131  & n8526 ;
  assign n9161 = ~\rEIP_reg[25]/NET0131  & ~n9160 ;
  assign n9162 = n5933 & n8525 ;
  assign n9163 = n8524 & ~n9162 ;
  assign n9164 = ~n9161 & n9163 ;
  assign n9168 = ~n9159 & ~n9164 ;
  assign n9169 = ~n9167 & n9168 ;
  assign n9175 = ~\rEIP_reg[14]/NET0131  & ~n8546 ;
  assign n9176 = n825 & ~n8547 ;
  assign n9177 = ~n9175 & n9176 ;
  assign n9170 = \Address[12]_pad  & ~n824 ;
  assign n9172 = ~n6544 & n8525 ;
  assign n9171 = ~\rEIP_reg[13]/NET0131  & ~n8525 ;
  assign n9173 = n8524 & ~n9171 ;
  assign n9174 = ~n9172 & n9173 ;
  assign n9178 = ~n9170 & ~n9174 ;
  assign n9179 = ~n9177 & n9178 ;
  assign n9181 = n5743 & n8624 ;
  assign n9182 = \rEIP_reg[21]/NET0131  & n9181 ;
  assign n9183 = ~\rEIP_reg[22]/NET0131  & ~n9182 ;
  assign n9184 = n825 & ~n8550 ;
  assign n9185 = ~n9183 & n9184 ;
  assign n9180 = \Address[20]_pad  & ~n824 ;
  assign n9186 = n5744 & n8525 ;
  assign n9188 = \rEIP_reg[21]/NET0131  & n9186 ;
  assign n9187 = ~\rEIP_reg[21]/NET0131  & ~n9186 ;
  assign n9189 = n8524 & ~n9187 ;
  assign n9190 = ~n9188 & n9189 ;
  assign n9191 = ~n9180 & ~n9190 ;
  assign n9192 = ~n9185 & n9191 ;
  assign n9198 = ~\rEIP_reg[10]/NET0131  & ~n8543 ;
  assign n9199 = n825 & ~n8544 ;
  assign n9200 = ~n9198 & n9199 ;
  assign n9193 = \Address[8]_pad  & ~n824 ;
  assign n9195 = ~n6398 & n8525 ;
  assign n9194 = ~\rEIP_reg[9]/NET0131  & ~n8525 ;
  assign n9196 = n8524 & ~n9194 ;
  assign n9197 = ~n9195 & n9196 ;
  assign n9201 = ~n9193 & ~n9197 ;
  assign n9202 = ~n9200 & n9201 ;
  assign n9208 = n3871 & n8838 ;
  assign n9209 = n3914 & n8841 ;
  assign n9210 = ~n9208 & ~n9209 ;
  assign n9211 = \DataWidth_reg[1]/NET0131  & ~n9210 ;
  assign n9203 = \Datai[0]_pad  & ~n3863 ;
  assign n9204 = \InstQueue_reg[0][0]/NET0131  & ~n3859 ;
  assign n9205 = ~n3862 & n9204 ;
  assign n9206 = ~n9203 & ~n9205 ;
  assign n9212 = ~n3919 & ~n9206 ;
  assign n9213 = ~n9211 & ~n9212 ;
  assign n9214 = n933 & ~n9213 ;
  assign n9215 = ~n508 & n3859 ;
  assign n9216 = ~n9204 & ~n9215 ;
  assign n9217 = n965 & ~n9216 ;
  assign n9207 = n1867 & ~n9206 ;
  assign n9218 = \InstQueue_reg[0][0]/NET0131  & ~n3929 ;
  assign n9219 = ~n9207 & ~n9218 ;
  assign n9220 = ~n9217 & n9219 ;
  assign n9221 = ~n9214 & n9220 ;
  assign n9227 = n3946 & n8841 ;
  assign n9228 = n3944 & n8838 ;
  assign n9229 = ~n9227 & ~n9228 ;
  assign n9230 = \DataWidth_reg[1]/NET0131  & ~n9229 ;
  assign n9222 = \Datai[0]_pad  & ~n3938 ;
  assign n9223 = \InstQueue_reg[10][0]/NET0131  & ~n3935 ;
  assign n9224 = ~n3937 & n9223 ;
  assign n9225 = ~n9222 & ~n9224 ;
  assign n9231 = ~n3951 & ~n9225 ;
  assign n9232 = ~n9230 & ~n9231 ;
  assign n9233 = n933 & ~n9232 ;
  assign n9234 = ~n508 & n3935 ;
  assign n9235 = ~n9223 & ~n9234 ;
  assign n9236 = n965 & ~n9235 ;
  assign n9226 = n1867 & ~n9225 ;
  assign n9237 = \InstQueue_reg[10][0]/NET0131  & ~n3929 ;
  assign n9238 = ~n9226 & ~n9237 ;
  assign n9239 = ~n9236 & n9238 ;
  assign n9240 = ~n9233 & n9239 ;
  assign n9246 = n3937 & n8838 ;
  assign n9247 = n3935 & n8841 ;
  assign n9248 = ~n9246 & ~n9247 ;
  assign n9249 = \DataWidth_reg[1]/NET0131  & ~n9248 ;
  assign n9241 = \Datai[0]_pad  & ~n3988 ;
  assign n9242 = \InstQueue_reg[12][0]/NET0131  & ~n3987 ;
  assign n9243 = ~n3963 & n9242 ;
  assign n9244 = ~n9241 & ~n9243 ;
  assign n9250 = ~n3998 & ~n9244 ;
  assign n9251 = ~n9249 & ~n9250 ;
  assign n9252 = n933 & ~n9251 ;
  assign n9253 = ~n508 & n3987 ;
  assign n9254 = ~n9242 & ~n9253 ;
  assign n9255 = n965 & ~n9254 ;
  assign n9245 = n1867 & ~n9244 ;
  assign n9256 = \InstQueue_reg[12][0]/NET0131  & ~n3929 ;
  assign n9257 = ~n9245 & ~n9256 ;
  assign n9258 = ~n9255 & n9257 ;
  assign n9259 = ~n9252 & n9258 ;
  assign n9265 = n3935 & n8838 ;
  assign n9266 = n3963 & n8841 ;
  assign n9267 = ~n9265 & ~n9266 ;
  assign n9268 = \DataWidth_reg[1]/NET0131  & ~n9267 ;
  assign n9260 = \Datai[0]_pad  & ~n4009 ;
  assign n9261 = \InstQueue_reg[13][0]/NET0131  & ~n3871 ;
  assign n9262 = ~n3987 & n9261 ;
  assign n9263 = ~n9260 & ~n9262 ;
  assign n9269 = ~n4019 & ~n9263 ;
  assign n9270 = ~n9268 & ~n9269 ;
  assign n9271 = n933 & ~n9270 ;
  assign n9272 = ~n508 & n3871 ;
  assign n9273 = ~n9261 & ~n9272 ;
  assign n9274 = n965 & ~n9273 ;
  assign n9264 = n1867 & ~n9263 ;
  assign n9275 = \InstQueue_reg[13][0]/NET0131  & ~n3929 ;
  assign n9276 = ~n9264 & ~n9275 ;
  assign n9277 = ~n9274 & n9276 ;
  assign n9278 = ~n9271 & n9277 ;
  assign n9284 = n3963 & n8838 ;
  assign n9285 = n3987 & n8841 ;
  assign n9286 = ~n9284 & ~n9285 ;
  assign n9287 = \DataWidth_reg[1]/NET0131  & ~n9286 ;
  assign n9279 = \Datai[0]_pad  & ~n3918 ;
  assign n9280 = \InstQueue_reg[14][0]/NET0131  & ~n3914 ;
  assign n9281 = ~n3871 & n9280 ;
  assign n9282 = ~n9279 & ~n9281 ;
  assign n9288 = ~n4039 & ~n9282 ;
  assign n9289 = ~n9287 & ~n9288 ;
  assign n9290 = n933 & ~n9289 ;
  assign n9291 = ~n508 & n3914 ;
  assign n9292 = ~n9280 & ~n9291 ;
  assign n9293 = n965 & ~n9292 ;
  assign n9283 = n1867 & ~n9282 ;
  assign n9294 = \InstQueue_reg[14][0]/NET0131  & ~n3929 ;
  assign n9295 = ~n9283 & ~n9294 ;
  assign n9296 = ~n9293 & n9295 ;
  assign n9297 = ~n9290 & n9296 ;
  assign n9303 = n3987 & n8838 ;
  assign n9304 = n3871 & n8841 ;
  assign n9305 = ~n9303 & ~n9304 ;
  assign n9306 = \DataWidth_reg[1]/NET0131  & ~n9305 ;
  assign n9298 = \Datai[0]_pad  & ~n4050 ;
  assign n9299 = \InstQueue_reg[15][0]/NET0131  & ~n3862 ;
  assign n9300 = ~n3914 & n9299 ;
  assign n9301 = ~n9298 & ~n9300 ;
  assign n9307 = ~n4060 & ~n9301 ;
  assign n9308 = ~n9306 & ~n9307 ;
  assign n9309 = n933 & ~n9308 ;
  assign n9310 = ~n508 & n3862 ;
  assign n9311 = ~n9299 & ~n9310 ;
  assign n9312 = n965 & ~n9311 ;
  assign n9302 = n1867 & ~n9301 ;
  assign n9313 = \InstQueue_reg[15][0]/NET0131  & ~n3929 ;
  assign n9314 = ~n9302 & ~n9313 ;
  assign n9315 = ~n9312 & n9314 ;
  assign n9316 = ~n9309 & n9315 ;
  assign n9322 = n3914 & n8838 ;
  assign n9323 = n3862 & n8841 ;
  assign n9324 = ~n9322 & ~n9323 ;
  assign n9325 = \DataWidth_reg[1]/NET0131  & ~n9324 ;
  assign n9317 = \Datai[0]_pad  & ~n4072 ;
  assign n9318 = \InstQueue_reg[1][0]/NET0131  & ~n4071 ;
  assign n9319 = ~n3859 & n9318 ;
  assign n9320 = ~n9317 & ~n9319 ;
  assign n9326 = ~n4082 & ~n9320 ;
  assign n9327 = ~n9325 & ~n9326 ;
  assign n9328 = n933 & ~n9327 ;
  assign n9329 = ~n508 & n4071 ;
  assign n9330 = ~n9318 & ~n9329 ;
  assign n9331 = n965 & ~n9330 ;
  assign n9321 = n1867 & ~n9320 ;
  assign n9332 = \InstQueue_reg[1][0]/NET0131  & ~n3929 ;
  assign n9333 = ~n9321 & ~n9332 ;
  assign n9334 = ~n9331 & n9333 ;
  assign n9335 = ~n9328 & n9334 ;
  assign n9341 = n3859 & n8841 ;
  assign n9342 = n3862 & n8838 ;
  assign n9343 = ~n9341 & ~n9342 ;
  assign n9344 = \DataWidth_reg[1]/NET0131  & ~n9343 ;
  assign n9336 = \Datai[0]_pad  & ~n4094 ;
  assign n9337 = \InstQueue_reg[2][0]/NET0131  & ~n4093 ;
  assign n9338 = ~n4071 & n9337 ;
  assign n9339 = ~n9336 & ~n9338 ;
  assign n9345 = ~n4104 & ~n9339 ;
  assign n9346 = ~n9344 & ~n9345 ;
  assign n9347 = n933 & ~n9346 ;
  assign n9348 = ~n508 & n4093 ;
  assign n9349 = ~n9337 & ~n9348 ;
  assign n9350 = n965 & ~n9349 ;
  assign n9340 = n1867 & ~n9339 ;
  assign n9351 = \InstQueue_reg[2][0]/NET0131  & ~n3929 ;
  assign n9352 = ~n9340 & ~n9351 ;
  assign n9353 = ~n9350 & n9352 ;
  assign n9354 = ~n9347 & n9353 ;
  assign n9360 = n4071 & n8838 ;
  assign n9361 = n4093 & n8841 ;
  assign n9362 = ~n9360 & ~n9361 ;
  assign n9363 = \DataWidth_reg[1]/NET0131  & ~n9362 ;
  assign n9355 = \Datai[0]_pad  & ~n4138 ;
  assign n9356 = \InstQueue_reg[4][0]/NET0131  & ~n4137 ;
  assign n9357 = ~n4115 & n9356 ;
  assign n9358 = ~n9355 & ~n9357 ;
  assign n9364 = ~n4148 & ~n9358 ;
  assign n9365 = ~n9363 & ~n9364 ;
  assign n9366 = n933 & ~n9365 ;
  assign n9367 = ~n508 & n4137 ;
  assign n9368 = ~n9356 & ~n9367 ;
  assign n9369 = n965 & ~n9368 ;
  assign n9359 = n1867 & ~n9358 ;
  assign n9370 = \InstQueue_reg[4][0]/NET0131  & ~n3929 ;
  assign n9371 = ~n9359 & ~n9370 ;
  assign n9372 = ~n9369 & n9371 ;
  assign n9373 = ~n9366 & n9372 ;
  assign n9379 = n4093 & n8838 ;
  assign n9380 = n4115 & n8841 ;
  assign n9381 = ~n9379 & ~n9380 ;
  assign n9382 = \DataWidth_reg[1]/NET0131  & ~n9381 ;
  assign n9374 = \Datai[0]_pad  & ~n4160 ;
  assign n9375 = \InstQueue_reg[5][0]/NET0131  & ~n4159 ;
  assign n9376 = ~n4137 & n9375 ;
  assign n9377 = ~n9374 & ~n9376 ;
  assign n9383 = ~n4170 & ~n9377 ;
  assign n9384 = ~n9382 & ~n9383 ;
  assign n9385 = n933 & ~n9384 ;
  assign n9386 = ~n508 & n4159 ;
  assign n9387 = ~n9375 & ~n9386 ;
  assign n9388 = n965 & ~n9387 ;
  assign n9378 = n1867 & ~n9377 ;
  assign n9389 = \InstQueue_reg[5][0]/NET0131  & ~n3929 ;
  assign n9390 = ~n9378 & ~n9389 ;
  assign n9391 = ~n9388 & n9390 ;
  assign n9392 = ~n9385 & n9391 ;
  assign n9398 = n4115 & n8838 ;
  assign n9399 = n4137 & n8841 ;
  assign n9400 = ~n9398 & ~n9399 ;
  assign n9401 = \DataWidth_reg[1]/NET0131  & ~n9400 ;
  assign n9393 = \Datai[0]_pad  & ~n4182 ;
  assign n9394 = \InstQueue_reg[6][0]/NET0131  & ~n4181 ;
  assign n9395 = ~n4159 & n9394 ;
  assign n9396 = ~n9393 & ~n9395 ;
  assign n9402 = ~n4192 & ~n9396 ;
  assign n9403 = ~n9401 & ~n9402 ;
  assign n9404 = n933 & ~n9403 ;
  assign n9405 = ~n508 & n4181 ;
  assign n9406 = ~n9394 & ~n9405 ;
  assign n9407 = n965 & ~n9406 ;
  assign n9397 = n1867 & ~n9396 ;
  assign n9408 = \InstQueue_reg[6][0]/NET0131  & ~n3929 ;
  assign n9409 = ~n9397 & ~n9408 ;
  assign n9410 = ~n9407 & n9409 ;
  assign n9411 = ~n9404 & n9410 ;
  assign n9417 = n4159 & n8838 ;
  assign n9418 = n4181 & n8841 ;
  assign n9419 = ~n9417 & ~n9418 ;
  assign n9420 = \DataWidth_reg[1]/NET0131  & ~n9419 ;
  assign n9412 = \Datai[0]_pad  & ~n3950 ;
  assign n9413 = \InstQueue_reg[8][0]/NET0131  & ~n3946 ;
  assign n9414 = ~n3944 & n9413 ;
  assign n9415 = ~n9412 & ~n9414 ;
  assign n9421 = ~n4233 & ~n9415 ;
  assign n9422 = ~n9420 & ~n9421 ;
  assign n9423 = n933 & ~n9422 ;
  assign n9424 = ~n508 & n3946 ;
  assign n9425 = ~n9413 & ~n9424 ;
  assign n9426 = n965 & ~n9425 ;
  assign n9416 = n1867 & ~n9415 ;
  assign n9427 = \InstQueue_reg[8][0]/NET0131  & ~n3929 ;
  assign n9428 = ~n9416 & ~n9427 ;
  assign n9429 = ~n9426 & n9428 ;
  assign n9430 = ~n9423 & n9429 ;
  assign n9436 = n4181 & n8838 ;
  assign n9437 = n3944 & n8841 ;
  assign n9438 = ~n9436 & ~n9437 ;
  assign n9439 = \DataWidth_reg[1]/NET0131  & ~n9438 ;
  assign n9431 = \Datai[0]_pad  & ~n3974 ;
  assign n9432 = \InstQueue_reg[9][0]/NET0131  & ~n3937 ;
  assign n9433 = ~n3946 & n9432 ;
  assign n9434 = ~n9431 & ~n9433 ;
  assign n9440 = ~n4253 & ~n9434 ;
  assign n9441 = ~n9439 & ~n9440 ;
  assign n9442 = n933 & ~n9441 ;
  assign n9443 = ~n508 & n3937 ;
  assign n9444 = ~n9432 & ~n9443 ;
  assign n9445 = n965 & ~n9444 ;
  assign n9435 = n1867 & ~n9434 ;
  assign n9446 = \InstQueue_reg[9][0]/NET0131  & ~n3929 ;
  assign n9447 = ~n9435 & ~n9446 ;
  assign n9448 = ~n9445 & n9447 ;
  assign n9449 = ~n9442 & n9448 ;
  assign n9455 = ~\rEIP_reg[6]/NET0131  & ~n8539 ;
  assign n9456 = n825 & ~n8540 ;
  assign n9457 = ~n9455 & n9456 ;
  assign n9450 = \Address[4]_pad  & ~n824 ;
  assign n9452 = ~n6265 & n8525 ;
  assign n9451 = ~\rEIP_reg[5]/NET0131  & ~n8525 ;
  assign n9453 = n8524 & ~n9451 ;
  assign n9454 = ~n9452 & n9453 ;
  assign n9458 = ~n9450 & ~n9454 ;
  assign n9459 = ~n9457 & n9458 ;
  assign n9464 = ~\rEIP_reg[29]/NET0131  & ~n8555 ;
  assign n9465 = n825 & ~n8556 ;
  assign n9466 = ~n9464 & n9465 ;
  assign n9460 = \Address[27]_pad  & ~n824 ;
  assign n9461 = ~\rEIP_reg[28]/NET0131  & ~n8528 ;
  assign n9462 = n8524 & ~n8529 ;
  assign n9463 = ~n9461 & n9462 ;
  assign n9467 = ~n9460 & ~n9463 ;
  assign n9468 = ~n9466 & n9467 ;
  assign n9474 = ~\rEIP_reg[17]/NET0131  & ~n8549 ;
  assign n9475 = n825 & ~n8625 ;
  assign n9476 = ~n9474 & n9475 ;
  assign n9469 = \Address[15]_pad  & ~n824 ;
  assign n9470 = n5737 & n8525 ;
  assign n9471 = ~\rEIP_reg[16]/NET0131  & ~n9470 ;
  assign n9472 = n8524 & ~n8619 ;
  assign n9473 = ~n9471 & n9472 ;
  assign n9477 = ~n9469 & ~n9473 ;
  assign n9478 = ~n9476 & n9477 ;
  assign n9483 = \rEIP_reg[24]/NET0131  & n8551 ;
  assign n9484 = ~\rEIP_reg[25]/NET0131  & ~n9483 ;
  assign n9485 = n825 & ~n8552 ;
  assign n9486 = ~n9484 & n9485 ;
  assign n9479 = \Address[23]_pad  & ~n824 ;
  assign n9480 = ~\rEIP_reg[24]/NET0131  & ~n8526 ;
  assign n9481 = n8524 & ~n9160 ;
  assign n9482 = ~n9480 & n9481 ;
  assign n9487 = ~n9479 & ~n9482 ;
  assign n9488 = ~n9486 & n9487 ;
  assign n9494 = \rEIP_reg[12]/NET0131  & n8545 ;
  assign n9495 = ~\rEIP_reg[13]/NET0131  & ~n9494 ;
  assign n9496 = n825 & ~n8546 ;
  assign n9497 = ~n9495 & n9496 ;
  assign n9489 = \Address[11]_pad  & ~n824 ;
  assign n9491 = ~n6508 & n8525 ;
  assign n9490 = ~\rEIP_reg[12]/NET0131  & ~n8525 ;
  assign n9492 = n8524 & ~n9490 ;
  assign n9493 = ~n9491 & n9492 ;
  assign n9498 = ~n9489 & ~n9493 ;
  assign n9499 = ~n9497 & n9498 ;
  assign n9508 = ~\rEIP_reg[5]/NET0131  & ~n8538 ;
  assign n9509 = n825 & ~n8539 ;
  assign n9510 = ~n9508 & n9509 ;
  assign n9500 = \Address[3]_pad  & ~n824 ;
  assign n9501 = \rEIP_reg[1]/NET0131  & n8525 ;
  assign n9502 = \rEIP_reg[2]/NET0131  & n9501 ;
  assign n9503 = \rEIP_reg[3]/NET0131  & n9502 ;
  assign n9505 = \rEIP_reg[4]/NET0131  & n9503 ;
  assign n9504 = ~\rEIP_reg[4]/NET0131  & ~n9503 ;
  assign n9506 = n8524 & ~n9504 ;
  assign n9507 = ~n9505 & n9506 ;
  assign n9511 = ~n9500 & ~n9507 ;
  assign n9512 = ~n9510 & n9511 ;
  assign n9518 = ~\rEIP_reg[21]/NET0131  & ~n9181 ;
  assign n9519 = n825 & ~n9182 ;
  assign n9520 = ~n9518 & n9519 ;
  assign n9513 = \Address[19]_pad  & ~n824 ;
  assign n9514 = n5741 & n8525 ;
  assign n9515 = ~\rEIP_reg[20]/NET0131  & ~n9514 ;
  assign n9516 = n8524 & ~n9186 ;
  assign n9517 = ~n9515 & n9516 ;
  assign n9521 = ~n9513 & ~n9517 ;
  assign n9522 = ~n9520 & n9521 ;
  assign n9528 = ~\rEIP_reg[9]/NET0131  & ~n8542 ;
  assign n9529 = n825 & ~n8543 ;
  assign n9530 = ~n9528 & n9529 ;
  assign n9523 = \Address[7]_pad  & ~n824 ;
  assign n9525 = ~n6361 & n8525 ;
  assign n9524 = ~\rEIP_reg[8]/NET0131  & ~n8525 ;
  assign n9526 = n8524 & ~n9524 ;
  assign n9527 = ~n9525 & n9526 ;
  assign n9531 = ~n9523 & ~n9527 ;
  assign n9532 = ~n9530 & n9531 ;
  assign n9540 = ~\rEIP_reg[16]/NET0131  & ~n8548 ;
  assign n9541 = n825 & ~n8549 ;
  assign n9542 = ~n9540 & n9541 ;
  assign n9533 = \Address[14]_pad  & ~n824 ;
  assign n9534 = n5732 & n8525 ;
  assign n9535 = \rEIP_reg[11]/NET0131  & n9534 ;
  assign n9536 = n5735 & n9535 ;
  assign n9537 = ~\rEIP_reg[15]/NET0131  & ~n9536 ;
  assign n9538 = n8524 & ~n9470 ;
  assign n9539 = ~n9537 & n9538 ;
  assign n9543 = ~n9533 & ~n9539 ;
  assign n9544 = ~n9542 & n9543 ;
  assign n9549 = ~\rEIP_reg[28]/NET0131  & ~n8554 ;
  assign n9550 = n825 & ~n8555 ;
  assign n9551 = ~n9549 & n9550 ;
  assign n9545 = \Address[26]_pad  & ~n824 ;
  assign n9546 = ~\rEIP_reg[27]/NET0131  & ~n8527 ;
  assign n9547 = n8524 & ~n8528 ;
  assign n9548 = ~n9546 & n9547 ;
  assign n9552 = ~n9545 & ~n9548 ;
  assign n9553 = ~n9551 & n9552 ;
  assign n9559 = ~\rEIP_reg[24]/NET0131  & ~n8551 ;
  assign n9560 = n825 & ~n9483 ;
  assign n9561 = ~n9559 & n9560 ;
  assign n9554 = \Address[22]_pad  & ~n824 ;
  assign n9555 = n5832 & n8525 ;
  assign n9556 = ~\rEIP_reg[23]/NET0131  & ~n9555 ;
  assign n9557 = n8524 & ~n8526 ;
  assign n9558 = ~n9556 & n9557 ;
  assign n9562 = ~n9554 & ~n9558 ;
  assign n9563 = ~n9561 & n9562 ;
  assign n9568 = ~\rEIP_reg[12]/NET0131  & ~n8545 ;
  assign n9569 = n825 & ~n9494 ;
  assign n9570 = ~n9568 & n9569 ;
  assign n9564 = \Address[10]_pad  & ~n824 ;
  assign n9565 = ~\rEIP_reg[11]/NET0131  & ~n9534 ;
  assign n9566 = n8524 & ~n9535 ;
  assign n9567 = ~n9565 & n9566 ;
  assign n9571 = ~n9564 & ~n9567 ;
  assign n9572 = ~n9570 & n9571 ;
  assign n9577 = ~\rEIP_reg[4]/NET0131  & ~n8537 ;
  assign n9578 = n825 & ~n8538 ;
  assign n9579 = ~n9577 & n9578 ;
  assign n9573 = \Address[2]_pad  & ~n824 ;
  assign n9574 = ~\rEIP_reg[3]/NET0131  & ~n9502 ;
  assign n9575 = n8524 & ~n9503 ;
  assign n9576 = ~n9574 & n9575 ;
  assign n9580 = ~n9573 & ~n9576 ;
  assign n9581 = ~n9579 & n9580 ;
  assign n9587 = \rEIP_reg[19]/NET0131  & n8624 ;
  assign n9588 = ~\rEIP_reg[20]/NET0131  & ~n9587 ;
  assign n9589 = n825 & ~n9181 ;
  assign n9590 = ~n9588 & n9589 ;
  assign n9582 = \Address[18]_pad  & ~n824 ;
  assign n9583 = n5739 & n8619 ;
  assign n9584 = ~\rEIP_reg[19]/NET0131  & ~n9583 ;
  assign n9585 = n8524 & ~n9514 ;
  assign n9586 = ~n9584 & n9585 ;
  assign n9591 = ~n9582 & ~n9586 ;
  assign n9592 = ~n9590 & n9591 ;
  assign n9598 = ~\rEIP_reg[8]/NET0131  & ~n8541 ;
  assign n9599 = n825 & ~n8542 ;
  assign n9600 = ~n9598 & n9599 ;
  assign n9593 = \Address[6]_pad  & ~n824 ;
  assign n9595 = ~n6328 & n8525 ;
  assign n9594 = ~\rEIP_reg[7]/NET0131  & ~n8525 ;
  assign n9596 = n8524 & ~n9594 ;
  assign n9597 = ~n9595 & n9596 ;
  assign n9601 = ~n9593 & ~n9597 ;
  assign n9602 = ~n9600 & n9601 ;
  assign n9607 = ~\rEIP_reg[27]/NET0131  & ~n8553 ;
  assign n9608 = n825 & ~n8554 ;
  assign n9609 = ~n9607 & n9608 ;
  assign n9603 = \Address[25]_pad  & ~n824 ;
  assign n9604 = ~\rEIP_reg[26]/NET0131  & ~n9162 ;
  assign n9605 = n8524 & ~n8527 ;
  assign n9606 = ~n9604 & n9605 ;
  assign n9610 = ~n9603 & ~n9606 ;
  assign n9611 = ~n9609 & n9610 ;
  assign n9620 = \rEIP_reg[31]/NET0131  & n8558 ;
  assign n9619 = ~\rEIP_reg[31]/NET0131  & ~n8558 ;
  assign n9621 = n825 & ~n9619 ;
  assign n9622 = ~n9620 & n9621 ;
  assign n9612 = \Address[29]_pad  & ~n824 ;
  assign n9614 = ~\rEIP_reg[30]/NET0131  & ~n6074 ;
  assign n9615 = ~n6152 & ~n9614 ;
  assign n9616 = n8525 & ~n9615 ;
  assign n9613 = ~\rEIP_reg[30]/NET0131  & ~n8525 ;
  assign n9617 = n8524 & ~n9613 ;
  assign n9618 = ~n9616 & n9617 ;
  assign n9623 = ~n9612 & ~n9618 ;
  assign n9624 = ~n9622 & n9623 ;
  assign n9630 = ~\rEIP_reg[15]/NET0131  & ~n8547 ;
  assign n9631 = n825 & ~n8548 ;
  assign n9632 = ~n9630 & n9631 ;
  assign n9625 = \Address[13]_pad  & ~n824 ;
  assign n9627 = ~n6579 & n8525 ;
  assign n9626 = ~\rEIP_reg[14]/NET0131  & ~n8525 ;
  assign n9628 = n8524 & ~n9626 ;
  assign n9629 = ~n9627 & n9628 ;
  assign n9633 = ~n9625 & ~n9629 ;
  assign n9634 = ~n9632 & n9633 ;
  assign n9640 = ~\rEIP_reg[11]/NET0131  & ~n8544 ;
  assign n9641 = n825 & ~n8545 ;
  assign n9642 = ~n9640 & n9641 ;
  assign n9635 = \Address[9]_pad  & ~n824 ;
  assign n9637 = ~n6437 & n8525 ;
  assign n9636 = ~\rEIP_reg[10]/NET0131  & ~n8525 ;
  assign n9638 = n8524 & ~n9636 ;
  assign n9639 = ~n9637 & n9638 ;
  assign n9643 = ~n9635 & ~n9639 ;
  assign n9644 = ~n9642 & n9643 ;
  assign n9650 = ~\rEIP_reg[23]/NET0131  & ~n8550 ;
  assign n9651 = n825 & ~n8551 ;
  assign n9652 = ~n9650 & n9651 ;
  assign n9646 = ~n5833 & n8525 ;
  assign n9645 = ~\rEIP_reg[22]/NET0131  & ~n8525 ;
  assign n9647 = n8524 & ~n9645 ;
  assign n9648 = ~n9646 & n9647 ;
  assign n9649 = \Address[21]_pad  & ~n824 ;
  assign n9653 = ~n9648 & ~n9649 ;
  assign n9654 = ~n9652 & n9653 ;
  assign n9655 = \DataWidth_reg[0]/NET0131  & \DataWidth_reg[1]/NET0131  ;
  assign n9656 = \ByteEnable_reg[2]/NET0131  & n9655 ;
  assign n9657 = ~\DataWidth_reg[1]/NET0131  & \rEIP_reg[1]/NET0131  ;
  assign n9658 = \DataWidth_reg[0]/NET0131  & ~n9657 ;
  assign n9659 = \rEIP_reg[0]/NET0131  & ~n9658 ;
  assign n9660 = ~n8534 & ~n9659 ;
  assign n9661 = ~n5692 & ~n9660 ;
  assign n9662 = ~n9656 & ~n9661 ;
  assign n9666 = ~HOLD_pad & \State_reg[0]/NET0131  ;
  assign n9667 = ~\State_reg[2]/NET0131  & ~n9666 ;
  assign n9668 = ~READY_n_pad & ~n9667 ;
  assign n9669 = \State_reg[1]/NET0131  & ~n9668 ;
  assign n9663 = HOLD_pad & \State_reg[2]/NET0131  ;
  assign n9664 = \RequestPending_reg/NET0131  & \State_reg[0]/NET0131  ;
  assign n9665 = ~n9663 & n9664 ;
  assign n9670 = ~n827 & ~n9665 ;
  assign n9671 = ~n9669 & n9670 ;
  assign n9674 = ~\DataWidth_reg[0]/NET0131  & ~\DataWidth_reg[1]/NET0131  ;
  assign n9675 = ~\rEIP_reg[0]/NET0131  & n9674 ;
  assign n9672 = \ByteEnable_reg[1]/NET0131  & n9655 ;
  assign n9673 = \rEIP_reg[1]/NET0131  & ~n9655 ;
  assign n9676 = ~n9672 & ~n9673 ;
  assign n9677 = ~n9675 & n9676 ;
  assign n9678 = ~READY_n_pad & \State_reg[0]/NET0131  ;
  assign n9679 = NA_n_pad & ~\State_reg[0]/NET0131  ;
  assign n9680 = \State_reg[2]/NET0131  & ~n9679 ;
  assign n9681 = ~n9678 & ~n9680 ;
  assign n9682 = ~HOLD_pad & ~n9681 ;
  assign n9683 = \State_reg[0]/NET0131  & ~\State_reg[1]/NET0131  ;
  assign n9684 = ~\State_reg[2]/NET0131  & n9683 ;
  assign n9685 = ~n9682 & ~n9684 ;
  assign n9686 = \RequestPending_reg/NET0131  & ~n9685 ;
  assign n9687 = ~n8524 & ~n9686 ;
  assign n9692 = ~\rEIP_reg[3]/NET0131  & ~n8536 ;
  assign n9693 = n825 & ~n8537 ;
  assign n9694 = ~n9692 & n9693 ;
  assign n9688 = \Address[1]_pad  & ~n824 ;
  assign n9689 = ~\rEIP_reg[2]/NET0131  & ~n9501 ;
  assign n9690 = n8524 & ~n9502 ;
  assign n9691 = ~n9689 & n9690 ;
  assign n9695 = ~n9688 & ~n9691 ;
  assign n9696 = ~n9694 & n9695 ;
  assign n9701 = ~\rEIP_reg[19]/NET0131  & ~n8624 ;
  assign n9702 = n825 & ~n9587 ;
  assign n9703 = ~n9701 & n9702 ;
  assign n9697 = \Address[17]_pad  & ~n824 ;
  assign n9698 = ~\rEIP_reg[18]/NET0131  & ~n8621 ;
  assign n9699 = n8524 & ~n9583 ;
  assign n9700 = ~n9698 & n9699 ;
  assign n9704 = ~n9697 & ~n9700 ;
  assign n9705 = ~n9703 & n9704 ;
  assign n9711 = ~\rEIP_reg[7]/NET0131  & ~n8540 ;
  assign n9712 = n825 & ~n8541 ;
  assign n9713 = ~n9711 & n9712 ;
  assign n9706 = \Address[5]_pad  & ~n824 ;
  assign n9708 = ~n6295 & n8525 ;
  assign n9707 = ~\rEIP_reg[6]/NET0131  & ~n8525 ;
  assign n9709 = n8524 & ~n9707 ;
  assign n9710 = ~n9708 & n9709 ;
  assign n9714 = ~n9706 & ~n9710 ;
  assign n9715 = ~n9713 & n9714 ;
  assign n9716 = \State_reg[0]/NET0131  & \State_reg[1]/NET0131  ;
  assign n9717 = ~\State_reg[2]/NET0131  & n9716 ;
  assign n9718 = ~HOLD_pad & ~\RequestPending_reg/NET0131  ;
  assign n9719 = READY_n_pad & ~n9718 ;
  assign n9720 = n9717 & n9719 ;
  assign n9721 = ~n827 & ~n9720 ;
  assign n9722 = ~NA_n_pad & ~n9721 ;
  assign n9723 = ~\RequestPending_reg/NET0131  & ~\State_reg[1]/NET0131  ;
  assign n9724 = ~\State_reg[2]/NET0131  & ~n9723 ;
  assign n9725 = HOLD_pad & \State_reg[0]/NET0131  ;
  assign n9726 = ~n9724 & n9725 ;
  assign n9727 = \State_reg[1]/NET0131  & \State_reg[2]/NET0131  ;
  assign n9728 = ~n9678 & n9727 ;
  assign n9729 = ~n9726 & ~n9728 ;
  assign n9730 = ~n9722 & n9729 ;
  assign n9731 = \ByteEnable_reg[3]/NET0131  & n9655 ;
  assign n9732 = \rEIP_reg[1]/NET0131  & ~n9675 ;
  assign n9733 = ~\DataWidth_reg[1]/NET0131  & ~n9732 ;
  assign n9734 = ~n9731 & ~n9733 ;
  assign n9739 = ~\rEIP_reg[2]/NET0131  & ~n8535 ;
  assign n9740 = n825 & ~n8536 ;
  assign n9741 = ~n9739 & n9740 ;
  assign n9735 = \Address[0]_pad  & ~n824 ;
  assign n9736 = ~\rEIP_reg[1]/NET0131  & ~n8525 ;
  assign n9737 = n8524 & ~n9501 ;
  assign n9738 = ~n9736 & n9737 ;
  assign n9742 = ~n9735 & ~n9738 ;
  assign n9743 = ~n9741 & n9742 ;
  assign n9744 = ~n827 & ~n9717 ;
  assign n9745 = ~\BS16_n_pad  & ~n9744 ;
  assign n9746 = ~n826 & ~n9717 ;
  assign n9747 = ~\DataWidth_reg[1]/NET0131  & n9746 ;
  assign n9748 = ~n9745 & ~n9747 ;
  assign n9749 = \BE_n[2]_pad  & ~n824 ;
  assign n9750 = \ByteEnable_reg[2]/NET0131  & n824 ;
  assign n9751 = ~n9749 & ~n9750 ;
  assign n9752 = ADS_n_pad & \State_reg[0]/NET0131  ;
  assign n9753 = n9746 & ~n9752 ;
  assign n9754 = \BE_n[0]_pad  & ~n824 ;
  assign n9755 = \ByteEnable_reg[0]/NET0131  & n824 ;
  assign n9756 = ~n9754 & ~n9755 ;
  assign n9757 = \BE_n[1]_pad  & ~n824 ;
  assign n9758 = \ByteEnable_reg[1]/NET0131  & n824 ;
  assign n9759 = ~n9757 & ~n9758 ;
  assign n9760 = \BE_n[3]_pad  & ~n824 ;
  assign n9761 = \ByteEnable_reg[3]/NET0131  & n824 ;
  assign n9762 = ~n9760 & ~n9761 ;
  assign n9763 = M_IO_n_pad & ~n824 ;
  assign n9764 = \MemoryFetch_reg/NET0131  & n824 ;
  assign n9765 = ~n9763 & ~n9764 ;
  assign n9766 = W_R_n_pad & ~n824 ;
  assign n9767 = ~\ReadRequest_reg/NET0131  & n824 ;
  assign n9768 = ~n9766 & ~n9767 ;
  assign n9769 = ~\State_reg[1]/NET0131  & \State_reg[2]/NET0131  ;
  assign n9770 = ~\State_reg[0]/NET0131  & ~n9769 ;
  assign n9771 = ~D_C_n_pad & ~n9770 ;
  assign n9772 = \CodeFetch_reg/NET0131  & n824 ;
  assign n9773 = ~n9771 & ~n9772 ;
  assign n9774 = \DataWidth_reg[0]/NET0131  & n9746 ;
  assign n9775 = ~n9745 & ~n9774 ;
  assign n9776 = \InstAddrPointer_reg[28]/NET0131  & n906 ;
  assign n9777 = ~n2335 & ~n9776 ;
  assign n9778 = n773 & ~n9777 ;
  assign n9780 = ~\InstAddrPointer_reg[28]/NET0131  & ~n765 ;
  assign n9781 = ~n740 & ~n9780 ;
  assign n9782 = n2340 & n9781 ;
  assign n9784 = ~n811 & n1391 ;
  assign n9779 = \InstAddrPointer_reg[28]/NET0131  & ~n1644 ;
  assign n9783 = ~n873 & n2322 ;
  assign n9785 = ~n9779 & ~n9783 ;
  assign n9786 = ~n9784 & n9785 ;
  assign n9787 = ~n9782 & n9786 ;
  assign n9788 = ~n2351 & n9787 ;
  assign n9789 = ~n9778 & n9788 ;
  assign n9790 = n929 & ~n9789 ;
  assign n9791 = \InstAddrPointer_reg[28]/NET0131  & n1661 ;
  assign n9792 = ~n2361 & ~n9791 ;
  assign n9793 = ~n9790 & n9792 ;
  assign n9795 = \PhyAddrPointer_reg[12]/NET0131  & n906 ;
  assign n9799 = ~n1460 & ~n2150 ;
  assign n9800 = ~n2151 & ~n9799 ;
  assign n9801 = n1014 & ~n9800 ;
  assign n9796 = n1312 & ~n2116 ;
  assign n9797 = ~n1014 & ~n2156 ;
  assign n9798 = ~n9796 & n9797 ;
  assign n9802 = ~n906 & ~n9798 ;
  assign n9803 = ~n9801 & n9802 ;
  assign n9804 = ~n9795 & ~n9803 ;
  assign n9805 = n773 & ~n9804 ;
  assign n9806 = \PhyAddrPointer_reg[12]/NET0131  & ~n1852 ;
  assign n9807 = \InstAddrPointer_reg[11]/NET0131  & n2170 ;
  assign n9809 = n1593 & n9807 ;
  assign n9808 = ~n1593 & ~n9807 ;
  assign n9810 = n899 & ~n9808 ;
  assign n9811 = ~n9809 & n9810 ;
  assign n9812 = ~n9806 & ~n9811 ;
  assign n9813 = ~n9805 & n9812 ;
  assign n9814 = n929 & ~n9813 ;
  assign n9818 = ~\DataWidth_reg[1]/NET0131  & ~n6494 ;
  assign n9815 = ~\PhyAddrPointer_reg[12]/NET0131  & ~n2465 ;
  assign n9816 = ~n2674 & ~n9815 ;
  assign n9817 = \DataWidth_reg[1]/NET0131  & ~n9816 ;
  assign n9819 = n933 & ~n9817 ;
  assign n9820 = ~n9818 & n9819 ;
  assign n9822 = n1867 & n6494 ;
  assign n9794 = \PhyAddrPointer_reg[12]/NET0131  & ~n1902 ;
  assign n9821 = \rEIP_reg[12]/NET0131  & n1655 ;
  assign n9823 = ~n9794 & ~n9821 ;
  assign n9824 = ~n9822 & n9823 ;
  assign n9825 = ~n9820 & n9824 ;
  assign n9826 = ~n9814 & n9825 ;
  assign n9828 = \InstAddrPointer_reg[17]/NET0131  & n906 ;
  assign n9829 = ~n2737 & ~n9828 ;
  assign n9830 = n773 & ~n9829 ;
  assign n9832 = \InstAddrPointer_reg[17]/NET0131  & ~n1816 ;
  assign n9831 = ~n873 & n2729 ;
  assign n9833 = n766 & n1586 ;
  assign n9834 = ~n811 & n1354 ;
  assign n9835 = ~n9833 & ~n9834 ;
  assign n9836 = ~n9831 & n9835 ;
  assign n9837 = ~n9832 & n9836 ;
  assign n9838 = ~n2744 & n9837 ;
  assign n9839 = ~n9830 & n9838 ;
  assign n9840 = n929 & ~n9839 ;
  assign n9827 = \InstAddrPointer_reg[17]/NET0131  & n1661 ;
  assign n9841 = ~n2755 & ~n9827 ;
  assign n9842 = ~n9840 & n9841 ;
  assign n9844 = \InstAddrPointer_reg[19]/NET0131  & n906 ;
  assign n9845 = ~n2522 & ~n9844 ;
  assign n9846 = n773 & ~n9845 ;
  assign n9848 = ~n836 & n1465 ;
  assign n9849 = n2216 & ~n9848 ;
  assign n9850 = \InstAddrPointer_reg[19]/NET0131  & ~n9849 ;
  assign n9852 = ~n873 & n1465 ;
  assign n9847 = n766 & n1619 ;
  assign n9851 = ~n811 & n1351 ;
  assign n9853 = ~n9847 & ~n9851 ;
  assign n9854 = ~n9852 & n9853 ;
  assign n9855 = ~n9850 & n9854 ;
  assign n9856 = ~n2529 & n9855 ;
  assign n9857 = ~n9846 & n9856 ;
  assign n9858 = n929 & ~n9857 ;
  assign n9843 = \InstAddrPointer_reg[19]/NET0131  & n1661 ;
  assign n9859 = ~n2505 & ~n9843 ;
  assign n9860 = ~n9858 & n9859 ;
  assign n9862 = \InstAddrPointer_reg[16]/NET0131  & n906 ;
  assign n9863 = ~n2699 & ~n9862 ;
  assign n9864 = n773 & ~n9863 ;
  assign n9865 = ~n873 & n2690 ;
  assign n9867 = \InstAddrPointer_reg[16]/NET0131  & ~n2073 ;
  assign n9861 = ~n811 & n1345 ;
  assign n9866 = n766 & n1799 ;
  assign n9868 = ~n9861 & ~n9866 ;
  assign n9869 = ~n9867 & n9868 ;
  assign n9870 = ~n9865 & n9869 ;
  assign n9871 = ~n2705 & n9870 ;
  assign n9872 = ~n9864 & n9871 ;
  assign n9873 = n929 & ~n9872 ;
  assign n9874 = \InstAddrPointer_reg[16]/NET0131  & n1661 ;
  assign n9875 = ~n2718 & ~n9874 ;
  assign n9876 = ~n9873 & n9875 ;
  assign n9878 = \InstAddrPointer_reg[20]/NET0131  & n906 ;
  assign n9882 = n1358 & n2695 ;
  assign n9884 = ~n1338 & n9882 ;
  assign n9883 = n1338 & ~n9882 ;
  assign n9885 = ~n1014 & ~n9883 ;
  assign n9886 = ~n9884 & n9885 ;
  assign n9879 = ~n1456 & ~n2015 ;
  assign n9880 = ~n1482 & ~n9879 ;
  assign n9881 = n1014 & ~n9880 ;
  assign n9887 = ~n906 & ~n9881 ;
  assign n9888 = ~n9886 & n9887 ;
  assign n9889 = ~n9878 & ~n9888 ;
  assign n9890 = n773 & ~n9889 ;
  assign n9891 = ~n2341 & ~n2343 ;
  assign n9892 = n899 & ~n2037 ;
  assign n9893 = ~n9891 & n9892 ;
  assign n9894 = ~READY_n_pad & ~n1456 ;
  assign n9895 = n840 & ~n9894 ;
  assign n9896 = ~n911 & ~n9895 ;
  assign n9897 = ~n862 & n9896 ;
  assign n9898 = \InstAddrPointer_reg[20]/NET0131  & ~n9897 ;
  assign n9877 = ~n811 & n1338 ;
  assign n9904 = ~\InstAddrPointer_reg[20]/NET0131  & READY_n_pad ;
  assign n9905 = ~n9894 & ~n9904 ;
  assign n9906 = ~n858 & n9905 ;
  assign n9899 = n788 & n1456 ;
  assign n9901 = n765 & ~n2343 ;
  assign n9900 = ~\InstAddrPointer_reg[20]/NET0131  & ~n765 ;
  assign n9902 = ~n740 & ~n9900 ;
  assign n9903 = ~n9901 & n9902 ;
  assign n9907 = ~n9899 & ~n9903 ;
  assign n9908 = ~n9906 & n9907 ;
  assign n9909 = ~n9877 & n9908 ;
  assign n9910 = ~n9898 & n9909 ;
  assign n9911 = ~n9893 & n9910 ;
  assign n9912 = ~n9890 & n9911 ;
  assign n9913 = n929 & ~n9912 ;
  assign n9914 = \rEIP_reg[20]/NET0131  & n1655 ;
  assign n9915 = \InstAddrPointer_reg[20]/NET0131  & n1661 ;
  assign n9916 = ~n9914 & ~n9915 ;
  assign n9917 = ~n9913 & n9916 ;
  assign n9919 = \InstAddrPointer_reg[18]/NET0131  & n906 ;
  assign n9920 = ~n2769 & ~n9919 ;
  assign n9921 = n773 & ~n9920 ;
  assign n9922 = \InstAddrPointer_reg[18]/NET0131  & ~n1816 ;
  assign n9923 = ~n873 & n1467 ;
  assign n9924 = n766 & n1608 ;
  assign n9925 = ~n811 & n1356 ;
  assign n9926 = ~n9924 & ~n9925 ;
  assign n9927 = ~n9923 & n9926 ;
  assign n9928 = ~n9922 & n9927 ;
  assign n9929 = ~n2775 & n9928 ;
  assign n9930 = ~n9921 & n9929 ;
  assign n9931 = n929 & ~n9930 ;
  assign n9918 = \InstAddrPointer_reg[18]/NET0131  & n1661 ;
  assign n9932 = ~n2785 & ~n9918 ;
  assign n9933 = ~n9931 & n9932 ;
  assign n9934 = \InstAddrPointer_reg[31]/NET0131  & n906 ;
  assign n9935 = ~n1849 & ~n9934 ;
  assign n9936 = n773 & ~n9935 ;
  assign n9941 = n766 & n1858 ;
  assign n9937 = ~n811 & n1843 ;
  assign n9938 = ~n836 & ~n1514 ;
  assign n9939 = n2216 & ~n9938 ;
  assign n9940 = \InstAddrPointer_reg[31]/NET0131  & ~n9939 ;
  assign n9942 = ~n873 & n1834 ;
  assign n9943 = ~n9940 & ~n9942 ;
  assign n9944 = ~n9937 & n9943 ;
  assign n9945 = ~n9941 & n9944 ;
  assign n9946 = ~n1862 & n9945 ;
  assign n9947 = ~n9936 & n9946 ;
  assign n9948 = n929 & ~n9947 ;
  assign n9949 = \InstAddrPointer_reg[31]/NET0131  & n1661 ;
  assign n9950 = ~n1866 & ~n9949 ;
  assign n9951 = ~n9948 & n9950 ;
  assign n9954 = \InstAddrPointer_reg[23]/NET0131  & n906 ;
  assign n9955 = ~n2283 & ~n9954 ;
  assign n9956 = n773 & ~n9955 ;
  assign n9958 = ~READY_n_pad & ~n1502 ;
  assign n9959 = ~\InstAddrPointer_reg[23]/NET0131  & READY_n_pad ;
  assign n9960 = ~n9958 & ~n9959 ;
  assign n9961 = ~n836 & n9960 ;
  assign n9962 = n1957 & ~n9961 ;
  assign n9963 = \InstAddrPointer_reg[23]/NET0131  & ~n9962 ;
  assign n9953 = n766 & n1807 ;
  assign n9964 = n788 & n1502 ;
  assign n9966 = ~n9953 & ~n9964 ;
  assign n9957 = ~n811 & n1368 ;
  assign n9965 = ~n858 & n9960 ;
  assign n9967 = ~n9957 & ~n9965 ;
  assign n9968 = n9966 & n9967 ;
  assign n9969 = ~n9963 & n9968 ;
  assign n9970 = ~n2289 & n9969 ;
  assign n9971 = ~n9956 & n9970 ;
  assign n9972 = n929 & ~n9971 ;
  assign n9952 = \InstAddrPointer_reg[23]/NET0131  & n1661 ;
  assign n9973 = ~n2272 & ~n9952 ;
  assign n9974 = ~n9972 & n9973 ;
  assign n9977 = \InstAddrPointer_reg[12]/NET0131  & n906 ;
  assign n9978 = ~n9803 & ~n9977 ;
  assign n9979 = n773 & ~n9978 ;
  assign n9980 = ~READY_n_pad & ~n1460 ;
  assign n9981 = ~\InstAddrPointer_reg[12]/NET0131  & READY_n_pad ;
  assign n9982 = ~n9980 & ~n9981 ;
  assign n9983 = ~n836 & n9982 ;
  assign n9984 = n1957 & ~n9983 ;
  assign n9985 = \InstAddrPointer_reg[12]/NET0131  & ~n9984 ;
  assign n9976 = ~n811 & n1312 ;
  assign n9986 = ~n858 & n9982 ;
  assign n9987 = n766 & n1593 ;
  assign n9988 = n788 & n1460 ;
  assign n9989 = ~n9987 & ~n9988 ;
  assign n9990 = ~n9986 & n9989 ;
  assign n9991 = ~n9976 & n9990 ;
  assign n9992 = ~n9985 & n9991 ;
  assign n9993 = ~n9811 & n9992 ;
  assign n9994 = ~n9979 & n9993 ;
  assign n9995 = n929 & ~n9994 ;
  assign n9975 = \InstAddrPointer_reg[12]/NET0131  & n1661 ;
  assign n9996 = ~n9821 & ~n9975 ;
  assign n9997 = ~n9995 & n9996 ;
  assign n9998 = \PhyAddrPointer_reg[20]/NET0131  & n906 ;
  assign n9999 = ~n9888 & ~n9998 ;
  assign n10000 = n773 & ~n9999 ;
  assign n10001 = \PhyAddrPointer_reg[20]/NET0131  & ~n1852 ;
  assign n10002 = ~n9893 & ~n10001 ;
  assign n10003 = ~n10000 & n10002 ;
  assign n10004 = n929 & ~n10003 ;
  assign n10008 = n2100 & n5705 ;
  assign n10005 = ~\PhyAddrPointer_reg[20]/NET0131  & ~n2508 ;
  assign n10006 = n969 & ~n2816 ;
  assign n10007 = ~n10005 & n10006 ;
  assign n10009 = \PhyAddrPointer_reg[20]/NET0131  & ~n1902 ;
  assign n10010 = ~n9914 & ~n10009 ;
  assign n10011 = ~n10007 & n10010 ;
  assign n10012 = ~n10008 & n10011 ;
  assign n10013 = ~n10004 & n10012 ;
  assign n10016 = \InstAddrPointer_reg[10]/NET0131  & n906 ;
  assign n10017 = ~n3205 & ~n10016 ;
  assign n10018 = n773 & ~n10017 ;
  assign n10019 = ~n873 & n1772 ;
  assign n10020 = \InstAddrPointer_reg[10]/NET0131  & ~n2073 ;
  assign n10015 = ~n811 & n1316 ;
  assign n10021 = n766 & n3210 ;
  assign n10022 = ~n10015 & ~n10021 ;
  assign n10023 = ~n10020 & n10022 ;
  assign n10024 = ~n10019 & n10023 ;
  assign n10025 = ~n3213 & n10024 ;
  assign n10026 = ~n10018 & n10025 ;
  assign n10027 = n929 & ~n10026 ;
  assign n10014 = \InstAddrPointer_reg[10]/NET0131  & n1661 ;
  assign n10028 = ~n3223 & ~n10014 ;
  assign n10029 = ~n10027 & n10028 ;
  assign n10047 = ~n1899 & ~n6169 ;
  assign n10049 = n2097 & ~n10047 ;
  assign n10048 = ~n2097 & n10047 ;
  assign n10050 = ~\DataWidth_reg[1]/NET0131  & ~n10048 ;
  assign n10051 = ~n10049 & n10050 ;
  assign n10046 = \DataWidth_reg[1]/NET0131  & ~\rEIP_reg[30]/NET0131  ;
  assign n10052 = n933 & ~n10046 ;
  assign n10053 = ~n10051 & n10052 ;
  assign n10032 = \EBX_reg[31]/NET0131  & ~n6148 ;
  assign n10033 = \EBX_reg[30]/NET0131  & ~n10032 ;
  assign n10031 = ~n6148 & n6149 ;
  assign n10034 = ~n5676 & ~n10031 ;
  assign n10035 = ~n10033 & n10034 ;
  assign n10030 = n5676 & ~n9615 ;
  assign n10036 = n3660 & ~n10030 ;
  assign n10037 = ~n10035 & n10036 ;
  assign n10038 = \rEIP_reg[30]/NET0131  & ~n5684 ;
  assign n10040 = n924 & ~n9615 ;
  assign n10039 = ~\EBX_reg[30]/NET0131  & ~n924 ;
  assign n10041 = n923 & ~n10039 ;
  assign n10042 = ~n10040 & n10041 ;
  assign n10043 = ~n10038 & ~n10042 ;
  assign n10044 = ~n10037 & n10043 ;
  assign n10045 = n929 & ~n10044 ;
  assign n10054 = \PhyAddrPointer_reg[30]/NET0131  & n953 ;
  assign n10055 = \rEIP_reg[30]/NET0131  & ~n5667 ;
  assign n10056 = ~n10054 & ~n10055 ;
  assign n10057 = ~n10045 & n10056 ;
  assign n10058 = ~n10053 & n10057 ;
  assign n10061 = \InstAddrPointer_reg[21]/NET0131  & n906 ;
  assign n10062 = ~n2799 & ~n10061 ;
  assign n10063 = n773 & ~n10062 ;
  assign n10064 = ~READY_n_pad & ~n1485 ;
  assign n10065 = ~\InstAddrPointer_reg[21]/NET0131  & READY_n_pad ;
  assign n10066 = ~n10064 & ~n10065 ;
  assign n10070 = ~n836 & n10066 ;
  assign n10071 = n1957 & ~n10070 ;
  assign n10072 = \InstAddrPointer_reg[21]/NET0131  & ~n10071 ;
  assign n10069 = ~n811 & n1335 ;
  assign n10068 = n766 & n1612 ;
  assign n10060 = n788 & n1485 ;
  assign n10067 = ~n858 & n10066 ;
  assign n10073 = ~n10060 & ~n10067 ;
  assign n10074 = ~n10068 & n10073 ;
  assign n10075 = ~n10069 & n10074 ;
  assign n10076 = ~n10072 & n10075 ;
  assign n10077 = ~n2806 & n10076 ;
  assign n10078 = ~n10063 & n10077 ;
  assign n10079 = n929 & ~n10078 ;
  assign n10059 = \InstAddrPointer_reg[21]/NET0131  & n1661 ;
  assign n10080 = ~n2814 & ~n10059 ;
  assign n10081 = ~n10079 & n10080 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g47406/_2_  = ~n946 ;
  assign \g47407/_2_  = ~n964 ;
  assign \g47411/_0_  = ~n966 ;
  assign \g47413/_0_  = ~n972 ;
  assign \g47424/_0_  = ~n1664 ;
  assign \g47434/_0_  = ~n1748 ;
  assign \g47437/_0_  = ~n1830 ;
  assign \g47447/_2_  = ~n1916 ;
  assign \g47448/_0_  = ~n1947 ;
  assign \g47451/_0_  = ~n1992 ;
  assign \g47452/_0_  = ~n2050 ;
  assign \g47453/_0_  = ~n2087 ;
  assign \g47465/_2_  = ~n2109 ;
  assign \g47466/_0_  = ~n2146 ;
  assign \g47467/_0_  = ~n2191 ;
  assign \g47471/_0_  = ~n2231 ;
  assign \g47485/_0_  = ~n2259 ;
  assign \g47486/_0_  = ~n2296 ;
  assign \g47487/_2_  = ~n2318 ;
  assign \g47488/_0_  = ~n2366 ;
  assign \g47489/_2_  = ~n2385 ;
  assign \g47491/_0_  = ~n2417 ;
  assign \g47494/_0_  = ~n2457 ;
  assign \g47510/_0_  = ~n2477 ;
  assign \g47511/_0_  = ~n2498 ;
  assign \g47512/_0_  = ~n2536 ;
  assign \g47515/_0_  = ~n2557 ;
  assign \g47516/_0_  = ~n2576 ;
  assign \g47517/_2_  = ~n2595 ;
  assign \g47524/_0_  = ~n2635 ;
  assign \g47525/_0_  = ~n2665 ;
  assign \g47550/_0_  = ~n2685 ;
  assign \g47551/_2_  = ~n2722 ;
  assign \g47552/_0_  = ~n2759 ;
  assign \g47554/_0_  = ~n2789 ;
  assign \g47555/_0_  = ~n2824 ;
  assign \g47556/_0_  = ~n2845 ;
  assign \g47558/_0_  = ~n2863 ;
  assign \g47563/_0_  = ~n2901 ;
  assign \g47564/_0_  = ~n2936 ;
  assign \g47565/_0_  = ~n3183 ;
  assign \g47584/_0_  = ~n3195 ;
  assign \g47592/_0_  = ~n3228 ;
  assign \g47597/_0_  = ~n3248 ;
  assign \g47598/_0_  = ~n3266 ;
  assign \g47601/_0_  = ~n3302 ;
  assign \g47602/_0_  = ~n3329 ;
  assign \g47603/_0_  = ~n3449 ;
  assign \g47604/_0_  = ~n3462 ;
  assign \g47606/_0_  = ~n3506 ;
  assign \g47630/_0_  = ~n3518 ;
  assign \g47636/_0_  = ~n3539 ;
  assign \g47641/_0_  = ~n3570 ;
  assign \g47642/_0_  = ~n3592 ;
  assign \g47643/_0_  = ~n3621 ;
  assign \g47644/_0_  = ~n3631 ;
  assign \g47645/_0_  = ~n3651 ;
  assign \g47646/_0_  = ~n3695 ;
  assign \g47648/_0_  = ~n3707 ;
  assign \g47679/_0_  = ~n3727 ;
  assign \g47680/_0_  = ~n3745 ;
  assign \g47681/_0_  = ~n3766 ;
  assign \g47683/_0_  = ~n3775 ;
  assign \g47687/_0_  = ~n3797 ;
  assign \g47690/_0_  = ~n3808 ;
  assign \g47746/_0_  = ~n3824 ;
  assign \g47747/_0_  = ~n3837 ;
  assign \g47754/_0_  = ~n3846 ;
  assign \g47756/_0_  = ~n3856 ;
  assign \g47804/_0_  = ~n3933 ;
  assign \g47805/_0_  = ~n3961 ;
  assign \g47806/_0_  = ~n3985 ;
  assign \g47807/_0_  = ~n4008 ;
  assign \g47809/_0_  = ~n4029 ;
  assign \g47810/_0_  = ~n4049 ;
  assign \g47812/_0_  = ~n4070 ;
  assign \g47813/_0_  = ~n4092 ;
  assign \g47814/_0_  = ~n4114 ;
  assign \g47815/_0_  = ~n4136 ;
  assign \g47816/_0_  = ~n4158 ;
  assign \g47817/_0_  = ~n4180 ;
  assign \g47818/_0_  = ~n4202 ;
  assign \g47819/_0_  = ~n4223 ;
  assign \g47820/_0_  = ~n4243 ;
  assign \g47821/_0_  = ~n4263 ;
  assign \g47836/_0_  = ~n4279 ;
  assign \g47848/_0_  = ~n4295 ;
  assign \g47851/_0_  = ~n4305 ;
  assign \g47852/_0_  = ~n4326 ;
  assign \g47943/_0_  = ~n4353 ;
  assign \g47944/_0_  = ~n4372 ;
  assign \g47945/_0_  = ~n4391 ;
  assign \g47946/_0_  = ~n4410 ;
  assign \g47947/_0_  = ~n4429 ;
  assign \g47949/_0_  = ~n4448 ;
  assign \g47950/_0_  = ~n4467 ;
  assign \g47952/_0_  = ~n4486 ;
  assign \g47953/_0_  = ~n4505 ;
  assign \g47954/_0_  = ~n4524 ;
  assign \g47955/_0_  = ~n4543 ;
  assign \g47956/_0_  = ~n4562 ;
  assign \g47957/_0_  = ~n4581 ;
  assign \g47958/_0_  = ~n4600 ;
  assign \g47959/_0_  = ~n4619 ;
  assign \g47960/_0_  = ~n4638 ;
  assign \g47999/_0_  = ~n4650 ;
  assign \g48/_0_  = ~n4660 ;
  assign \g48005/_0_  = ~n4669 ;
  assign \g48006/_0_  = ~n4682 ;
  assign \g48007/_0_  = ~n4723 ;
  assign \g48008/_0_  = ~n4764 ;
  assign \g48009/_0_  = ~n4807 ;
  assign \g48010/_0_  = ~n4849 ;
  assign \g48011/_0_  = ~n4861 ;
  assign \g48012/_0_  = ~n4907 ;
  assign \g48013/_0_  = ~n4951 ;
  assign \g48014/_0_  = ~n4994 ;
  assign \g48015/_0_  = ~n5038 ;
  assign \g48057/_0_  = ~n5061 ;
  assign \g48058/_0_  = ~n5084 ;
  assign \g48059/_0_  = ~n5103 ;
  assign \g48060/_0_  = ~n5122 ;
  assign \g48061/_0_  = ~n5141 ;
  assign \g48062/_0_  = ~n5160 ;
  assign \g48063/_0_  = ~n5179 ;
  assign \g48064/_0_  = ~n5198 ;
  assign \g48066/_0_  = ~n5217 ;
  assign \g48067/_0_  = ~n5236 ;
  assign \g48068/_0_  = ~n5255 ;
  assign \g48069/_0_  = ~n5274 ;
  assign \g48070/_0_  = ~n5293 ;
  assign \g48071/_0_  = ~n5312 ;
  assign \g48073/_0_  = ~n5331 ;
  assign \g48074/_0_  = ~n5350 ;
  assign \g48075/_0_  = ~n5369 ;
  assign \g48076/_0_  = ~n5388 ;
  assign \g48077/_0_  = ~n5407 ;
  assign \g48078/_0_  = ~n5426 ;
  assign \g48079/_0_  = ~n5445 ;
  assign \g48080/_0_  = ~n5464 ;
  assign \g48081/_0_  = ~n5483 ;
  assign \g48082/_0_  = ~n5502 ;
  assign \g48084/_0_  = ~n5521 ;
  assign \g48085/_0_  = ~n5540 ;
  assign \g48086/_0_  = ~n5559 ;
  assign \g48087/_0_  = ~n5578 ;
  assign \g48089/_0_  = ~n5597 ;
  assign \g48090/_0_  = ~n5616 ;
  assign \g48091/_0_  = ~n5635 ;
  assign \g48093/_0_  = ~n5654 ;
  assign \g48094/_0_  = ~n5665 ;
  assign \g48119/_0_  = ~n5702 ;
  assign \g48120/_0_  = ~n5782 ;
  assign \g48121/_0_  = ~n5817 ;
  assign \g48122/_0_  = ~n5854 ;
  assign \g48123/_0_  = ~n5889 ;
  assign \g48124/_0_  = ~n5928 ;
  assign \g48125/_0_  = ~n5966 ;
  assign \g48126/_0_  = ~n6004 ;
  assign \g48127/_0_  = ~n6038 ;
  assign \g48128/_0_  = ~n6072 ;
  assign \g48129/_0_  = ~n6110 ;
  assign \g48130/_0_  = ~n6145 ;
  assign \g48131/_0_  = ~n6179 ;
  assign \g48132/_0_  = ~n6214 ;
  assign \g48133/_0_  = ~n6247 ;
  assign \g48134/_0_  = ~n6281 ;
  assign \g48135/_0_  = ~n6314 ;
  assign \g48136/_0_  = ~n6348 ;
  assign \g48137/_0_  = ~n6380 ;
  assign \g48138/_0_  = ~n6414 ;
  assign \g48140/_0_  = ~n6423 ;
  assign \g48144/_0_  = ~n6457 ;
  assign \g48145/_0_  = ~n6491 ;
  assign \g48146/_0_  = ~n6529 ;
  assign \g48147/_0_  = ~n6564 ;
  assign \g48148/_0_  = ~n6599 ;
  assign \g48150/_0_  = ~n6633 ;
  assign \g48151/_0_  = ~n6668 ;
  assign \g48152/_0_  = ~n6705 ;
  assign \g48153/_0_  = ~n6739 ;
  assign \g48154/_0_  = ~n6772 ;
  assign \g48176/_0_  = ~n6785 ;
  assign \g48189/_0_  = ~n6799 ;
  assign \g48192/_0_  = ~n6813 ;
  assign \g48193/_0_  = ~n6824 ;
  assign \g48194/_0_  = ~n6834 ;
  assign \g48195/_0_  = ~n6843 ;
  assign \g48196/_0_  = ~n6853 ;
  assign \g48197/_0_  = ~n6863 ;
  assign \g48198/_0_  = ~n6874 ;
  assign \g48199/_0_  = ~n6884 ;
  assign \g48200/_0_  = ~n6898 ;
  assign \g48263/_0_  = ~n6904 ;
  assign \g48265/_0_  = ~n6910 ;
  assign \g48273/_0_  = ~n6929 ;
  assign \g48313/_0_  = ~n6945 ;
  assign \g48318/_0_  = ~n6965 ;
  assign \g48319/_0_  = ~n6973 ;
  assign \g48321/_0_  = ~n6980 ;
  assign \g48323/_0_  = ~n6990 ;
  assign \g48324/_0_  = ~n7040 ;
  assign \g48325/_0_  = ~n7089 ;
  assign \g48326/_0_  = ~n7138 ;
  assign \g48327/_0_  = ~n7188 ;
  assign \g48328/_0_  = ~n7191 ;
  assign \g48329/_0_  = ~n7241 ;
  assign \g48330/_0_  = ~n7290 ;
  assign \g48331/_0_  = ~n7337 ;
  assign \g48332/_0_  = ~n7358 ;
  assign \g48333/_0_  = ~n7379 ;
  assign \g48472/_0_  = ~n7390 ;
  assign \g48519/_0_  = ~n7402 ;
  assign \g48520/_0_  = ~n7408 ;
  assign \g48521/_0_  = ~n7420 ;
  assign \g48522/_0_  = ~n7432 ;
  assign \g48523/_0_  = ~n7444 ;
  assign \g48524/_0_  = ~n7457 ;
  assign \g48525/_0_  = ~n7465 ;
  assign \g48527/_0_  = ~n7475 ;
  assign \g48529/_0_  = ~n7485 ;
  assign \g48530/_0_  = ~n7495 ;
  assign \g48531/_0_  = ~n7505 ;
  assign \g48532/_0_  = ~n7515 ;
  assign \g48533/_0_  = ~n7525 ;
  assign \g48534/_0_  = ~n7535 ;
  assign \g48535/_0_  = ~n7545 ;
  assign \g48536/_0_  = ~n7555 ;
  assign \g48537/_0_  = ~n7565 ;
  assign \g48538/_0_  = ~n7575 ;
  assign \g48539/_0_  = ~n7586 ;
  assign \g48540/_0_  = ~n7597 ;
  assign \g48541/_0_  = ~n7608 ;
  assign \g48542/_0_  = ~n7618 ;
  assign \g48543/_0_  = ~n7627 ;
  assign \g48545/_0_  = ~n7637 ;
  assign \g48546/_0_  = ~n7647 ;
  assign \g48547/_0_  = ~n7650 ;
  assign \g48639/_0_  = ~n7673 ;
  assign \g48642/_0_  = ~n7692 ;
  assign \g48645/_0_  = ~n7711 ;
  assign \g48648/_0_  = ~n7730 ;
  assign \g48652/_0_  = ~n7749 ;
  assign \g48655/_0_  = ~n7768 ;
  assign \g48658/_0_  = ~n7787 ;
  assign \g48661/_0_  = ~n7806 ;
  assign \g48664/_0_  = ~n7825 ;
  assign \g48667/_0_  = ~n7844 ;
  assign \g48670/_0_  = ~n7863 ;
  assign \g48673/_0_  = ~n7882 ;
  assign \g48678/_0_  = ~n7901 ;
  assign \g48681/_0_  = ~n7920 ;
  assign \g48684/_0_  = ~n7939 ;
  assign \g48688/_0_  = ~n7958 ;
  assign \g48793/_0_  = ~n7966 ;
  assign \g48812/_0_  = ~n7972 ;
  assign \g48813/_0_  = ~n7980 ;
  assign \g48814/_0_  = ~n7991 ;
  assign \g48824/_0_  = ~n7999 ;
  assign \g48825/_0_  = ~n8011 ;
  assign \g48826/_0_  = ~n8021 ;
  assign \g48827/_0_  = ~n8031 ;
  assign \g48828/_0_  = ~n8041 ;
  assign \g48829/_0_  = ~n8051 ;
  assign \g48830/_0_  = ~n8061 ;
  assign \g48831/_0_  = ~n8071 ;
  assign \g48833/_0_  = ~n8081 ;
  assign \g48834/_0_  = ~n8087 ;
  assign \g48835/_0_  = ~n8097 ;
  assign \g48836/_0_  = ~n8102 ;
  assign \g48837/_0_  = ~n8112 ;
  assign \g48838/_0_  = ~n8117 ;
  assign \g48839/_0_  = ~n8127 ;
  assign \g48840/_0_  = ~n8137 ;
  assign \g48841/_0_  = ~n8147 ;
  assign \g48842/_0_  = ~n8157 ;
  assign \g48843/_0_  = ~n8167 ;
  assign \g48844/_0_  = ~n8177 ;
  assign \g48845/_0_  = ~n8188 ;
  assign \g48846/_0_  = ~n8198 ;
  assign \g48847/_0_  = ~n8204 ;
  assign \g48848/_0_  = ~n8214 ;
  assign \g48908/_0_  = ~n8237 ;
  assign \g48909/_0_  = ~n8256 ;
  assign \g48910/_0_  = ~n8275 ;
  assign \g48912/_0_  = ~n8294 ;
  assign \g48913/_0_  = ~n8313 ;
  assign \g48915/_0_  = ~n8332 ;
  assign \g48917/_0_  = ~n8351 ;
  assign \g48932/_0_  = ~n8370 ;
  assign \g48933/_0_  = ~n8389 ;
  assign \g48935/_0_  = ~n8408 ;
  assign \g48937/_0_  = ~n8427 ;
  assign \g48938/_0_  = ~n8446 ;
  assign \g48939/_0_  = ~n8465 ;
  assign \g48940/_0_  = ~n8484 ;
  assign \g48942/_0_  = ~n8503 ;
  assign \g48945/_0_  = ~n8522 ;
  assign \g48971/_0_  = ~n8562 ;
  assign \g49007/_0_  = ~n8573 ;
  assign \g49047/_0_  = ~n8581 ;
  assign \g49048/_0_  = ~n8592 ;
  assign \g49050/_0_  = ~n8600 ;
  assign \g49182/_0_  = ~n8617 ;
  assign \g49280/_0_  = ~n8630 ;
  assign \g49332/_0_  = ~n8638 ;
  assign \g49335/_0_  = ~n8646 ;
  assign \g49336/_0_  = ~n8654 ;
  assign \g49337/_0_  = ~n8662 ;
  assign \g49338/_0_  = ~n8670 ;
  assign \g49339/_0_  = ~n8678 ;
  assign \g49340/_0_  = ~n8686 ;
  assign \g49341/_0_  = ~n8694 ;
  assign \g49342/_0_  = ~n8702 ;
  assign \g49343/_0_  = ~n8710 ;
  assign \g49344/_0_  = ~n8718 ;
  assign \g49345/_0_  = ~n8726 ;
  assign \g49346/_0_  = ~n8734 ;
  assign \g49347/_0_  = ~n8742 ;
  assign \g49348/_0_  = ~n8750 ;
  assign \g49349/_0_  = ~n8758 ;
  assign \g49356/_0_  = ~n8773 ;
  assign \g49375/_0_  = ~n8783 ;
  assign \g49396/_0_  = ~n8789 ;
  assign \g49397/_0_  = ~n8812 ;
  assign \g49400/_0_  = ~n8831 ;
  assign \g49404/_0_  = ~n8854 ;
  assign \g49406/_0_  = ~n8873 ;
  assign \g49414/_0_  = ~n8892 ;
  assign \g49422/_0_  = ~n8911 ;
  assign \g49426/_0_  = ~n8930 ;
  assign \g49430/_0_  = ~n8949 ;
  assign \g49434/_0_  = ~n8968 ;
  assign \g49437/_0_  = ~n8987 ;
  assign \g49440/_0_  = ~n9006 ;
  assign \g49441/_0_  = ~n9025 ;
  assign \g49444/_0_  = ~n9044 ;
  assign \g49448/_0_  = ~n9063 ;
  assign \g49451/_0_  = ~n9082 ;
  assign \g49455/_0_  = ~n9101 ;
  assign \g49456/_0_  = ~n9120 ;
  assign \g49460/_0_  = ~n9139 ;
  assign \g49466/_0_  = ~n9158 ;
  assign \g49563/_0_  = ~n9169 ;
  assign \g49592/_0_  = ~n9179 ;
  assign \g49915/_0_  = ~n9192 ;
  assign \g49941/_0_  = ~n9202 ;
  assign \g50023/_0_  = ~n9221 ;
  assign \g50026/_0_  = ~n9240 ;
  assign \g50029/_0_  = ~n9259 ;
  assign \g50031/_0_  = ~n9278 ;
  assign \g50033/_0_  = ~n9297 ;
  assign \g50035/_0_  = ~n9316 ;
  assign \g50037/_0_  = ~n9335 ;
  assign \g50040/_0_  = ~n9354 ;
  assign \g50050/_0_  = ~n9373 ;
  assign \g50056/_0_  = ~n9392 ;
  assign \g50059/_0_  = ~n9411 ;
  assign \g50065/_0_  = ~n9430 ;
  assign \g50067/_0_  = ~n9449 ;
  assign \g50150/_0_  = ~n9459 ;
  assign \g50283/_0_  = ~n9468 ;
  assign \g50284/_0_  = ~n9478 ;
  assign \g50501/_0_  = ~n9488 ;
  assign \g50594/_0_  = ~n9499 ;
  assign \g50807/_0_  = ~n9512 ;
  assign \g50866/_0_  = ~n9522 ;
  assign \g50875/_0_  = ~n9532 ;
  assign \g51449/_0_  = ~n9544 ;
  assign \g51510/_0_  = ~n9553 ;
  assign \g51534/_0_  = ~n9563 ;
  assign \g52310/_0_  = ~n9572 ;
  assign \g53066/_0_  = ~n9581 ;
  assign \g53087/_0_  = ~n9592 ;
  assign \g53151/_0_  = ~n9602 ;
  assign \g53608/_0_  = ~n9611 ;
  assign \g53634/_0_  = ~n9624 ;
  assign \g54053/_0_  = ~n9634 ;
  assign \g54091/_0_  = ~n9644 ;
  assign \g54103/_0_  = ~n9654 ;
  assign \g54268/_0_  = ~n9662 ;
  assign \g54277/_0_  = ~n9671 ;
  assign \g54287/_0_  = ~n9677 ;
  assign \g54294/_0_  = n9687 ;
  assign \g54449/_0_  = ~n9696 ;
  assign \g54453/_0_  = ~n9705 ;
  assign \g54484/_0_  = ~n9715 ;
  assign \g54528/_0_  = ~n9730 ;
  assign \g54582/_0_  = ~n9734 ;
  assign \g55448/_0_  = ~n9743 ;
  assign \g55693/_1_  = ~n9655 ;
  assign \g55874/_0_  = n9748 ;
  assign \g56203/_0_  = ~n9751 ;
  assign \g56303/_0_  = ~n9753 ;
  assign \g56329/_0_  = ~n9756 ;
  assign \g56336/_0_  = ~n9759 ;
  assign \g56345/_0_  = ~n9762 ;
  assign \g56367/_0_  = ~n9765 ;
  assign \g56411/_0_  = ~n9768 ;
  assign \g56529/_0_  = n9773 ;
  assign \g56858/_0_  = ~n9775 ;
  assign \g60443/_1_  = ~n8534 ;
  assign \g63395/_0_  = ~n9793 ;
  assign \g63442/_0_  = ~n9826 ;
  assign \g63595/_0_  = ~n9842 ;
  assign \g63996/_0_  = ~n9860 ;
  assign \g64048/_0_  = ~n9876 ;
  assign \g64071/_0_  = ~n9917 ;
  assign \g64085/_0_  = ~n9933 ;
  assign \g64096/_0_  = ~n9951 ;
  assign \g64119/_0_  = ~n9974 ;
  assign \g64216/_0_  = ~n9997 ;
  assign \g64513/_0_  = ~n10013 ;
  assign \g64566/_0_  = ~n10029 ;
  assign \g64694/_0_  = ~n10058 ;
  assign \g64913/_0_  = ~n10081 ;
endmodule
