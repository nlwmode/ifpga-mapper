module top (\a0_pad , \a1_pad , \a2_pad , \a3_pad , \a4_pad , \b0_pad , \b1_pad , \b2_pad , \b3_pad , \b4_pad , \b5_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \c3_pad , \c4_pad , \c5_pad , c_pad, \d0_pad , \d1_pad , \d2_pad , \d3_pad , \d4_pad , \d5_pad , d_pad, \e0_pad , \e2_pad , \e3_pad , \e4_pad , \e5_pad , e_pad, \f0_pad , \f1_pad , \f2_pad , \f3_pad , \f4_pad , \f5_pad , f_pad, \g0_pad , \g1_pad , \g2_pad , \g3_pad , \g4_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , \h3_pad , \h4_pad , \h5_pad , h_pad, \i0_pad , \i10_pad , \i1_pad , \i2_pad , \i3_pad , \i4_pad , \i5_pad , i_pad, \j0_pad , \j2_pad , \j3_pad , \j4_pad , \j5_pad , j_pad, \k0_pad , \k1_pad , \k2_pad , \k3_pad , \k4_pad , \k5_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , \l3_pad , \l4_pad , \l5_pad , \l6_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , \m3_pad , \m4_pad , \m5_pad , \m6_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , \n3_pad , \n4_pad , \n5_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , \o3_pad , \o4_pad , \o5_pad , o_pad, \p0_pad , \p10_pad , \p1_pad , \p2_pad , \p3_pad , \p4_pad , \p5_pad , p_pad, \q0_pad , \q1_pad , \q2_pad , \q3_pad , \q4_pad , \q5_pad , q_pad, \r0_pad , \r1_pad , \r2_pad , \r3_pad , \r4_pad , \r5_pad , \r6_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , \s3_pad , \s4_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , \t3_pad , \t4_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , \u3_pad , \u4_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , \v3_pad , \v4_pad , v_pad, \w0_pad , \w1_pad , \w2_pad , \w3_pad , \w4_pad , w_pad, \x0_pad , \x1_pad , \x2_pad , \x3_pad , \x4_pad , \y0_pad , \y1_pad , \y2_pad , \y3_pad , \y4_pad , \z0_pad , \z1_pad , \z2_pad , \z3_pad , \z4_pad , z_pad, \a10_pad , \a6_pad , \a7_pad , \a8_pad , \a9_pad , \b10_pad , \b6_pad , \b7_pad , \b8_pad , \b9_pad , \c10_pad , \c53 , \c6_pad , \c7_pad , \c8_pad , \c9_pad , \d10_pad , \d6_pad , \d7_pad , \d8_pad , \d9_pad , \e10_pad , \e6_pad , \e7_pad , \e8_pad , \e9_pad , \f10_pad , \f22 , \f6_pad , \f7_pad , \f8_pad , \f9_pad , \g10_pad , \g6_pad , \g7_pad , \g8_pad , \g9_pad , \h6_pad , \h7_pad , \h8_pad , \h9_pad , \i6_pad , \i7_pad , \i8_pad , \i9_pad , \j10_pad , \j6_pad , \j7_pad , \j8_pad , \j9_pad , \k10_pad , \k53 , \k6_pad , \k7_pad , \k8_pad , \k9_pad , \l10_pad , \l7_pad , \l8_pad , \l9_pad , \m10_pad , \m7_pad , \m8_pad , \m9_pad , \n10_pad , \n6_pad , \n7_pad , \n8_pad , \n9_pad , \o10_pad , \o6_pad , \o7_pad , \o8_pad , \o9_pad , \p6_pad , \p7_pad , \p8_pad , \p9_pad , \q10_pad , \q6_pad , \q7_pad , \q8_pad , \q9_pad , \r10_pad , \r7_pad , \r8_pad , \r9_pad , \s5_pad , \s7_pad , \s8_pad , \s9_pad , \t10_pad , \t5_pad , \t6_pad , \t7_pad , \t8_pad , \t9_pad , \u5_pad , \u7_pad , \u8_pad , \u9_pad , \v10_pad , \v5_pad , \v6_pad , \v7_pad , \v8_pad , \v9_pad , \w10_pad , \w5_pad , \w6_pad , \w7_pad , \w8_pad , \w9_pad , \x10_pad , \x21 , \x5_pad , \x6_pad , \x7_pad , \x8_pad , \x9_pad , \y10_pad , \y5_pad , \y6_pad , \y7_pad , \y8_pad , \y9_pad , \z5_pad , \z6_pad , \z7_pad , \z8_pad , \z9_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input \a3_pad  ;
	input \a4_pad  ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input \b3_pad  ;
	input \b4_pad  ;
	input \b5_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \c3_pad  ;
	input \c4_pad  ;
	input \c5_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \d3_pad  ;
	input \d4_pad  ;
	input \d5_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input \e2_pad  ;
	input \e3_pad  ;
	input \e4_pad  ;
	input \e5_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \f3_pad  ;
	input \f4_pad  ;
	input \f5_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input \g3_pad  ;
	input \g4_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input \h3_pad  ;
	input \h4_pad  ;
	input \h5_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i10_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input \i3_pad  ;
	input \i4_pad  ;
	input \i5_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input \j2_pad  ;
	input \j3_pad  ;
	input \j4_pad  ;
	input \j5_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input \k3_pad  ;
	input \k4_pad  ;
	input \k5_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input \l3_pad  ;
	input \l4_pad  ;
	input \l5_pad  ;
	input \l6_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input \m3_pad  ;
	input \m4_pad  ;
	input \m5_pad  ;
	input \m6_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input \n3_pad  ;
	input \n4_pad  ;
	input \n5_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input \o3_pad  ;
	input \o4_pad  ;
	input \o5_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input \p10_pad  ;
	input \p1_pad  ;
	input \p2_pad  ;
	input \p3_pad  ;
	input \p4_pad  ;
	input \p5_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input \q1_pad  ;
	input \q2_pad  ;
	input \q3_pad  ;
	input \q4_pad  ;
	input \q5_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input \r1_pad  ;
	input \r2_pad  ;
	input \r3_pad  ;
	input \r4_pad  ;
	input \r5_pad  ;
	input \r6_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input \s3_pad  ;
	input \s4_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input \t3_pad  ;
	input \t4_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input \u3_pad  ;
	input \u4_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input \w2_pad  ;
	input \w3_pad  ;
	input \w4_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input \x2_pad  ;
	input \x3_pad  ;
	input \x4_pad  ;
	input \y0_pad  ;
	input \y1_pad  ;
	input \y2_pad  ;
	input \y3_pad  ;
	input \y4_pad  ;
	input \z0_pad  ;
	input \z1_pad  ;
	input \z2_pad  ;
	input \z3_pad  ;
	input \z4_pad  ;
	input z_pad ;
	output \a10_pad  ;
	output \a6_pad  ;
	output \a7_pad  ;
	output \a8_pad  ;
	output \a9_pad  ;
	output \b10_pad  ;
	output \b6_pad  ;
	output \b7_pad  ;
	output \b8_pad  ;
	output \b9_pad  ;
	output \c10_pad  ;
	output \c53  ;
	output \c6_pad  ;
	output \c7_pad  ;
	output \c8_pad  ;
	output \c9_pad  ;
	output \d10_pad  ;
	output \d6_pad  ;
	output \d7_pad  ;
	output \d8_pad  ;
	output \d9_pad  ;
	output \e10_pad  ;
	output \e6_pad  ;
	output \e7_pad  ;
	output \e8_pad  ;
	output \e9_pad  ;
	output \f10_pad  ;
	output \f22  ;
	output \f6_pad  ;
	output \f7_pad  ;
	output \f8_pad  ;
	output \f9_pad  ;
	output \g10_pad  ;
	output \g6_pad  ;
	output \g7_pad  ;
	output \g8_pad  ;
	output \g9_pad  ;
	output \h6_pad  ;
	output \h7_pad  ;
	output \h8_pad  ;
	output \h9_pad  ;
	output \i6_pad  ;
	output \i7_pad  ;
	output \i8_pad  ;
	output \i9_pad  ;
	output \j10_pad  ;
	output \j6_pad  ;
	output \j7_pad  ;
	output \j8_pad  ;
	output \j9_pad  ;
	output \k10_pad  ;
	output \k53  ;
	output \k6_pad  ;
	output \k7_pad  ;
	output \k8_pad  ;
	output \k9_pad  ;
	output \l10_pad  ;
	output \l7_pad  ;
	output \l8_pad  ;
	output \l9_pad  ;
	output \m10_pad  ;
	output \m7_pad  ;
	output \m8_pad  ;
	output \m9_pad  ;
	output \n10_pad  ;
	output \n6_pad  ;
	output \n7_pad  ;
	output \n8_pad  ;
	output \n9_pad  ;
	output \o10_pad  ;
	output \o6_pad  ;
	output \o7_pad  ;
	output \o8_pad  ;
	output \o9_pad  ;
	output \p6_pad  ;
	output \p7_pad  ;
	output \p8_pad  ;
	output \p9_pad  ;
	output \q10_pad  ;
	output \q6_pad  ;
	output \q7_pad  ;
	output \q8_pad  ;
	output \q9_pad  ;
	output \r10_pad  ;
	output \r7_pad  ;
	output \r8_pad  ;
	output \r9_pad  ;
	output \s5_pad  ;
	output \s7_pad  ;
	output \s8_pad  ;
	output \s9_pad  ;
	output \t10_pad  ;
	output \t5_pad  ;
	output \t6_pad  ;
	output \t7_pad  ;
	output \t8_pad  ;
	output \t9_pad  ;
	output \u5_pad  ;
	output \u7_pad  ;
	output \u8_pad  ;
	output \u9_pad  ;
	output \v10_pad  ;
	output \v5_pad  ;
	output \v6_pad  ;
	output \v7_pad  ;
	output \v8_pad  ;
	output \v9_pad  ;
	output \w10_pad  ;
	output \w5_pad  ;
	output \w6_pad  ;
	output \w7_pad  ;
	output \w8_pad  ;
	output \w9_pad  ;
	output \x10_pad  ;
	output \x21  ;
	output \x5_pad  ;
	output \x6_pad  ;
	output \x7_pad  ;
	output \x8_pad  ;
	output \x9_pad  ;
	output \y10_pad  ;
	output \y5_pad  ;
	output \y6_pad  ;
	output \y7_pad  ;
	output \y8_pad  ;
	output \y9_pad  ;
	output \z5_pad  ;
	output \z6_pad  ;
	output \z7_pad  ;
	output \z8_pad  ;
	output \z9_pad  ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	LUT4 #(
		.INIT('h0008)
	) name0 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\r5_pad ,
		_w174_,
		_w175_
	);
	LUT3 #(
		.INIT('h40)
	) name2 (
		\i5_pad ,
		\o5_pad ,
		\p10_pad ,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\b5_pad ,
		\i10_pad ,
		_w177_
	);
	LUT4 #(
		.INIT('h0100)
	) name4 (
		\b5_pad ,
		\d5_pad ,
		\e5_pad ,
		\i10_pad ,
		_w178_
	);
	LUT3 #(
		.INIT('hba)
	) name5 (
		\e5_pad ,
		_w176_,
		_w178_,
		_w179_
	);
	LUT4 #(
		.INIT('h1011)
	) name6 (
		\c5_pad ,
		\e5_pad ,
		_w176_,
		_w178_,
		_w180_
	);
	LUT4 #(
		.INIT('h0203)
	) name7 (
		\b5_pad ,
		\d5_pad ,
		\e5_pad ,
		\i10_pad ,
		_w181_
	);
	LUT3 #(
		.INIT('h15)
	) name8 (
		\d5_pad ,
		_w176_,
		_w181_,
		_w182_
	);
	LUT3 #(
		.INIT('h40)
	) name9 (
		_w175_,
		_w180_,
		_w182_,
		_w183_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name10 (
		\r4_pad ,
		_w175_,
		_w180_,
		_w182_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\s4_pad ,
		_w184_,
		_w185_
	);
	LUT3 #(
		.INIT('h80)
	) name12 (
		\r4_pad ,
		\r5_pad ,
		_w174_,
		_w186_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\l5_pad ,
		\m5_pad ,
		_w187_
	);
	LUT4 #(
		.INIT('h0020)
	) name14 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w188_
	);
	LUT4 #(
		.INIT('h00df)
	) name15 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w189_
	);
	LUT3 #(
		.INIT('h01)
	) name16 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		_w190_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name17 (
		_w189_,
		_w180_,
		_w182_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		_w186_,
		_w191_,
		_w192_
	);
	LUT3 #(
		.INIT('h80)
	) name19 (
		\s4_pad ,
		\t4_pad ,
		_w184_,
		_w193_
	);
	LUT3 #(
		.INIT('h48)
	) name20 (
		\t4_pad ,
		_w192_,
		_w185_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\m4_pad ,
		\q0_pad ,
		_w195_
	);
	LUT4 #(
		.INIT('h0777)
	) name22 (
		\f3_pad ,
		\m0_pad ,
		\n0_pad ,
		\p5_pad ,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT4 #(
		.INIT('h153f)
	) name24 (
		\h4_pad ,
		\m5_pad ,
		\p0_pad ,
		\r0_pad ,
		_w198_
	);
	LUT4 #(
		.INIT('h153f)
	) name25 (
		\k0_pad ,
		\l0_pad ,
		\m3_pad ,
		\q3_pad ,
		_w199_
	);
	LUT4 #(
		.INIT('h135f)
	) name26 (
		\o0_pad ,
		\r4_pad ,
		\r5_pad ,
		\u0_pad ,
		_w200_
	);
	LUT4 #(
		.INIT('h0777)
	) name27 (
		\d4_pad ,
		\s0_pad ,
		\t0_pad ,
		\w4_pad ,
		_w201_
	);
	LUT4 #(
		.INIT('h8000)
	) name28 (
		_w200_,
		_w201_,
		_w198_,
		_w199_,
		_w202_
	);
	LUT2 #(
		.INIT('h7)
	) name29 (
		_w197_,
		_w202_,
		_w203_
	);
	LUT3 #(
		.INIT('h40)
	) name30 (
		\k1_pad ,
		\o1_pad ,
		\r6_pad ,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\f1_pad ,
		\m6_pad ,
		_w205_
	);
	LUT4 #(
		.INIT('h0100)
	) name32 (
		\f1_pad ,
		\h1_pad ,
		\i1_pad ,
		\m6_pad ,
		_w206_
	);
	LUT3 #(
		.INIT('hba)
	) name33 (
		\i1_pad ,
		_w204_,
		_w206_,
		_w207_
	);
	LUT4 #(
		.INIT('h1011)
	) name34 (
		\g1_pad ,
		\i1_pad ,
		_w204_,
		_w206_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		i_pad,
		_w208_,
		_w209_
	);
	LUT3 #(
		.INIT('h23)
	) name36 (
		i_pad,
		\s1_pad ,
		_w208_,
		_w210_
	);
	LUT3 #(
		.INIT('h01)
	) name37 (
		\a1_pad ,
		\b1_pad ,
		\c1_pad ,
		_w211_
	);
	LUT4 #(
		.INIT('h0100)
	) name38 (
		\a1_pad ,
		\b1_pad ,
		\c1_pad ,
		\r1_pad ,
		_w212_
	);
	LUT4 #(
		.INIT('h5051)
	) name39 (
		\p1_pad ,
		\q1_pad ,
		\z0_pad ,
		_w212_,
		_w213_
	);
	LUT3 #(
		.INIT('h01)
	) name40 (
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w214_
	);
	LUT4 #(
		.INIT('h5554)
	) name41 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w215_
	);
	LUT4 #(
		.INIT('haaab)
	) name42 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\v0_pad ,
		_w215_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\x0_pad ,
		\y0_pad ,
		_w218_
	);
	LUT3 #(
		.INIT('h02)
	) name45 (
		\w0_pad ,
		\x0_pad ,
		\y0_pad ,
		_w219_
	);
	LUT3 #(
		.INIT('h10)
	) name46 (
		\v0_pad ,
		_w215_,
		_w219_,
		_w220_
	);
	LUT3 #(
		.INIT('h45)
	) name47 (
		h_pad,
		_w213_,
		_w220_,
		_w221_
	);
	LUT3 #(
		.INIT('h06)
	) name48 (
		\s1_pad ,
		_w209_,
		_w221_,
		_w222_
	);
	LUT3 #(
		.INIT('h04)
	) name49 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		_w223_
	);
	LUT4 #(
		.INIT('h0004)
	) name50 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w224_
	);
	LUT3 #(
		.INIT('h01)
	) name51 (
		\d1_pad ,
		\w0_pad ,
		\z0_pad ,
		_w225_
	);
	LUT3 #(
		.INIT('h80)
	) name52 (
		_w211_,
		_w218_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\v0_pad ,
		_w215_,
		_w227_
	);
	LUT3 #(
		.INIT('h15)
	) name54 (
		_w224_,
		_w226_,
		_w227_,
		_w228_
	);
	LUT4 #(
		.INIT('h5444)
	) name55 (
		\x2_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		b_pad,
		_w229_,
		_w230_
	);
	LUT4 #(
		.INIT('h7b00)
	) name57 (
		\t1_pad ,
		_w228_,
		_w222_,
		_w230_,
		_w231_
	);
	LUT3 #(
		.INIT('h54)
	) name58 (
		g_pad,
		_w215_,
		_w208_,
		_w232_
	);
	LUT4 #(
		.INIT('h0010)
	) name59 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w233_
	);
	LUT4 #(
		.INIT('h5545)
	) name60 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w234_
	);
	LUT4 #(
		.INIT('h00ab)
	) name61 (
		g_pad,
		_w215_,
		_w208_,
		_w234_,
		_w235_
	);
	LUT4 #(
		.INIT('h0203)
	) name62 (
		\f1_pad ,
		\h1_pad ,
		\i1_pad ,
		\m6_pad ,
		_w236_
	);
	LUT3 #(
		.INIT('h15)
	) name63 (
		\h1_pad ,
		_w204_,
		_w236_,
		_w237_
	);
	LUT4 #(
		.INIT('h20a0)
	) name64 (
		_w226_,
		_w208_,
		_w217_,
		_w237_,
		_w238_
	);
	LUT4 #(
		.INIT('h0040)
	) name65 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w239_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\r1_pad ,
		\v0_pad ,
		_w240_
	);
	LUT3 #(
		.INIT('h51)
	) name67 (
		f_pad,
		_w239_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w238_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		j_pad,
		\q1_pad ,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\q2_pad ,
		\r2_pad ,
		_w244_
	);
	LUT3 #(
		.INIT('h07)
	) name71 (
		_w239_,
		_w243_,
		_w244_,
		_w245_
	);
	LUT4 #(
		.INIT('haa80)
	) name72 (
		\s2_pad ,
		_w239_,
		_w243_,
		_w244_,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		j_pad,
		\p1_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w239_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w246_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\q2_pad ,
		\r2_pad ,
		_w250_
	);
	LUT3 #(
		.INIT('h07)
	) name77 (
		_w239_,
		_w243_,
		_w250_,
		_w251_
	);
	LUT4 #(
		.INIT('h5540)
	) name78 (
		\s2_pad ,
		_w239_,
		_w243_,
		_w250_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w248_,
		_w252_,
		_w253_
	);
	LUT3 #(
		.INIT('h1b)
	) name80 (
		_w232_,
		_w249_,
		_w253_,
		_w254_
	);
	LUT4 #(
		.INIT('h8488)
	) name81 (
		\t2_pad ,
		_w234_,
		_w242_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('he)
	) name82 (
		_w235_,
		_w255_,
		_w256_
	);
	LUT4 #(
		.INIT('h00fe)
	) name83 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w257_
	);
	LUT4 #(
		.INIT('hff01)
	) name84 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w258_
	);
	LUT3 #(
		.INIT('h54)
	) name85 (
		\e0_pad ,
		_w180_,
		_w257_,
		_w259_
	);
	LUT4 #(
		.INIT('h0004)
	) name86 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w260_
	);
	LUT4 #(
		.INIT('h00fb)
	) name87 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w261_
	);
	LUT4 #(
		.INIT('h00ab)
	) name88 (
		\e0_pad ,
		_w180_,
		_w257_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\f3_pad ,
		\g3_pad ,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\h0_pad ,
		\q5_pad ,
		_w264_
	);
	LUT3 #(
		.INIT('h13)
	) name91 (
		_w174_,
		_w263_,
		_w264_,
		_w265_
	);
	LUT4 #(
		.INIT('h5450)
	) name92 (
		\h3_pad ,
		_w174_,
		_w263_,
		_w264_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		\h0_pad ,
		\p5_pad ,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w174_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w266_,
		_w268_,
		_w269_
	);
	LUT3 #(
		.INIT('h54)
	) name96 (
		\i3_pad ,
		_w266_,
		_w268_,
		_w270_
	);
	LUT4 #(
		.INIT('h4445)
	) name97 (
		\h0_pad ,
		\i3_pad ,
		_w266_,
		_w268_,
		_w271_
	);
	LUT4 #(
		.INIT('h5155)
	) name98 (
		\h0_pad ,
		\j3_pad ,
		\p3_pad ,
		_w270_,
		_w272_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name99 (
		\q3_pad ,
		\r3_pad ,
		_w259_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\q3_pad ,
		\r3_pad ,
		_w274_
	);
	LUT4 #(
		.INIT('h00ab)
	) name101 (
		\e0_pad ,
		_w180_,
		_w257_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		\t4_pad ,
		\u4_pad ,
		_w276_
	);
	LUT4 #(
		.INIT('h0001)
	) name103 (
		\v4_pad ,
		\w4_pad ,
		\x4_pad ,
		\y4_pad ,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\s4_pad ,
		\z4_pad ,
		_w278_
	);
	LUT4 #(
		.INIT('h4000)
	) name105 (
		_w257_,
		_w276_,
		_w277_,
		_w278_,
		_w279_
	);
	LUT4 #(
		.INIT('h1500)
	) name106 (
		\r4_pad ,
		_w180_,
		_w182_,
		_w279_,
		_w280_
	);
	LUT4 #(
		.INIT('h4044)
	) name107 (
		\j5_pad ,
		\k5_pad ,
		\r4_pad ,
		\r5_pad ,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\d0_pad ,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w280_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\f3_pad ,
		\g3_pad ,
		_w284_
	);
	LUT3 #(
		.INIT('h07)
	) name111 (
		_w174_,
		_w264_,
		_w284_,
		_w285_
	);
	LUT4 #(
		.INIT('haa80)
	) name112 (
		\h3_pad ,
		_w174_,
		_w264_,
		_w284_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w268_,
		_w286_,
		_w287_
	);
	LUT4 #(
		.INIT('h1115)
	) name114 (
		\h0_pad ,
		\i3_pad ,
		_w268_,
		_w286_,
		_w288_
	);
	LUT4 #(
		.INIT('h2223)
	) name115 (
		\e0_pad ,
		\h0_pad ,
		_w180_,
		_w257_,
		_w289_
	);
	LUT4 #(
		.INIT('hf700)
	) name116 (
		\k3_pad ,
		\p3_pad ,
		_w288_,
		_w289_,
		_w290_
	);
	LUT3 #(
		.INIT('h01)
	) name117 (
		_w275_,
		_w283_,
		_w290_,
		_w291_
	);
	LUT4 #(
		.INIT('h999c)
	) name118 (
		\e0_pad ,
		\s3_pad ,
		_w180_,
		_w257_,
		_w292_
	);
	LUT3 #(
		.INIT('h40)
	) name119 (
		_w273_,
		_w291_,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name120 (
		\t3_pad ,
		_w261_,
		_w262_,
		_w293_,
		_w294_
	);
	LUT4 #(
		.INIT('h8000)
	) name121 (
		\s4_pad ,
		\t4_pad ,
		\u4_pad ,
		_w184_,
		_w295_
	);
	LUT3 #(
		.INIT('h48)
	) name122 (
		\u4_pad ,
		_w192_,
		_w193_,
		_w296_
	);
	LUT3 #(
		.INIT('h20)
	) name123 (
		\s0_pad ,
		_w280_,
		_w282_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		\j0_pad ,
		\q5_pad ,
		_w298_
	);
	LUT3 #(
		.INIT('h80)
	) name125 (
		\d4_pad ,
		\e4_pad ,
		\f4_pad ,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\j0_pad ,
		\p5_pad ,
		_w300_
	);
	LUT4 #(
		.INIT('h5700)
	) name127 (
		\i4_pad ,
		_w298_,
		_w299_,
		_w300_,
		_w301_
	);
	LUT3 #(
		.INIT('h08)
	) name128 (
		\g4_pad ,
		\p4_pad ,
		_w301_,
		_w302_
	);
	LUT4 #(
		.INIT('h0080)
	) name129 (
		\g4_pad ,
		\p4_pad ,
		\q0_pad ,
		_w301_,
		_w303_
	);
	LUT3 #(
		.INIT('h80)
	) name130 (
		\p3_pad ,
		\s3_pad ,
		\t3_pad ,
		_w304_
	);
	LUT3 #(
		.INIT('h80)
	) name131 (
		\m0_pad ,
		_w274_,
		_w304_,
		_w305_
	);
	LUT4 #(
		.INIT('h0777)
	) name132 (
		\l0_pad ,
		\l3_pad ,
		\n5_pad ,
		\p0_pad ,
		_w306_
	);
	LUT4 #(
		.INIT('h135f)
	) name133 (
		\g4_pad ,
		\l5_pad ,
		\r0_pad ,
		\u0_pad ,
		_w307_
	);
	LUT4 #(
		.INIT('h0777)
	) name134 (
		\n0_pad ,
		\q5_pad ,
		\t0_pad ,
		\v4_pad ,
		_w308_
	);
	LUT3 #(
		.INIT('h80)
	) name135 (
		_w306_,
		_w307_,
		_w308_,
		_w309_
	);
	LUT3 #(
		.INIT('h01)
	) name136 (
		\r3_pad ,
		\s3_pad ,
		\t3_pad ,
		_w310_
	);
	LUT4 #(
		.INIT('h0002)
	) name137 (
		\n3_pad ,
		\o3_pad ,
		\p3_pad ,
		\q3_pad ,
		_w311_
	);
	LUT3 #(
		.INIT('h80)
	) name138 (
		\k0_pad ,
		_w310_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\o0_pad ,
		_w261_,
		_w313_
	);
	LUT4 #(
		.INIT('h0100)
	) name140 (
		_w305_,
		_w312_,
		_w313_,
		_w309_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		_w303_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('hb)
	) name142 (
		_w297_,
		_w315_,
		_w316_
	);
	LUT4 #(
		.INIT('h5c0c)
	) name143 (
		i_pad,
		\s1_pad ,
		\t1_pad ,
		_w208_,
		_w317_
	);
	LUT3 #(
		.INIT('h01)
	) name144 (
		_w210_,
		_w221_,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('h5444)
	) name145 (
		\y2_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		b_pad,
		_w319_,
		_w320_
	);
	LUT4 #(
		.INIT('h7b00)
	) name147 (
		\u1_pad ,
		_w228_,
		_w318_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\w2_pad ,
		\x2_pad ,
		_w322_
	);
	LUT4 #(
		.INIT('h0001)
	) name149 (
		\w2_pad ,
		\x2_pad ,
		\y2_pad ,
		\z2_pad ,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		_w234_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w235_,
		_w324_,
		_w325_
	);
	LUT4 #(
		.INIT('h0002)
	) name152 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w326_
	);
	LUT3 #(
		.INIT('h07)
	) name153 (
		\r4_pad ,
		_w279_,
		_w326_,
		_w327_
	);
	LUT3 #(
		.INIT('h51)
	) name154 (
		\p5_pad ,
		\q5_pad ,
		\v4_pad ,
		_w328_
	);
	LUT4 #(
		.INIT('h7f00)
	) name155 (
		\r5_pad ,
		_w276_,
		_w277_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('h0004)
	) name156 (
		\r4_pad ,
		\s4_pad ,
		\t4_pad ,
		\u4_pad ,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		_w257_,
		_w330_,
		_w331_
	);
	LUT3 #(
		.INIT('h45)
	) name158 (
		\f0_pad ,
		_w329_,
		_w331_,
		_w332_
	);
	LUT4 #(
		.INIT('h6366)
	) name159 (
		\f0_pad ,
		\u3_pad ,
		_w329_,
		_w331_,
		_w333_
	);
	LUT4 #(
		.INIT('h3202)
	) name160 (
		\l3_pad ,
		z_pad,
		_w327_,
		_w333_,
		_w334_
	);
	LUT3 #(
		.INIT('h48)
	) name161 (
		\v4_pad ,
		_w192_,
		_w295_,
		_w335_
	);
	LUT4 #(
		.INIT('h0010)
	) name162 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w336_
	);
	LUT4 #(
		.INIT('h007f)
	) name163 (
		_w174_,
		_w310_,
		_w311_,
		_w336_,
		_w337_
	);
	LUT4 #(
		.INIT('h8000)
	) name164 (
		_w174_,
		_w177_,
		_w274_,
		_w304_,
		_w338_
	);
	LUT4 #(
		.INIT('h0080)
	) name165 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w339_
	);
	LUT4 #(
		.INIT('hff7d)
	) name166 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w340_
	);
	LUT3 #(
		.INIT('hdf)
	) name167 (
		_w337_,
		_w338_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\r1_pad ,
		_w239_,
		_w342_
	);
	LUT3 #(
		.INIT('h08)
	) name169 (
		_w208_,
		_w237_,
		_w342_,
		_w343_
	);
	LUT4 #(
		.INIT('h0400)
	) name170 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w344_
	);
	LUT4 #(
		.INIT('h5155)
	) name171 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w345_
	);
	LUT4 #(
		.INIT('h7f00)
	) name172 (
		_w214_,
		_w208_,
		_w237_,
		_w345_,
		_w346_
	);
	LUT4 #(
		.INIT('haa2a)
	) name173 (
		\v0_pad ,
		_w208_,
		_w237_,
		_w342_,
		_w347_
	);
	LUT3 #(
		.INIT('h84)
	) name174 (
		\v0_pad ,
		_w346_,
		_w343_,
		_w348_
	);
	LUT4 #(
		.INIT('h1555)
	) name175 (
		k_pad,
		\s1_pad ,
		\t1_pad ,
		\u1_pad ,
		_w349_
	);
	LUT4 #(
		.INIT('h5554)
	) name176 (
		k_pad,
		\s1_pad ,
		\t1_pad ,
		\u1_pad ,
		_w350_
	);
	LUT4 #(
		.INIT('h0b4f)
	) name177 (
		i_pad,
		_w208_,
		_w349_,
		_w350_,
		_w351_
	);
	LUT4 #(
		.INIT('h8488)
	) name178 (
		\v1_pad ,
		_w228_,
		_w221_,
		_w351_,
		_w352_
	);
	LUT4 #(
		.INIT('ha888)
	) name179 (
		\z2_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		b_pad,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('hb)
	) name181 (
		_w352_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\w2_pad ,
		\x2_pad ,
		_w356_
	);
	LUT4 #(
		.INIT('h8000)
	) name183 (
		\w2_pad ,
		\x2_pad ,
		\y2_pad ,
		\z2_pad ,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w234_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		\g0_pad ,
		_w180_,
		_w359_
	);
	LUT3 #(
		.INIT('h23)
	) name186 (
		\g0_pad ,
		\u3_pad ,
		_w180_,
		_w360_
	);
	LUT3 #(
		.INIT('h12)
	) name187 (
		\u3_pad ,
		_w332_,
		_w359_,
		_w361_
	);
	LUT4 #(
		.INIT('h5540)
	) name188 (
		\m3_pad ,
		\r4_pad ,
		_w279_,
		_w326_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		z_pad,
		_w362_,
		_w363_
	);
	LUT4 #(
		.INIT('h7b00)
	) name190 (
		\v3_pad ,
		_w327_,
		_w361_,
		_w363_,
		_w364_
	);
	LUT4 #(
		.INIT('h60c0)
	) name191 (
		\v4_pad ,
		\w4_pad ,
		_w192_,
		_w295_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\w0_pad ,
		_w347_,
		_w366_
	);
	LUT3 #(
		.INIT('h80)
	) name193 (
		\r1_pad ,
		\v0_pad ,
		_w239_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		_w346_,
		_w367_,
		_w368_
	);
	LUT4 #(
		.INIT('h0048)
	) name195 (
		\w0_pad ,
		_w346_,
		_w347_,
		_w367_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		\v1_pad ,
		_w350_,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		\v1_pad ,
		_w349_,
		_w371_
	);
	LUT4 #(
		.INIT('hfb40)
	) name198 (
		i_pad,
		_w208_,
		_w370_,
		_w371_,
		_w372_
	);
	LUT4 #(
		.INIT('h8488)
	) name199 (
		\w1_pad ,
		_w228_,
		_w221_,
		_w372_,
		_w373_
	);
	LUT4 #(
		.INIT('ha888)
	) name200 (
		\a3_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		b_pad,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('hb)
	) name202 (
		_w373_,
		_w375_,
		_w376_
	);
	LUT3 #(
		.INIT('h54)
	) name203 (
		\t2_pad ,
		_w248_,
		_w252_,
		_w377_
	);
	LUT4 #(
		.INIT('h4445)
	) name204 (
		j_pad,
		\t2_pad ,
		_w248_,
		_w252_,
		_w378_
	);
	LUT4 #(
		.INIT('h1115)
	) name205 (
		j_pad,
		\t2_pad ,
		_w246_,
		_w248_,
		_w379_
	);
	LUT3 #(
		.INIT('hd8)
	) name206 (
		_w232_,
		_w378_,
		_w379_,
		_w380_
	);
	LUT4 #(
		.INIT('h8884)
	) name207 (
		\w2_pad ,
		_w234_,
		_w242_,
		_w380_,
		_w381_
	);
	LUT4 #(
		.INIT('h5c0c)
	) name208 (
		\g0_pad ,
		\u3_pad ,
		\v3_pad ,
		_w180_,
		_w382_
	);
	LUT3 #(
		.INIT('h01)
	) name209 (
		_w332_,
		_w360_,
		_w382_,
		_w383_
	);
	LUT4 #(
		.INIT('h5540)
	) name210 (
		\n3_pad ,
		\r4_pad ,
		_w279_,
		_w326_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		z_pad,
		_w384_,
		_w385_
	);
	LUT4 #(
		.INIT('h7b00)
	) name212 (
		\w3_pad ,
		_w327_,
		_w383_,
		_w385_,
		_w386_
	);
	LUT4 #(
		.INIT('h070f)
	) name213 (
		\v4_pad ,
		\w4_pad ,
		\x4_pad ,
		_w295_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\w4_pad ,
		\x4_pad ,
		_w388_
	);
	LUT3 #(
		.INIT('h80)
	) name215 (
		\v4_pad ,
		_w295_,
		_w388_,
		_w389_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name216 (
		\v4_pad ,
		_w192_,
		_w295_,
		_w388_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w387_,
		_w390_,
		_w391_
	);
	LUT3 #(
		.INIT('h80)
	) name218 (
		\w0_pad ,
		\x0_pad ,
		_w347_,
		_w392_
	);
	LUT3 #(
		.INIT('h48)
	) name219 (
		\x0_pad ,
		_w368_,
		_w366_,
		_w393_
	);
	LUT3 #(
		.INIT('h01)
	) name220 (
		\v1_pad ,
		\w1_pad ,
		_w350_,
		_w394_
	);
	LUT3 #(
		.INIT('h08)
	) name221 (
		\v1_pad ,
		\w1_pad ,
		_w349_,
		_w395_
	);
	LUT4 #(
		.INIT('hfb40)
	) name222 (
		i_pad,
		_w208_,
		_w394_,
		_w395_,
		_w396_
	);
	LUT4 #(
		.INIT('h8488)
	) name223 (
		\x1_pad ,
		_w228_,
		_w221_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('ha888)
	) name224 (
		\b3_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		b_pad,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('hb)
	) name226 (
		_w397_,
		_w399_,
		_w400_
	);
	LUT3 #(
		.INIT('h51)
	) name227 (
		\w2_pad ,
		_w232_,
		_w378_,
		_w401_
	);
	LUT3 #(
		.INIT('ha8)
	) name228 (
		\w2_pad ,
		_w232_,
		_w379_,
		_w402_
	);
	LUT3 #(
		.INIT('h01)
	) name229 (
		_w242_,
		_w402_,
		_w401_,
		_w403_
	);
	LUT3 #(
		.INIT('h48)
	) name230 (
		\x2_pad ,
		_w234_,
		_w403_,
		_w404_
	);
	LUT3 #(
		.INIT('h01)
	) name231 (
		\u3_pad ,
		\v3_pad ,
		\w3_pad ,
		_w405_
	);
	LUT4 #(
		.INIT('h0010)
	) name232 (
		\g0_pad ,
		\i0_pad ,
		_w180_,
		_w405_,
		_w406_
	);
	LUT4 #(
		.INIT('h1555)
	) name233 (
		\i0_pad ,
		\u3_pad ,
		\v3_pad ,
		\w3_pad ,
		_w407_
	);
	LUT3 #(
		.INIT('hb0)
	) name234 (
		\g0_pad ,
		_w180_,
		_w407_,
		_w408_
	);
	LUT3 #(
		.INIT('h01)
	) name235 (
		_w332_,
		_w406_,
		_w408_,
		_w409_
	);
	LUT4 #(
		.INIT('haa80)
	) name236 (
		\o3_pad ,
		\r4_pad ,
		_w279_,
		_w326_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		z_pad,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('h48ff)
	) name238 (
		\x3_pad ,
		_w327_,
		_w409_,
		_w411_,
		_w412_
	);
	LUT4 #(
		.INIT('h8000)
	) name239 (
		\v4_pad ,
		\y4_pad ,
		_w295_,
		_w388_,
		_w413_
	);
	LUT3 #(
		.INIT('h48)
	) name240 (
		\y4_pad ,
		_w192_,
		_w389_,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		\c3_pad ,
		\d3_pad ,
		_w415_
	);
	LUT3 #(
		.INIT('h80)
	) name242 (
		\c3_pad ,
		\d3_pad ,
		\e3_pad ,
		_w416_
	);
	LUT3 #(
		.INIT('h4c)
	) name243 (
		_w205_,
		_w239_,
		_w416_,
		_w417_
	);
	LUT3 #(
		.INIT('h15)
	) name244 (
		_w224_,
		_w205_,
		_w233_,
		_w418_
	);
	LUT2 #(
		.INIT('hb)
	) name245 (
		_w417_,
		_w418_,
		_w419_
	);
	LUT3 #(
		.INIT('h48)
	) name246 (
		\y0_pad ,
		_w368_,
		_w392_,
		_w420_
	);
	LUT4 #(
		.INIT('h0080)
	) name247 (
		\v1_pad ,
		\w1_pad ,
		\x1_pad ,
		_w349_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		k_pad,
		_w421_,
		_w422_
	);
	LUT4 #(
		.INIT('h0023)
	) name249 (
		i_pad,
		k_pad,
		_w208_,
		_w421_,
		_w423_
	);
	LUT4 #(
		.INIT('h0001)
	) name250 (
		\v1_pad ,
		\w1_pad ,
		\x1_pad ,
		_w350_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		k_pad,
		_w424_,
		_w425_
	);
	LUT4 #(
		.INIT('h0010)
	) name252 (
		i_pad,
		k_pad,
		_w208_,
		_w424_,
		_w426_
	);
	LUT3 #(
		.INIT('h01)
	) name253 (
		_w221_,
		_w426_,
		_w423_,
		_w427_
	);
	LUT4 #(
		.INIT('h5444)
	) name254 (
		\c3_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		b_pad,
		_w428_,
		_w429_
	);
	LUT4 #(
		.INIT('h7b00)
	) name256 (
		\y1_pad ,
		_w228_,
		_w427_,
		_w429_,
		_w430_
	);
	LUT3 #(
		.INIT('h08)
	) name257 (
		_w232_,
		_w322_,
		_w378_,
		_w431_
	);
	LUT3 #(
		.INIT('h04)
	) name258 (
		_w232_,
		_w356_,
		_w379_,
		_w432_
	);
	LUT3 #(
		.INIT('h54)
	) name259 (
		_w242_,
		_w431_,
		_w432_,
		_w433_
	);
	LUT3 #(
		.INIT('h48)
	) name260 (
		\y2_pad ,
		_w234_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		\x3_pad ,
		_w407_,
		_w435_
	);
	LUT3 #(
		.INIT('h0b)
	) name262 (
		\g0_pad ,
		_w180_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('h5554)
	) name263 (
		\i0_pad ,
		\u3_pad ,
		\v3_pad ,
		\w3_pad ,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		\x3_pad ,
		_w437_,
		_w438_
	);
	LUT3 #(
		.INIT('h04)
	) name265 (
		\g0_pad ,
		_w180_,
		_w438_,
		_w439_
	);
	LUT3 #(
		.INIT('h01)
	) name266 (
		_w332_,
		_w439_,
		_w436_,
		_w440_
	);
	LUT4 #(
		.INIT('haa80)
	) name267 (
		\p3_pad ,
		\r4_pad ,
		_w279_,
		_w326_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		z_pad,
		_w441_,
		_w442_
	);
	LUT4 #(
		.INIT('h48ff)
	) name269 (
		\y3_pad ,
		_w327_,
		_w440_,
		_w442_,
		_w443_
	);
	LUT3 #(
		.INIT('h48)
	) name270 (
		\z4_pad ,
		_w192_,
		_w413_,
		_w444_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		\y0_pad ,
		\z0_pad ,
		_w445_
	);
	LUT4 #(
		.INIT('h8000)
	) name272 (
		\w0_pad ,
		\x0_pad ,
		_w347_,
		_w445_,
		_w446_
	);
	LUT4 #(
		.INIT('h60c0)
	) name273 (
		\y0_pad ,
		\z0_pad ,
		_w368_,
		_w392_,
		_w447_
	);
	LUT3 #(
		.INIT('h8c)
	) name274 (
		i_pad,
		\y1_pad ,
		_w208_,
		_w448_
	);
	LUT3 #(
		.INIT('h10)
	) name275 (
		i_pad,
		\y1_pad ,
		_w208_,
		_w449_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name276 (
		\y1_pad ,
		_w209_,
		_w425_,
		_w422_,
		_w450_
	);
	LUT4 #(
		.INIT('h8884)
	) name277 (
		\z1_pad ,
		_w228_,
		_w221_,
		_w450_,
		_w451_
	);
	LUT4 #(
		.INIT('ha888)
	) name278 (
		\d3_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		b_pad,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('hb)
	) name280 (
		_w451_,
		_w453_,
		_w454_
	);
	LUT4 #(
		.INIT('haa8a)
	) name281 (
		\y2_pad ,
		_w232_,
		_w356_,
		_w379_,
		_w455_
	);
	LUT4 #(
		.INIT('h5515)
	) name282 (
		\y2_pad ,
		_w232_,
		_w322_,
		_w378_,
		_w456_
	);
	LUT3 #(
		.INIT('h01)
	) name283 (
		_w242_,
		_w456_,
		_w455_,
		_w457_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name284 (
		\z2_pad ,
		_w234_,
		_w235_,
		_w457_,
		_w458_
	);
	LUT3 #(
		.INIT('h08)
	) name285 (
		\x3_pad ,
		\y3_pad ,
		_w407_,
		_w459_
	);
	LUT3 #(
		.INIT('h0b)
	) name286 (
		\g0_pad ,
		_w180_,
		_w459_,
		_w460_
	);
	LUT3 #(
		.INIT('h01)
	) name287 (
		\x3_pad ,
		\y3_pad ,
		_w437_,
		_w461_
	);
	LUT3 #(
		.INIT('h04)
	) name288 (
		\g0_pad ,
		_w180_,
		_w461_,
		_w462_
	);
	LUT3 #(
		.INIT('h01)
	) name289 (
		_w332_,
		_w462_,
		_w460_,
		_w463_
	);
	LUT4 #(
		.INIT('haa80)
	) name290 (
		\q3_pad ,
		\r4_pad ,
		_w279_,
		_w326_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		z_pad,
		_w464_,
		_w465_
	);
	LUT4 #(
		.INIT('h48ff)
	) name292 (
		\z3_pad ,
		_w327_,
		_w463_,
		_w465_,
		_w466_
	);
	LUT3 #(
		.INIT('h48)
	) name293 (
		\a1_pad ,
		_w368_,
		_w446_,
		_w467_
	);
	LUT3 #(
		.INIT('h8a)
	) name294 (
		\z1_pad ,
		_w422_,
		_w448_,
		_w468_
	);
	LUT4 #(
		.INIT('h2322)
	) name295 (
		\z1_pad ,
		_w221_,
		_w425_,
		_w449_,
		_w469_
	);
	LUT4 #(
		.INIT('h8488)
	) name296 (
		\a2_pad ,
		_w228_,
		_w468_,
		_w469_,
		_w470_
	);
	LUT4 #(
		.INIT('ha888)
	) name297 (
		\e3_pad ,
		_w224_,
		_w226_,
		_w227_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		b_pad,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('hb)
	) name299 (
		_w470_,
		_w472_,
		_w473_
	);
	LUT3 #(
		.INIT('h31)
	) name300 (
		\v2_pad ,
		_w232_,
		_w379_,
		_w474_
	);
	LUT3 #(
		.INIT('hc4)
	) name301 (
		\u2_pad ,
		_w232_,
		_w378_,
		_w475_
	);
	LUT3 #(
		.INIT('h01)
	) name302 (
		_w242_,
		_w475_,
		_w474_,
		_w476_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name303 (
		\a3_pad ,
		_w234_,
		_w235_,
		_w476_,
		_w477_
	);
	LUT4 #(
		.INIT('h0080)
	) name304 (
		\x3_pad ,
		\y3_pad ,
		\z3_pad ,
		_w407_,
		_w478_
	);
	LUT4 #(
		.INIT('h0023)
	) name305 (
		\g0_pad ,
		\i0_pad ,
		_w180_,
		_w478_,
		_w479_
	);
	LUT4 #(
		.INIT('h0001)
	) name306 (
		\x3_pad ,
		\y3_pad ,
		\z3_pad ,
		_w437_,
		_w480_
	);
	LUT4 #(
		.INIT('h0010)
	) name307 (
		\g0_pad ,
		\i0_pad ,
		_w180_,
		_w480_,
		_w481_
	);
	LUT4 #(
		.INIT('haaa9)
	) name308 (
		\a4_pad ,
		_w332_,
		_w481_,
		_w479_,
		_w482_
	);
	LUT4 #(
		.INIT('h5540)
	) name309 (
		\r3_pad ,
		\r4_pad ,
		_w279_,
		_w326_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		z_pad,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('hd0)
	) name311 (
		_w327_,
		_w482_,
		_w484_,
		_w485_
	);
	LUT3 #(
		.INIT('h80)
	) name312 (
		\a1_pad ,
		\b1_pad ,
		_w446_,
		_w486_
	);
	LUT4 #(
		.INIT('h60c0)
	) name313 (
		\a1_pad ,
		\b1_pad ,
		_w368_,
		_w446_,
		_w487_
	);
	LUT2 #(
		.INIT('hd)
	) name314 (
		\b2_pad ,
		b_pad,
		_w488_
	);
	LUT4 #(
		.INIT('h2333)
	) name315 (
		\a3_pad ,
		j_pad,
		\u2_pad ,
		_w377_,
		_w489_
	);
	LUT4 #(
		.INIT('h2223)
	) name316 (
		g_pad,
		j_pad,
		_w215_,
		_w208_,
		_w490_
	);
	LUT4 #(
		.INIT('hf700)
	) name317 (
		\a3_pad ,
		\v2_pad ,
		_w379_,
		_w490_,
		_w491_
	);
	LUT4 #(
		.INIT('h0013)
	) name318 (
		_w232_,
		_w242_,
		_w489_,
		_w491_,
		_w492_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name319 (
		\b3_pad ,
		_w234_,
		_w235_,
		_w492_,
		_w493_
	);
	LUT3 #(
		.INIT('h9a)
	) name320 (
		\a4_pad ,
		\g0_pad ,
		_w180_,
		_w494_
	);
	LUT4 #(
		.INIT('h0100)
	) name321 (
		_w332_,
		_w481_,
		_w479_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('hcc80)
	) name322 (
		\r4_pad ,
		\s3_pad ,
		_w279_,
		_w326_,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		z_pad,
		_w496_,
		_w497_
	);
	LUT4 #(
		.INIT('h48ff)
	) name324 (
		\b4_pad ,
		_w327_,
		_w495_,
		_w497_,
		_w498_
	);
	LUT4 #(
		.INIT('h8000)
	) name325 (
		\a1_pad ,
		\b1_pad ,
		\c1_pad ,
		_w446_,
		_w499_
	);
	LUT3 #(
		.INIT('h48)
	) name326 (
		\c1_pad ,
		_w368_,
		_w486_,
		_w500_
	);
	LUT3 #(
		.INIT('hde)
	) name327 (
		\b2_pad ,
		b_pad,
		\c2_pad ,
		_w501_
	);
	LUT3 #(
		.INIT('hc8)
	) name328 (
		\b3_pad ,
		_w232_,
		_w489_,
		_w502_
	);
	LUT4 #(
		.INIT('h4445)
	) name329 (
		\b3_pad ,
		g_pad,
		_w215_,
		_w208_,
		_w503_
	);
	LUT3 #(
		.INIT('h01)
	) name330 (
		_w242_,
		_w491_,
		_w503_,
		_w504_
	);
	LUT4 #(
		.INIT('h8488)
	) name331 (
		\c3_pad ,
		_w234_,
		_w502_,
		_w504_,
		_w505_
	);
	LUT3 #(
		.INIT('h9a)
	) name332 (
		\b4_pad ,
		\g0_pad ,
		_w180_,
		_w506_
	);
	LUT4 #(
		.INIT('h4888)
	) name333 (
		\c4_pad ,
		_w327_,
		_w495_,
		_w506_,
		_w507_
	);
	LUT4 #(
		.INIT('hcc80)
	) name334 (
		\r4_pad ,
		\t3_pad ,
		_w279_,
		_w326_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		z_pad,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('hb)
	) name336 (
		_w507_,
		_w509_,
		_w510_
	);
	LUT3 #(
		.INIT('h8c)
	) name337 (
		\b5_pad ,
		\d5_pad ,
		\i10_pad ,
		_w511_
	);
	LUT4 #(
		.INIT('heac0)
	) name338 (
		_w189_,
		_w176_,
		_w181_,
		_w511_,
		_w512_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name339 (
		_w174_,
		_w177_,
		_w274_,
		_w304_,
		_w513_
	);
	LUT3 #(
		.INIT('h07)
	) name340 (
		_w177_,
		_w260_,
		_w326_,
		_w514_
	);
	LUT2 #(
		.INIT('hb)
	) name341 (
		_w513_,
		_w514_,
		_w515_
	);
	LUT3 #(
		.INIT('h48)
	) name342 (
		\d1_pad ,
		_w368_,
		_w499_,
		_w516_
	);
	LUT3 #(
		.INIT('h80)
	) name343 (
		\b2_pad ,
		\c2_pad ,
		\d2_pad ,
		_w517_
	);
	LUT4 #(
		.INIT('hdfec)
	) name344 (
		\b2_pad ,
		b_pad,
		\c2_pad ,
		\d2_pad ,
		_w518_
	);
	LUT4 #(
		.INIT('h999a)
	) name345 (
		\c3_pad ,
		g_pad,
		_w215_,
		_w208_,
		_w519_
	);
	LUT3 #(
		.INIT('h40)
	) name346 (
		_w502_,
		_w504_,
		_w519_,
		_w520_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name347 (
		\d3_pad ,
		_w234_,
		_w235_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('hd)
	) name348 (
		\d4_pad ,
		z_pad,
		_w522_
	);
	LUT4 #(
		.INIT('h0f08)
	) name349 (
		\e5_pad ,
		_w189_,
		_w176_,
		_w178_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		l_pad,
		\q1_pad ,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		l_pad,
		\p1_pad ,
		_w525_
	);
	LUT4 #(
		.INIT('h5700)
	) name352 (
		\g2_pad ,
		_w517_,
		_w524_,
		_w525_,
		_w526_
	);
	LUT3 #(
		.INIT('h08)
	) name353 (
		\e2_pad ,
		\n2_pad ,
		_w526_,
		_w527_
	);
	LUT4 #(
		.INIT('h0f07)
	) name354 (
		\e2_pad ,
		\n2_pad ,
		_w344_,
		_w526_,
		_w528_
	);
	LUT4 #(
		.INIT('h0a05)
	) name355 (
		\e2_pad ,
		\n2_pad ,
		_w344_,
		_w526_,
		_w529_
	);
	LUT4 #(
		.INIT('hffae)
	) name356 (
		b_pad,
		\s1_pad ,
		_w528_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\c3_pad ,
		\d3_pad ,
		_w531_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name358 (
		\b3_pad ,
		_w232_,
		_w489_,
		_w531_,
		_w532_
	);
	LUT4 #(
		.INIT('h00ab)
	) name359 (
		g_pad,
		_w215_,
		_w208_,
		_w415_,
		_w533_
	);
	LUT4 #(
		.INIT('h0001)
	) name360 (
		_w242_,
		_w491_,
		_w503_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('h8488)
	) name361 (
		\e3_pad ,
		_w234_,
		_w532_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('he)
	) name362 (
		_w235_,
		_w535_,
		_w536_
	);
	LUT3 #(
		.INIT('hf6)
	) name363 (
		\d4_pad ,
		\e4_pad ,
		z_pad,
		_w537_
	);
	LUT4 #(
		.INIT('h3132)
	) name364 (
		\h5_pad ,
		z_pad,
		_w187_,
		_w302_,
		_w538_
	);
	LUT4 #(
		.INIT('h1110)
	) name365 (
		\h5_pad ,
		z_pad,
		_w187_,
		_w302_,
		_w539_
	);
	LUT4 #(
		.INIT('h010a)
	) name366 (
		\f5_pad ,
		\p10_pad ,
		_w187_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('he)
	) name367 (
		z_pad,
		_w540_,
		_w541_
	);
	LUT3 #(
		.INIT('hc6)
	) name368 (
		\e2_pad ,
		\f2_pad ,
		_w526_,
		_w542_
	);
	LUT4 #(
		.INIT('hfeae)
	) name369 (
		b_pad,
		\t1_pad ,
		_w528_,
		_w542_,
		_w543_
	);
	LUT4 #(
		.INIT('h4844)
	) name370 (
		\f3_pad ,
		_w261_,
		_w280_,
		_w282_,
		_w544_
	);
	LUT4 #(
		.INIT('hff78)
	) name371 (
		\d4_pad ,
		\e4_pad ,
		\f4_pad ,
		z_pad,
		_w545_
	);
	LUT4 #(
		.INIT('h0503)
	) name372 (
		\f5_pad ,
		\p10_pad ,
		_w187_,
		_w539_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		z_pad,
		_w546_,
		_w547_
	);
	LUT4 #(
		.INIT('hbbbe)
	) name374 (
		b_pad,
		\g2_pad ,
		_w517_,
		_w524_,
		_w548_
	);
	LUT4 #(
		.INIT('h6066)
	) name375 (
		\f3_pad ,
		_w259_,
		_w280_,
		_w282_,
		_w549_
	);
	LUT3 #(
		.INIT('h48)
	) name376 (
		\g3_pad ,
		_w261_,
		_w549_,
		_w550_
	);
	LUT4 #(
		.INIT('h0f07)
	) name377 (
		\g4_pad ,
		\p4_pad ,
		_w188_,
		_w301_,
		_w551_
	);
	LUT4 #(
		.INIT('h0a05)
	) name378 (
		\g4_pad ,
		\p4_pad ,
		_w188_,
		_w301_,
		_w552_
	);
	LUT4 #(
		.INIT('hffce)
	) name379 (
		\u3_pad ,
		z_pad,
		_w551_,
		_w552_,
		_w553_
	);
	LUT3 #(
		.INIT('h8c)
	) name380 (
		\f1_pad ,
		\h1_pad ,
		\m6_pad ,
		_w554_
	);
	LUT4 #(
		.INIT('hf888)
	) name381 (
		_w204_,
		_w236_,
		_w345_,
		_w554_,
		_w555_
	);
	LUT4 #(
		.INIT('h0f07)
	) name382 (
		\e2_pad ,
		\f2_pad ,
		\h2_pad ,
		_w526_,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		\f2_pad ,
		\h2_pad ,
		_w557_
	);
	LUT3 #(
		.INIT('h20)
	) name384 (
		\e2_pad ,
		_w526_,
		_w557_,
		_w558_
	);
	LUT3 #(
		.INIT('h02)
	) name385 (
		_w528_,
		_w556_,
		_w558_,
		_w559_
	);
	LUT3 #(
		.INIT('h51)
	) name386 (
		b_pad,
		\u1_pad ,
		_w528_,
		_w560_
	);
	LUT2 #(
		.INIT('hb)
	) name387 (
		_w559_,
		_w560_,
		_w561_
	);
	LUT4 #(
		.INIT('hab00)
	) name388 (
		\e0_pad ,
		_w180_,
		_w257_,
		_w285_,
		_w562_
	);
	LUT4 #(
		.INIT('h5400)
	) name389 (
		\e0_pad ,
		_w180_,
		_w257_,
		_w265_,
		_w563_
	);
	LUT4 #(
		.INIT('h000b)
	) name390 (
		_w280_,
		_w282_,
		_w563_,
		_w562_,
		_w564_
	);
	LUT3 #(
		.INIT('h48)
	) name391 (
		\h3_pad ,
		_w261_,
		_w564_,
		_w565_
	);
	LUT3 #(
		.INIT('hc6)
	) name392 (
		\g4_pad ,
		\h4_pad ,
		_w301_,
		_w566_
	);
	LUT4 #(
		.INIT('hfece)
	) name393 (
		\v3_pad ,
		z_pad,
		_w551_,
		_w566_,
		_w567_
	);
	LUT4 #(
		.INIT('h3230)
	) name394 (
		\i1_pad ,
		_w204_,
		_w206_,
		_w345_,
		_w568_
	);
	LUT4 #(
		.INIT('h0800)
	) name395 (
		\e2_pad ,
		\i2_pad ,
		_w526_,
		_w557_,
		_w569_
	);
	LUT3 #(
		.INIT('h48)
	) name396 (
		\i2_pad ,
		_w528_,
		_w558_,
		_w570_
	);
	LUT3 #(
		.INIT('h51)
	) name397 (
		b_pad,
		\v1_pad ,
		_w528_,
		_w571_
	);
	LUT2 #(
		.INIT('hb)
	) name398 (
		_w570_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		_w259_,
		_w287_,
		_w573_
	);
	LUT4 #(
		.INIT('h7077)
	) name400 (
		_w259_,
		_w269_,
		_w280_,
		_w282_,
		_w574_
	);
	LUT4 #(
		.INIT('h8488)
	) name401 (
		\i3_pad ,
		_w261_,
		_w573_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('he)
	) name402 (
		_w262_,
		_w575_,
		_w576_
	);
	LUT4 #(
		.INIT('hddde)
	) name403 (
		\i4_pad ,
		z_pad,
		_w298_,
		_w299_,
		_w577_
	);
	LUT3 #(
		.INIT('h0b)
	) name404 (
		\j5_pad ,
		\k5_pad ,
		z_pad,
		_w578_
	);
	LUT3 #(
		.INIT('h60)
	) name405 (
		\j5_pad ,
		_w174_,
		_w578_,
		_w579_
	);
	LUT4 #(
		.INIT('h0080)
	) name406 (
		\e2_pad ,
		\n2_pad ,
		\r6_pad ,
		_w526_,
		_w580_
	);
	LUT4 #(
		.INIT('hf1f4)
	) name407 (
		b_pad,
		\r6_pad ,
		_w223_,
		_w527_,
		_w581_
	);
	LUT4 #(
		.INIT('h8000)
	) name408 (
		\f2_pad ,
		\h2_pad ,
		\i2_pad ,
		\j2_pad ,
		_w582_
	);
	LUT3 #(
		.INIT('h20)
	) name409 (
		\e2_pad ,
		_w526_,
		_w582_,
		_w583_
	);
	LUT4 #(
		.INIT('h00c8)
	) name410 (
		\j2_pad ,
		_w528_,
		_w569_,
		_w583_,
		_w584_
	);
	LUT3 #(
		.INIT('h51)
	) name411 (
		b_pad,
		\w1_pad ,
		_w528_,
		_w585_
	);
	LUT2 #(
		.INIT('hb)
	) name412 (
		_w584_,
		_w585_,
		_w586_
	);
	LUT4 #(
		.INIT('h0001)
	) name413 (
		\l3_pad ,
		\m3_pad ,
		\n3_pad ,
		\o3_pad ,
		_w587_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		_w261_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w262_,
		_w588_,
		_w589_
	);
	LUT4 #(
		.INIT('h0f07)
	) name416 (
		\g4_pad ,
		\h4_pad ,
		\j4_pad ,
		_w301_,
		_w590_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\h4_pad ,
		\j4_pad ,
		_w591_
	);
	LUT3 #(
		.INIT('h20)
	) name418 (
		\g4_pad ,
		_w301_,
		_w591_,
		_w592_
	);
	LUT3 #(
		.INIT('h02)
	) name419 (
		_w551_,
		_w590_,
		_w592_,
		_w593_
	);
	LUT3 #(
		.INIT('h31)
	) name420 (
		\w3_pad ,
		z_pad,
		_w551_,
		_w594_
	);
	LUT2 #(
		.INIT('hb)
	) name421 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT4 #(
		.INIT('h0208)
	) name422 (
		\j5_pad ,
		\k5_pad ,
		z_pad,
		_w174_,
		_w596_
	);
	LUT4 #(
		.INIT('h3133)
	) name423 (
		\e2_pad ,
		l_pad,
		_w526_,
		_w582_,
		_w597_
	);
	LUT3 #(
		.INIT('h84)
	) name424 (
		\k2_pad ,
		_w528_,
		_w597_,
		_w598_
	);
	LUT3 #(
		.INIT('h51)
	) name425 (
		b_pad,
		\x1_pad ,
		_w528_,
		_w599_
	);
	LUT2 #(
		.INIT('hb)
	) name426 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT4 #(
		.INIT('h8000)
	) name427 (
		\l3_pad ,
		\m3_pad ,
		\n3_pad ,
		\o3_pad ,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		_w261_,
		_w601_,
		_w602_
	);
	LUT4 #(
		.INIT('h0800)
	) name429 (
		\g4_pad ,
		\k4_pad ,
		_w301_,
		_w591_,
		_w603_
	);
	LUT3 #(
		.INIT('h48)
	) name430 (
		\k4_pad ,
		_w551_,
		_w592_,
		_w604_
	);
	LUT3 #(
		.INIT('h31)
	) name431 (
		\x3_pad ,
		z_pad,
		_w551_,
		_w605_
	);
	LUT2 #(
		.INIT('hb)
	) name432 (
		_w604_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		\o2_pad ,
		s_pad,
		_w607_
	);
	LUT4 #(
		.INIT('h135f)
	) name434 (
		o_pad,
		r_pad,
		\t2_pad ,
		\u1_pad ,
		_w608_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		_w607_,
		_w608_,
		_w609_
	);
	LUT4 #(
		.INIT('h135f)
	) name436 (
		\j2_pad ,
		q_pad,
		t_pad,
		\x1_pad ,
		_w610_
	);
	LUT4 #(
		.INIT('h153f)
	) name437 (
		\a3_pad ,
		\e3_pad ,
		m_pad,
		n_pad,
		_w611_
	);
	LUT4 #(
		.INIT('h0777)
	) name438 (
		\a2_pad ,
		p_pad,
		w_pad,
		\y0_pad ,
		_w612_
	);
	LUT4 #(
		.INIT('h153f)
	) name439 (
		\d1_pad ,
		\g2_pad ,
		u_pad,
		v_pad,
		_w613_
	);
	LUT4 #(
		.INIT('h8000)
	) name440 (
		_w612_,
		_w613_,
		_w610_,
		_w611_,
		_w614_
	);
	LUT2 #(
		.INIT('h7)
	) name441 (
		_w609_,
		_w614_,
		_w615_
	);
	LUT3 #(
		.INIT('h08)
	) name442 (
		\k2_pad ,
		\l2_pad ,
		_w597_,
		_w616_
	);
	LUT4 #(
		.INIT('hc060)
	) name443 (
		\k2_pad ,
		\l2_pad ,
		_w528_,
		_w597_,
		_w617_
	);
	LUT3 #(
		.INIT('h51)
	) name444 (
		b_pad,
		\y1_pad ,
		_w528_,
		_w618_
	);
	LUT2 #(
		.INIT('hb)
	) name445 (
		_w617_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		_w259_,
		_w271_,
		_w620_
	);
	LUT4 #(
		.INIT('h8acf)
	) name447 (
		_w259_,
		_w280_,
		_w282_,
		_w288_,
		_w621_
	);
	LUT4 #(
		.INIT('h8488)
	) name448 (
		\l3_pad ,
		_w261_,
		_w620_,
		_w621_,
		_w622_
	);
	LUT4 #(
		.INIT('h8000)
	) name449 (
		\h4_pad ,
		\j4_pad ,
		\k4_pad ,
		\l4_pad ,
		_w623_
	);
	LUT3 #(
		.INIT('h20)
	) name450 (
		\g4_pad ,
		_w301_,
		_w623_,
		_w624_
	);
	LUT4 #(
		.INIT('h00c8)
	) name451 (
		\l4_pad ,
		_w551_,
		_w603_,
		_w624_,
		_w625_
	);
	LUT3 #(
		.INIT('h31)
	) name452 (
		\y3_pad ,
		z_pad,
		_w551_,
		_w626_
	);
	LUT2 #(
		.INIT('hb)
	) name453 (
		_w625_,
		_w626_,
		_w627_
	);
	LUT4 #(
		.INIT('h0545)
	) name454 (
		\a0_pad ,
		\r5_pad ,
		\z4_pad ,
		_w413_,
		_w628_
	);
	LUT4 #(
		.INIT('h0222)
	) name455 (
		_w174_,
		_w177_,
		_w310_,
		_w311_,
		_w629_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name456 (
		\l5_pad ,
		\m5_pad ,
		\n5_pad ,
		z_pad,
		_w630_
	);
	LUT3 #(
		.INIT('h20)
	) name457 (
		_w337_,
		_w629_,
		_w630_,
		_w631_
	);
	LUT4 #(
		.INIT('h0455)
	) name458 (
		z_pad,
		_w190_,
		_w628_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		\m2_pad ,
		s_pad,
		_w633_
	);
	LUT4 #(
		.INIT('h135f)
	) name460 (
		o_pad,
		q_pad,
		\s2_pad ,
		\w1_pad ,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT4 #(
		.INIT('h153f)
	) name462 (
		\i2_pad ,
		r_pad,
		\t1_pad ,
		t_pad,
		_w636_
	);
	LUT4 #(
		.INIT('h0777)
	) name463 (
		\d3_pad ,
		m_pad,
		n_pad,
		\z2_pad ,
		_w637_
	);
	LUT4 #(
		.INIT('h153f)
	) name464 (
		p_pad,
		w_pad,
		\x0_pad ,
		\z1_pad ,
		_w638_
	);
	LUT4 #(
		.INIT('h153f)
	) name465 (
		\c1_pad ,
		\d2_pad ,
		u_pad,
		v_pad,
		_w639_
	);
	LUT4 #(
		.INIT('h8000)
	) name466 (
		_w638_,
		_w639_,
		_w636_,
		_w637_,
		_w640_
	);
	LUT2 #(
		.INIT('h7)
	) name467 (
		_w635_,
		_w640_,
		_w641_
	);
	LUT4 #(
		.INIT('h1151)
	) name468 (
		c_pad,
		\d1_pad ,
		\r1_pad ,
		_w499_,
		_w642_
	);
	LUT3 #(
		.INIT('h04)
	) name469 (
		\e3_pad ,
		\y2_pad ,
		\z2_pad ,
		_w643_
	);
	LUT4 #(
		.INIT('h0001)
	) name470 (
		\a3_pad ,
		\b3_pad ,
		\c3_pad ,
		\d3_pad ,
		_w644_
	);
	LUT4 #(
		.INIT('h0444)
	) name471 (
		_w205_,
		_w239_,
		_w643_,
		_w644_,
		_w645_
	);
	LUT4 #(
		.INIT('h0100)
	) name472 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w646_
	);
	LUT4 #(
		.INIT('h007f)
	) name473 (
		_w239_,
		_w643_,
		_w644_,
		_w646_,
		_w647_
	);
	LUT4 #(
		.INIT('h0fef)
	) name474 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w648_
	);
	LUT3 #(
		.INIT('h20)
	) name475 (
		_w647_,
		_w645_,
		_w648_,
		_w649_
	);
	LUT4 #(
		.INIT('h0455)
	) name476 (
		b_pad,
		_w214_,
		_w642_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('h0080)
	) name477 (
		\k2_pad ,
		\l2_pad ,
		\m2_pad ,
		_w597_,
		_w651_
	);
	LUT3 #(
		.INIT('h51)
	) name478 (
		b_pad,
		\z1_pad ,
		_w528_,
		_w652_
	);
	LUT4 #(
		.INIT('h48ff)
	) name479 (
		\m2_pad ,
		_w528_,
		_w616_,
		_w652_,
		_w653_
	);
	LUT4 #(
		.INIT('h999c)
	) name480 (
		\e0_pad ,
		\l3_pad ,
		_w180_,
		_w257_,
		_w654_
	);
	LUT3 #(
		.INIT('h40)
	) name481 (
		_w620_,
		_w621_,
		_w654_,
		_w655_
	);
	LUT3 #(
		.INIT('h48)
	) name482 (
		\m3_pad ,
		_w261_,
		_w655_,
		_w656_
	);
	LUT4 #(
		.INIT('h3133)
	) name483 (
		\g4_pad ,
		\j0_pad ,
		_w301_,
		_w623_,
		_w657_
	);
	LUT3 #(
		.INIT('h84)
	) name484 (
		\m4_pad ,
		_w551_,
		_w657_,
		_w658_
	);
	LUT3 #(
		.INIT('h31)
	) name485 (
		\z3_pad ,
		z_pad,
		_w551_,
		_w659_
	);
	LUT2 #(
		.INIT('hb)
	) name486 (
		_w658_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		\l2_pad ,
		s_pad,
		_w661_
	);
	LUT4 #(
		.INIT('h135f)
	) name488 (
		o_pad,
		q_pad,
		\r2_pad ,
		\v1_pad ,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		_w661_,
		_w662_,
		_w663_
	);
	LUT4 #(
		.INIT('h153f)
	) name490 (
		\h2_pad ,
		r_pad,
		\s1_pad ,
		t_pad,
		_w664_
	);
	LUT4 #(
		.INIT('h0777)
	) name491 (
		\c3_pad ,
		m_pad,
		n_pad,
		\y2_pad ,
		_w665_
	);
	LUT4 #(
		.INIT('h153f)
	) name492 (
		p_pad,
		\w0_pad ,
		w_pad,
		\y1_pad ,
		_w666_
	);
	LUT4 #(
		.INIT('h153f)
	) name493 (
		\b1_pad ,
		\c2_pad ,
		u_pad,
		v_pad,
		_w667_
	);
	LUT4 #(
		.INIT('h8000)
	) name494 (
		_w666_,
		_w667_,
		_w664_,
		_w665_,
		_w668_
	);
	LUT2 #(
		.INIT('h7)
	) name495 (
		_w663_,
		_w668_,
		_w669_
	);
	LUT4 #(
		.INIT('h8000)
	) name496 (
		\k2_pad ,
		\l2_pad ,
		\m2_pad ,
		\o2_pad ,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w582_,
		_w670_,
		_w671_
	);
	LUT3 #(
		.INIT('he0)
	) name498 (
		b_pad,
		_w528_,
		_w671_,
		_w672_
	);
	LUT4 #(
		.INIT('h999c)
	) name499 (
		\e0_pad ,
		\m3_pad ,
		_w180_,
		_w257_,
		_w673_
	);
	LUT4 #(
		.INIT('h4000)
	) name500 (
		_w620_,
		_w621_,
		_w654_,
		_w673_,
		_w674_
	);
	LUT3 #(
		.INIT('h48)
	) name501 (
		\n3_pad ,
		_w261_,
		_w674_,
		_w675_
	);
	LUT3 #(
		.INIT('h08)
	) name502 (
		\m4_pad ,
		\n4_pad ,
		_w657_,
		_w676_
	);
	LUT4 #(
		.INIT('hc060)
	) name503 (
		\m4_pad ,
		\n4_pad ,
		_w551_,
		_w657_,
		_w677_
	);
	LUT3 #(
		.INIT('h31)
	) name504 (
		\a4_pad ,
		z_pad,
		_w551_,
		_w678_
	);
	LUT2 #(
		.INIT('hb)
	) name505 (
		_w677_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		\k2_pad ,
		s_pad,
		_w680_
	);
	LUT4 #(
		.INIT('h153f)
	) name507 (
		\m1_pad ,
		o_pad,
		\q2_pad ,
		r_pad,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name508 (
		_w680_,
		_w681_,
		_w682_
	);
	LUT4 #(
		.INIT('h153f)
	) name509 (
		\f2_pad ,
		q_pad,
		\r1_pad ,
		t_pad,
		_w683_
	);
	LUT4 #(
		.INIT('h0777)
	) name510 (
		\b3_pad ,
		m_pad,
		n_pad,
		\x2_pad ,
		_w684_
	);
	LUT4 #(
		.INIT('h0777)
	) name511 (
		\p1_pad ,
		p_pad,
		\v0_pad ,
		w_pad,
		_w685_
	);
	LUT4 #(
		.INIT('h153f)
	) name512 (
		\a1_pad ,
		\b2_pad ,
		u_pad,
		v_pad,
		_w686_
	);
	LUT4 #(
		.INIT('h8000)
	) name513 (
		_w685_,
		_w686_,
		_w683_,
		_w684_,
		_w687_
	);
	LUT2 #(
		.INIT('h7)
	) name514 (
		_w682_,
		_w687_,
		_w688_
	);
	LUT3 #(
		.INIT('h8a)
	) name515 (
		_w528_,
		_w597_,
		_w670_,
		_w689_
	);
	LUT3 #(
		.INIT('h31)
	) name516 (
		\a2_pad ,
		b_pad,
		_w528_,
		_w690_
	);
	LUT4 #(
		.INIT('he0ff)
	) name517 (
		\o2_pad ,
		_w651_,
		_w689_,
		_w690_,
		_w691_
	);
	LUT4 #(
		.INIT('h999c)
	) name518 (
		\e0_pad ,
		\n3_pad ,
		_w180_,
		_w257_,
		_w692_
	);
	LUT4 #(
		.INIT('h4888)
	) name519 (
		\o3_pad ,
		_w261_,
		_w674_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('he)
	) name520 (
		_w262_,
		_w693_,
		_w694_
	);
	LUT4 #(
		.INIT('h0080)
	) name521 (
		\m4_pad ,
		\n4_pad ,
		\o4_pad ,
		_w657_,
		_w695_
	);
	LUT3 #(
		.INIT('h31)
	) name522 (
		\b4_pad ,
		z_pad,
		_w551_,
		_w696_
	);
	LUT4 #(
		.INIT('h48ff)
	) name523 (
		\o4_pad ,
		_w551_,
		_w676_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		\b0_pad ,
		_w336_,
		_w698_
	);
	LUT3 #(
		.INIT('h04)
	) name525 (
		\c0_pad ,
		\p5_pad ,
		_w339_,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT4 #(
		.INIT('h0016)
	) name527 (
		\p5_pad ,
		\q5_pad ,
		\r5_pad ,
		z_pad,
		_w701_
	);
	LUT3 #(
		.INIT('hc8)
	) name528 (
		\c0_pad ,
		\r5_pad ,
		_w339_,
		_w702_
	);
	LUT3 #(
		.INIT('hc8)
	) name529 (
		\b0_pad ,
		\q5_pad ,
		_w336_,
		_w703_
	);
	LUT3 #(
		.INIT('h10)
	) name530 (
		_w702_,
		_w703_,
		_w701_,
		_w704_
	);
	LUT2 #(
		.INIT('hb)
	) name531 (
		_w700_,
		_w704_,
		_w705_
	);
	LUT3 #(
		.INIT('h20)
	) name532 (
		u_pad,
		_w238_,
		_w241_,
		_w706_
	);
	LUT4 #(
		.INIT('h0080)
	) name533 (
		\e2_pad ,
		\n2_pad ,
		s_pad,
		_w526_,
		_w707_
	);
	LUT2 #(
		.INIT('h2)
	) name534 (
		q_pad,
		_w234_,
		_w708_
	);
	LUT3 #(
		.INIT('h80)
	) name535 (
		m_pad,
		_w643_,
		_w644_,
		_w709_
	);
	LUT4 #(
		.INIT('h8000)
	) name536 (
		\c3_pad ,
		\d3_pad ,
		\e3_pad ,
		o_pad,
		_w710_
	);
	LUT4 #(
		.INIT('h153f)
	) name537 (
		\e2_pad ,
		p_pad,
		\q1_pad ,
		t_pad,
		_w711_
	);
	LUT4 #(
		.INIT('h135f)
	) name538 (
		\l1_pad ,
		v_pad,
		w_pad,
		\z0_pad ,
		_w712_
	);
	LUT4 #(
		.INIT('h135f)
	) name539 (
		\n1_pad ,
		n_pad,
		r_pad,
		\w2_pad ,
		_w713_
	);
	LUT4 #(
		.INIT('h4000)
	) name540 (
		_w710_,
		_w711_,
		_w712_,
		_w713_,
		_w714_
	);
	LUT3 #(
		.INIT('h10)
	) name541 (
		_w708_,
		_w709_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w707_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('hb)
	) name543 (
		_w706_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		d_pad,
		_w646_,
		_w718_
	);
	LUT4 #(
		.INIT('h4000)
	) name545 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w719_
	);
	LUT3 #(
		.INIT('h04)
	) name546 (
		e_pad,
		\p1_pad ,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		_w718_,
		_w720_,
		_w721_
	);
	LUT4 #(
		.INIT('h0114)
	) name548 (
		b_pad,
		\p1_pad ,
		\q1_pad ,
		\r1_pad ,
		_w722_
	);
	LUT3 #(
		.INIT('hc8)
	) name549 (
		e_pad,
		\r1_pad ,
		_w719_,
		_w723_
	);
	LUT3 #(
		.INIT('hc8)
	) name550 (
		d_pad,
		\q1_pad ,
		_w646_,
		_w724_
	);
	LUT3 #(
		.INIT('h10)
	) name551 (
		_w723_,
		_w724_,
		_w722_,
		_w725_
	);
	LUT2 #(
		.INIT('hb)
	) name552 (
		_w721_,
		_w725_,
		_w726_
	);
	LUT3 #(
		.INIT('h5c)
	) name553 (
		\l6_pad ,
		\p2_pad ,
		_w580_,
		_w727_
	);
	LUT3 #(
		.INIT('hc4)
	) name554 (
		\j3_pad ,
		_w259_,
		_w271_,
		_w728_
	);
	LUT3 #(
		.INIT('h31)
	) name555 (
		\k3_pad ,
		_w259_,
		_w288_,
		_w729_
	);
	LUT3 #(
		.INIT('h01)
	) name556 (
		_w283_,
		_w729_,
		_w728_,
		_w730_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name557 (
		\p3_pad ,
		_w261_,
		_w262_,
		_w730_,
		_w731_
	);
	LUT4 #(
		.INIT('h8000)
	) name558 (
		\m4_pad ,
		\n4_pad ,
		\o4_pad ,
		\q4_pad ,
		_w732_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w623_,
		_w732_,
		_w733_
	);
	LUT3 #(
		.INIT('he0)
	) name560 (
		z_pad,
		_w551_,
		_w733_,
		_w734_
	);
	LUT3 #(
		.INIT('h04)
	) name561 (
		\c0_pad ,
		\q5_pad ,
		_w339_,
		_w735_
	);
	LUT3 #(
		.INIT('hc8)
	) name562 (
		\c0_pad ,
		\p5_pad ,
		_w339_,
		_w736_
	);
	LUT4 #(
		.INIT('h010d)
	) name563 (
		\r5_pad ,
		_w698_,
		_w736_,
		_w735_,
		_w737_
	);
	LUT2 #(
		.INIT('h2)
	) name564 (
		_w701_,
		_w737_,
		_w738_
	);
	LUT4 #(
		.INIT('hbffb)
	) name565 (
		b_pad,
		\l1_pad ,
		\m1_pad ,
		\n1_pad ,
		_w739_
	);
	LUT4 #(
		.INIT('h7f00)
	) name566 (
		_w205_,
		_w239_,
		_w416_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h7)
	) name567 (
		_w647_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		\q0_pad ,
		\q4_pad ,
		_w742_
	);
	LUT4 #(
		.INIT('h0777)
	) name569 (
		\i3_pad ,
		\m0_pad ,
		\p0_pad ,
		\w3_pad ,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name570 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT4 #(
		.INIT('h135f)
	) name571 (
		\l4_pad ,
		\o0_pad ,
		\r0_pad ,
		\z3_pad ,
		_w745_
	);
	LUT4 #(
		.INIT('h153f)
	) name572 (
		\k0_pad ,
		\l0_pad ,
		\p3_pad ,
		\t3_pad ,
		_w746_
	);
	LUT4 #(
		.INIT('h0777)
	) name573 (
		\c4_pad ,
		\n0_pad ,
		\u0_pad ,
		\u4_pad ,
		_w747_
	);
	LUT4 #(
		.INIT('h0777)
	) name574 (
		\i4_pad ,
		\s0_pad ,
		\t0_pad ,
		\z4_pad ,
		_w748_
	);
	LUT4 #(
		.INIT('h8000)
	) name575 (
		_w747_,
		_w748_,
		_w745_,
		_w746_,
		_w749_
	);
	LUT2 #(
		.INIT('h7)
	) name576 (
		_w744_,
		_w749_,
		_w750_
	);
	LUT3 #(
		.INIT('h04)
	) name577 (
		e_pad,
		\q1_pad ,
		_w719_,
		_w751_
	);
	LUT3 #(
		.INIT('hc8)
	) name578 (
		e_pad,
		\p1_pad ,
		_w719_,
		_w752_
	);
	LUT4 #(
		.INIT('h010d)
	) name579 (
		\r1_pad ,
		_w718_,
		_w752_,
		_w751_,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		_w722_,
		_w753_,
		_w754_
	);
	LUT4 #(
		.INIT('h4844)
	) name581 (
		\q2_pad ,
		_w234_,
		_w238_,
		_w241_,
		_w755_
	);
	LUT4 #(
		.INIT('h0007)
	) name582 (
		_w259_,
		_w272_,
		_w283_,
		_w290_,
		_w756_
	);
	LUT4 #(
		.INIT('hf4f8)
	) name583 (
		\q3_pad ,
		_w261_,
		_w262_,
		_w756_,
		_w757_
	);
	LUT3 #(
		.INIT('h8a)
	) name584 (
		_w551_,
		_w657_,
		_w732_,
		_w758_
	);
	LUT3 #(
		.INIT('h31)
	) name585 (
		\c4_pad ,
		z_pad,
		_w551_,
		_w759_
	);
	LUT4 #(
		.INIT('he0ff)
	) name586 (
		\q4_pad ,
		_w695_,
		_w758_,
		_w759_,
		_w760_
	);
	LUT3 #(
		.INIT('h04)
	) name587 (
		\c0_pad ,
		\r5_pad ,
		_w339_,
		_w761_
	);
	LUT3 #(
		.INIT('hc8)
	) name588 (
		\c0_pad ,
		\q5_pad ,
		_w339_,
		_w762_
	);
	LUT4 #(
		.INIT('h010d)
	) name589 (
		\p5_pad ,
		_w698_,
		_w762_,
		_w761_,
		_w763_
	);
	LUT2 #(
		.INIT('h2)
	) name590 (
		_w701_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		\o4_pad ,
		\q0_pad ,
		_w765_
	);
	LUT4 #(
		.INIT('h0777)
	) name592 (
		\h3_pad ,
		\m0_pad ,
		\p0_pad ,
		\v3_pad ,
		_w766_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w765_,
		_w766_,
		_w767_
	);
	LUT4 #(
		.INIT('h135f)
	) name594 (
		\k4_pad ,
		\o0_pad ,
		\r0_pad ,
		\y3_pad ,
		_w768_
	);
	LUT4 #(
		.INIT('h153f)
	) name595 (
		\k0_pad ,
		\l0_pad ,
		\o3_pad ,
		\s3_pad ,
		_w769_
	);
	LUT4 #(
		.INIT('h0777)
	) name596 (
		\b4_pad ,
		\n0_pad ,
		\t4_pad ,
		\u0_pad ,
		_w770_
	);
	LUT4 #(
		.INIT('h0777)
	) name597 (
		\f4_pad ,
		\s0_pad ,
		\t0_pad ,
		\y4_pad ,
		_w771_
	);
	LUT4 #(
		.INIT('h8000)
	) name598 (
		_w770_,
		_w771_,
		_w768_,
		_w769_,
		_w772_
	);
	LUT2 #(
		.INIT('h7)
	) name599 (
		_w767_,
		_w772_,
		_w773_
	);
	LUT3 #(
		.INIT('h04)
	) name600 (
		e_pad,
		\r1_pad ,
		_w719_,
		_w774_
	);
	LUT3 #(
		.INIT('hc8)
	) name601 (
		e_pad,
		\q1_pad ,
		_w719_,
		_w775_
	);
	LUT4 #(
		.INIT('h010d)
	) name602 (
		\p1_pad ,
		_w718_,
		_w775_,
		_w774_,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name603 (
		_w722_,
		_w776_,
		_w777_
	);
	LUT4 #(
		.INIT('h6066)
	) name604 (
		\q2_pad ,
		_w232_,
		_w238_,
		_w241_,
		_w778_
	);
	LUT3 #(
		.INIT('h48)
	) name605 (
		\r2_pad ,
		_w234_,
		_w778_,
		_w779_
	);
	LUT3 #(
		.INIT('hc8)
	) name606 (
		\q3_pad ,
		_w259_,
		_w272_,
		_w780_
	);
	LUT4 #(
		.INIT('h2223)
	) name607 (
		\e0_pad ,
		\q3_pad ,
		_w180_,
		_w257_,
		_w781_
	);
	LUT3 #(
		.INIT('h01)
	) name608 (
		_w283_,
		_w290_,
		_w781_,
		_w782_
	);
	LUT4 #(
		.INIT('h8488)
	) name609 (
		\r3_pad ,
		_w261_,
		_w780_,
		_w782_,
		_w783_
	);
	LUT3 #(
		.INIT('h84)
	) name610 (
		\r4_pad ,
		_w191_,
		_w183_,
		_w784_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		\n4_pad ,
		\q0_pad ,
		_w785_
	);
	LUT4 #(
		.INIT('h0777)
	) name612 (
		\g3_pad ,
		\m0_pad ,
		\p0_pad ,
		\u3_pad ,
		_w786_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT4 #(
		.INIT('h135f)
	) name614 (
		\j4_pad ,
		\o0_pad ,
		\r0_pad ,
		\x3_pad ,
		_w788_
	);
	LUT4 #(
		.INIT('h153f)
	) name615 (
		\k0_pad ,
		\l0_pad ,
		\n3_pad ,
		\r3_pad ,
		_w789_
	);
	LUT4 #(
		.INIT('h0777)
	) name616 (
		\a4_pad ,
		\n0_pad ,
		\s4_pad ,
		\u0_pad ,
		_w790_
	);
	LUT4 #(
		.INIT('h0777)
	) name617 (
		\e4_pad ,
		\s0_pad ,
		\t0_pad ,
		\x4_pad ,
		_w791_
	);
	LUT4 #(
		.INIT('h8000)
	) name618 (
		_w790_,
		_w791_,
		_w788_,
		_w789_,
		_w792_
	);
	LUT2 #(
		.INIT('h7)
	) name619 (
		_w787_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('h6366)
	) name620 (
		h_pad,
		\s1_pad ,
		_w213_,
		_w220_,
		_w794_
	);
	LUT4 #(
		.INIT('h5404)
	) name621 (
		b_pad,
		\w2_pad ,
		_w228_,
		_w794_,
		_w795_
	);
	LUT4 #(
		.INIT('hab00)
	) name622 (
		g_pad,
		_w215_,
		_w208_,
		_w245_,
		_w796_
	);
	LUT4 #(
		.INIT('h5400)
	) name623 (
		g_pad,
		_w215_,
		_w208_,
		_w251_,
		_w797_
	);
	LUT4 #(
		.INIT('h000b)
	) name624 (
		_w238_,
		_w241_,
		_w797_,
		_w796_,
		_w798_
	);
	LUT3 #(
		.INIT('h48)
	) name625 (
		\s2_pad ,
		_w234_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('h8488)
	) name626 (
		\s3_pad ,
		_w261_,
		_w273_,
		_w291_,
		_w800_
	);
	LUT2 #(
		.INIT('he)
	) name627 (
		_w262_,
		_w800_,
		_w801_
	);
	LUT4 #(
		.INIT('h1020)
	) name628 (
		\s4_pad ,
		_w186_,
		_w191_,
		_w184_,
		_w802_
	);
	assign \a10_pad  = _w194_ ;
	assign \a6_pad  = _w203_ ;
	assign \a7_pad  = _w231_ ;
	assign \a8_pad  = _w256_ ;
	assign \a9_pad  = _w294_ ;
	assign \b10_pad  = _w296_ ;
	assign \b6_pad  = _w316_ ;
	assign \b7_pad  = _w321_ ;
	assign \b8_pad  = _w325_ ;
	assign \b9_pad  = _w334_ ;
	assign \c10_pad  = _w335_ ;
	assign \c53  = _w341_ ;
	assign \c6_pad  = _w348_ ;
	assign \c7_pad  = _w355_ ;
	assign \c8_pad  = _w358_ ;
	assign \c9_pad  = _w364_ ;
	assign \d10_pad  = _w365_ ;
	assign \d6_pad  = _w369_ ;
	assign \d7_pad  = _w376_ ;
	assign \d8_pad  = _w381_ ;
	assign \d9_pad  = _w386_ ;
	assign \e10_pad  = _w391_ ;
	assign \e6_pad  = _w393_ ;
	assign \e7_pad  = _w400_ ;
	assign \e8_pad  = _w404_ ;
	assign \e9_pad  = _w412_ ;
	assign \f10_pad  = _w414_ ;
	assign \f22  = _w419_ ;
	assign \f6_pad  = _w420_ ;
	assign \f7_pad  = _w430_ ;
	assign \f8_pad  = _w434_ ;
	assign \f9_pad  = _w443_ ;
	assign \g10_pad  = _w444_ ;
	assign \g6_pad  = _w447_ ;
	assign \g7_pad  = _w454_ ;
	assign \g8_pad  = _w458_ ;
	assign \g9_pad  = _w466_ ;
	assign \h6_pad  = _w467_ ;
	assign \h7_pad  = _w473_ ;
	assign \h8_pad  = _w477_ ;
	assign \h9_pad  = _w485_ ;
	assign \i6_pad  = _w487_ ;
	assign \i7_pad  = _w488_ ;
	assign \i8_pad  = _w493_ ;
	assign \i9_pad  = _w498_ ;
	assign \j10_pad  = _w179_ ;
	assign \j6_pad  = _w500_ ;
	assign \j7_pad  = _w501_ ;
	assign \j8_pad  = _w505_ ;
	assign \j9_pad  = _w510_ ;
	assign \k10_pad  = _w512_ ;
	assign \k53  = _w515_ ;
	assign \k6_pad  = _w516_ ;
	assign \k7_pad  = _w518_ ;
	assign \k8_pad  = _w521_ ;
	assign \k9_pad  = _w522_ ;
	assign \l10_pad  = _w523_ ;
	assign \l7_pad  = _w530_ ;
	assign \l8_pad  = _w536_ ;
	assign \l9_pad  = _w537_ ;
	assign \m10_pad  = _w541_ ;
	assign \m7_pad  = _w543_ ;
	assign \m8_pad  = _w544_ ;
	assign \m9_pad  = _w545_ ;
	assign \n10_pad  = _w547_ ;
	assign \n6_pad  = _w207_ ;
	assign \n7_pad  = _w548_ ;
	assign \n8_pad  = _w550_ ;
	assign \n9_pad  = _w553_ ;
	assign \o10_pad  = _w538_ ;
	assign \o6_pad  = _w555_ ;
	assign \o7_pad  = _w561_ ;
	assign \o8_pad  = _w565_ ;
	assign \o9_pad  = _w567_ ;
	assign \p6_pad  = _w568_ ;
	assign \p7_pad  = _w572_ ;
	assign \p8_pad  = _w576_ ;
	assign \p9_pad  = _w577_ ;
	assign \q10_pad  = _w579_ ;
	assign \q6_pad  = _w581_ ;
	assign \q7_pad  = _w586_ ;
	assign \q8_pad  = _w589_ ;
	assign \q9_pad  = _w595_ ;
	assign \r10_pad  = _w596_ ;
	assign \r7_pad  = _w600_ ;
	assign \r8_pad  = _w602_ ;
	assign \r9_pad  = _w606_ ;
	assign \s5_pad  = _w615_ ;
	assign \s7_pad  = _w619_ ;
	assign \s8_pad  = _w622_ ;
	assign \s9_pad  = _w627_ ;
	assign \t10_pad  = _w632_ ;
	assign \t5_pad  = _w641_ ;
	assign \t6_pad  = _w650_ ;
	assign \t7_pad  = _w653_ ;
	assign \t8_pad  = _w656_ ;
	assign \t9_pad  = _w660_ ;
	assign \u5_pad  = _w669_ ;
	assign \u7_pad  = _w672_ ;
	assign \u8_pad  = _w675_ ;
	assign \u9_pad  = _w679_ ;
	assign \v10_pad  = _w258_ ;
	assign \v5_pad  = _w688_ ;
	assign \v6_pad  = _w216_ ;
	assign \v7_pad  = _w691_ ;
	assign \v8_pad  = _w694_ ;
	assign \v9_pad  = _w697_ ;
	assign \w10_pad  = _w705_ ;
	assign \w5_pad  = _w717_ ;
	assign \w6_pad  = _w726_ ;
	assign \w7_pad  = _w727_ ;
	assign \w8_pad  = _w731_ ;
	assign \w9_pad  = _w734_ ;
	assign \x10_pad  = _w738_ ;
	assign \x21  = _w741_ ;
	assign \x5_pad  = _w750_ ;
	assign \x6_pad  = _w754_ ;
	assign \x7_pad  = _w755_ ;
	assign \x8_pad  = _w757_ ;
	assign \x9_pad  = _w760_ ;
	assign \y10_pad  = _w764_ ;
	assign \y5_pad  = _w773_ ;
	assign \y6_pad  = _w777_ ;
	assign \y7_pad  = _w779_ ;
	assign \y8_pad  = _w783_ ;
	assign \y9_pad  = _w784_ ;
	assign \z5_pad  = _w793_ ;
	assign \z6_pad  = _w795_ ;
	assign \z7_pad  = _w799_ ;
	assign \z8_pad  = _w801_ ;
	assign \z9_pad  = _w802_ ;
endmodule;