module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G1_pad , \G2_pad , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G288_pad , \G290_pad , \G296_pad , \G302_pad , \G310_pad , \G312_pad , \G315_pad , \G327_pad , \G45_pad , \G47_pad , \G49_pad , \G53_pad , \G55_pad , \_al_n0 , \_al_n1 , \g1452/_0_ , \g1456/_1_ , \g1462/_0_ , \g1463/_0_ , \g1504/_3_ , \g1524/_1_ , \g1524/_2_ , \g1527/_3_ , \g31/_0_ , \g45/_1_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G1_pad  ;
	input \G2_pad  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G288_pad  ;
	output \G290_pad  ;
	output \G296_pad  ;
	output \G302_pad  ;
	output \G310_pad  ;
	output \G312_pad  ;
	output \G315_pad  ;
	output \G327_pad  ;
	output \G45_pad  ;
	output \G47_pad  ;
	output \G49_pad  ;
	output \G53_pad  ;
	output \G55_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1452/_0_  ;
	output \g1456/_1_  ;
	output \g1462/_0_  ;
	output \g1463/_0_  ;
	output \g1504/_3_  ;
	output \g1524/_1_  ;
	output \g1524/_2_  ;
	output \g1527/_3_  ;
	output \g31/_0_  ;
	output \g45/_1_  ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\G40_reg/NET0131 ,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w24_,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w28_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\G39_reg/NET0131 ,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w28_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\G42_reg/NET0131 ,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w25_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\G16_pad ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w35_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\G16_pad ,
		\G4_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\G40_reg/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\G16_pad ,
		\G40_reg/NET0131 ,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\G1_pad ,
		_w24_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w41_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		_w39_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\G38_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\G42_reg/NET0131 ,
		_w47_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w40_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\G38_reg/NET0131 ,
		_w24_,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\G40_reg/NET0131 ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w53_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w38_,
		_w51_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w46_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w26_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\G38_reg/NET0131 ,
		_w36_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\G16_pad ,
		_w61_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w62_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w24_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\G40_reg/NET0131 ,
		_w36_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\G39_reg/NET0131 ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w66_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\G38_reg/NET0131 ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w30_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\G10_pad ,
		\G11_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\G12_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w33_,
		_w40_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\G10_pad ,
		\G11_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\G15_pad ,
		_w39_,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w74_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w75_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\G5_pad ,
		_w27_,
		_w81_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w61_,
		_w65_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w52_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w82_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w50_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\G41_reg/NET0131 ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w39_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\G5_pad ,
		_w27_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\G13_pad ,
		\G15_pad ,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\G42_reg/NET0131 ,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		\G38_reg/NET0131 ,
		_w28_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		\G40_reg/NET0131 ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\G39_reg/NET0131 ,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\G6_pad ,
		\G7_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\G8_pad ,
		\G9_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w97_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\G40_reg/NET0131 ,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\G41_reg/NET0131 ,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w102_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w96_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		\G1_pad ,
		_w29_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\G42_reg/NET0131 ,
		\G6_pad ,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\G7_pad ,
		\G8_pad ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\G9_pad ,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w109_,
		_w110_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w112_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w107_,
		_w108_,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		_w39_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w28_,
		_w108_,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\G39_reg/NET0131 ,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\G39_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\G42_reg/NET0131 ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w119_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\G40_reg/NET0131 ,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w117_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w106_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\G16_pad ,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\G41_reg/NET0131 ,
		\G5_pad ,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\G42_reg/NET0131 ,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\G1_pad ,
		\G3_pad ,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w59_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		\G2_pad ,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w128_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		_w61_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\G40_reg/NET0131 ,
		_w36_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		\G4_pad ,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\G14_pad ,
		\G15_pad ,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w88_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w135_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\G39_reg/NET0131 ,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w133_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\G38_reg/NET0131 ,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w142_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\G0_pad ,
		\G38_reg/NET0131 ,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\G39_reg/NET0131 ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w142_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w67_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w55_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w141_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w126_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\G18_pad ,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		\G40_reg/NET0131 ,
		_w62_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\G38_reg/NET0131 ,
		_w36_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\G42_reg/NET0131 ,
		_w76_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\G15_pad ,
		_w32_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w154_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\G16_pad ,
		_w103_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w153_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w152_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w151_,
		_w156_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w99_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\G16_pad ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		\G4_pad ,
		_w35_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w36_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		_w164_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		\G0_pad ,
		_w36_,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		\G4_pad ,
		_w24_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\G38_reg/NET0131 ,
		_w168_,
		_w170_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w169_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\G38_reg/NET0131 ,
		_w128_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w130_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		_w61_,
		_w171_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w173_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\G2_pad ,
		_w129_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\G16_pad ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\G41_reg/NET0131 ,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		\G14_pad ,
		\G15_pad ,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\G41_reg/NET0131 ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name157 (
		_w87_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w39_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w178_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w161_,
		_w167_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w183_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w175_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		\G18_pad ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w37_,
		_w165_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w74_,
		_w154_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		\G38_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w40_,
		_w48_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		_w109_,
		_w190_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w189_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\G38_reg/NET0131 ,
		_w66_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w177_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w188_,
		_w194_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w196_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w175_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\G18_pad ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\G16_pad ,
		\G1_pad ,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		\G38_reg/NET0131 ,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		\G0_pad ,
		_w190_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\G16_pad ,
		\G38_reg/NET0131 ,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\G42_reg/NET0131 ,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		_w29_,
		_w202_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w203_,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\G10_pad ,
		\G12_pad ,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\G11_pad ,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w75_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w208_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\G39_reg/NET0131 ,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		\G1_pad ,
		\G38_reg/NET0131 ,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		\G41_reg/NET0131 ,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\G42_reg/NET0131 ,
		_w61_,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		\G41_reg/NET0131 ,
		_w143_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		_w217_,
		_w218_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		_w219_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		\G4_pad ,
		_w65_,
		_w222_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w120_,
		_w204_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w222_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w33_,
		_w218_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w221_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w215_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		\G18_pad ,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w61_,
		_w87_,
		_w230_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		\G39_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		\G41_reg/NET0131 ,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		_w216_,
		_w230_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\G15_pad ,
		_w89_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w39_,
		_w137_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\G3_pad ,
		_w66_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		_w202_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\G41_reg/NET0131 ,
		\G5_pad ,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		\G16_pad ,
		\G39_reg/NET0131 ,
		_w240_
	);
	LUT2 #(
		.INIT('h2)
	) name217 (
		\G42_reg/NET0131 ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		\G40_reg/NET0131 ,
		_w142_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		_w239_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w232_,
		_w241_,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w243_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w42_,
		_w83_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w176_,
		_w232_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w246_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		_w59_,
		_w109_,
		_w249_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		\G16_pad ,
		_w87_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w249_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\G39_reg/NET0131 ,
		_w135_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w181_,
		_w251_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w252_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w245_,
		_w248_,
		_w255_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		_w254_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\G38_reg/NET0131 ,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\G16_pad ,
		_w91_,
		_w258_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		_w153_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w144_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		_w67_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\G16_pad ,
		\G41_reg/NET0131 ,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w71_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		_w36_,
		_w165_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		\G39_reg/NET0131 ,
		_w71_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w99_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name244 (
		\G15_pad ,
		_w25_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\G41_reg/NET0131 ,
		_w82_,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w268_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w267_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\G40_reg/NET0131 ,
		_w40_,
		_w272_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w261_,
		_w265_,
		_w274_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w273_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w257_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		\G18_pad ,
		_w276_,
		_w277_
	);
	assign \G288_pad  = _w27_ ;
	assign \G290_pad  = _w31_ ;
	assign \G296_pad  = _w34_ ;
	assign \G302_pad  = _w58_ ;
	assign \G310_pad  = _w60_ ;
	assign \G312_pad  = _w64_ ;
	assign \G315_pad  = _w70_ ;
	assign \G327_pad  = _w72_ ;
	assign \G45_pad  = _w80_ ;
	assign \G47_pad  = _w81_ ;
	assign \G49_pad  = _w86_ ;
	assign \G53_pad  = _w89_ ;
	assign \G55_pad  = _w90_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1452/_0_  = _w150_ ;
	assign \g1456/_1_  = _w187_ ;
	assign \g1462/_0_  = _w200_ ;
	assign \g1463/_0_  = _w229_ ;
	assign \g1504/_3_  = _w234_ ;
	assign \g1524/_1_  = _w235_ ;
	assign \g1524/_2_  = _w236_ ;
	assign \g1527/_3_  = _w238_ ;
	assign \g31/_0_  = _w277_ ;
	assign \g45/_1_  = _w167_ ;
endmodule;