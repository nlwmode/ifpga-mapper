module top( \cont1_reg[0]/NET0131  , \cont1_reg[1]/NET0131  , \cont1_reg[2]/NET0131  , \cont1_reg[3]/NET0131  , \cont1_reg[4]/NET0131  , \cont1_reg[5]/NET0131  , \cont1_reg[6]/NET0131  , \cont1_reg[7]/NET0131  , \cont1_reg[8]/NET0131  , \cont_reg[0]/NET0131  , \cont_reg[1]/NET0131  , \cont_reg[2]/NET0131  , \cont_reg[3]/NET0131  , \cont_reg[4]/NET0131  , \r_in_reg[0]/NET0131  , \r_in_reg[1]/NET0131  , \r_in_reg[2]/NET0131  , \r_in_reg[3]/NET0131  , \r_in_reg[4]/NET0131  , \r_in_reg[5]/NET0131  , \stato_reg[0]/NET0131  , \stato_reg[1]/NET0131  , \stato_reg[2]/NET0131  , \stato_reg[3]/NET0131  , stbi_pad , \x_in[0]_pad  , \x_in[1]_pad  , \x_in[2]_pad  , \x_in[3]_pad  , \x_in[4]_pad  , \x_in[5]_pad  , \x_out[0]_pad  , \x_out[1]_pad  , \x_out[2]_pad  , \x_out[3]_pad  , \x_out[4]_pad  , \x_out[5]_pad  , \_al_n0  , \_al_n1  , \g2420/_0_  , \g2432/_0_  , \g2433/_0_  , \g2442/_0_  , \g2449/_0_  , \g2469/_0_  , \g2489/_0_  , \g2492/_0_  , \g2531/_0_  , \g2532/_0_  , \g2533/_0_  , \g2534/_0_  , \g2536/_0_  , \g2542/_0_  , \g2619/_0_  , \g2620/_0_  , \g2662/_0_  , \g2663/_0_  , \g2665/_0_  , \g2666/_0_  , \g2667/_0_  , \g2668/_0_  , \g2712/_0_  , \g3382/_0_  , \g34/_0_  , \g3435/_0_  , \g3443/_0_  , \g3735/_0_  , \g4020/_0_  , \g64/_0_  );
  input \cont1_reg[0]/NET0131  ;
  input \cont1_reg[1]/NET0131  ;
  input \cont1_reg[2]/NET0131  ;
  input \cont1_reg[3]/NET0131  ;
  input \cont1_reg[4]/NET0131  ;
  input \cont1_reg[5]/NET0131  ;
  input \cont1_reg[6]/NET0131  ;
  input \cont1_reg[7]/NET0131  ;
  input \cont1_reg[8]/NET0131  ;
  input \cont_reg[0]/NET0131  ;
  input \cont_reg[1]/NET0131  ;
  input \cont_reg[2]/NET0131  ;
  input \cont_reg[3]/NET0131  ;
  input \cont_reg[4]/NET0131  ;
  input \r_in_reg[0]/NET0131  ;
  input \r_in_reg[1]/NET0131  ;
  input \r_in_reg[2]/NET0131  ;
  input \r_in_reg[3]/NET0131  ;
  input \r_in_reg[4]/NET0131  ;
  input \r_in_reg[5]/NET0131  ;
  input \stato_reg[0]/NET0131  ;
  input \stato_reg[1]/NET0131  ;
  input \stato_reg[2]/NET0131  ;
  input \stato_reg[3]/NET0131  ;
  input stbi_pad ;
  input \x_in[0]_pad  ;
  input \x_in[1]_pad  ;
  input \x_in[2]_pad  ;
  input \x_in[3]_pad  ;
  input \x_in[4]_pad  ;
  input \x_in[5]_pad  ;
  input \x_out[0]_pad  ;
  input \x_out[1]_pad  ;
  input \x_out[2]_pad  ;
  input \x_out[3]_pad  ;
  input \x_out[4]_pad  ;
  input \x_out[5]_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g2420/_0_  ;
  output \g2432/_0_  ;
  output \g2433/_0_  ;
  output \g2442/_0_  ;
  output \g2449/_0_  ;
  output \g2469/_0_  ;
  output \g2489/_0_  ;
  output \g2492/_0_  ;
  output \g2531/_0_  ;
  output \g2532/_0_  ;
  output \g2533/_0_  ;
  output \g2534/_0_  ;
  output \g2536/_0_  ;
  output \g2542/_0_  ;
  output \g2619/_0_  ;
  output \g2620/_0_  ;
  output \g2662/_0_  ;
  output \g2663/_0_  ;
  output \g2665/_0_  ;
  output \g2666/_0_  ;
  output \g2667/_0_  ;
  output \g2668/_0_  ;
  output \g2712/_0_  ;
  output \g3382/_0_  ;
  output \g34/_0_  ;
  output \g3435/_0_  ;
  output \g3443/_0_  ;
  output \g3735/_0_  ;
  output \g4020/_0_  ;
  output \g64/_0_  ;
  wire n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 ;
  assign n38 = \cont1_reg[2]/NET0131  & \r_in_reg[2]/NET0131  ;
  assign n39 = ~\cont1_reg[1]/NET0131  & ~\r_in_reg[1]/NET0131  ;
  assign n40 = \cont1_reg[1]/NET0131  & \r_in_reg[1]/NET0131  ;
  assign n41 = \cont1_reg[0]/NET0131  & \r_in_reg[0]/NET0131  ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = ~n39 & ~n42 ;
  assign n44 = ~n38 & ~n43 ;
  assign n45 = ~\cont1_reg[4]/NET0131  & ~\r_in_reg[4]/NET0131  ;
  assign n46 = ~\cont1_reg[2]/NET0131  & ~\r_in_reg[2]/NET0131  ;
  assign n47 = ~\cont1_reg[3]/NET0131  & ~\r_in_reg[3]/NET0131  ;
  assign n48 = ~n46 & ~n47 ;
  assign n49 = ~n45 & n48 ;
  assign n50 = ~n44 & n49 ;
  assign n51 = \cont1_reg[5]/NET0131  & \r_in_reg[5]/NET0131  ;
  assign n52 = \cont1_reg[4]/NET0131  & \r_in_reg[4]/NET0131  ;
  assign n53 = \cont1_reg[3]/NET0131  & \r_in_reg[3]/NET0131  ;
  assign n54 = ~n45 & n53 ;
  assign n55 = ~n52 & ~n54 ;
  assign n56 = ~n51 & n55 ;
  assign n57 = ~n50 & n56 ;
  assign n58 = ~\cont1_reg[5]/NET0131  & ~\r_in_reg[5]/NET0131  ;
  assign n59 = \cont1_reg[6]/NET0131  & \r_in_reg[1]/NET0131  ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~n57 & n60 ;
  assign n62 = ~\cont1_reg[2]/NET0131  & \r_in_reg[2]/NET0131  ;
  assign n63 = \cont1_reg[2]/NET0131  & ~\r_in_reg[2]/NET0131  ;
  assign n64 = ~n62 & n63 ;
  assign n65 = \cont1_reg[1]/NET0131  & ~\r_in_reg[1]/NET0131  ;
  assign n66 = \cont1_reg[0]/NET0131  & ~\r_in_reg[0]/NET0131  ;
  assign n67 = ~n65 & ~n66 ;
  assign n68 = ~\cont1_reg[1]/NET0131  & \r_in_reg[1]/NET0131  ;
  assign n69 = ~n62 & ~n68 ;
  assign n70 = ~n67 & n69 ;
  assign n71 = ~n64 & ~n70 ;
  assign n72 = \cont1_reg[5]/NET0131  & ~\r_in_reg[5]/NET0131  ;
  assign n73 = ~\cont1_reg[6]/NET0131  & ~n72 ;
  assign n74 = \cont1_reg[4]/NET0131  & ~\r_in_reg[4]/NET0131  ;
  assign n75 = \cont1_reg[3]/NET0131  & ~\r_in_reg[3]/NET0131  ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = n73 & n76 ;
  assign n78 = n71 & n77 ;
  assign n79 = ~\r_in_reg[1]/NET0131  & ~n73 ;
  assign n80 = ~\cont1_reg[4]/NET0131  & \r_in_reg[4]/NET0131  ;
  assign n81 = ~\cont1_reg[3]/NET0131  & \r_in_reg[3]/NET0131  ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = ~n74 & ~n82 ;
  assign n84 = ~\cont1_reg[5]/NET0131  & \r_in_reg[5]/NET0131  ;
  assign n85 = ~\r_in_reg[1]/NET0131  & ~n84 ;
  assign n86 = ~n83 & n85 ;
  assign n87 = ~n79 & ~n86 ;
  assign n88 = ~n78 & ~n87 ;
  assign n89 = ~\cont1_reg[7]/NET0131  & ~n88 ;
  assign n90 = ~n61 & n89 ;
  assign n91 = ~\stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n92 = ~\stato_reg[0]/NET0131  & ~\stato_reg[3]/NET0131  ;
  assign n93 = n91 & n92 ;
  assign n94 = \cont1_reg[7]/NET0131  & n88 ;
  assign n95 = \cont1_reg[7]/NET0131  & n60 ;
  assign n96 = ~n57 & n95 ;
  assign n97 = ~n94 & ~n96 ;
  assign n98 = n93 & n97 ;
  assign n99 = ~n90 & n98 ;
  assign n100 = ~\cont1_reg[0]/NET0131  & ~\cont1_reg[1]/NET0131  ;
  assign n101 = ~\cont1_reg[2]/NET0131  & n100 ;
  assign n102 = \cont1_reg[3]/NET0131  & \cont1_reg[4]/NET0131  ;
  assign n103 = \cont1_reg[5]/NET0131  & \cont1_reg[6]/NET0131  ;
  assign n104 = n102 & n103 ;
  assign n105 = ~n101 & n104 ;
  assign n106 = ~\cont1_reg[7]/NET0131  & ~n105 ;
  assign n107 = ~\r_in_reg[2]/NET0131  & \r_in_reg[3]/NET0131  ;
  assign n108 = ~n101 & n102 ;
  assign n109 = \cont1_reg[6]/NET0131  & \cont1_reg[7]/NET0131  ;
  assign n110 = \cont1_reg[5]/NET0131  & n109 ;
  assign n111 = n108 & n110 ;
  assign n112 = n107 & ~n111 ;
  assign n113 = ~n106 & n112 ;
  assign n114 = ~\cont1_reg[2]/NET0131  & ~\cont1_reg[3]/NET0131  ;
  assign n115 = ~\cont1_reg[4]/NET0131  & n114 ;
  assign n116 = n103 & ~n115 ;
  assign n117 = ~\cont1_reg[7]/NET0131  & ~n116 ;
  assign n118 = \r_in_reg[2]/NET0131  & \r_in_reg[3]/NET0131  ;
  assign n119 = n110 & ~n115 ;
  assign n120 = n118 & ~n119 ;
  assign n121 = ~n117 & n120 ;
  assign n122 = \cont1_reg[2]/NET0131  & \cont1_reg[4]/NET0131  ;
  assign n123 = ~n100 & n122 ;
  assign n124 = ~n102 & ~n123 ;
  assign n125 = ~\r_in_reg[2]/NET0131  & ~\r_in_reg[3]/NET0131  ;
  assign n126 = ~\cont1_reg[6]/NET0131  & ~\cont1_reg[7]/NET0131  ;
  assign n127 = ~\cont1_reg[5]/NET0131  & n126 ;
  assign n128 = n125 & n127 ;
  assign n129 = n124 & n128 ;
  assign n130 = ~n121 & ~n129 ;
  assign n131 = ~n113 & n130 ;
  assign n132 = \cont1_reg[4]/NET0131  & \cont1_reg[5]/NET0131  ;
  assign n133 = ~\cont1_reg[1]/NET0131  & ~\cont1_reg[2]/NET0131  ;
  assign n134 = \cont1_reg[3]/NET0131  & \cont1_reg[5]/NET0131  ;
  assign n135 = ~n133 & n134 ;
  assign n136 = ~n132 & ~n135 ;
  assign n137 = ~\cont1_reg[6]/NET0131  & n136 ;
  assign n138 = \r_in_reg[2]/NET0131  & ~\r_in_reg[3]/NET0131  ;
  assign n139 = \cont1_reg[7]/NET0131  & n138 ;
  assign n140 = ~n137 & n139 ;
  assign n141 = ~\cont1_reg[7]/NET0131  & n138 ;
  assign n142 = n137 & n141 ;
  assign n143 = ~n140 & ~n142 ;
  assign n144 = ~\cont1_reg[5]/NET0131  & ~\cont1_reg[6]/NET0131  ;
  assign n145 = n124 & n144 ;
  assign n146 = \cont1_reg[7]/NET0131  & n125 ;
  assign n147 = ~n145 & n146 ;
  assign n148 = n143 & ~n147 ;
  assign n149 = n131 & n148 ;
  assign n150 = \stato_reg[0]/NET0131  & ~\stato_reg[3]/NET0131  ;
  assign n151 = \stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n152 = n150 & n151 ;
  assign n153 = ~n149 & n152 ;
  assign n154 = n91 & n150 ;
  assign n155 = ~\cont1_reg[8]/NET0131  & ~n127 ;
  assign n156 = n102 & ~n133 ;
  assign n157 = ~\cont1_reg[0]/NET0131  & ~\cont1_reg[2]/NET0131  ;
  assign n158 = ~\cont1_reg[8]/NET0131  & ~n157 ;
  assign n159 = n156 & n158 ;
  assign n160 = ~n155 & ~n159 ;
  assign n161 = ~\cont1_reg[5]/NET0131  & ~n156 ;
  assign n162 = ~\cont1_reg[6]/NET0131  & n161 ;
  assign n163 = ~n160 & n162 ;
  assign n164 = n154 & ~n163 ;
  assign n165 = \stato_reg[1]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n166 = n92 & n165 ;
  assign n167 = ~\r_in_reg[0]/NET0131  & ~\r_in_reg[1]/NET0131  ;
  assign n168 = ~\r_in_reg[4]/NET0131  & ~\r_in_reg[5]/NET0131  ;
  assign n169 = n167 & n168 ;
  assign n170 = n125 & n169 ;
  assign n171 = \r_in_reg[0]/NET0131  & \r_in_reg[1]/NET0131  ;
  assign n172 = \r_in_reg[4]/NET0131  & \r_in_reg[5]/NET0131  ;
  assign n173 = n118 & n172 ;
  assign n174 = n171 & n173 ;
  assign n175 = ~n170 & ~n174 ;
  assign n176 = n166 & n175 ;
  assign n177 = ~\stato_reg[1]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n178 = \stato_reg[0]/NET0131  & \stato_reg[3]/NET0131  ;
  assign n179 = n177 & ~n178 ;
  assign n180 = \cont1_reg[7]/NET0131  & ~n179 ;
  assign n181 = ~n176 & n180 ;
  assign n182 = ~n164 & n181 ;
  assign n183 = ~\cont1_reg[6]/NET0131  & n154 ;
  assign n184 = n161 & n183 ;
  assign n185 = ~n160 & n184 ;
  assign n186 = ~\cont1_reg[7]/NET0131  & ~n185 ;
  assign n187 = ~n182 & ~n186 ;
  assign n188 = ~\cont1_reg[3]/NET0131  & ~\cont1_reg[4]/NET0131  ;
  assign n189 = \cont1_reg[1]/NET0131  & \cont1_reg[2]/NET0131  ;
  assign n190 = n188 & ~n189 ;
  assign n191 = \cont1_reg[5]/NET0131  & ~\cont1_reg[8]/NET0131  ;
  assign n192 = ~n126 & n191 ;
  assign n193 = ~n190 & n192 ;
  assign n194 = \cont1_reg[6]/NET0131  & n193 ;
  assign n195 = ~\cont1_reg[7]/NET0131  & ~n194 ;
  assign n196 = ~\cont1_reg[8]/NET0131  & ~n126 ;
  assign n197 = ~n190 & n196 ;
  assign n198 = n110 & n197 ;
  assign n199 = n92 & n151 ;
  assign n200 = ~n198 & n199 ;
  assign n201 = ~n195 & n200 ;
  assign n202 = ~n187 & ~n201 ;
  assign n203 = ~n153 & n202 ;
  assign n204 = ~n99 & n203 ;
  assign n205 = n154 & n160 ;
  assign n206 = ~n196 & n199 ;
  assign n207 = ~n179 & ~n206 ;
  assign n208 = ~\cont1_reg[0]/NET0131  & \r_in_reg[1]/NET0131  ;
  assign n209 = ~n66 & ~n208 ;
  assign n210 = n93 & n209 ;
  assign n211 = \cont1_reg[1]/NET0131  & ~n210 ;
  assign n212 = n207 & n211 ;
  assign n213 = ~n205 & n212 ;
  assign n214 = n154 & ~n160 ;
  assign n215 = n93 & ~n209 ;
  assign n216 = n196 & n199 ;
  assign n217 = ~\cont1_reg[1]/NET0131  & ~n216 ;
  assign n218 = ~n215 & n217 ;
  assign n219 = ~n214 & n218 ;
  assign n220 = ~n213 & ~n219 ;
  assign n221 = n166 & n174 ;
  assign n222 = \cont1_reg[1]/NET0131  & n166 ;
  assign n223 = ~n170 & n222 ;
  assign n224 = ~n221 & ~n223 ;
  assign n225 = n150 & n165 ;
  assign n226 = ~\cont_reg[1]/NET0131  & ~\r_in_reg[0]/NET0131  ;
  assign n227 = ~\cont_reg[0]/NET0131  & \r_in_reg[0]/NET0131  ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = n225 & n228 ;
  assign n230 = ~\cont1_reg[0]/NET0131  & ~\r_in_reg[2]/NET0131  ;
  assign n231 = ~n138 & ~n230 ;
  assign n232 = ~\cont1_reg[1]/NET0131  & n231 ;
  assign n233 = \cont1_reg[1]/NET0131  & ~n231 ;
  assign n234 = n152 & ~n233 ;
  assign n235 = ~n232 & n234 ;
  assign n236 = ~n229 & ~n235 ;
  assign n237 = n224 & n236 ;
  assign n238 = ~n220 & n237 ;
  assign n239 = \cont1_reg[2]/NET0131  & \r_in_reg[3]/NET0131  ;
  assign n240 = ~\r_in_reg[2]/NET0131  & ~n100 ;
  assign n241 = n239 & n240 ;
  assign n242 = \r_in_reg[3]/NET0131  & n62 ;
  assign n243 = ~\cont1_reg[2]/NET0131  & \r_in_reg[3]/NET0131  ;
  assign n244 = n100 & n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = ~n241 & n245 ;
  assign n247 = n152 & ~n246 ;
  assign n248 = ~n133 & ~n189 ;
  assign n249 = \r_in_reg[2]/NET0131  & n248 ;
  assign n250 = ~\r_in_reg[3]/NET0131  & ~n249 ;
  assign n251 = n63 & ~n100 ;
  assign n252 = n46 & n100 ;
  assign n253 = ~n251 & ~n252 ;
  assign n254 = n152 & n253 ;
  assign n255 = n250 & n254 ;
  assign n256 = ~n247 & ~n255 ;
  assign n257 = ~n160 & ~n248 ;
  assign n258 = n127 & ~n156 ;
  assign n259 = ~\cont1_reg[8]/NET0131  & ~n258 ;
  assign n260 = \cont1_reg[2]/NET0131  & ~n259 ;
  assign n261 = ~n257 & ~n260 ;
  assign n262 = n154 & ~n261 ;
  assign n263 = n166 & ~n170 ;
  assign n264 = ~\cont1_reg[2]/NET0131  & ~n174 ;
  assign n265 = n263 & ~n264 ;
  assign n266 = ~\cont_reg[2]/NET0131  & ~\r_in_reg[0]/NET0131  ;
  assign n267 = ~\cont_reg[1]/NET0131  & \r_in_reg[0]/NET0131  ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = n225 & n268 ;
  assign n270 = n216 & n248 ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = ~n265 & n271 ;
  assign n273 = ~n41 & n68 ;
  assign n274 = n39 & ~n66 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = ~n38 & ~n46 ;
  assign n277 = n93 & ~n276 ;
  assign n278 = n275 & n277 ;
  assign n279 = n93 & n276 ;
  assign n280 = ~n275 & n279 ;
  assign n281 = ~n278 & ~n280 ;
  assign n282 = \cont1_reg[2]/NET0131  & ~n207 ;
  assign n283 = n281 & ~n282 ;
  assign n284 = n272 & n283 ;
  assign n285 = ~n262 & n284 ;
  assign n286 = n256 & n285 ;
  assign n287 = \r_in_reg[3]/NET0131  & \r_in_reg[4]/NET0131  ;
  assign n288 = ~\r_in_reg[5]/NET0131  & ~n287 ;
  assign n289 = ~\r_in_reg[2]/NET0131  & ~\r_in_reg[5]/NET0131  ;
  assign n290 = ~n171 & n289 ;
  assign n291 = ~n288 & ~n290 ;
  assign n292 = n166 & ~n291 ;
  assign n293 = n175 & n292 ;
  assign n294 = \stato_reg[2]/NET0131  & n92 ;
  assign n295 = \r_in_reg[1]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n296 = n294 & ~n295 ;
  assign n297 = n150 & n177 ;
  assign n298 = ~stbi_pad & n297 ;
  assign n299 = ~n296 & ~n298 ;
  assign n300 = ~n205 & n299 ;
  assign n301 = ~n293 & n300 ;
  assign n302 = ~\stato_reg[0]/NET0131  & n177 ;
  assign n303 = ~n154 & ~n302 ;
  assign n304 = ~n206 & n303 ;
  assign n305 = \r_in_reg[1]/NET0131  & n93 ;
  assign n306 = stbi_pad & n297 ;
  assign n307 = ~n305 & ~n306 ;
  assign n308 = n304 & n307 ;
  assign n309 = ~n176 & n308 ;
  assign n310 = ~\stato_reg[3]/NET0131  & \x_out[3]_pad  ;
  assign n311 = ~n302 & n310 ;
  assign n312 = n100 & n114 ;
  assign n313 = \cont1_reg[8]/NET0131  & n312 ;
  assign n314 = \cont1_reg[3]/NET0131  & \cont1_reg[8]/NET0131  ;
  assign n315 = ~n101 & n314 ;
  assign n316 = ~n313 & ~n315 ;
  assign n317 = ~\stato_reg[0]/NET0131  & \stato_reg[3]/NET0131  ;
  assign n318 = n177 & n317 ;
  assign n319 = ~\cont1_reg[3]/NET0131  & ~\cont1_reg[8]/NET0131  ;
  assign n320 = n318 & ~n319 ;
  assign n321 = n316 & n320 ;
  assign n322 = ~n311 & ~n321 ;
  assign n323 = ~\stato_reg[3]/NET0131  & \x_out[4]_pad  ;
  assign n324 = ~n302 & n323 ;
  assign n325 = \cont1_reg[8]/NET0131  & ~n312 ;
  assign n326 = ~\cont1_reg[4]/NET0131  & ~n325 ;
  assign n327 = \cont1_reg[4]/NET0131  & \cont1_reg[8]/NET0131  ;
  assign n328 = ~n312 & n327 ;
  assign n329 = n318 & ~n328 ;
  assign n330 = ~n326 & n329 ;
  assign n331 = ~n324 & ~n330 ;
  assign n332 = ~\stato_reg[3]/NET0131  & \x_out[5]_pad  ;
  assign n333 = ~n302 & n332 ;
  assign n334 = ~\cont1_reg[5]/NET0131  & ~\cont1_reg[8]/NET0131  ;
  assign n335 = ~\cont1_reg[5]/NET0131  & n188 ;
  assign n336 = n101 & n335 ;
  assign n337 = ~n334 & ~n336 ;
  assign n338 = n101 & n188 ;
  assign n339 = \cont1_reg[5]/NET0131  & \cont1_reg[8]/NET0131  ;
  assign n340 = ~n338 & n339 ;
  assign n341 = n318 & ~n340 ;
  assign n342 = n337 & n341 ;
  assign n343 = ~n333 & ~n342 ;
  assign n344 = \stato_reg[2]/NET0131  & ~\stato_reg[3]/NET0131  ;
  assign n345 = ~n150 & ~n344 ;
  assign n346 = ~n318 & n345 ;
  assign n347 = \cont_reg[1]/NET0131  & ~n346 ;
  assign n348 = \cont_reg[1]/NET0131  & n166 ;
  assign n349 = n175 & n348 ;
  assign n350 = ~n347 & ~n349 ;
  assign n351 = ~\cont_reg[0]/NET0131  & ~\cont_reg[1]/NET0131  ;
  assign n352 = ~\cont_reg[2]/NET0131  & n351 ;
  assign n353 = \cont_reg[3]/NET0131  & \cont_reg[4]/NET0131  ;
  assign n354 = ~n352 & n353 ;
  assign n355 = \cont_reg[0]/NET0131  & \cont_reg[1]/NET0131  ;
  assign n356 = ~n351 & ~n355 ;
  assign n357 = n166 & n356 ;
  assign n358 = ~n354 & n357 ;
  assign n359 = ~n175 & n358 ;
  assign n360 = n350 & ~n359 ;
  assign n361 = \cont_reg[2]/NET0131  & ~n346 ;
  assign n362 = \cont_reg[2]/NET0131  & n166 ;
  assign n363 = n175 & n362 ;
  assign n364 = ~n361 & ~n363 ;
  assign n365 = n166 & ~n354 ;
  assign n366 = ~n175 & n365 ;
  assign n367 = ~\cont_reg[2]/NET0131  & ~n355 ;
  assign n368 = \cont_reg[2]/NET0131  & n355 ;
  assign n369 = ~n367 & ~n368 ;
  assign n370 = n366 & n369 ;
  assign n371 = n364 & ~n370 ;
  assign n372 = ~n176 & n346 ;
  assign n373 = \cont_reg[2]/NET0131  & \cont_reg[3]/NET0131  ;
  assign n374 = n355 & n373 ;
  assign n375 = n166 & ~n374 ;
  assign n376 = ~n354 & n375 ;
  assign n377 = ~n175 & n376 ;
  assign n378 = n372 & ~n377 ;
  assign n379 = \cont_reg[3]/NET0131  & ~n378 ;
  assign n380 = n368 & n377 ;
  assign n381 = ~n379 & ~n380 ;
  assign n382 = ~\cont_reg[4]/NET0131  & n374 ;
  assign n383 = n166 & n382 ;
  assign n384 = ~n175 & n383 ;
  assign n385 = ~\cont_reg[4]/NET0131  & ~n384 ;
  assign n386 = ~n377 & ~n384 ;
  assign n387 = n372 & n386 ;
  assign n388 = ~n385 & ~n387 ;
  assign n389 = ~\stato_reg[3]/NET0131  & \x_out[2]_pad  ;
  assign n390 = ~n302 & n389 ;
  assign n391 = \cont1_reg[2]/NET0131  & \cont1_reg[8]/NET0131  ;
  assign n392 = ~n100 & n391 ;
  assign n393 = ~\cont1_reg[2]/NET0131  & \cont1_reg[8]/NET0131  ;
  assign n394 = n100 & n393 ;
  assign n395 = ~n392 & ~n394 ;
  assign n396 = ~\cont1_reg[2]/NET0131  & ~\cont1_reg[8]/NET0131  ;
  assign n397 = n318 & ~n396 ;
  assign n398 = n395 & n397 ;
  assign n399 = ~n390 & ~n398 ;
  assign n400 = \cont_reg[0]/NET0131  & ~n346 ;
  assign n401 = \cont_reg[0]/NET0131  & n166 ;
  assign n402 = n175 & n401 ;
  assign n403 = ~n400 & ~n402 ;
  assign n404 = ~\cont_reg[0]/NET0131  & n166 ;
  assign n405 = ~n354 & n404 ;
  assign n406 = ~n175 & n405 ;
  assign n407 = n403 & ~n406 ;
  assign n408 = \cont1_reg[0]/NET0131  & n318 ;
  assign n409 = ~\stato_reg[3]/NET0131  & \x_out[0]_pad  ;
  assign n410 = ~n302 & n409 ;
  assign n411 = ~n408 & ~n410 ;
  assign n412 = ~\stato_reg[3]/NET0131  & \x_out[1]_pad  ;
  assign n413 = ~n302 & n412 ;
  assign n414 = \cont1_reg[0]/NET0131  & \cont1_reg[8]/NET0131  ;
  assign n415 = \cont1_reg[1]/NET0131  & n414 ;
  assign n416 = ~\cont1_reg[1]/NET0131  & ~n414 ;
  assign n417 = ~n415 & ~n416 ;
  assign n418 = n318 & n417 ;
  assign n419 = ~n413 & ~n418 ;
  assign n420 = ~\stato_reg[3]/NET0131  & \x_in[3]_pad  ;
  assign n421 = n177 & n420 ;
  assign n422 = ~\stato_reg[3]/NET0131  & ~n177 ;
  assign n423 = ~n318 & ~n422 ;
  assign n424 = \r_in_reg[3]/NET0131  & ~n423 ;
  assign n425 = ~n421 & ~n424 ;
  assign n426 = ~\stato_reg[3]/NET0131  & \x_in[5]_pad  ;
  assign n427 = n177 & n426 ;
  assign n428 = \r_in_reg[5]/NET0131  & ~n423 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = ~\stato_reg[3]/NET0131  & \x_in[0]_pad  ;
  assign n431 = n177 & n430 ;
  assign n432 = \r_in_reg[0]/NET0131  & ~n423 ;
  assign n433 = ~n431 & ~n432 ;
  assign n434 = ~\stato_reg[3]/NET0131  & \x_in[1]_pad  ;
  assign n435 = n177 & n434 ;
  assign n436 = \r_in_reg[1]/NET0131  & ~n423 ;
  assign n437 = ~n435 & ~n436 ;
  assign n438 = ~\stato_reg[3]/NET0131  & \x_in[2]_pad  ;
  assign n439 = n177 & n438 ;
  assign n440 = \r_in_reg[2]/NET0131  & ~n423 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~\stato_reg[3]/NET0131  & \x_in[4]_pad  ;
  assign n443 = n177 & n442 ;
  assign n444 = \r_in_reg[4]/NET0131  & ~n423 ;
  assign n445 = ~n443 & ~n444 ;
  assign n446 = n166 & ~n175 ;
  assign n447 = ~n152 & ~n446 ;
  assign n448 = n38 & ~n46 ;
  assign n449 = ~n39 & ~n46 ;
  assign n450 = ~n42 & n449 ;
  assign n451 = ~n448 & ~n450 ;
  assign n452 = ~n47 & ~n53 ;
  assign n453 = \r_in_reg[1]/NET0131  & ~n452 ;
  assign n454 = n451 & n453 ;
  assign n455 = ~\r_in_reg[1]/NET0131  & ~n452 ;
  assign n456 = n71 & n455 ;
  assign n457 = ~n454 & ~n456 ;
  assign n458 = \r_in_reg[1]/NET0131  & n452 ;
  assign n459 = ~n451 & n458 ;
  assign n460 = ~\r_in_reg[1]/NET0131  & n452 ;
  assign n461 = ~n71 & n460 ;
  assign n462 = ~n459 & ~n461 ;
  assign n463 = n93 & n462 ;
  assign n464 = n457 & n463 ;
  assign n465 = \cont1_reg[3]/NET0131  & n179 ;
  assign n466 = \cont1_reg[3]/NET0131  & n166 ;
  assign n467 = n175 & n466 ;
  assign n468 = ~n465 & ~n467 ;
  assign n469 = ~n189 & n196 ;
  assign n470 = \cont1_reg[3]/NET0131  & n199 ;
  assign n471 = ~n469 & n470 ;
  assign n472 = ~\cont1_reg[3]/NET0131  & n199 ;
  assign n473 = n469 & n472 ;
  assign n474 = ~n471 & ~n473 ;
  assign n475 = \r_in_reg[3]/NET0131  & n166 ;
  assign n476 = ~n175 & n475 ;
  assign n477 = ~\cont_reg[3]/NET0131  & ~\r_in_reg[0]/NET0131  ;
  assign n478 = ~\cont_reg[2]/NET0131  & \r_in_reg[0]/NET0131  ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = n225 & n479 ;
  assign n481 = ~n476 & ~n480 ;
  assign n482 = n474 & n481 ;
  assign n483 = n468 & n482 ;
  assign n484 = \cont1_reg[3]/NET0131  & ~n133 ;
  assign n485 = ~\cont1_reg[3]/NET0131  & n133 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = n138 & n486 ;
  assign n488 = \cont1_reg[2]/NET0131  & \cont1_reg[3]/NET0131  ;
  assign n489 = ~n114 & ~n488 ;
  assign n490 = n118 & ~n489 ;
  assign n491 = ~n487 & ~n490 ;
  assign n492 = \cont1_reg[3]/NET0131  & ~n101 ;
  assign n493 = n107 & ~n312 ;
  assign n494 = ~n492 & n493 ;
  assign n495 = ~n100 & n488 ;
  assign n496 = n125 & n495 ;
  assign n497 = \cont1_reg[2]/NET0131  & ~n100 ;
  assign n498 = ~\cont1_reg[3]/NET0131  & n125 ;
  assign n499 = ~n497 & n498 ;
  assign n500 = ~n496 & ~n499 ;
  assign n501 = ~n494 & n500 ;
  assign n502 = n491 & n501 ;
  assign n503 = n152 & ~n502 ;
  assign n504 = ~n160 & ~n486 ;
  assign n505 = ~\cont1_reg[3]/NET0131  & n160 ;
  assign n506 = n154 & ~n505 ;
  assign n507 = ~n504 & n506 ;
  assign n508 = ~n503 & ~n507 ;
  assign n509 = n483 & n508 ;
  assign n510 = ~n464 & n509 ;
  assign n511 = \r_in_reg[1]/NET0131  & ~n109 ;
  assign n512 = ~n45 & ~n58 ;
  assign n513 = ~n38 & ~n53 ;
  assign n514 = ~n47 & ~n513 ;
  assign n515 = n512 & n514 ;
  assign n516 = n52 & ~n58 ;
  assign n517 = ~n51 & ~n516 ;
  assign n518 = ~n515 & n517 ;
  assign n519 = n48 & n512 ;
  assign n520 = n43 & n519 ;
  assign n521 = \r_in_reg[1]/NET0131  & ~n520 ;
  assign n522 = n518 & n521 ;
  assign n523 = ~n511 & ~n522 ;
  assign n524 = ~n72 & ~n74 ;
  assign n525 = n126 & n524 ;
  assign n526 = ~n80 & ~n84 ;
  assign n527 = ~n72 & n126 ;
  assign n528 = ~n526 & n527 ;
  assign n529 = ~n525 & ~n528 ;
  assign n530 = ~n67 & ~n68 ;
  assign n531 = ~n63 & ~n75 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = n62 & ~n75 ;
  assign n534 = ~n81 & ~n533 ;
  assign n535 = ~n528 & n534 ;
  assign n536 = ~n532 & n535 ;
  assign n537 = ~n529 & ~n536 ;
  assign n538 = ~\r_in_reg[1]/NET0131  & n537 ;
  assign n539 = n523 & ~n538 ;
  assign n540 = \cont1_reg[8]/NET0131  & n93 ;
  assign n541 = ~n539 & n540 ;
  assign n542 = ~\cont1_reg[8]/NET0131  & n93 ;
  assign n543 = n539 & n542 ;
  assign n544 = ~n541 & ~n543 ;
  assign n545 = \cont1_reg[8]/NET0131  & n120 ;
  assign n546 = \cont1_reg[8]/NET0131  & n107 ;
  assign n547 = ~n111 & n546 ;
  assign n548 = ~n545 & ~n547 ;
  assign n549 = n107 & n110 ;
  assign n550 = n108 & n549 ;
  assign n551 = n118 & n119 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = ~\cont1_reg[8]/NET0131  & ~n552 ;
  assign n554 = n548 & ~n553 ;
  assign n555 = n126 & n136 ;
  assign n556 = ~\cont1_reg[8]/NET0131  & ~n555 ;
  assign n557 = ~\cont1_reg[6]/NET0131  & \cont1_reg[8]/NET0131  ;
  assign n558 = ~\cont1_reg[7]/NET0131  & n557 ;
  assign n559 = n136 & n558 ;
  assign n560 = n138 & ~n559 ;
  assign n561 = ~n556 & n560 ;
  assign n562 = \cont1_reg[8]/NET0131  & n127 ;
  assign n563 = n124 & n562 ;
  assign n564 = \cont1_reg[8]/NET0131  & n125 ;
  assign n565 = ~n129 & ~n564 ;
  assign n566 = ~n563 & ~n565 ;
  assign n567 = ~n561 & ~n566 ;
  assign n568 = n554 & n567 ;
  assign n569 = n152 & ~n568 ;
  assign n570 = ~n154 & ~n179 ;
  assign n571 = ~n176 & n570 ;
  assign n572 = \cont1_reg[8]/NET0131  & ~n571 ;
  assign n573 = n110 & ~n190 ;
  assign n574 = ~\cont1_reg[8]/NET0131  & ~n573 ;
  assign n575 = n199 & ~n574 ;
  assign n576 = ~n572 & ~n575 ;
  assign n577 = ~n569 & n576 ;
  assign n578 = n544 & n577 ;
  assign n579 = \r_in_reg[1]/NET0131  & n55 ;
  assign n580 = ~n50 & n579 ;
  assign n581 = ~\r_in_reg[1]/NET0131  & n83 ;
  assign n582 = ~\r_in_reg[1]/NET0131  & n76 ;
  assign n583 = n71 & n582 ;
  assign n584 = ~n581 & ~n583 ;
  assign n585 = ~n580 & n584 ;
  assign n586 = ~n72 & ~n84 ;
  assign n587 = n93 & ~n586 ;
  assign n588 = ~n585 & n587 ;
  assign n589 = n93 & n586 ;
  assign n590 = n585 & n589 ;
  assign n591 = ~n588 & ~n590 ;
  assign n592 = ~\cont1_reg[5]/NET0131  & ~n102 ;
  assign n593 = ~\cont1_reg[2]/NET0131  & ~\cont1_reg[5]/NET0131  ;
  assign n594 = n100 & n593 ;
  assign n595 = ~n592 & ~n594 ;
  assign n596 = \cont1_reg[5]/NET0131  & n102 ;
  assign n597 = ~n101 & n596 ;
  assign n598 = n107 & ~n597 ;
  assign n599 = n595 & n598 ;
  assign n600 = \cont1_reg[5]/NET0131  & ~n115 ;
  assign n601 = ~\cont1_reg[4]/NET0131  & ~\cont1_reg[5]/NET0131  ;
  assign n602 = n114 & n601 ;
  assign n603 = n118 & ~n602 ;
  assign n604 = ~n600 & n603 ;
  assign n605 = ~n599 & ~n604 ;
  assign n606 = ~\cont1_reg[5]/NET0131  & n125 ;
  assign n607 = n124 & n606 ;
  assign n608 = \cont1_reg[5]/NET0131  & n125 ;
  assign n609 = ~n124 & n608 ;
  assign n610 = ~n607 & ~n609 ;
  assign n611 = ~n484 & n601 ;
  assign n612 = n136 & n138 ;
  assign n613 = ~n611 & n612 ;
  assign n614 = n610 & ~n613 ;
  assign n615 = n605 & n614 ;
  assign n616 = n152 & ~n615 ;
  assign n617 = ~n160 & n161 ;
  assign n618 = n155 & ~n156 ;
  assign n619 = \cont1_reg[5]/NET0131  & ~n618 ;
  assign n620 = ~n617 & ~n619 ;
  assign n621 = n154 & ~n620 ;
  assign n622 = ~\cont1_reg[5]/NET0131  & ~n197 ;
  assign n623 = ~n193 & n199 ;
  assign n624 = ~n622 & n623 ;
  assign n625 = \cont1_reg[5]/NET0131  & n166 ;
  assign n626 = ~n170 & n625 ;
  assign n627 = ~n221 & ~n626 ;
  assign n628 = \cont1_reg[5]/NET0131  & n179 ;
  assign n629 = \cont_reg[4]/NET0131  & \r_in_reg[0]/NET0131  ;
  assign n630 = n225 & n629 ;
  assign n631 = ~n628 & ~n630 ;
  assign n632 = n627 & n631 ;
  assign n633 = ~n624 & n632 ;
  assign n634 = ~n621 & n633 ;
  assign n635 = ~n616 & n634 ;
  assign n636 = n591 & n635 ;
  assign n637 = n518 & ~n520 ;
  assign n638 = \r_in_reg[1]/NET0131  & ~n637 ;
  assign n639 = n524 & ~n534 ;
  assign n640 = n524 & n531 ;
  assign n641 = ~n530 & n640 ;
  assign n642 = ~n639 & ~n641 ;
  assign n643 = ~n72 & ~n526 ;
  assign n644 = ~\r_in_reg[1]/NET0131  & ~n643 ;
  assign n645 = n642 & n644 ;
  assign n646 = ~\cont1_reg[6]/NET0131  & ~n645 ;
  assign n647 = ~n638 & n646 ;
  assign n648 = \cont1_reg[6]/NET0131  & n645 ;
  assign n649 = n59 & ~n637 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = n93 & n650 ;
  assign n652 = ~n647 & n651 ;
  assign n653 = ~\cont1_reg[5]/NET0131  & n124 ;
  assign n654 = \cont1_reg[6]/NET0131  & n125 ;
  assign n655 = ~n653 & n654 ;
  assign n656 = ~\cont1_reg[6]/NET0131  & n125 ;
  assign n657 = n653 & n656 ;
  assign n658 = ~n655 & ~n657 ;
  assign n659 = ~\cont1_reg[6]/NET0131  & ~n597 ;
  assign n660 = ~n105 & n107 ;
  assign n661 = ~n659 & n660 ;
  assign n662 = ~\cont1_reg[6]/NET0131  & n138 ;
  assign n663 = n136 & n662 ;
  assign n664 = \cont1_reg[6]/NET0131  & n138 ;
  assign n665 = ~n136 & n664 ;
  assign n666 = ~n663 & ~n665 ;
  assign n667 = ~\cont1_reg[4]/NET0131  & ~\cont1_reg[6]/NET0131  ;
  assign n668 = n114 & n667 ;
  assign n669 = ~n144 & ~n668 ;
  assign n670 = ~n116 & n118 ;
  assign n671 = n669 & n670 ;
  assign n672 = n666 & ~n671 ;
  assign n673 = ~n661 & n672 ;
  assign n674 = n658 & n673 ;
  assign n675 = n152 & ~n674 ;
  assign n676 = n154 & n161 ;
  assign n677 = ~n160 & n676 ;
  assign n678 = n193 & n199 ;
  assign n679 = ~\cont1_reg[6]/NET0131  & ~n678 ;
  assign n680 = ~n677 & n679 ;
  assign n681 = n154 & ~n617 ;
  assign n682 = \cont1_reg[6]/NET0131  & ~n179 ;
  assign n683 = ~n623 & n682 ;
  assign n684 = ~n176 & n683 ;
  assign n685 = ~n681 & n684 ;
  assign n686 = ~n680 & ~n685 ;
  assign n687 = ~n675 & ~n686 ;
  assign n688 = ~n652 & n687 ;
  assign n689 = \cont1_reg[0]/NET0131  & n166 ;
  assign n690 = ~n170 & n689 ;
  assign n691 = ~n221 & ~n690 ;
  assign n692 = ~\stato_reg[1]/NET0131  & n150 ;
  assign n693 = ~n302 & ~n692 ;
  assign n694 = ~n199 & n693 ;
  assign n695 = \cont1_reg[0]/NET0131  & ~n694 ;
  assign n696 = ~\cont1_reg[0]/NET0131  & ~\r_in_reg[0]/NET0131  ;
  assign n697 = ~n41 & ~n696 ;
  assign n698 = n93 & n697 ;
  assign n699 = \cont1_reg[0]/NET0131  & \r_in_reg[2]/NET0131  ;
  assign n700 = ~n230 & ~n699 ;
  assign n701 = n152 & ~n700 ;
  assign n702 = \cont_reg[0]/NET0131  & ~\r_in_reg[0]/NET0131  ;
  assign n703 = n225 & n702 ;
  assign n704 = ~n701 & ~n703 ;
  assign n705 = ~n698 & n704 ;
  assign n706 = ~n695 & n705 ;
  assign n707 = n691 & n706 ;
  assign n708 = \stato_reg[0]/NET0131  & ~n151 ;
  assign n709 = n422 & n708 ;
  assign n710 = ~n294 & ~n709 ;
  assign n711 = \r_in_reg[1]/NET0131  & n514 ;
  assign n712 = \r_in_reg[1]/NET0131  & n48 ;
  assign n713 = n43 & n712 ;
  assign n714 = ~n711 & ~n713 ;
  assign n715 = ~\r_in_reg[1]/NET0131  & n534 ;
  assign n716 = ~n532 & n715 ;
  assign n717 = n714 & ~n716 ;
  assign n718 = ~n74 & ~n80 ;
  assign n719 = n93 & n718 ;
  assign n720 = ~n717 & n719 ;
  assign n721 = n93 & ~n718 ;
  assign n722 = n717 & n721 ;
  assign n723 = ~n720 & ~n722 ;
  assign n724 = n154 & n484 ;
  assign n725 = ~n160 & n724 ;
  assign n726 = ~\cont1_reg[3]/NET0131  & ~n189 ;
  assign n727 = n196 & n726 ;
  assign n728 = n199 & n727 ;
  assign n729 = ~\cont1_reg[4]/NET0131  & ~n728 ;
  assign n730 = ~n725 & n729 ;
  assign n731 = ~n160 & n484 ;
  assign n732 = n154 & ~n731 ;
  assign n733 = n199 & ~n727 ;
  assign n734 = \cont1_reg[4]/NET0131  & ~n179 ;
  assign n735 = ~n263 & n734 ;
  assign n736 = ~n733 & n735 ;
  assign n737 = ~n732 & n736 ;
  assign n738 = ~n730 & ~n737 ;
  assign n739 = ~\cont_reg[4]/NET0131  & ~\r_in_reg[0]/NET0131  ;
  assign n740 = ~\cont_reg[3]/NET0131  & \r_in_reg[0]/NET0131  ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = n225 & n741 ;
  assign n743 = ~n221 & ~n742 ;
  assign n744 = ~n152 & n743 ;
  assign n745 = n188 & ~n497 ;
  assign n746 = n125 & ~n745 ;
  assign n747 = n124 & n746 ;
  assign n748 = n107 & ~n108 ;
  assign n749 = ~\cont1_reg[2]/NET0131  & ~\cont1_reg[4]/NET0131  ;
  assign n750 = n100 & n749 ;
  assign n751 = ~n188 & ~n750 ;
  assign n752 = n748 & n751 ;
  assign n753 = ~n747 & ~n752 ;
  assign n754 = ~\cont1_reg[4]/NET0131  & n138 ;
  assign n755 = ~n484 & n754 ;
  assign n756 = n138 & n156 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = \cont1_reg[4]/NET0131  & ~n114 ;
  assign n759 = ~n115 & ~n758 ;
  assign n760 = n118 & ~n759 ;
  assign n761 = n757 & ~n760 ;
  assign n762 = n743 & n761 ;
  assign n763 = n753 & n762 ;
  assign n764 = ~n744 & ~n763 ;
  assign n765 = ~n738 & ~n764 ;
  assign n766 = n723 & n765 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g2420/_0_  = ~n204 ;
  assign \g2432/_0_  = ~n238 ;
  assign \g2433/_0_  = ~n286 ;
  assign \g2442/_0_  = ~n301 ;
  assign \g2449/_0_  = ~n309 ;
  assign \g2469/_0_  = ~n322 ;
  assign \g2489/_0_  = ~n331 ;
  assign \g2492/_0_  = ~n343 ;
  assign \g2531/_0_  = ~n360 ;
  assign \g2532/_0_  = ~n371 ;
  assign \g2533/_0_  = ~n381 ;
  assign \g2534/_0_  = n388 ;
  assign \g2536/_0_  = ~n399 ;
  assign \g2542/_0_  = ~n407 ;
  assign \g2619/_0_  = ~n411 ;
  assign \g2620/_0_  = ~n419 ;
  assign \g2662/_0_  = ~n425 ;
  assign \g2663/_0_  = ~n429 ;
  assign \g2665/_0_  = ~n433 ;
  assign \g2666/_0_  = ~n437 ;
  assign \g2667/_0_  = ~n441 ;
  assign \g2668/_0_  = ~n445 ;
  assign \g2712/_0_  = ~n447 ;
  assign \g3382/_0_  = ~n510 ;
  assign \g34/_0_  = ~n578 ;
  assign \g3435/_0_  = ~n636 ;
  assign \g3443/_0_  = ~n688 ;
  assign \g3735/_0_  = ~n707 ;
  assign \g4020/_0_  = ~n710 ;
  assign \g64/_0_  = ~n766 ;
endmodule
