module top( \C_0_pad  , \C_10_pad  , \C_11_pad  , \C_12_pad  , \C_13_pad  , \C_14_pad  , \C_15_pad  , \C_16_pad  , \C_1_pad  , \C_2_pad  , \C_3_pad  , \C_4_pad  , \C_5_pad  , \C_6_pad  , \C_7_pad  , \C_8_pad  , \C_9_pad  , \P_0_pad  , \X_10_reg/NET0131  , \X_11_reg/NET0131  , \X_12_reg/NET0131  , \X_13_reg/NET0131  , \X_14_reg/NET0131  , \X_15_reg/NET0131  , \X_16_reg/P0002  , \X_1_reg/NET0131  , \X_2_reg/NET0131  , \X_3_reg/NET0131  , \X_4_reg/NET0131  , \X_5_reg/NET0131  , \X_6_reg/NET0131  , \X_7_reg/NET0131  , \X_8_reg/NET0131  , \X_9_reg/NET0131  , \X_12_reg/P0001  , \X_13_reg/P0001  , \X_14_reg/P0001  , \X_15_reg/P0001  , \X_16_reg/P0000  , \X_9_reg/P0001  , Z_pad , \_al_n0  , \_al_n1  , \g1160/_3_  , \g1169/_0_  , \g1185/_0_  , \g1212/_2_  , \g1218/_0_  , \g1234/_0_  , \g16/_1_  , \g17/_0_  , \g27/_2_  , \g29/_3_  , \g669/_1__syn_2  , \g714/_0_  , \g721/_0_  , \g734/_0_  , \g743/_0_  , \g763/_0_  );
  input \C_0_pad  ;
  input \C_10_pad  ;
  input \C_11_pad  ;
  input \C_12_pad  ;
  input \C_13_pad  ;
  input \C_14_pad  ;
  input \C_15_pad  ;
  input \C_16_pad  ;
  input \C_1_pad  ;
  input \C_2_pad  ;
  input \C_3_pad  ;
  input \C_4_pad  ;
  input \C_5_pad  ;
  input \C_6_pad  ;
  input \C_7_pad  ;
  input \C_8_pad  ;
  input \C_9_pad  ;
  input \P_0_pad  ;
  input \X_10_reg/NET0131  ;
  input \X_11_reg/NET0131  ;
  input \X_12_reg/NET0131  ;
  input \X_13_reg/NET0131  ;
  input \X_14_reg/NET0131  ;
  input \X_15_reg/NET0131  ;
  input \X_16_reg/P0002  ;
  input \X_1_reg/NET0131  ;
  input \X_2_reg/NET0131  ;
  input \X_3_reg/NET0131  ;
  input \X_4_reg/NET0131  ;
  input \X_5_reg/NET0131  ;
  input \X_6_reg/NET0131  ;
  input \X_7_reg/NET0131  ;
  input \X_8_reg/NET0131  ;
  input \X_9_reg/NET0131  ;
  output \X_12_reg/P0001  ;
  output \X_13_reg/P0001  ;
  output \X_14_reg/P0001  ;
  output \X_15_reg/P0001  ;
  output \X_16_reg/P0000  ;
  output \X_9_reg/P0001  ;
  output Z_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1160/_3_  ;
  output \g1169/_0_  ;
  output \g1185/_0_  ;
  output \g1212/_2_  ;
  output \g1218/_0_  ;
  output \g1234/_0_  ;
  output \g16/_1_  ;
  output \g17/_0_  ;
  output \g27/_2_  ;
  output \g29/_3_  ;
  output \g669/_1__syn_2  ;
  output \g714/_0_  ;
  output \g721/_0_  ;
  output \g734/_0_  ;
  output \g743/_0_  ;
  output \g763/_0_  ;
  wire n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 ;
  assign n35 = \C_13_pad  & \X_13_reg/NET0131  ;
  assign n36 = \C_14_pad  & ~\X_13_reg/NET0131  ;
  assign n37 = \X_14_reg/NET0131  & n36 ;
  assign n38 = ~n35 & ~n37 ;
  assign n39 = \P_0_pad  & ~n38 ;
  assign n40 = \C_15_pad  & \X_15_reg/NET0131  ;
  assign n41 = \C_16_pad  & ~\X_15_reg/NET0131  ;
  assign n42 = \X_16_reg/P0002  & n41 ;
  assign n43 = ~n40 & ~n42 ;
  assign n44 = \P_0_pad  & ~\X_13_reg/NET0131  ;
  assign n45 = ~\X_14_reg/NET0131  & n44 ;
  assign n46 = ~n43 & n45 ;
  assign n47 = ~n39 & ~n46 ;
  assign n48 = ~\X_10_reg/NET0131  & ~\X_11_reg/NET0131  ;
  assign n49 = ~\X_12_reg/NET0131  & ~\X_9_reg/NET0131  ;
  assign n50 = n48 & n49 ;
  assign n51 = ~n47 & n50 ;
  assign n52 = \P_0_pad  & ~\X_9_reg/NET0131  ;
  assign n53 = ~\X_10_reg/NET0131  & n52 ;
  assign n54 = \C_11_pad  & \X_11_reg/NET0131  ;
  assign n55 = n53 & n54 ;
  assign n56 = \C_10_pad  & \X_10_reg/NET0131  ;
  assign n57 = n52 & n56 ;
  assign n58 = ~n55 & ~n57 ;
  assign n59 = ~n51 & n58 ;
  assign n60 = ~\X_1_reg/NET0131  & ~\X_2_reg/NET0131  ;
  assign n61 = ~\X_3_reg/NET0131  & ~\X_4_reg/NET0131  ;
  assign n62 = n60 & n61 ;
  assign n63 = ~\X_6_reg/NET0131  & n62 ;
  assign n64 = ~\X_7_reg/NET0131  & ~\X_8_reg/NET0131  ;
  assign n65 = ~\X_5_reg/NET0131  & n64 ;
  assign n66 = n63 & n65 ;
  assign n67 = ~n59 & n66 ;
  assign n73 = \C_3_pad  & \X_3_reg/NET0131  ;
  assign n74 = \C_4_pad  & ~\X_3_reg/NET0131  ;
  assign n75 = \X_4_reg/NET0131  & n74 ;
  assign n76 = ~n73 & ~n75 ;
  assign n77 = n60 & ~n76 ;
  assign n68 = \C_5_pad  & \X_5_reg/NET0131  ;
  assign n69 = \C_6_pad  & ~\X_5_reg/NET0131  ;
  assign n70 = \X_6_reg/NET0131  & n69 ;
  assign n71 = ~n68 & ~n70 ;
  assign n72 = n62 & ~n71 ;
  assign n79 = \C_2_pad  & ~\X_1_reg/NET0131  ;
  assign n80 = \X_2_reg/NET0131  & n79 ;
  assign n78 = \C_1_pad  & \X_1_reg/NET0131  ;
  assign n81 = ~\C_0_pad  & ~n78 ;
  assign n82 = ~n80 & n81 ;
  assign n83 = ~n72 & n82 ;
  assign n84 = ~n77 & n83 ;
  assign n85 = \P_0_pad  & ~n84 ;
  assign n86 = \C_9_pad  & \P_0_pad  ;
  assign n87 = \X_9_reg/NET0131  & n86 ;
  assign n88 = \C_12_pad  & ~\X_11_reg/NET0131  ;
  assign n89 = \X_12_reg/NET0131  & n88 ;
  assign n90 = n53 & n89 ;
  assign n91 = ~n87 & ~n90 ;
  assign n92 = n66 & ~n91 ;
  assign n93 = \C_7_pad  & \X_7_reg/NET0131  ;
  assign n94 = \C_8_pad  & ~\X_7_reg/NET0131  ;
  assign n95 = \X_8_reg/NET0131  & n94 ;
  assign n96 = ~n93 & ~n95 ;
  assign n97 = \P_0_pad  & ~\X_5_reg/NET0131  ;
  assign n98 = n63 & n97 ;
  assign n99 = ~n96 & n98 ;
  assign n100 = ~n92 & ~n99 ;
  assign n101 = ~n85 & n100 ;
  assign n102 = ~n67 & n101 ;
  assign n103 = \X_7_reg/NET0131  & \X_8_reg/NET0131  ;
  assign n104 = \P_0_pad  & \X_1_reg/NET0131  ;
  assign n105 = \X_2_reg/NET0131  & n104 ;
  assign n106 = \X_3_reg/NET0131  & n105 ;
  assign n107 = \X_4_reg/NET0131  & n106 ;
  assign n108 = \X_5_reg/NET0131  & \X_6_reg/NET0131  ;
  assign n109 = n107 & n108 ;
  assign n110 = n103 & n109 ;
  assign n111 = \X_10_reg/NET0131  & \X_4_reg/NET0131  ;
  assign n112 = \X_9_reg/NET0131  & n111 ;
  assign n113 = n103 & n108 ;
  assign n114 = n112 & n113 ;
  assign n115 = n106 & n114 ;
  assign n116 = \X_11_reg/NET0131  & n115 ;
  assign n117 = ~\X_11_reg/NET0131  & ~n115 ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = \X_7_reg/NET0131  & ~n109 ;
  assign n120 = ~n64 & ~n103 ;
  assign n121 = ~n119 & ~n120 ;
  assign n122 = n119 & n120 ;
  assign n123 = ~n121 & ~n122 ;
  assign n124 = \X_12_reg/NET0131  & n116 ;
  assign n125 = \X_13_reg/NET0131  & n124 ;
  assign n126 = ~\X_2_reg/NET0131  & ~n104 ;
  assign n127 = ~n105 & ~n126 ;
  assign n128 = \X_9_reg/NET0131  & n110 ;
  assign n129 = ~\X_10_reg/NET0131  & ~n128 ;
  assign n130 = ~n115 & ~n129 ;
  assign n131 = \X_14_reg/NET0131  & n125 ;
  assign n132 = \X_5_reg/NET0131  & n107 ;
  assign n133 = ~\X_6_reg/NET0131  & ~n132 ;
  assign n134 = ~n109 & ~n133 ;
  assign n135 = \X_15_reg/NET0131  & n131 ;
  assign n136 = ~\X_4_reg/NET0131  & ~n106 ;
  assign n137 = ~n107 & ~n136 ;
  assign n138 = ~\X_7_reg/NET0131  & n109 ;
  assign n139 = ~n119 & ~n138 ;
  assign n140 = ~\X_5_reg/NET0131  & ~n107 ;
  assign n141 = ~n132 & ~n140 ;
  assign n142 = ~\X_3_reg/NET0131  & ~n105 ;
  assign n143 = ~n106 & ~n142 ;
  assign n144 = ~\P_0_pad  & ~\X_1_reg/NET0131  ;
  assign n145 = ~n104 & ~n144 ;
  assign \X_12_reg/P0001  = ~\X_12_reg/NET0131  ;
  assign \X_13_reg/P0001  = ~\X_13_reg/NET0131  ;
  assign \X_14_reg/P0001  = ~\X_14_reg/NET0131  ;
  assign \X_15_reg/P0001  = ~\X_15_reg/NET0131  ;
  assign \X_16_reg/P0000  = ~\X_16_reg/P0002  ;
  assign \X_9_reg/P0001  = ~\X_9_reg/NET0131  ;
  assign Z_pad = ~n102 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1160/_3_  = n110 ;
  assign \g1169/_0_  = n118 ;
  assign \g1185/_0_  = n123 ;
  assign \g1212/_2_  = n125 ;
  assign \g1218/_0_  = n127 ;
  assign \g1234/_0_  = n130 ;
  assign \g16/_1_  = n131 ;
  assign \g17/_0_  = n134 ;
  assign \g27/_2_  = n124 ;
  assign \g29/_3_  = n116 ;
  assign \g669/_1__syn_2  = n135 ;
  assign \g714/_0_  = n137 ;
  assign \g721/_0_  = ~n139 ;
  assign \g734/_0_  = n141 ;
  assign \g743/_0_  = n143 ;
  assign \g763/_0_  = n145 ;
endmodule
