module top( a_pad , b_pad , c_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , \a0_pad  , \b0_pad  , \c0_pad  , \d0_pad  , \e0_pad  , \f0_pad  , \g0_pad  , \h0_pad  , \i0_pad  , \j0_pad  , \k0_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  , \t0_pad  , z_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  output \a0_pad  ;
  output \b0_pad  ;
  output \c0_pad  ;
  output \d0_pad  ;
  output \e0_pad  ;
  output \f0_pad  ;
  output \g0_pad  ;
  output \h0_pad  ;
  output \i0_pad  ;
  output \j0_pad  ;
  output \k0_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  output \t0_pad  ;
  output z_pad ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 ;
  assign n37 = ~t_pad & ~u_pad ;
  assign n38 = v_pad & ~n37 ;
  assign n39 = f_pad & n38 ;
  assign n27 = ~v_pad & ~y_pad ;
  assign n31 = ~s_pad & ~t_pad ;
  assign n32 = ~n27 & n31 ;
  assign n33 = u_pad & ~v_pad ;
  assign n34 = ~u_pad & v_pad ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = n32 & ~n35 ;
  assign n40 = ~w_pad & ~n36 ;
  assign n41 = ~n39 & n40 ;
  assign n25 = v_pad & ~w_pad ;
  assign n26 = q_pad & ~n25 ;
  assign n28 = s_pad & ~t_pad ;
  assign n29 = n27 & n28 ;
  assign n30 = u_pad & n29 ;
  assign n42 = ~n26 & ~n30 ;
  assign n43 = ~n41 & n42 ;
  assign n46 = y_pad & n31 ;
  assign n47 = u_pad & ~n46 ;
  assign n48 = ~v_pad & ~n47 ;
  assign n44 = g_pad & ~n37 ;
  assign n45 = v_pad & ~n44 ;
  assign n49 = w_pad & ~n29 ;
  assign n50 = ~n45 & ~n49 ;
  assign n51 = ~n48 & n50 ;
  assign n52 = q_pad & n32 ;
  assign n53 = ~u_pad & ~w_pad ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = ~v_pad & ~n54 ;
  assign n56 = ~h_pad & ~n33 ;
  assign n57 = n30 & n56 ;
  assign n58 = q_pad & ~n57 ;
  assign n59 = w_pad & ~n58 ;
  assign n60 = ~n37 & n56 ;
  assign n61 = s_pad & n37 ;
  assign n62 = ~n49 & ~n61 ;
  assign n63 = ~n60 & n62 ;
  assign n64 = ~n59 & ~n63 ;
  assign n65 = ~n55 & ~n64 ;
  assign n68 = t_pad & ~u_pad ;
  assign n69 = s_pad & n68 ;
  assign n70 = ~v_pad & ~n69 ;
  assign n66 = i_pad & ~n37 ;
  assign n67 = v_pad & ~n66 ;
  assign n71 = ~w_pad & ~n67 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = ~s_pad & ~v_pad ;
  assign n74 = ~n28 & ~n73 ;
  assign n75 = ~u_pad & ~n74 ;
  assign n76 = j_pad & n38 ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = ~w_pad & ~n77 ;
  assign n79 = ~a_pad & ~k_pad ;
  assign n80 = l_pad & n79 ;
  assign n82 = ~m_pad & n_pad ;
  assign n81 = k_pad & ~l_pad ;
  assign n83 = ~a_pad & n81 ;
  assign n84 = ~n82 & n83 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = k_pad & l_pad ;
  assign n88 = ~m_pad & ~n86 ;
  assign n87 = m_pad & n86 ;
  assign n89 = ~a_pad & ~n87 ;
  assign n90 = ~n88 & n89 ;
  assign n93 = ~n_pad & ~n87 ;
  assign n92 = n_pad & n87 ;
  assign n91 = ~m_pad & n81 ;
  assign n94 = ~a_pad & ~n91 ;
  assign n95 = ~n92 & n94 ;
  assign n96 = ~n93 & n95 ;
  assign n97 = n81 & n82 ;
  assign n98 = ~x_pad & ~n97 ;
  assign n100 = ~o_pad & n98 ;
  assign n99 = o_pad & ~n98 ;
  assign n101 = ~a_pad & ~n99 ;
  assign n102 = ~n100 & n101 ;
  assign n104 = ~q_pad & r_pad ;
  assign n105 = n99 & ~n104 ;
  assign n106 = ~p_pad & ~n105 ;
  assign n103 = p_pad & n99 ;
  assign n107 = ~a_pad & ~n103 ;
  assign n108 = ~n106 & n107 ;
  assign n110 = q_pad & n103 ;
  assign n109 = ~q_pad & ~n103 ;
  assign n111 = ~a_pad & ~n109 ;
  assign n112 = ~n110 & n111 ;
  assign n118 = ~r_pad & ~n110 ;
  assign n113 = ~p_pad & ~q_pad ;
  assign n114 = p_pad & q_pad ;
  assign n115 = r_pad & n114 ;
  assign n116 = ~n113 & ~n115 ;
  assign n117 = n99 & ~n116 ;
  assign n119 = ~a_pad & ~n117 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = ~p_pad & n104 ;
  assign n122 = n99 & n121 ;
  assign n124 = s_pad & n122 ;
  assign n123 = ~s_pad & ~n122 ;
  assign n125 = ~a_pad & ~n123 ;
  assign n126 = ~n124 & n125 ;
  assign n128 = ~n34 & n124 ;
  assign n129 = ~t_pad & ~n128 ;
  assign n127 = t_pad & n124 ;
  assign n130 = ~a_pad & ~n127 ;
  assign n131 = ~n129 & n130 ;
  assign n132 = u_pad & ~n127 ;
  assign n133 = n69 & n122 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = ~a_pad & ~n134 ;
  assign n136 = ~t_pad & u_pad ;
  assign n137 = ~n68 & ~n136 ;
  assign n138 = n124 & n137 ;
  assign n139 = v_pad & ~n138 ;
  assign n140 = n33 & n127 ;
  assign n141 = ~n139 & ~n140 ;
  assign n142 = ~a_pad & ~n141 ;
  assign n143 = y_pad & n73 ;
  assign n144 = n136 & n143 ;
  assign n145 = ~w_pad & ~n144 ;
  assign n146 = ~a_pad & ~n30 ;
  assign n147 = ~n145 & n146 ;
  assign n148 = b_pad & ~x_pad ;
  assign n149 = ~b_pad & x_pad ;
  assign n150 = ~n148 & ~n149 ;
  assign n151 = ~a_pad & ~n150 ;
  assign n152 = c_pad & ~y_pad ;
  assign n153 = ~c_pad & y_pad ;
  assign n154 = ~n152 & ~n153 ;
  assign n155 = ~a_pad & ~n154 ;
  assign n156 = e_pad & ~n37 ;
  assign n157 = v_pad & ~n61 ;
  assign n158 = ~n156 & n157 ;
  assign n159 = ~w_pad & ~n33 ;
  assign n160 = ~n158 & n159 ;
  assign \a0_pad  = n43 ;
  assign \b0_pad  = n51 ;
  assign \c0_pad  = n65 ;
  assign \d0_pad  = n72 ;
  assign \e0_pad  = n78 ;
  assign \f0_pad  = n79 ;
  assign \g0_pad  = ~n85 ;
  assign \h0_pad  = n90 ;
  assign \i0_pad  = n96 ;
  assign \j0_pad  = n102 ;
  assign \k0_pad  = n108 ;
  assign \l0_pad  = n112 ;
  assign \m0_pad  = n120 ;
  assign \n0_pad  = n126 ;
  assign \o0_pad  = n131 ;
  assign \p0_pad  = n135 ;
  assign \q0_pad  = n142 ;
  assign \r0_pad  = n147 ;
  assign \s0_pad  = n151 ;
  assign \t0_pad  = n155 ;
  assign z_pad = n160 ;
endmodule
