module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  output v_pad ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n55 = ~c_pad & ~s_pad ;
  assign n54 = ~a_pad & s_pad ;
  assign n56 = t_pad & ~n54 ;
  assign n57 = ~n55 & n56 ;
  assign n59 = ~b_pad & s_pad ;
  assign n58 = ~d_pad & ~s_pad ;
  assign n60 = ~t_pad & ~n58 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = ~n57 & ~n61 ;
  assign n63 = r_pad & ~n62 ;
  assign n45 = ~h_pad & ~s_pad ;
  assign n44 = ~f_pad & s_pad ;
  assign n46 = ~t_pad & ~n44 ;
  assign n47 = ~n45 & n46 ;
  assign n49 = ~e_pad & s_pad ;
  assign n48 = ~g_pad & ~s_pad ;
  assign n50 = t_pad & ~n48 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = ~n47 & ~n51 ;
  assign n53 = ~r_pad & ~n52 ;
  assign n64 = q_pad & ~n53 ;
  assign n65 = ~n63 & n64 ;
  assign n33 = ~i_pad & s_pad ;
  assign n32 = ~k_pad & ~s_pad ;
  assign n34 = t_pad & ~n32 ;
  assign n35 = ~n33 & n34 ;
  assign n37 = ~l_pad & ~s_pad ;
  assign n36 = ~j_pad & s_pad ;
  assign n38 = ~t_pad & ~n36 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = ~n35 & ~n39 ;
  assign n41 = r_pad & ~n40 ;
  assign n23 = ~p_pad & ~s_pad ;
  assign n22 = ~n_pad & s_pad ;
  assign n24 = ~t_pad & ~n22 ;
  assign n25 = ~n23 & n24 ;
  assign n27 = ~m_pad & s_pad ;
  assign n26 = ~o_pad & ~s_pad ;
  assign n28 = t_pad & ~n26 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = ~r_pad & ~n30 ;
  assign n42 = ~q_pad & ~n31 ;
  assign n43 = ~n41 & n42 ;
  assign n66 = u_pad & ~n43 ;
  assign n67 = ~n65 & n66 ;
  assign v_pad = n67 ;
endmodule
