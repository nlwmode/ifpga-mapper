module top( ctr_pad , \cts_reg/NET0131  , g_button_pad , key_pad , \last_g_reg/NET0131  , \last_r_reg/NET0131  , r_button_pad , rtr_pad , rts_pad , \sign_reg[3]/NET0131  , start_pad , \stato_reg[0]/NET0131  , \stato_reg[1]/NET0131  , \stato_reg[2]/NET0131  , \stato_reg[3]/NET0131  , test_pad , \v_in[0]_pad  , \v_in[1]_pad  , \v_in[2]_pad  , \v_in[3]_pad  , \v_out_reg[0]/NET0131  , \v_out_reg[1]/NET0131  , \v_out_reg[2]/NET0131  , \v_out_reg[3]/NET0131  , \voto0_reg/NET0131  , \voto1_reg/NET0131  , \voto2_reg/NET0131  , \voto3_reg/NET0131  , \_al_n0  , \_al_n1  , \g1181/_2_  , \g1199/_0_  , \g1200/_0_  , \g1201/_0_  , \g1202/_0_  , \g1205/_0_  , \g1208/_0_  , \g1209/_0_  , \g1210/_0_  , \g1211/_0_  , \g1212/_0_  , \g1216/_0_  , \g1217/_0_  , \g1218/_0_  , \g1219/_0_  , \g1579/_0_  , \g36/_0_  );
  input ctr_pad ;
  input \cts_reg/NET0131  ;
  input g_button_pad ;
  input key_pad ;
  input \last_g_reg/NET0131  ;
  input \last_r_reg/NET0131  ;
  input r_button_pad ;
  input rtr_pad ;
  input rts_pad ;
  input \sign_reg[3]/NET0131  ;
  input start_pad ;
  input \stato_reg[0]/NET0131  ;
  input \stato_reg[1]/NET0131  ;
  input \stato_reg[2]/NET0131  ;
  input \stato_reg[3]/NET0131  ;
  input test_pad ;
  input \v_in[0]_pad  ;
  input \v_in[1]_pad  ;
  input \v_in[2]_pad  ;
  input \v_in[3]_pad  ;
  input \v_out_reg[0]/NET0131  ;
  input \v_out_reg[1]/NET0131  ;
  input \v_out_reg[2]/NET0131  ;
  input \v_out_reg[3]/NET0131  ;
  input \voto0_reg/NET0131  ;
  input \voto1_reg/NET0131  ;
  input \voto2_reg/NET0131  ;
  input \voto3_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1181/_2_  ;
  output \g1199/_0_  ;
  output \g1200/_0_  ;
  output \g1201/_0_  ;
  output \g1202/_0_  ;
  output \g1205/_0_  ;
  output \g1208/_0_  ;
  output \g1209/_0_  ;
  output \g1210/_0_  ;
  output \g1211/_0_  ;
  output \g1212/_0_  ;
  output \g1216/_0_  ;
  output \g1217/_0_  ;
  output \g1218/_0_  ;
  output \g1219/_0_  ;
  output \g1579/_0_  ;
  output \g36/_0_  ;
  wire n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 ;
  assign n35 = ~\stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n38 = ~\stato_reg[3]/NET0131  & n35 ;
  assign n39 = ~\stato_reg[0]/NET0131  & n38 ;
  assign n40 = \voto1_reg/NET0131  & \voto2_reg/NET0131  ;
  assign n41 = rtr_pad & ~\voto0_reg/NET0131  ;
  assign n42 = ~\voto3_reg/NET0131  & n41 ;
  assign n43 = n40 & n42 ;
  assign n44 = n39 & ~n43 ;
  assign n45 = ~rtr_pad & ~\stato_reg[2]/NET0131  ;
  assign n46 = n44 & ~n45 ;
  assign n29 = \stato_reg[1]/NET0131  & \stato_reg[2]/NET0131  ;
  assign n30 = ~\stato_reg[3]/NET0131  & n29 ;
  assign n31 = \stato_reg[1]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n32 = ~\stato_reg[0]/NET0131  & \stato_reg[3]/NET0131  ;
  assign n33 = n31 & n32 ;
  assign n34 = ~n30 & ~n33 ;
  assign n36 = \stato_reg[0]/NET0131  & ~\stato_reg[3]/NET0131  ;
  assign n37 = n35 & n36 ;
  assign n47 = n31 & n36 ;
  assign n48 = ~n37 & ~n47 ;
  assign n49 = n34 & n48 ;
  assign n50 = ~n46 & n49 ;
  assign n51 = ~\stato_reg[1]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n52 = n36 & n51 ;
  assign n53 = ~start_pad & n52 ;
  assign n54 = n29 & n36 ;
  assign n55 = ~n53 & ~n54 ;
  assign n56 = ~n33 & n55 ;
  assign n57 = ~\stato_reg[0]/NET0131  & ~\stato_reg[3]/NET0131  ;
  assign n58 = n31 & n57 ;
  assign n59 = ~start_pad & n58 ;
  assign n60 = n32 & n51 ;
  assign n61 = ~n38 & ~n60 ;
  assign n62 = ~n59 & n61 ;
  assign n63 = n56 & n62 ;
  assign n64 = \voto1_reg/NET0131  & ~n63 ;
  assign n67 = n29 & n57 ;
  assign n71 = ~rts_pad & n67 ;
  assign n72 = ~n47 & ~n71 ;
  assign n73 = \voto1_reg/NET0131  & ~n72 ;
  assign n65 = \stato_reg[3]/NET0131  & n51 ;
  assign n66 = \stato_reg[0]/NET0131  & n65 ;
  assign n68 = rts_pad & n67 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = \v_in[1]_pad  & ~n69 ;
  assign n74 = key_pad & start_pad ;
  assign n75 = n58 & n74 ;
  assign n76 = g_button_pad & ~\last_g_reg/NET0131  ;
  assign n77 = ~\voto1_reg/NET0131  & ~n76 ;
  assign n78 = \voto1_reg/NET0131  & n76 ;
  assign n79 = ~n77 & ~n78 ;
  assign n80 = n75 & n79 ;
  assign n81 = ~n70 & ~n80 ;
  assign n82 = ~n73 & n81 ;
  assign n83 = ~n64 & n82 ;
  assign n92 = ~\last_r_reg/NET0131  & r_button_pad ;
  assign n93 = n75 & n92 ;
  assign n94 = ~\voto2_reg/NET0131  & ~n93 ;
  assign n95 = n75 & ~n92 ;
  assign n96 = \voto2_reg/NET0131  & n61 ;
  assign n97 = ~n95 & n96 ;
  assign n98 = ~n94 & ~n97 ;
  assign n84 = \voto2_reg/NET0131  & ~n56 ;
  assign n86 = \voto2_reg/NET0131  & n59 ;
  assign n85 = \v_in[2]_pad  & n66 ;
  assign n87 = \voto2_reg/NET0131  & n47 ;
  assign n88 = rts_pad & ~\v_in[2]_pad  ;
  assign n89 = ~rts_pad & ~\voto2_reg/NET0131  ;
  assign n90 = ~n88 & ~n89 ;
  assign n91 = n67 & n90 ;
  assign n99 = ~n87 & ~n91 ;
  assign n100 = ~n85 & n99 ;
  assign n101 = ~n86 & n100 ;
  assign n102 = ~n84 & n101 ;
  assign n103 = ~n98 & n102 ;
  assign n106 = n39 & n43 ;
  assign n104 = ~rtr_pad & ~\stato_reg[0]/NET0131  ;
  assign n105 = n65 & ~n104 ;
  assign n107 = n51 & n57 ;
  assign n108 = ~test_pad & n107 ;
  assign n109 = ~n105 & ~n108 ;
  assign n110 = ~n106 & n109 ;
  assign n113 = \v_in[0]_pad  & \v_in[1]_pad  ;
  assign n114 = \v_in[2]_pad  & \v_in[3]_pad  ;
  assign n115 = n113 & n114 ;
  assign n116 = n66 & n115 ;
  assign n111 = rtr_pad & n54 ;
  assign n112 = \stato_reg[1]/NET0131  & n57 ;
  assign n119 = ~n111 & ~n112 ;
  assign n117 = start_pad & n52 ;
  assign n118 = ~rts_pad & n37 ;
  assign n120 = ~n117 & ~n118 ;
  assign n121 = n119 & n120 ;
  assign n122 = ~n116 & n121 ;
  assign n123 = ~n36 & ~n112 ;
  assign n124 = ~n29 & ~n123 ;
  assign n125 = n34 & ~n51 ;
  assign n126 = ~n124 & n125 ;
  assign n127 = ~rtr_pad & n39 ;
  assign n128 = n126 & ~n127 ;
  assign n129 = \v_out_reg[3]/NET0131  & ~n128 ;
  assign n130 = rtr_pad & \voto3_reg/NET0131  ;
  assign n131 = n39 & n130 ;
  assign n132 = ~n129 & ~n131 ;
  assign n133 = ~\stato_reg[0]/NET0131  & ~\stato_reg[2]/NET0131  ;
  assign n134 = \stato_reg[3]/NET0131  & ~n133 ;
  assign n135 = \sign_reg[3]/NET0131  & ~n134 ;
  assign n136 = ~n108 & n135 ;
  assign n137 = ~n66 & ~n136 ;
  assign n138 = \v_out_reg[0]/NET0131  & ~n128 ;
  assign n139 = rtr_pad & \voto0_reg/NET0131  ;
  assign n140 = n39 & n139 ;
  assign n141 = ~n138 & ~n140 ;
  assign n142 = \v_out_reg[1]/NET0131  & ~n128 ;
  assign n143 = rtr_pad & \voto1_reg/NET0131  ;
  assign n144 = n39 & n143 ;
  assign n145 = ~n142 & ~n144 ;
  assign n146 = \v_out_reg[2]/NET0131  & ~n126 ;
  assign n147 = ~rtr_pad & ~\v_out_reg[2]/NET0131  ;
  assign n148 = rtr_pad & ~\voto2_reg/NET0131  ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n39 & n149 ;
  assign n151 = ~n146 & ~n150 ;
  assign n152 = ~key_pad & start_pad ;
  assign n153 = n58 & ~n152 ;
  assign n154 = n61 & ~n153 ;
  assign n155 = n56 & n154 ;
  assign n156 = \voto3_reg/NET0131  & ~n155 ;
  assign n159 = ~\voto1_reg/NET0131  & ~\voto2_reg/NET0131  ;
  assign n160 = ~n40 & ~n159 ;
  assign n162 = ~\voto0_reg/NET0131  & ~n160 ;
  assign n161 = \voto0_reg/NET0131  & n160 ;
  assign n163 = n47 & ~n161 ;
  assign n164 = ~n162 & n163 ;
  assign n157 = \v_in[3]_pad  & ~n69 ;
  assign n158 = \voto3_reg/NET0131  & n71 ;
  assign n165 = ~n157 & ~n158 ;
  assign n166 = ~n164 & n165 ;
  assign n167 = ~n156 & n166 ;
  assign n174 = ~n38 & ~n47 ;
  assign n175 = ~n112 & n174 ;
  assign n176 = ~n66 & n175 ;
  assign n177 = \cts_reg/NET0131  & ~n176 ;
  assign n168 = ~n54 & ~n60 ;
  assign n169 = rtr_pad & ~n168 ;
  assign n170 = ~n33 & ~n169 ;
  assign n171 = \cts_reg/NET0131  & ~n170 ;
  assign n172 = ~n39 & ~n52 ;
  assign n173 = rtr_pad & ~n172 ;
  assign n178 = ~n171 & ~n173 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = ~\stato_reg[0]/NET0131  & n31 ;
  assign n181 = \stato_reg[3]/NET0131  & ~n51 ;
  assign n182 = ~n180 & n181 ;
  assign n183 = ~n58 & ~n182 ;
  assign n184 = \last_g_reg/NET0131  & n183 ;
  assign n186 = ~g_button_pad & n74 ;
  assign n185 = ~\last_g_reg/NET0131  & ~n74 ;
  assign n187 = n58 & ~n185 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = ~n184 & ~n188 ;
  assign n190 = \last_r_reg/NET0131  & n183 ;
  assign n192 = ~r_button_pad & n74 ;
  assign n191 = ~\last_r_reg/NET0131  & ~n74 ;
  assign n193 = n58 & ~n191 ;
  assign n194 = ~n192 & n193 ;
  assign n195 = ~n190 & ~n194 ;
  assign n196 = n61 & ~n71 ;
  assign n197 = n55 & n196 ;
  assign n198 = \voto0_reg/NET0131  & ~n197 ;
  assign n199 = \v_in[0]_pad  & ~n69 ;
  assign n200 = ~start_pad & ~\voto0_reg/NET0131  ;
  assign n201 = n153 & ~n200 ;
  assign n202 = ~\sign_reg[3]/NET0131  & n33 ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = ~n199 & n203 ;
  assign n205 = ~n198 & n204 ;
  assign n206 = ~n36 & ~n65 ;
  assign n207 = ~n180 & n206 ;
  assign n208 = ~n39 & ~n71 ;
  assign n209 = n207 & n208 ;
  assign n210 = ctr_pad & ~n209 ;
  assign n211 = ~n118 & ~n210 ;
  assign n212 = ~n44 & ~n54 ;
  assign n213 = rtr_pad & ~n212 ;
  assign n216 = \stato_reg[0]/NET0131  & ~n115 ;
  assign n217 = ~n104 & ~n216 ;
  assign n218 = n65 & ~n217 ;
  assign n214 = ~n37 & ~n67 ;
  assign n215 = rts_pad & ~n214 ;
  assign n219 = ~n53 & ~n107 ;
  assign n220 = ~n59 & n219 ;
  assign n221 = ~n215 & n220 ;
  assign n222 = ~n218 & n221 ;
  assign n223 = ~n213 & n222 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1181/_2_  = ~n50 ;
  assign \g1199/_0_  = ~n83 ;
  assign \g1200/_0_  = ~n103 ;
  assign \g1201/_0_  = ~n110 ;
  assign \g1202/_0_  = ~n122 ;
  assign \g1205/_0_  = ~n132 ;
  assign \g1208/_0_  = ~n137 ;
  assign \g1209/_0_  = ~n141 ;
  assign \g1210/_0_  = ~n145 ;
  assign \g1211/_0_  = ~n151 ;
  assign \g1212/_0_  = ~n167 ;
  assign \g1216/_0_  = ~n179 ;
  assign \g1217/_0_  = ~n189 ;
  assign \g1218/_0_  = ~n195 ;
  assign \g1219/_0_  = ~n205 ;
  assign \g1579/_0_  = ~n211 ;
  assign \g36/_0_  = ~n223 ;
endmodule
