module top (\102GAT(31)_pad , \105GAT(32)_pad , \108GAT(33)_pad , \112GAT(34)_pad , \115GAT(35)_pad , \11GAT(3)_pad , \14GAT(4)_pad , \17GAT(5)_pad , \1GAT(0)_pad , \21GAT(6)_pad , \24GAT(7)_pad , \27GAT(8)_pad , \30GAT(9)_pad , \34GAT(10)_pad , \37GAT(11)_pad , \40GAT(12)_pad , \43GAT(13)_pad , \47GAT(14)_pad , \4GAT(1)_pad , \50GAT(15)_pad , \53GAT(16)_pad , \56GAT(17)_pad , \60GAT(18)_pad , \63GAT(19)_pad , \66GAT(20)_pad , \69GAT(21)_pad , \73GAT(22)_pad , \76GAT(23)_pad , \79GAT(24)_pad , \82GAT(25)_pad , \86GAT(26)_pad , \89GAT(27)_pad , \8GAT(2)_pad , \92GAT(28)_pad , \95GAT(29)_pad , \99GAT(30)_pad , \203GAT(82) , \309GAT(131) , \360GAT(162) , \421GAT(188)_pad , \430GAT(193)_pad , \431GAT(194)_pad , \432GAT(195)_pad );
	input \102GAT(31)_pad  ;
	input \105GAT(32)_pad  ;
	input \108GAT(33)_pad  ;
	input \112GAT(34)_pad  ;
	input \115GAT(35)_pad  ;
	input \11GAT(3)_pad  ;
	input \14GAT(4)_pad  ;
	input \17GAT(5)_pad  ;
	input \1GAT(0)_pad  ;
	input \21GAT(6)_pad  ;
	input \24GAT(7)_pad  ;
	input \27GAT(8)_pad  ;
	input \30GAT(9)_pad  ;
	input \34GAT(10)_pad  ;
	input \37GAT(11)_pad  ;
	input \40GAT(12)_pad  ;
	input \43GAT(13)_pad  ;
	input \47GAT(14)_pad  ;
	input \4GAT(1)_pad  ;
	input \50GAT(15)_pad  ;
	input \53GAT(16)_pad  ;
	input \56GAT(17)_pad  ;
	input \60GAT(18)_pad  ;
	input \63GAT(19)_pad  ;
	input \66GAT(20)_pad  ;
	input \69GAT(21)_pad  ;
	input \73GAT(22)_pad  ;
	input \76GAT(23)_pad  ;
	input \79GAT(24)_pad  ;
	input \82GAT(25)_pad  ;
	input \86GAT(26)_pad  ;
	input \89GAT(27)_pad  ;
	input \8GAT(2)_pad  ;
	input \92GAT(28)_pad  ;
	input \95GAT(29)_pad  ;
	input \99GAT(30)_pad  ;
	output \203GAT(82)  ;
	output \309GAT(131)  ;
	output \360GAT(162)  ;
	output \421GAT(188)_pad  ;
	output \430GAT(193)_pad  ;
	output \431GAT(194)_pad  ;
	output \432GAT(195)_pad  ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\50GAT(15)_pad ,
		\56GAT(17)_pad ,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\24GAT(7)_pad ,
		\30GAT(9)_pad ,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\63GAT(19)_pad ,
		\69GAT(21)_pad ,
		_w39_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\102GAT(31)_pad ,
		\108GAT(33)_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\76GAT(23)_pad ,
		\82GAT(25)_pad ,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\37GAT(11)_pad ,
		\43GAT(13)_pad ,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\11GAT(3)_pad ,
		\17GAT(5)_pad ,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\1GAT(0)_pad ,
		\4GAT(1)_pad ,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\89GAT(27)_pad ,
		\95GAT(29)_pad ,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w37_,
		_w38_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w39_,
		_w40_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w41_,
		_w42_,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w43_,
		_w44_,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w45_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w47_,
		_w48_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w46_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w50_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\1GAT(0)_pad ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\4GAT(1)_pad ,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\8GAT(2)_pad ,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\50GAT(15)_pad ,
		_w53_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\56GAT(17)_pad ,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\60GAT(18)_pad ,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\89GAT(27)_pad ,
		_w53_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\95GAT(29)_pad ,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\99GAT(30)_pad ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\24GAT(7)_pad ,
		_w53_,
		_w63_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\30GAT(9)_pad ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\34GAT(10)_pad ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\11GAT(3)_pad ,
		_w53_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\17GAT(5)_pad ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\21GAT(6)_pad ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\102GAT(31)_pad ,
		_w53_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\108GAT(33)_pad ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\112GAT(34)_pad ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\37GAT(11)_pad ,
		_w53_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\43GAT(13)_pad ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\47GAT(14)_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\63GAT(19)_pad ,
		_w53_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\69GAT(21)_pad ,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\73GAT(22)_pad ,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\76GAT(23)_pad ,
		_w53_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\76GAT(23)_pad ,
		_w53_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\82GAT(25)_pad ,
		\86GAT(26)_pad ,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w56_,
		_w59_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w62_,
		_w65_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w68_,
		_w71_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w74_,
		_w77_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w82_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w84_,
		_w85_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w83_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w87_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\34GAT(10)_pad ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		_w64_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		\40GAT(12)_pad ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\21GAT(6)_pad ,
		_w90_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		_w67_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\27GAT(8)_pad ,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\73GAT(22)_pad ,
		_w90_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		_w76_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\79GAT(24)_pad ,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\112GAT(34)_pad ,
		_w90_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		_w70_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\115GAT(35)_pad ,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\47GAT(14)_pad ,
		_w90_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		_w73_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		\53GAT(16)_pad ,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\8GAT(2)_pad ,
		_w90_,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		_w55_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		\14GAT(4)_pad ,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\99GAT(30)_pad ,
		_w90_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		_w61_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\105GAT(32)_pad ,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		\60GAT(18)_pad ,
		_w90_,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		_w58_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		\66GAT(20)_pad ,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\86GAT(26)_pad ,
		_w90_,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\82GAT(25)_pad ,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w82_,
		_w90_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		\92GAT(28)_pad ,
		_w80_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w116_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w93_,
		_w96_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w99_,
		_w102_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w105_,
		_w108_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w111_,
		_w114_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w120_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w122_,
		_w123_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w121_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w125_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\66GAT(20)_pad ,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		_w113_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\53GAT(16)_pad ,
		_w128_,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w104_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w130_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\40GAT(12)_pad ,
		_w128_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w92_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\27GAT(8)_pad ,
		_w128_,
		_w136_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		_w95_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w135_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w133_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\105GAT(32)_pad ,
		_w128_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		_w110_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\115GAT(35)_pad ,
		_w128_,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		_w101_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\92GAT(28)_pad ,
		_w128_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w78_,
		_w116_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w144_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name110 (
		\79GAT(24)_pad ,
		_w128_,
		_w147_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		_w98_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w141_,
		_w143_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w146_,
		_w148_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w139_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\14GAT(4)_pad ,
		_w128_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		_w107_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w152_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		_w135_,
		_w148_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w146_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		_w133_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w138_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		_w141_,
		_w146_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w132_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w135_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w133_,
		_w156_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w137_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w162_,
		_w164_,
		_w165_
	);
	assign \203GAT(82)  = _w53_ ;
	assign \309GAT(131)  = _w90_ ;
	assign \360GAT(162)  = _w128_ ;
	assign \421GAT(188)_pad  = _w155_ ;
	assign \430GAT(193)_pad  = _w139_ ;
	assign \431GAT(194)_pad  = _w159_ ;
	assign \432GAT(195)_pad  = _w165_ ;
endmodule;