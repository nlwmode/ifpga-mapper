module top( \ccyc_addr_in[0]_pad  , \ccyc_addr_in[11]_pad  , \ccyc_addr_in[12]_pad  , \ccyc_addr_in[13]_pad  , \ccyc_addr_in[14]_pad  , \ccyc_addr_in[15]_pad  , \ccyc_addr_in[16]_pad  , \ccyc_addr_in[17]_pad  , \ccyc_addr_in[18]_pad  , \ccyc_addr_in[19]_pad  , \ccyc_addr_in[20]_pad  , \ccyc_addr_in[21]_pad  , \ccyc_addr_in[22]_pad  , \ccyc_addr_in[23]_pad  , \ccyc_addr_in[24]_pad  , \ccyc_addr_in[25]_pad  , \ccyc_addr_in[26]_pad  , \ccyc_addr_in[27]_pad  , \ccyc_addr_in[28]_pad  , \ccyc_addr_in[29]_pad  , \ccyc_addr_in[30]_pad  , \ccyc_addr_in[31]_pad  , \ccyc_addr_out[11]_pad  , \ccyc_addr_out[12]_pad  , \ccyc_addr_out[13]_pad  , \ccyc_addr_out[14]_pad  , \ccyc_addr_out[15]_pad  , \ccyc_addr_out[16]_pad  , \ccyc_addr_out[17]_pad  , \ccyc_addr_out[18]_pad  , \ccyc_addr_out[19]_pad  , \ccyc_addr_out[20]_pad  , \ccyc_addr_out[21]_pad  , \ccyc_addr_out[22]_pad  , \ccyc_addr_out[23]_pad  , \ccyc_addr_out[24]_pad  , \ccyc_addr_out[25]_pad  , \ccyc_addr_out[26]_pad  , \ccyc_addr_out[27]_pad  , \ccyc_addr_out[28]_pad  , \ccyc_addr_out[29]_pad  , \ccyc_addr_out[30]_pad  , \ccyc_addr_out[31]_pad  );
  input \ccyc_addr_in[0]_pad  ;
  input \ccyc_addr_in[11]_pad  ;
  input \ccyc_addr_in[12]_pad  ;
  input \ccyc_addr_in[13]_pad  ;
  input \ccyc_addr_in[14]_pad  ;
  input \ccyc_addr_in[15]_pad  ;
  input \ccyc_addr_in[16]_pad  ;
  input \ccyc_addr_in[17]_pad  ;
  input \ccyc_addr_in[18]_pad  ;
  input \ccyc_addr_in[19]_pad  ;
  input \ccyc_addr_in[20]_pad  ;
  input \ccyc_addr_in[21]_pad  ;
  input \ccyc_addr_in[22]_pad  ;
  input \ccyc_addr_in[23]_pad  ;
  input \ccyc_addr_in[24]_pad  ;
  input \ccyc_addr_in[25]_pad  ;
  input \ccyc_addr_in[26]_pad  ;
  input \ccyc_addr_in[27]_pad  ;
  input \ccyc_addr_in[28]_pad  ;
  input \ccyc_addr_in[29]_pad  ;
  input \ccyc_addr_in[30]_pad  ;
  input \ccyc_addr_in[31]_pad  ;
  output \ccyc_addr_out[11]_pad  ;
  output \ccyc_addr_out[12]_pad  ;
  output \ccyc_addr_out[13]_pad  ;
  output \ccyc_addr_out[14]_pad  ;
  output \ccyc_addr_out[15]_pad  ;
  output \ccyc_addr_out[16]_pad  ;
  output \ccyc_addr_out[17]_pad  ;
  output \ccyc_addr_out[18]_pad  ;
  output \ccyc_addr_out[19]_pad  ;
  output \ccyc_addr_out[20]_pad  ;
  output \ccyc_addr_out[21]_pad  ;
  output \ccyc_addr_out[22]_pad  ;
  output \ccyc_addr_out[23]_pad  ;
  output \ccyc_addr_out[24]_pad  ;
  output \ccyc_addr_out[25]_pad  ;
  output \ccyc_addr_out[26]_pad  ;
  output \ccyc_addr_out[27]_pad  ;
  output \ccyc_addr_out[28]_pad  ;
  output \ccyc_addr_out[29]_pad  ;
  output \ccyc_addr_out[30]_pad  ;
  output \ccyc_addr_out[31]_pad  ;
  wire n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 ;
  assign n23 = ~\ccyc_addr_in[14]_pad  & ~\ccyc_addr_in[15]_pad  ;
  assign n24 = ~\ccyc_addr_in[12]_pad  & ~\ccyc_addr_in[13]_pad  ;
  assign n25 = n23 & n24 ;
  assign n26 = ~\ccyc_addr_in[0]_pad  & ~n25 ;
  assign n27 = ~\ccyc_addr_in[0]_pad  & ~\ccyc_addr_in[11]_pad  ;
  assign n28 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[11]_pad  ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = ~n26 & ~n29 ;
  assign n31 = ~\ccyc_addr_in[0]_pad  & \ccyc_addr_in[11]_pad  ;
  assign n32 = ~\ccyc_addr_in[12]_pad  & ~n31 ;
  assign n33 = ~n26 & ~n32 ;
  assign n34 = \ccyc_addr_in[12]_pad  & ~\ccyc_addr_in[13]_pad  ;
  assign n35 = n23 & n34 ;
  assign n36 = n27 & n35 ;
  assign n37 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[13]_pad  ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = n31 & n35 ;
  assign n40 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[14]_pad  ;
  assign n41 = ~n39 & ~n40 ;
  assign n42 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[15]_pad  ;
  assign n43 = ~\ccyc_addr_in[12]_pad  & \ccyc_addr_in[13]_pad  ;
  assign n44 = n23 & n43 ;
  assign n45 = n27 & n44 ;
  assign n46 = ~n42 & ~n45 ;
  assign n47 = n31 & n44 ;
  assign n48 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[16]_pad  ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = \ccyc_addr_in[12]_pad  & \ccyc_addr_in[13]_pad  ;
  assign n51 = n23 & n50 ;
  assign n52 = n27 & n51 ;
  assign n53 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[17]_pad  ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = n31 & n51 ;
  assign n56 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[18]_pad  ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = \ccyc_addr_in[14]_pad  & ~\ccyc_addr_in[15]_pad  ;
  assign n59 = n24 & n58 ;
  assign n60 = n27 & n59 ;
  assign n61 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[19]_pad  ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = n31 & n59 ;
  assign n64 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[20]_pad  ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = n34 & n58 ;
  assign n67 = n27 & n66 ;
  assign n68 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[21]_pad  ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = n31 & n66 ;
  assign n71 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[22]_pad  ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[23]_pad  ;
  assign n74 = n43 & n58 ;
  assign n75 = n27 & n74 ;
  assign n76 = ~n73 & ~n75 ;
  assign n77 = n31 & n74 ;
  assign n78 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[24]_pad  ;
  assign n79 = ~n77 & ~n78 ;
  assign n80 = n50 & n58 ;
  assign n81 = n27 & n80 ;
  assign n82 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[25]_pad  ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = n31 & n80 ;
  assign n85 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[26]_pad  ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = ~\ccyc_addr_in[14]_pad  & \ccyc_addr_in[15]_pad  ;
  assign n88 = n24 & n87 ;
  assign n89 = n27 & n88 ;
  assign n90 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[27]_pad  ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = n31 & n88 ;
  assign n93 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[28]_pad  ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = n34 & n87 ;
  assign n96 = n27 & n95 ;
  assign n97 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[29]_pad  ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = n31 & n95 ;
  assign n100 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[30]_pad  ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = \ccyc_addr_in[0]_pad  & \ccyc_addr_in[31]_pad  ;
  assign n103 = n27 & n43 ;
  assign n104 = n87 & n103 ;
  assign n105 = ~n102 & ~n104 ;
  assign \ccyc_addr_out[11]_pad  = n30 ;
  assign \ccyc_addr_out[12]_pad  = n33 ;
  assign \ccyc_addr_out[13]_pad  = ~n38 ;
  assign \ccyc_addr_out[14]_pad  = ~n41 ;
  assign \ccyc_addr_out[15]_pad  = ~n46 ;
  assign \ccyc_addr_out[16]_pad  = ~n49 ;
  assign \ccyc_addr_out[17]_pad  = ~n54 ;
  assign \ccyc_addr_out[18]_pad  = ~n57 ;
  assign \ccyc_addr_out[19]_pad  = ~n62 ;
  assign \ccyc_addr_out[20]_pad  = ~n65 ;
  assign \ccyc_addr_out[21]_pad  = ~n69 ;
  assign \ccyc_addr_out[22]_pad  = ~n72 ;
  assign \ccyc_addr_out[23]_pad  = ~n76 ;
  assign \ccyc_addr_out[24]_pad  = ~n79 ;
  assign \ccyc_addr_out[25]_pad  = ~n83 ;
  assign \ccyc_addr_out[26]_pad  = ~n86 ;
  assign \ccyc_addr_out[27]_pad  = ~n91 ;
  assign \ccyc_addr_out[28]_pad  = ~n94 ;
  assign \ccyc_addr_out[29]_pad  = ~n98 ;
  assign \ccyc_addr_out[30]_pad  = ~n101 ;
  assign \ccyc_addr_out[31]_pad  = ~n105 ;
endmodule
