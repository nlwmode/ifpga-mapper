module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, \j0_pad , j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u0_pad , \v0_pad , \w0_pad , \x0_pad , \y0_pad , \z0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u0_pad  ;
	output \v0_pad  ;
	output \w0_pad  ;
	output \x0_pad  ;
	output \y0_pad  ;
	output \z0_pad  ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	LUT3 #(
		.INIT('h82)
	) name0 (
		q_pad,
		r_pad,
		u_pad,
		_w37_
	);
	LUT3 #(
		.INIT('h0e)
	) name1 (
		p_pad,
		q_pad,
		s_pad,
		_w38_
	);
	LUT2 #(
		.INIT('hb)
	) name2 (
		_w37_,
		_w38_,
		_w39_
	);
	LUT4 #(
		.INIT('h57fd)
	) name3 (
		q_pad,
		r_pad,
		u_pad,
		v_pad,
		_w40_
	);
	LUT3 #(
		.INIT('h0e)
	) name4 (
		o_pad,
		q_pad,
		s_pad,
		_w41_
	);
	LUT2 #(
		.INIT('h7)
	) name5 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		r_pad,
		u_pad,
		v_pad,
		_w43_
	);
	LUT3 #(
		.INIT('h0e)
	) name7 (
		n_pad,
		q_pad,
		s_pad,
		_w44_
	);
	LUT4 #(
		.INIT('h28ff)
	) name8 (
		q_pad,
		w_pad,
		_w43_,
		_w44_,
		_w45_
	);
	LUT4 #(
		.INIT('h0001)
	) name9 (
		r_pad,
		u_pad,
		v_pad,
		w_pad,
		_w46_
	);
	LUT3 #(
		.INIT('h0e)
	) name10 (
		m_pad,
		q_pad,
		s_pad,
		_w47_
	);
	LUT4 #(
		.INIT('h28ff)
	) name11 (
		q_pad,
		x_pad,
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		q_pad,
		y_pad,
		_w49_
	);
	LUT3 #(
		.INIT('hb0)
	) name13 (
		x_pad,
		_w46_,
		_w49_,
		_w50_
	);
	LUT3 #(
		.INIT('h02)
	) name14 (
		q_pad,
		x_pad,
		y_pad,
		_w51_
	);
	LUT3 #(
		.INIT('h0e)
	) name15 (
		l_pad,
		q_pad,
		s_pad,
		_w52_
	);
	LUT3 #(
		.INIT('h70)
	) name16 (
		_w46_,
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('hb)
	) name17 (
		_w50_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		x_pad,
		y_pad,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		q_pad,
		z_pad,
		_w56_
	);
	LUT3 #(
		.INIT('h70)
	) name20 (
		_w46_,
		_w55_,
		_w56_,
		_w57_
	);
	LUT4 #(
		.INIT('h0002)
	) name21 (
		q_pad,
		x_pad,
		y_pad,
		z_pad,
		_w58_
	);
	LUT3 #(
		.INIT('h0e)
	) name22 (
		k_pad,
		q_pad,
		s_pad,
		_w59_
	);
	LUT3 #(
		.INIT('h70)
	) name23 (
		_w46_,
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('hb)
	) name24 (
		_w57_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h01)
	) name25 (
		x_pad,
		y_pad,
		z_pad,
		_w62_
	);
	LUT4 #(
		.INIT('h00ac)
	) name26 (
		\a0_pad ,
		j_pad,
		q_pad,
		s_pad,
		_w63_
	);
	LUT4 #(
		.INIT('h005c)
	) name27 (
		\a0_pad ,
		j_pad,
		q_pad,
		s_pad,
		_w64_
	);
	LUT4 #(
		.INIT('h087f)
	) name28 (
		_w46_,
		_w62_,
		_w63_,
		_w64_,
		_w65_
	);
	LUT4 #(
		.INIT('h0001)
	) name29 (
		\a0_pad ,
		x_pad,
		y_pad,
		z_pad,
		_w66_
	);
	LUT4 #(
		.INIT('h00ac)
	) name30 (
		\b0_pad ,
		i_pad,
		q_pad,
		s_pad,
		_w67_
	);
	LUT4 #(
		.INIT('h005c)
	) name31 (
		\b0_pad ,
		i_pad,
		q_pad,
		s_pad,
		_w68_
	);
	LUT4 #(
		.INIT('h087f)
	) name32 (
		_w46_,
		_w66_,
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\a0_pad ,
		\b0_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\c0_pad ,
		q_pad,
		_w71_
	);
	LUT4 #(
		.INIT('h7f00)
	) name35 (
		_w46_,
		_w62_,
		_w70_,
		_w71_,
		_w72_
	);
	LUT4 #(
		.INIT('h0100)
	) name36 (
		\a0_pad ,
		\b0_pad ,
		\c0_pad ,
		q_pad,
		_w73_
	);
	LUT3 #(
		.INIT('h0e)
	) name37 (
		h_pad,
		q_pad,
		s_pad,
		_w74_
	);
	LUT4 #(
		.INIT('h7f00)
	) name38 (
		_w46_,
		_w62_,
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('hb)
	) name39 (
		_w72_,
		_w75_,
		_w76_
	);
	LUT3 #(
		.INIT('h01)
	) name40 (
		\a0_pad ,
		\b0_pad ,
		\c0_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\d0_pad ,
		q_pad,
		_w78_
	);
	LUT4 #(
		.INIT('h7f00)
	) name42 (
		_w46_,
		_w62_,
		_w77_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\d0_pad ,
		q_pad,
		_w80_
	);
	LUT4 #(
		.INIT('h8000)
	) name44 (
		_w46_,
		_w62_,
		_w77_,
		_w80_,
		_w81_
	);
	LUT3 #(
		.INIT('h0e)
	) name45 (
		g_pad,
		q_pad,
		s_pad,
		_w82_
	);
	LUT3 #(
		.INIT('hef)
	) name46 (
		_w79_,
		_w81_,
		_w82_,
		_w83_
	);
	LUT4 #(
		.INIT('h0001)
	) name47 (
		\a0_pad ,
		\b0_pad ,
		\c0_pad ,
		\d0_pad ,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\e0_pad ,
		q_pad,
		_w85_
	);
	LUT4 #(
		.INIT('h7f00)
	) name49 (
		_w46_,
		_w62_,
		_w84_,
		_w85_,
		_w86_
	);
	LUT3 #(
		.INIT('h10)
	) name50 (
		\d0_pad ,
		\e0_pad ,
		q_pad,
		_w87_
	);
	LUT4 #(
		.INIT('h8000)
	) name51 (
		_w46_,
		_w62_,
		_w77_,
		_w87_,
		_w88_
	);
	LUT3 #(
		.INIT('h0e)
	) name52 (
		f_pad,
		q_pad,
		s_pad,
		_w89_
	);
	LUT3 #(
		.INIT('hef)
	) name53 (
		_w86_,
		_w88_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\d0_pad ,
		\e0_pad ,
		_w91_
	);
	LUT4 #(
		.INIT('h8000)
	) name55 (
		_w46_,
		_w62_,
		_w77_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\f0_pad ,
		q_pad,
		_w93_
	);
	LUT4 #(
		.INIT('h0100)
	) name57 (
		\d0_pad ,
		\e0_pad ,
		\f0_pad ,
		q_pad,
		_w94_
	);
	LUT4 #(
		.INIT('h8000)
	) name58 (
		_w46_,
		_w62_,
		_w77_,
		_w94_,
		_w95_
	);
	LUT3 #(
		.INIT('h0e)
	) name59 (
		e_pad,
		q_pad,
		s_pad,
		_w96_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name60 (
		_w92_,
		_w93_,
		_w95_,
		_w96_,
		_w97_
	);
	LUT3 #(
		.INIT('h01)
	) name61 (
		\d0_pad ,
		\e0_pad ,
		\f0_pad ,
		_w98_
	);
	LUT4 #(
		.INIT('h8000)
	) name62 (
		_w46_,
		_w62_,
		_w77_,
		_w98_,
		_w99_
	);
	LUT4 #(
		.INIT('h00ca)
	) name63 (
		d_pad,
		\g0_pad ,
		q_pad,
		s_pad,
		_w100_
	);
	LUT4 #(
		.INIT('h003a)
	) name64 (
		d_pad,
		\g0_pad ,
		q_pad,
		s_pad,
		_w101_
	);
	LUT3 #(
		.INIT('h27)
	) name65 (
		_w99_,
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\h0_pad ,
		q_pad,
		_w103_
	);
	LUT3 #(
		.INIT('hb0)
	) name67 (
		\g0_pad ,
		_w99_,
		_w103_,
		_w104_
	);
	LUT3 #(
		.INIT('h10)
	) name68 (
		\g0_pad ,
		\h0_pad ,
		q_pad,
		_w105_
	);
	LUT3 #(
		.INIT('h0e)
	) name69 (
		c_pad,
		q_pad,
		s_pad,
		_w106_
	);
	LUT3 #(
		.INIT('h70)
	) name70 (
		_w99_,
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('hb)
	) name71 (
		_w104_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\g0_pad ,
		\h0_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\i0_pad ,
		q_pad,
		_w110_
	);
	LUT3 #(
		.INIT('h70)
	) name74 (
		_w99_,
		_w109_,
		_w110_,
		_w111_
	);
	LUT4 #(
		.INIT('h0100)
	) name75 (
		\g0_pad ,
		\h0_pad ,
		\i0_pad ,
		q_pad,
		_w112_
	);
	LUT3 #(
		.INIT('h0e)
	) name76 (
		b_pad,
		q_pad,
		s_pad,
		_w113_
	);
	LUT3 #(
		.INIT('h70)
	) name77 (
		_w99_,
		_w112_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('hb)
	) name78 (
		_w111_,
		_w114_,
		_w115_
	);
	LUT3 #(
		.INIT('h01)
	) name79 (
		\g0_pad ,
		\h0_pad ,
		\i0_pad ,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\j0_pad ,
		q_pad,
		_w117_
	);
	LUT3 #(
		.INIT('h70)
	) name81 (
		_w99_,
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\j0_pad ,
		q_pad,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w116_,
		_w119_,
		_w120_
	);
	LUT3 #(
		.INIT('h0e)
	) name84 (
		a_pad,
		q_pad,
		s_pad,
		_w121_
	);
	LUT3 #(
		.INIT('h70)
	) name85 (
		_w99_,
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('hb)
	) name86 (
		_w118_,
		_w122_,
		_w123_
	);
	assign \k0_pad  = _w39_ ;
	assign \l0_pad  = _w42_ ;
	assign \m0_pad  = _w45_ ;
	assign \n0_pad  = _w48_ ;
	assign \o0_pad  = _w54_ ;
	assign \p0_pad  = _w61_ ;
	assign \q0_pad  = _w65_ ;
	assign \r0_pad  = _w69_ ;
	assign \s0_pad  = _w76_ ;
	assign \t0_pad  = _w83_ ;
	assign \u0_pad  = _w90_ ;
	assign \v0_pad  = _w97_ ;
	assign \w0_pad  = _w102_ ;
	assign \x0_pad  = _w108_ ;
	assign \y0_pad  = _w115_ ;
	assign \z0_pad  = _w123_ ;
endmodule;