module top (\cont1_reg[0]/NET0131 , \cont1_reg[1]/NET0131 , \cont1_reg[2]/NET0131 , \cont1_reg[3]/NET0131 , \cont1_reg[4]/NET0131 , \cont1_reg[5]/NET0131 , \cont1_reg[6]/NET0131 , \cont1_reg[7]/NET0131 , \cont1_reg[8]/NET0131 , \cont_reg[0]/NET0131 , \cont_reg[1]/NET0131 , \cont_reg[2]/NET0131 , \cont_reg[3]/NET0131 , \cont_reg[4]/NET0131 , \r_in_reg[0]/NET0131 , \r_in_reg[1]/NET0131 , \r_in_reg[2]/NET0131 , \r_in_reg[3]/NET0131 , \r_in_reg[4]/NET0131 , \r_in_reg[5]/NET0131 , \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , \stato_reg[2]/NET0131 , \stato_reg[3]/NET0131 , stbi_pad, \x_in[0]_pad , \x_in[1]_pad , \x_in[2]_pad , \x_in[3]_pad , \x_in[4]_pad , \x_in[5]_pad , \x_out[0]_pad , \x_out[1]_pad , \x_out[2]_pad , \x_out[3]_pad , \x_out[4]_pad , \x_out[5]_pad , \_al_n0 , \_al_n1 , \g2420/_0_ , \g2432/_0_ , \g2433/_0_ , \g2442/_0_ , \g2449/_0_ , \g2469/_0_ , \g2489/_0_ , \g2492/_0_ , \g2531/_0_ , \g2532/_0_ , \g2533/_0_ , \g2534/_0_ , \g2536/_0_ , \g2542/_0_ , \g2619/_0_ , \g2620/_0_ , \g2662/_0_ , \g2663/_0_ , \g2665/_0_ , \g2666/_0_ , \g2667/_0_ , \g2668/_0_ , \g2712/_0_ , \g3382/_0_ , \g34/_0_ , \g3435/_0_ , \g3443/_0_ , \g3735/_0_ , \g4020/_0_ , \g64/_0_ );
	input \cont1_reg[0]/NET0131  ;
	input \cont1_reg[1]/NET0131  ;
	input \cont1_reg[2]/NET0131  ;
	input \cont1_reg[3]/NET0131  ;
	input \cont1_reg[4]/NET0131  ;
	input \cont1_reg[5]/NET0131  ;
	input \cont1_reg[6]/NET0131  ;
	input \cont1_reg[7]/NET0131  ;
	input \cont1_reg[8]/NET0131  ;
	input \cont_reg[0]/NET0131  ;
	input \cont_reg[1]/NET0131  ;
	input \cont_reg[2]/NET0131  ;
	input \cont_reg[3]/NET0131  ;
	input \cont_reg[4]/NET0131  ;
	input \r_in_reg[0]/NET0131  ;
	input \r_in_reg[1]/NET0131  ;
	input \r_in_reg[2]/NET0131  ;
	input \r_in_reg[3]/NET0131  ;
	input \r_in_reg[4]/NET0131  ;
	input \r_in_reg[5]/NET0131  ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	input \stato_reg[2]/NET0131  ;
	input \stato_reg[3]/NET0131  ;
	input stbi_pad ;
	input \x_in[0]_pad  ;
	input \x_in[1]_pad  ;
	input \x_in[2]_pad  ;
	input \x_in[3]_pad  ;
	input \x_in[4]_pad  ;
	input \x_in[5]_pad  ;
	input \x_out[0]_pad  ;
	input \x_out[1]_pad  ;
	input \x_out[2]_pad  ;
	input \x_out[3]_pad  ;
	input \x_out[4]_pad  ;
	input \x_out[5]_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g2420/_0_  ;
	output \g2432/_0_  ;
	output \g2433/_0_  ;
	output \g2442/_0_  ;
	output \g2449/_0_  ;
	output \g2469/_0_  ;
	output \g2489/_0_  ;
	output \g2492/_0_  ;
	output \g2531/_0_  ;
	output \g2532/_0_  ;
	output \g2533/_0_  ;
	output \g2534/_0_  ;
	output \g2536/_0_  ;
	output \g2542/_0_  ;
	output \g2619/_0_  ;
	output \g2620/_0_  ;
	output \g2662/_0_  ;
	output \g2663/_0_  ;
	output \g2665/_0_  ;
	output \g2666/_0_  ;
	output \g2667/_0_  ;
	output \g2668/_0_  ;
	output \g2712/_0_  ;
	output \g3382/_0_  ;
	output \g34/_0_  ;
	output \g3435/_0_  ;
	output \g3443/_0_  ;
	output \g3735/_0_  ;
	output \g4020/_0_  ;
	output \g64/_0_  ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w39_
	);
	LUT4 #(
		.INIT('h135f)
	) name1 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w40_
	);
	LUT4 #(
		.INIT('hec80)
	) name2 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w42_
	);
	LUT4 #(
		.INIT('hfac8)
	) name4 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w43_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5 (
		_w39_,
		_w41_,
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w45_
	);
	LUT4 #(
		.INIT('h137f)
	) name7 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\cont1_reg[6]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w48_
	);
	LUT4 #(
		.INIT('hc080)
	) name10 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w49_
	);
	LUT3 #(
		.INIT('hb0)
	) name11 (
		_w44_,
		_w47_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w51_
	);
	LUT4 #(
		.INIT('hf531)
	) name13 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w52_
	);
	LUT4 #(
		.INIT('h8caf)
	) name14 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w53_
	);
	LUT3 #(
		.INIT('h45)
	) name15 (
		_w51_,
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w55_
	);
	LUT3 #(
		.INIT('h31)
	) name17 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w57_
	);
	LUT4 #(
		.INIT('hf531)
	) name19 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w56_,
		_w58_,
		_w59_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name21 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w60_
	);
	LUT4 #(
		.INIT('h7310)
	) name22 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w61_
	);
	LUT3 #(
		.INIT('h23)
	) name23 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w62_
	);
	LUT3 #(
		.INIT('h45)
	) name24 (
		_w60_,
		_w61_,
		_w62_,
		_w63_
	);
	LUT4 #(
		.INIT('h5540)
	) name25 (
		\cont1_reg[7]/NET0131 ,
		_w54_,
		_w59_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w50_,
		_w64_,
		_w65_
	);
	LUT4 #(
		.INIT('h0010)
	) name27 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w66_
	);
	LUT4 #(
		.INIT('h002a)
	) name28 (
		\cont1_reg[7]/NET0131 ,
		_w54_,
		_w59_,
		_w63_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\cont1_reg[7]/NET0131 ,
		_w49_,
		_w68_
	);
	LUT3 #(
		.INIT('hb0)
	) name30 (
		_w44_,
		_w47_,
		_w68_,
		_w69_
	);
	LUT3 #(
		.INIT('h02)
	) name31 (
		_w66_,
		_w67_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		_w71_
	);
	LUT3 #(
		.INIT('h01)
	) name33 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		_w74_
	);
	LUT4 #(
		.INIT('h8000)
	) name36 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		_w75_
	);
	LUT3 #(
		.INIT('h45)
	) name37 (
		\cont1_reg[7]/NET0131 ,
		_w72_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w77_
	);
	LUT3 #(
		.INIT('h80)
	) name39 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name40 (
		_w72_,
		_w73_,
		_w77_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w76_,
		_w79_,
		_w80_
	);
	LUT3 #(
		.INIT('h01)
	) name42 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w81_
	);
	LUT3 #(
		.INIT('h51)
	) name43 (
		\cont1_reg[7]/NET0131 ,
		_w74_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w83_
	);
	LUT3 #(
		.INIT('hd0)
	) name45 (
		_w78_,
		_w81_,
		_w83_,
		_w84_
	);
	LUT4 #(
		.INIT('he000)
	) name46 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w73_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		_w88_
	);
	LUT3 #(
		.INIT('h01)
	) name50 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		_w89_
	);
	LUT4 #(
		.INIT('h1000)
	) name51 (
		_w73_,
		_w85_,
		_w87_,
		_w89_,
		_w90_
	);
	LUT3 #(
		.INIT('h0b)
	) name52 (
		_w82_,
		_w84_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w93_
	);
	LUT4 #(
		.INIT('he000)
	) name55 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w95_
	);
	LUT3 #(
		.INIT('h08)
	) name57 (
		\cont1_reg[7]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w96_
	);
	LUT4 #(
		.INIT('hfe00)
	) name58 (
		\cont1_reg[6]/NET0131 ,
		_w92_,
		_w94_,
		_w96_,
		_w97_
	);
	LUT3 #(
		.INIT('h04)
	) name59 (
		\cont1_reg[7]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w98_
	);
	LUT4 #(
		.INIT('h0100)
	) name60 (
		\cont1_reg[6]/NET0131 ,
		_w92_,
		_w94_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		_w100_
	);
	LUT3 #(
		.INIT('h02)
	) name62 (
		\cont1_reg[7]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w101_
	);
	LUT4 #(
		.INIT('hef00)
	) name63 (
		_w73_,
		_w85_,
		_w100_,
		_w101_,
		_w102_
	);
	LUT3 #(
		.INIT('h01)
	) name64 (
		_w97_,
		_w99_,
		_w102_,
		_w103_
	);
	LUT4 #(
		.INIT('h0080)
	) name65 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w104_
	);
	LUT4 #(
		.INIT('hbf00)
	) name66 (
		_w80_,
		_w91_,
		_w103_,
		_w104_,
		_w105_
	);
	LUT4 #(
		.INIT('h0020)
	) name67 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w106_
	);
	LUT4 #(
		.INIT('h00fe)
	) name68 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w107_
	);
	LUT4 #(
		.INIT('he000)
	) name69 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w108_
	);
	LUT3 #(
		.INIT('h0e)
	) name70 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w109_
	);
	LUT3 #(
		.INIT('h15)
	) name71 (
		_w107_,
		_w108_,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('h01)
	) name72 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		_w108_,
		_w111_
	);
	LUT3 #(
		.INIT('h8a)
	) name73 (
		_w106_,
		_w110_,
		_w111_,
		_w112_
	);
	LUT4 #(
		.INIT('h0004)
	) name74 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w113_
	);
	LUT4 #(
		.INIT('h0001)
	) name75 (
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w115_
	);
	LUT4 #(
		.INIT('h8000)
	) name77 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w116_
	);
	LUT4 #(
		.INIT('h0777)
	) name78 (
		_w87_,
		_w114_,
		_w115_,
		_w116_,
		_w117_
	);
	LUT4 #(
		.INIT('h0103)
	) name79 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\cont1_reg[7]/NET0131 ,
		_w118_,
		_w119_
	);
	LUT3 #(
		.INIT('h70)
	) name81 (
		_w113_,
		_w117_,
		_w119_,
		_w120_
	);
	LUT4 #(
		.INIT('h0010)
	) name82 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		_w106_,
		_w108_,
		_w121_
	);
	LUT3 #(
		.INIT('h45)
	) name83 (
		\cont1_reg[7]/NET0131 ,
		_w110_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w124_
	);
	LUT4 #(
		.INIT('h0007)
	) name86 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w126_
	);
	LUT4 #(
		.INIT('h00a8)
	) name88 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w127_
	);
	LUT4 #(
		.INIT('h3133)
	) name89 (
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		_w125_,
		_w126_,
		_w128_
	);
	LUT3 #(
		.INIT('h0e)
	) name90 (
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w129_
	);
	LUT4 #(
		.INIT('h0040)
	) name91 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w130_
	);
	LUT4 #(
		.INIT('hdf00)
	) name92 (
		_w78_,
		_w125_,
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w128_,
		_w131_,
		_w132_
	);
	LUT4 #(
		.INIT('h00f4)
	) name94 (
		_w112_,
		_w120_,
		_w122_,
		_w132_,
		_w133_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name95 (
		_w65_,
		_w70_,
		_w105_,
		_w133_,
		_w134_
	);
	LUT4 #(
		.INIT('h0222)
	) name96 (
		_w106_,
		_w107_,
		_w108_,
		_w109_,
		_w135_
	);
	LUT3 #(
		.INIT('h45)
	) name97 (
		_w118_,
		_w129_,
		_w130_,
		_w136_
	);
	LUT3 #(
		.INIT('h8d)
	) name98 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w137_
	);
	LUT3 #(
		.INIT('h2a)
	) name99 (
		\cont1_reg[1]/NET0131 ,
		_w66_,
		_w137_,
		_w138_
	);
	LUT3 #(
		.INIT('h40)
	) name100 (
		_w135_,
		_w136_,
		_w138_,
		_w139_
	);
	LUT4 #(
		.INIT('ha888)
	) name101 (
		_w106_,
		_w107_,
		_w108_,
		_w109_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w66_,
		_w137_,
		_w141_
	);
	LUT3 #(
		.INIT('h15)
	) name103 (
		\cont1_reg[1]/NET0131 ,
		_w129_,
		_w130_,
		_w142_
	);
	LUT3 #(
		.INIT('h10)
	) name104 (
		_w140_,
		_w141_,
		_w142_,
		_w143_
	);
	LUT3 #(
		.INIT('h80)
	) name105 (
		_w113_,
		_w115_,
		_w116_,
		_w144_
	);
	LUT4 #(
		.INIT('h20a0)
	) name106 (
		\cont1_reg[1]/NET0131 ,
		_w87_,
		_w113_,
		_w114_,
		_w145_
	);
	LUT4 #(
		.INIT('h0008)
	) name107 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w146_
	);
	LUT3 #(
		.INIT('hac)
	) name108 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w146_,
		_w147_,
		_w148_
	);
	LUT3 #(
		.INIT('he2)
	) name110 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w149_
	);
	LUT3 #(
		.INIT('h84)
	) name111 (
		\cont1_reg[1]/NET0131 ,
		_w104_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h0001)
	) name112 (
		_w144_,
		_w145_,
		_w148_,
		_w150_,
		_w151_
	);
	LUT3 #(
		.INIT('h1f)
	) name113 (
		_w139_,
		_w143_,
		_w151_,
		_w152_
	);
	LUT4 #(
		.INIT('haf9f)
	) name114 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w71_,
		_w153_
	);
	LUT2 #(
		.INIT('h6)
	) name115 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w154_
	);
	LUT4 #(
		.INIT('h009f)
	) name116 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w155_
	);
	LUT4 #(
		.INIT('hff1e)
	) name117 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w156_
	);
	LUT3 #(
		.INIT('h80)
	) name118 (
		_w104_,
		_w155_,
		_w156_,
		_w157_
	);
	LUT3 #(
		.INIT('h0d)
	) name119 (
		_w104_,
		_w153_,
		_w157_,
		_w158_
	);
	LUT4 #(
		.INIT('h00ea)
	) name120 (
		_w107_,
		_w108_,
		_w109_,
		_w154_,
		_w159_
	);
	LUT4 #(
		.INIT('h88a8)
	) name121 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w89_,
		_w108_,
		_w160_
	);
	LUT3 #(
		.INIT('ha8)
	) name122 (
		_w106_,
		_w159_,
		_w160_,
		_w161_
	);
	LUT3 #(
		.INIT('h4c)
	) name123 (
		_w87_,
		_w113_,
		_w114_,
		_w162_
	);
	LUT3 #(
		.INIT('h15)
	) name124 (
		\cont1_reg[2]/NET0131 ,
		_w115_,
		_w116_,
		_w163_
	);
	LUT3 #(
		.INIT('hac)
	) name125 (
		\cont_reg[1]/NET0131 ,
		\cont_reg[2]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w146_,
		_w164_,
		_w165_
	);
	LUT3 #(
		.INIT('h80)
	) name127 (
		_w129_,
		_w130_,
		_w154_,
		_w166_
	);
	LUT4 #(
		.INIT('h000d)
	) name128 (
		_w162_,
		_w163_,
		_w165_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('hecce)
	) name129 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w168_
	);
	LUT2 #(
		.INIT('h6)
	) name130 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w169_
	);
	LUT3 #(
		.INIT('hd7)
	) name131 (
		_w66_,
		_w168_,
		_w169_,
		_w170_
	);
	LUT4 #(
		.INIT('h8a88)
	) name132 (
		\cont1_reg[2]/NET0131 ,
		_w118_,
		_w129_,
		_w130_,
		_w171_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT4 #(
		.INIT('hdfff)
	) name134 (
		_w158_,
		_w161_,
		_w167_,
		_w172_,
		_w173_
	);
	LUT3 #(
		.INIT('h07)
	) name135 (
		\r_in_reg[3]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w174_
	);
	LUT4 #(
		.INIT('h0007)
	) name136 (
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w175_
	);
	LUT3 #(
		.INIT('ha8)
	) name137 (
		_w113_,
		_w174_,
		_w175_,
		_w176_
	);
	LUT3 #(
		.INIT('h04)
	) name138 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\r_in_reg[1]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w178_
	);
	LUT4 #(
		.INIT('h0002)
	) name140 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w179_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name141 (
		stbi_pad,
		_w177_,
		_w178_,
		_w179_,
		_w180_
	);
	LUT4 #(
		.INIT('hecff)
	) name142 (
		_w117_,
		_w135_,
		_w176_,
		_w180_,
		_w181_
	);
	LUT3 #(
		.INIT('h01)
	) name143 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w182_
	);
	LUT4 #(
		.INIT('hfede)
	) name144 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w183_
	);
	LUT3 #(
		.INIT('hb0)
	) name145 (
		_w129_,
		_w130_,
		_w183_,
		_w184_
	);
	LUT4 #(
		.INIT('h135f)
	) name146 (
		\r_in_reg[1]/NET0131 ,
		stbi_pad,
		_w66_,
		_w179_,
		_w185_
	);
	LUT4 #(
		.INIT('h8fff)
	) name147 (
		_w113_,
		_w117_,
		_w184_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\stato_reg[3]/NET0131 ,
		\x_out[3]_pad ,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w182_,
		_w187_,
		_w188_
	);
	LUT4 #(
		.INIT('h0001)
	) name150 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w189_
	);
	LUT4 #(
		.INIT('h6f3f)
	) name151 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w71_,
		_w190_
	);
	LUT4 #(
		.INIT('h0100)
	) name152 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w192_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT3 #(
		.INIT('hea)
	) name155 (
		_w188_,
		_w190_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\stato_reg[3]/NET0131 ,
		\x_out[4]_pad ,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		_w182_,
		_w195_,
		_w196_
	);
	LUT4 #(
		.INIT('ha600)
	) name158 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w189_,
		_w191_,
		_w197_
	);
	LUT2 #(
		.INIT('he)
	) name159 (
		_w196_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\stato_reg[3]/NET0131 ,
		\x_out[5]_pad ,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w182_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w201_
	);
	LUT3 #(
		.INIT('h01)
	) name163 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w202_
	);
	LUT3 #(
		.INIT('h13)
	) name164 (
		_w72_,
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w204_
	);
	LUT4 #(
		.INIT('h80f0)
	) name166 (
		_w72_,
		_w123_,
		_w191_,
		_w204_,
		_w205_
	);
	LUT3 #(
		.INIT('hea)
	) name167 (
		_w200_,
		_w203_,
		_w205_,
		_w206_
	);
	LUT4 #(
		.INIT('hfe05)
	) name168 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w207_
	);
	LUT2 #(
		.INIT('h2)
	) name169 (
		\cont_reg[1]/NET0131 ,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\cont_reg[1]/NET0131 ,
		_w113_,
		_w209_
	);
	LUT3 #(
		.INIT('h01)
	) name171 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		\cont_reg[2]/NET0131 ,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\cont_reg[3]/NET0131 ,
		\cont_reg[4]/NET0131 ,
		_w211_
	);
	LUT2 #(
		.INIT('h6)
	) name173 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		_w212_
	);
	LUT4 #(
		.INIT('h8a00)
	) name174 (
		_w113_,
		_w210_,
		_w211_,
		_w212_,
		_w213_
	);
	LUT4 #(
		.INIT('hfdec)
	) name175 (
		_w117_,
		_w208_,
		_w209_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\cont_reg[2]/NET0131 ,
		_w207_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\cont_reg[2]/NET0131 ,
		_w113_,
		_w216_
	);
	LUT3 #(
		.INIT('h13)
	) name178 (
		_w117_,
		_w215_,
		_w216_,
		_w217_
	);
	LUT3 #(
		.INIT('h8a)
	) name179 (
		_w113_,
		_w210_,
		_w211_,
		_w218_
	);
	LUT3 #(
		.INIT('h80)
	) name180 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		\cont_reg[2]/NET0131 ,
		_w219_
	);
	LUT3 #(
		.INIT('h78)
	) name181 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		\cont_reg[2]/NET0131 ,
		_w220_
	);
	LUT3 #(
		.INIT('h40)
	) name182 (
		_w117_,
		_w218_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('hd)
	) name183 (
		_w217_,
		_w221_,
		_w222_
	);
	LUT3 #(
		.INIT('h70)
	) name184 (
		_w113_,
		_w117_,
		_w207_,
		_w223_
	);
	LUT4 #(
		.INIT('h8000)
	) name185 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		\cont_reg[2]/NET0131 ,
		\cont_reg[3]/NET0131 ,
		_w224_
	);
	LUT4 #(
		.INIT('h008a)
	) name186 (
		_w113_,
		_w210_,
		_w211_,
		_w224_,
		_w225_
	);
	LUT4 #(
		.INIT('h4070)
	) name187 (
		_w113_,
		_w117_,
		_w207_,
		_w225_,
		_w226_
	);
	LUT3 #(
		.INIT('h40)
	) name188 (
		_w117_,
		_w219_,
		_w225_,
		_w227_
	);
	LUT3 #(
		.INIT('hf2)
	) name189 (
		\cont_reg[3]/NET0131 ,
		_w226_,
		_w227_,
		_w228_
	);
	LUT3 #(
		.INIT('h40)
	) name190 (
		\cont_reg[4]/NET0131 ,
		_w113_,
		_w224_,
		_w229_
	);
	LUT3 #(
		.INIT('h45)
	) name191 (
		\cont_reg[4]/NET0131 ,
		_w117_,
		_w229_,
		_w230_
	);
	LUT3 #(
		.INIT('hab)
	) name192 (
		_w117_,
		_w225_,
		_w229_,
		_w231_
	);
	LUT3 #(
		.INIT('h13)
	) name193 (
		_w223_,
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		\stato_reg[3]/NET0131 ,
		\x_out[2]_pad ,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w182_,
		_w233_,
		_w234_
	);
	LUT4 #(
		.INIT('h1eff)
	) name196 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w236_
	);
	LUT3 #(
		.INIT('h08)
	) name198 (
		_w191_,
		_w235_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('he)
	) name199 (
		_w234_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		\cont_reg[0]/NET0131 ,
		_w207_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\cont_reg[0]/NET0131 ,
		_w113_,
		_w240_
	);
	LUT4 #(
		.INIT('h4044)
	) name202 (
		\cont_reg[0]/NET0131 ,
		_w113_,
		_w210_,
		_w211_,
		_w241_
	);
	LUT4 #(
		.INIT('hfdec)
	) name203 (
		_w117_,
		_w239_,
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		\stato_reg[3]/NET0131 ,
		\x_out[0]_pad ,
		_w243_
	);
	LUT4 #(
		.INIT('hb3a0)
	) name205 (
		\cont1_reg[0]/NET0131 ,
		_w182_,
		_w191_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		\stato_reg[3]/NET0131 ,
		\x_out[1]_pad ,
		_w245_
	);
	LUT3 #(
		.INIT('h6c)
	) name207 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w246_
	);
	LUT4 #(
		.INIT('hdc50)
	) name208 (
		_w182_,
		_w191_,
		_w245_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h0100)
	) name209 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		\x_in[3]_pad ,
		_w248_
	);
	LUT4 #(
		.INIT('hfe03)
	) name210 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w249_
	);
	LUT3 #(
		.INIT('hce)
	) name211 (
		\r_in_reg[3]/NET0131 ,
		_w248_,
		_w249_,
		_w250_
	);
	LUT4 #(
		.INIT('h0100)
	) name212 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		\x_in[5]_pad ,
		_w251_
	);
	LUT3 #(
		.INIT('hf2)
	) name213 (
		\r_in_reg[5]/NET0131 ,
		_w249_,
		_w251_,
		_w252_
	);
	LUT4 #(
		.INIT('h0100)
	) name214 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		\x_in[0]_pad ,
		_w253_
	);
	LUT3 #(
		.INIT('hf2)
	) name215 (
		\r_in_reg[0]/NET0131 ,
		_w249_,
		_w253_,
		_w254_
	);
	LUT4 #(
		.INIT('h0100)
	) name216 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		\x_in[1]_pad ,
		_w255_
	);
	LUT3 #(
		.INIT('hf2)
	) name217 (
		\r_in_reg[1]/NET0131 ,
		_w249_,
		_w255_,
		_w256_
	);
	LUT4 #(
		.INIT('h0100)
	) name218 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		\x_in[2]_pad ,
		_w257_
	);
	LUT3 #(
		.INIT('hf2)
	) name219 (
		\r_in_reg[2]/NET0131 ,
		_w249_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('h0100)
	) name220 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		\x_in[4]_pad ,
		_w259_
	);
	LUT3 #(
		.INIT('hf2)
	) name221 (
		\r_in_reg[4]/NET0131 ,
		_w249_,
		_w259_,
		_w260_
	);
	LUT3 #(
		.INIT('hae)
	) name222 (
		_w104_,
		_w113_,
		_w117_,
		_w261_
	);
	LUT4 #(
		.INIT('hfac8)
	) name223 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w262_
	);
	LUT3 #(
		.INIT('h84)
	) name224 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w263_
	);
	LUT4 #(
		.INIT('h2300)
	) name225 (
		_w40_,
		_w39_,
		_w262_,
		_w263_,
		_w264_
	);
	LUT3 #(
		.INIT('h21)
	) name226 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w265_
	);
	LUT4 #(
		.INIT('h4500)
	) name227 (
		_w51_,
		_w52_,
		_w53_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w264_,
		_w266_,
		_w267_
	);
	LUT3 #(
		.INIT('h48)
	) name229 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w268_
	);
	LUT4 #(
		.INIT('hdc00)
	) name230 (
		_w40_,
		_w39_,
		_w262_,
		_w268_,
		_w269_
	);
	LUT3 #(
		.INIT('h12)
	) name231 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w270_
	);
	LUT4 #(
		.INIT('hba00)
	) name232 (
		_w51_,
		_w52_,
		_w53_,
		_w270_,
		_w271_
	);
	LUT3 #(
		.INIT('h02)
	) name233 (
		_w66_,
		_w269_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w267_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\cont1_reg[3]/NET0131 ,
		_w118_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		\cont1_reg[3]/NET0131 ,
		_w113_,
		_w275_
	);
	LUT3 #(
		.INIT('h13)
	) name237 (
		_w117_,
		_w274_,
		_w275_,
		_w276_
	);
	LUT4 #(
		.INIT('h65ff)
	) name238 (
		\cont1_reg[3]/NET0131 ,
		_w124_,
		_w129_,
		_w130_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		\r_in_reg[3]/NET0131 ,
		_w113_,
		_w278_
	);
	LUT3 #(
		.INIT('hac)
	) name240 (
		\cont_reg[2]/NET0131 ,
		\cont_reg[3]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w146_,
		_w279_,
		_w280_
	);
	LUT4 #(
		.INIT('h008c)
	) name242 (
		_w117_,
		_w277_,
		_w278_,
		_w280_,
		_w281_
	);
	LUT3 #(
		.INIT('he0)
	) name243 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w282_
	);
	LUT3 #(
		.INIT('h1e)
	) name244 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w283_
	);
	LUT4 #(
		.INIT('h9000)
	) name245 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w284_
	);
	LUT3 #(
		.INIT('h07)
	) name246 (
		_w95_,
		_w283_,
		_w284_,
		_w285_
	);
	LUT4 #(
		.INIT('hfe00)
	) name247 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w286_
	);
	LUT3 #(
		.INIT('h02)
	) name248 (
		_w77_,
		_w189_,
		_w286_,
		_w287_
	);
	LUT3 #(
		.INIT('he0)
	) name249 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w288_
	);
	LUT4 #(
		.INIT('hc6ff)
	) name250 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w71_,
		_w87_,
		_w289_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name251 (
		_w104_,
		_w285_,
		_w287_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h00ea)
	) name252 (
		_w107_,
		_w108_,
		_w109_,
		_w283_,
		_w291_
	);
	LUT4 #(
		.INIT('h0111)
	) name253 (
		\cont1_reg[3]/NET0131 ,
		_w107_,
		_w108_,
		_w109_,
		_w292_
	);
	LUT3 #(
		.INIT('h02)
	) name254 (
		_w106_,
		_w291_,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('h0008)
	) name255 (
		_w276_,
		_w281_,
		_w290_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('hb)
	) name256 (
		_w273_,
		_w294_,
		_w295_
	);
	LUT3 #(
		.INIT('h70)
	) name257 (
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w296_
	);
	LUT4 #(
		.INIT('hfac8)
	) name258 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w297_
	);
	LUT4 #(
		.INIT('hec80)
	) name259 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w298_
	);
	LUT4 #(
		.INIT('h137f)
	) name260 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w299_
	);
	LUT3 #(
		.INIT('h70)
	) name261 (
		_w297_,
		_w298_,
		_w299_,
		_w300_
	);
	LUT3 #(
		.INIT('h80)
	) name262 (
		_w41_,
		_w43_,
		_w297_,
		_w301_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name263 (
		\r_in_reg[1]/NET0131 ,
		_w41_,
		_w43_,
		_w297_,
		_w302_
	);
	LUT3 #(
		.INIT('h15)
	) name264 (
		_w296_,
		_w300_,
		_w302_,
		_w303_
	);
	LUT4 #(
		.INIT('hf531)
	) name265 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w304_
	);
	LUT4 #(
		.INIT('h8caf)
	) name266 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w305_
	);
	LUT4 #(
		.INIT('h0301)
	) name267 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w306_
	);
	LUT4 #(
		.INIT('hefaf)
	) name268 (
		_w55_,
		_w57_,
		_w88_,
		_w305_,
		_w307_
	);
	LUT4 #(
		.INIT('h08ce)
	) name269 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w308_
	);
	LUT4 #(
		.INIT('hf531)
	) name270 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name271 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT4 #(
		.INIT('h8cef)
	) name272 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w311_
	);
	LUT3 #(
		.INIT('hb0)
	) name273 (
		_w305_,
		_w306_,
		_w311_,
		_w312_
	);
	LUT4 #(
		.INIT('h1011)
	) name274 (
		\r_in_reg[1]/NET0131 ,
		_w307_,
		_w310_,
		_w312_,
		_w313_
	);
	LUT4 #(
		.INIT('h77b7)
	) name275 (
		\cont1_reg[8]/NET0131 ,
		_w66_,
		_w303_,
		_w313_,
		_w314_
	);
	LUT4 #(
		.INIT('ha200)
	) name276 (
		\cont1_reg[8]/NET0131 ,
		_w78_,
		_w81_,
		_w83_,
		_w315_
	);
	LUT3 #(
		.INIT('h20)
	) name277 (
		\cont1_reg[8]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w316_
	);
	LUT4 #(
		.INIT('hbf00)
	) name278 (
		_w72_,
		_w73_,
		_w78_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w315_,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('h4000)
	) name280 (
		_w72_,
		_w73_,
		_w77_,
		_w78_,
		_w319_
	);
	LUT3 #(
		.INIT('h20)
	) name281 (
		_w78_,
		_w81_,
		_w83_,
		_w320_
	);
	LUT3 #(
		.INIT('h54)
	) name282 (
		\cont1_reg[8]/NET0131 ,
		_w319_,
		_w320_,
		_w321_
	);
	LUT4 #(
		.INIT('h5551)
	) name283 (
		\cont1_reg[8]/NET0131 ,
		_w88_,
		_w92_,
		_w94_,
		_w322_
	);
	LUT3 #(
		.INIT('h10)
	) name284 (
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w323_
	);
	LUT4 #(
		.INIT('he0f0)
	) name285 (
		_w92_,
		_w94_,
		_w95_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w322_,
		_w324_,
		_w325_
	);
	LUT4 #(
		.INIT('h0100)
	) name287 (
		\cont1_reg[5]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w326_
	);
	LUT3 #(
		.INIT('h10)
	) name288 (
		_w73_,
		_w85_,
		_w326_,
		_w327_
	);
	LUT3 #(
		.INIT('h02)
	) name289 (
		\cont1_reg[8]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w328_
	);
	LUT3 #(
		.INIT('h32)
	) name290 (
		_w90_,
		_w327_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('h0002)
	) name291 (
		_w318_,
		_w321_,
		_w325_,
		_w329_,
		_w330_
	);
	LUT4 #(
		.INIT('hfedc)
	) name292 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w331_
	);
	LUT4 #(
		.INIT('h80aa)
	) name293 (
		\cont1_reg[8]/NET0131 ,
		_w113_,
		_w117_,
		_w331_,
		_w332_
	);
	LUT4 #(
		.INIT('hae00)
	) name294 (
		\cont1_reg[8]/NET0131 ,
		_w78_,
		_w125_,
		_w130_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w332_,
		_w333_,
		_w334_
	);
	LUT4 #(
		.INIT('h3bff)
	) name296 (
		_w104_,
		_w314_,
		_w330_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\r_in_reg[1]/NET0131 ,
		_w46_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w44_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		\r_in_reg[1]/NET0131 ,
		_w61_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		\r_in_reg[1]/NET0131 ,
		_w58_,
		_w339_
	);
	LUT3 #(
		.INIT('h13)
	) name301 (
		_w54_,
		_w338_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h9)
	) name302 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w341_
	);
	LUT4 #(
		.INIT('hdf75)
	) name303 (
		_w66_,
		_w337_,
		_w340_,
		_w341_,
		_w342_
	);
	LUT3 #(
		.INIT('h07)
	) name304 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w343_
	);
	LUT4 #(
		.INIT('h0001)
	) name305 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT3 #(
		.INIT('h80)
	) name307 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w346_
	);
	LUT3 #(
		.INIT('h8c)
	) name308 (
		_w72_,
		_w77_,
		_w346_,
		_w347_
	);
	LUT4 #(
		.INIT('hfe00)
	) name309 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w349_
	);
	LUT4 #(
		.INIT('h0001)
	) name311 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		_w350_
	);
	LUT3 #(
		.INIT('h02)
	) name312 (
		_w83_,
		_w348_,
		_w350_,
		_w351_
	);
	LUT3 #(
		.INIT('h07)
	) name313 (
		_w345_,
		_w347_,
		_w351_,
		_w352_
	);
	LUT4 #(
		.INIT('h56ff)
	) name314 (
		\cont1_reg[5]/NET0131 ,
		_w73_,
		_w85_,
		_w87_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w282_,
		_w349_,
		_w354_
	);
	LUT3 #(
		.INIT('h10)
	) name316 (
		_w92_,
		_w94_,
		_w95_,
		_w355_
	);
	LUT3 #(
		.INIT('h8a)
	) name317 (
		_w353_,
		_w354_,
		_w355_,
		_w356_
	);
	LUT3 #(
		.INIT('h2a)
	) name318 (
		_w104_,
		_w352_,
		_w356_,
		_w357_
	);
	LUT4 #(
		.INIT('h0404)
	) name319 (
		\cont1_reg[5]/NET0131 ,
		_w107_,
		_w108_,
		_w109_,
		_w358_
	);
	LUT4 #(
		.INIT('h5959)
	) name320 (
		\cont1_reg[5]/NET0131 ,
		_w107_,
		_w108_,
		_w109_,
		_w359_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		_w106_,
		_w359_,
		_w360_
	);
	LUT3 #(
		.INIT('h45)
	) name322 (
		\cont1_reg[5]/NET0131 ,
		_w125_,
		_w129_,
		_w361_
	);
	LUT3 #(
		.INIT('hb0)
	) name323 (
		_w125_,
		_w127_,
		_w130_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		_w361_,
		_w362_,
		_w363_
	);
	LUT4 #(
		.INIT('h20a0)
	) name325 (
		\cont1_reg[5]/NET0131 ,
		_w87_,
		_w113_,
		_w114_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\cont_reg[4]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w365_
	);
	LUT4 #(
		.INIT('h0777)
	) name327 (
		\cont1_reg[5]/NET0131 ,
		_w118_,
		_w146_,
		_w365_,
		_w366_
	);
	LUT3 #(
		.INIT('h10)
	) name328 (
		_w144_,
		_w364_,
		_w366_,
		_w367_
	);
	LUT3 #(
		.INIT('h10)
	) name329 (
		_w360_,
		_w363_,
		_w367_,
		_w368_
	);
	LUT3 #(
		.INIT('hdf)
	) name330 (
		_w342_,
		_w357_,
		_w368_,
		_w369_
	);
	LUT3 #(
		.INIT('ha2)
	) name331 (
		\r_in_reg[1]/NET0131 ,
		_w300_,
		_w301_,
		_w370_
	);
	LUT4 #(
		.INIT('hdf55)
	) name332 (
		_w304_,
		_w308_,
		_w309_,
		_w311_,
		_w371_
	);
	LUT4 #(
		.INIT('h7310)
	) name333 (
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		\r_in_reg[1]/NET0131 ,
		_w372_,
		_w373_
	);
	LUT3 #(
		.INIT('h15)
	) name335 (
		\cont1_reg[6]/NET0131 ,
		_w371_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w370_,
		_w374_,
		_w375_
	);
	LUT3 #(
		.INIT('h80)
	) name337 (
		\cont1_reg[6]/NET0131 ,
		_w371_,
		_w373_,
		_w376_
	);
	LUT3 #(
		.INIT('ha2)
	) name338 (
		_w48_,
		_w300_,
		_w301_,
		_w377_
	);
	LUT3 #(
		.INIT('h02)
	) name339 (
		_w66_,
		_w376_,
		_w377_,
		_w378_
	);
	LUT3 #(
		.INIT('h02)
	) name340 (
		\cont1_reg[6]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w379_
	);
	LUT4 #(
		.INIT('hfe00)
	) name341 (
		\cont1_reg[5]/NET0131 ,
		_w73_,
		_w85_,
		_w379_,
		_w380_
	);
	LUT3 #(
		.INIT('h01)
	) name342 (
		\cont1_reg[6]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w381_
	);
	LUT4 #(
		.INIT('h0100)
	) name343 (
		\cont1_reg[5]/NET0131 ,
		_w73_,
		_w85_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w380_,
		_w382_,
		_w383_
	);
	LUT3 #(
		.INIT('h45)
	) name345 (
		\cont1_reg[6]/NET0131 ,
		_w72_,
		_w346_,
		_w384_
	);
	LUT3 #(
		.INIT('hb0)
	) name346 (
		_w72_,
		_w75_,
		_w77_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name347 (
		_w384_,
		_w385_,
		_w386_
	);
	LUT4 #(
		.INIT('h56ff)
	) name348 (
		\cont1_reg[6]/NET0131 ,
		_w92_,
		_w94_,
		_w95_,
		_w387_
	);
	LUT4 #(
		.INIT('h0001)
	) name349 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		\cont1_reg[6]/NET0131 ,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w100_,
		_w388_,
		_w389_
	);
	LUT3 #(
		.INIT('hd0)
	) name351 (
		_w74_,
		_w81_,
		_w83_,
		_w390_
	);
	LUT3 #(
		.INIT('h2a)
	) name352 (
		_w387_,
		_w389_,
		_w390_,
		_w391_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name353 (
		_w104_,
		_w383_,
		_w386_,
		_w391_,
		_w392_
	);
	LUT3 #(
		.INIT('h04)
	) name354 (
		\cont1_reg[5]/NET0131 ,
		_w106_,
		_w108_,
		_w393_
	);
	LUT4 #(
		.INIT('h4555)
	) name355 (
		\cont1_reg[6]/NET0131 ,
		_w125_,
		_w127_,
		_w130_,
		_w394_
	);
	LUT3 #(
		.INIT('hb0)
	) name356 (
		_w110_,
		_w393_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		_w106_,
		_w358_,
		_w396_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\cont1_reg[6]/NET0131 ,
		_w118_,
		_w397_
	);
	LUT4 #(
		.INIT('h0700)
	) name359 (
		_w113_,
		_w117_,
		_w362_,
		_w397_,
		_w398_
	);
	LUT3 #(
		.INIT('h45)
	) name360 (
		_w395_,
		_w396_,
		_w398_,
		_w399_
	);
	LUT4 #(
		.INIT('hfff4)
	) name361 (
		_w375_,
		_w378_,
		_w392_,
		_w399_,
		_w400_
	);
	LUT4 #(
		.INIT('h20a0)
	) name362 (
		\cont1_reg[0]/NET0131 ,
		_w87_,
		_w113_,
		_w114_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w144_,
		_w401_,
		_w402_
	);
	LUT4 #(
		.INIT('hfe9c)
	) name364 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		\cont1_reg[0]/NET0131 ,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h6)
	) name366 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		_w66_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h6)
	) name368 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		\cont_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w408_
	);
	LUT4 #(
		.INIT('h31f5)
	) name370 (
		_w104_,
		_w146_,
		_w407_,
		_w408_,
		_w409_
	);
	LUT3 #(
		.INIT('h10)
	) name371 (
		_w404_,
		_w406_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h7)
	) name372 (
		_w402_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('h0078)
	) name373 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w412_
	);
	LUT4 #(
		.INIT('h557f)
	) name374 (
		\r_in_reg[1]/NET0131 ,
		_w41_,
		_w43_,
		_w298_,
		_w413_
	);
	LUT4 #(
		.INIT('h4500)
	) name375 (
		\r_in_reg[1]/NET0131 ,
		_w308_,
		_w309_,
		_w311_,
		_w414_
	);
	LUT2 #(
		.INIT('h9)
	) name376 (
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w415_
	);
	LUT4 #(
		.INIT('h5df7)
	) name377 (
		_w66_,
		_w413_,
		_w414_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w106_,
		_w282_,
		_w417_
	);
	LUT3 #(
		.INIT('h07)
	) name379 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w418_
	);
	LUT4 #(
		.INIT('h1555)
	) name380 (
		\cont1_reg[4]/NET0131 ,
		_w129_,
		_w130_,
		_w418_,
		_w419_
	);
	LUT3 #(
		.INIT('hb0)
	) name381 (
		_w110_,
		_w417_,
		_w419_,
		_w420_
	);
	LUT4 #(
		.INIT('hea00)
	) name382 (
		_w107_,
		_w108_,
		_w109_,
		_w282_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		_w106_,
		_w421_,
		_w422_
	);
	LUT3 #(
		.INIT('h4c)
	) name384 (
		_w129_,
		_w130_,
		_w418_,
		_w423_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		\cont1_reg[4]/NET0131 ,
		_w118_,
		_w424_
	);
	LUT3 #(
		.INIT('h10)
	) name386 (
		_w162_,
		_w423_,
		_w424_,
		_w425_
	);
	LUT3 #(
		.INIT('h45)
	) name387 (
		_w420_,
		_w422_,
		_w425_,
		_w426_
	);
	LUT3 #(
		.INIT('hac)
	) name388 (
		\cont_reg[3]/NET0131 ,
		\cont_reg[4]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w146_,
		_w427_,
		_w428_
	);
	LUT3 #(
		.INIT('h01)
	) name390 (
		_w104_,
		_w144_,
		_w428_,
		_w429_
	);
	LUT3 #(
		.INIT('ha2)
	) name391 (
		_w87_,
		_w123_,
		_w288_,
		_w430_
	);
	LUT3 #(
		.INIT('hb0)
	) name392 (
		_w72_,
		_w73_,
		_w77_,
		_w431_
	);
	LUT4 #(
		.INIT('h0001)
	) name393 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w123_,
		_w432_,
		_w433_
	);
	LUT4 #(
		.INIT('h0777)
	) name395 (
		_w86_,
		_w430_,
		_w431_,
		_w433_,
		_w434_
	);
	LUT4 #(
		.INIT('hc6ff)
	) name396 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w93_,
		_w95_,
		_w435_
	);
	LUT3 #(
		.INIT('h1e)
	) name397 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w436_
	);
	LUT2 #(
		.INIT('h2)
	) name398 (
		_w83_,
		_w436_,
		_w437_
	);
	LUT4 #(
		.INIT('h0010)
	) name399 (
		_w144_,
		_w428_,
		_w435_,
		_w437_,
		_w438_
	);
	LUT3 #(
		.INIT('h15)
	) name400 (
		_w429_,
		_w434_,
		_w438_,
		_w439_
	);
	LUT3 #(
		.INIT('hfd)
	) name401 (
		_w416_,
		_w426_,
		_w439_,
		_w440_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g2420/_0_  = _w134_ ;
	assign \g2432/_0_  = _w152_ ;
	assign \g2433/_0_  = _w173_ ;
	assign \g2442/_0_  = _w181_ ;
	assign \g2449/_0_  = _w186_ ;
	assign \g2469/_0_  = _w194_ ;
	assign \g2489/_0_  = _w198_ ;
	assign \g2492/_0_  = _w206_ ;
	assign \g2531/_0_  = _w214_ ;
	assign \g2532/_0_  = _w222_ ;
	assign \g2533/_0_  = _w228_ ;
	assign \g2534/_0_  = _w232_ ;
	assign \g2536/_0_  = _w238_ ;
	assign \g2542/_0_  = _w242_ ;
	assign \g2619/_0_  = _w244_ ;
	assign \g2620/_0_  = _w247_ ;
	assign \g2662/_0_  = _w250_ ;
	assign \g2663/_0_  = _w252_ ;
	assign \g2665/_0_  = _w254_ ;
	assign \g2666/_0_  = _w256_ ;
	assign \g2667/_0_  = _w258_ ;
	assign \g2668/_0_  = _w260_ ;
	assign \g2712/_0_  = _w261_ ;
	assign \g3382/_0_  = _w295_ ;
	assign \g34/_0_  = _w335_ ;
	assign \g3435/_0_  = _w369_ ;
	assign \g3443/_0_  = _w400_ ;
	assign \g3735/_0_  = _w411_ ;
	assign \g4020/_0_  = _w412_ ;
	assign \g64/_0_  = _w440_ ;
endmodule;