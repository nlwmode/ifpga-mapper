module top (CLR_pad, \v0_pad , \v10_reg/NET0131 , \v11_reg/NET0131 , \v12_reg/NET0131 , \v1_pad , \v2_pad , \v3_pad , \v4_pad , \v5_pad , \v6_pad , \v7_reg/NET0131 , \v8_reg/NET0131 , \v9_reg/NET0131 , \_al_n0 , \_al_n1 , \g1759/_1_ , \g1762/_1_ , \g1764/_1_ , \g1765/_0_ , \g1786/_2_ , \g1791/_3_ , \g1808/_3_ , \g1822/_2_ , \g1929/_3_ , \g2713/_1_ , \g2744/_0_ , \v13_D_11_pad , \v13_D_12_pad , \v13_D_13_pad , \v13_D_14_pad , \v13_D_16_pad , \v13_D_18_pad , \v13_D_19_pad , \v13_D_21_pad , \v13_D_22_pad , \v13_D_23_pad , \v13_D_24_pad , \v13_D_7_pad , \v13_D_8_pad , \v13_D_9_pad );
	input CLR_pad ;
	input \v0_pad  ;
	input \v10_reg/NET0131  ;
	input \v11_reg/NET0131  ;
	input \v12_reg/NET0131  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input \v5_pad  ;
	input \v6_pad  ;
	input \v7_reg/NET0131  ;
	input \v8_reg/NET0131  ;
	input \v9_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1759/_1_  ;
	output \g1762/_1_  ;
	output \g1764/_1_  ;
	output \g1765/_0_  ;
	output \g1786/_2_  ;
	output \g1791/_3_  ;
	output \g1808/_3_  ;
	output \g1822/_2_  ;
	output \g1929/_3_  ;
	output \g2713/_1_  ;
	output \g2744/_0_  ;
	output \v13_D_11_pad  ;
	output \v13_D_12_pad  ;
	output \v13_D_13_pad  ;
	output \v13_D_14_pad  ;
	output \v13_D_16_pad  ;
	output \v13_D_18_pad  ;
	output \v13_D_19_pad  ;
	output \v13_D_21_pad  ;
	output \v13_D_22_pad  ;
	output \v13_D_23_pad  ;
	output \v13_D_24_pad  ;
	output \v13_D_7_pad  ;
	output \v13_D_8_pad  ;
	output \v13_D_9_pad  ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		_w16_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\v4_pad ,
		\v5_pad ,
		_w18_
	);
	LUT4 #(
		.INIT('h0040)
	) name3 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w19_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w20_
	);
	LUT3 #(
		.INIT('h80)
	) name5 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w21_
	);
	LUT3 #(
		.INIT('h40)
	) name6 (
		\v1_pad ,
		\v3_pad ,
		\v6_pad ,
		_w22_
	);
	LUT4 #(
		.INIT('ha888)
	) name7 (
		_w16_,
		_w19_,
		_w21_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\v6_pad ,
		\v8_reg/NET0131 ,
		_w24_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w25_
	);
	LUT4 #(
		.INIT('h0010)
	) name10 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w26_
	);
	LUT3 #(
		.INIT('h08)
	) name11 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w27_
	);
	LUT4 #(
		.INIT('h0800)
	) name12 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w28_
	);
	LUT4 #(
		.INIT('h0002)
	) name13 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w29_
	);
	LUT4 #(
		.INIT('h0015)
	) name14 (
		_w28_,
		_w24_,
		_w26_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w33_
	);
	LUT4 #(
		.INIT('h8a00)
	) name18 (
		\v10_reg/NET0131 ,
		\v1_pad ,
		\v6_pad ,
		\v8_reg/NET0131 ,
		_w34_
	);
	LUT3 #(
		.INIT('h01)
	) name19 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w35_
	);
	LUT4 #(
		.INIT('h0001)
	) name20 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w36_
	);
	LUT4 #(
		.INIT('haa80)
	) name21 (
		_w31_,
		_w32_,
		_w34_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w38_
	);
	LUT4 #(
		.INIT('h0222)
	) name23 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		\v4_pad ,
		\v5_pad ,
		_w39_
	);
	LUT3 #(
		.INIT('hc8)
	) name24 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w40_
	);
	LUT4 #(
		.INIT('h5d00)
	) name25 (
		\v9_reg/NET0131 ,
		_w38_,
		_w39_,
		_w40_,
		_w41_
	);
	LUT4 #(
		.INIT('h0100)
	) name26 (
		_w23_,
		_w37_,
		_w41_,
		_w30_,
		_w42_
	);
	LUT4 #(
		.INIT('h0800)
	) name27 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\v7_reg/NET0131 ,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w45_
	);
	LUT3 #(
		.INIT('h08)
	) name30 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w46_
	);
	LUT4 #(
		.INIT('h0020)
	) name31 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w47_
	);
	LUT3 #(
		.INIT('h07)
	) name32 (
		_w45_,
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w50_
	);
	LUT4 #(
		.INIT('hadbd)
	) name35 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		_w49_,
		_w51_,
		_w52_
	);
	LUT3 #(
		.INIT('h10)
	) name37 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w54_
	);
	LUT4 #(
		.INIT('h0020)
	) name39 (
		\v1_pad ,
		\v2_pad ,
		\v6_pad ,
		\v8_reg/NET0131 ,
		_w55_
	);
	LUT3 #(
		.INIT('h80)
	) name40 (
		_w54_,
		_w53_,
		_w55_,
		_w56_
	);
	LUT4 #(
		.INIT('h0100)
	) name41 (
		_w44_,
		_w52_,
		_w56_,
		_w48_,
		_w57_
	);
	LUT4 #(
		.INIT('h02aa)
	) name42 (
		CLR_pad,
		\v7_reg/NET0131 ,
		_w42_,
		_w57_,
		_w58_
	);
	LUT3 #(
		.INIT('h02)
	) name43 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w59_
	);
	LUT4 #(
		.INIT('hfd00)
	) name44 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w60_
	);
	LUT3 #(
		.INIT('h60)
	) name45 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w61_
	);
	LUT3 #(
		.INIT('h02)
	) name46 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v6_pad ,
		_w62_
	);
	LUT4 #(
		.INIT('h0004)
	) name47 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v6_pad ,
		_w63_
	);
	LUT3 #(
		.INIT('h01)
	) name48 (
		_w61_,
		_w63_,
		_w60_,
		_w64_
	);
	LUT3 #(
		.INIT('h40)
	) name49 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w65_
	);
	LUT3 #(
		.INIT('hbc)
	) name50 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w66_
	);
	LUT4 #(
		.INIT('h00f7)
	) name51 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w67_
	);
	LUT4 #(
		.INIT('hf351)
	) name52 (
		\v2_pad ,
		_w65_,
		_w66_,
		_w67_,
		_w68_
	);
	LUT4 #(
		.INIT('h00ef)
	) name53 (
		\v10_reg/NET0131 ,
		\v1_pad ,
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w69_
	);
	LUT4 #(
		.INIT('h0010)
	) name54 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w70_
	);
	LUT3 #(
		.INIT('h0d)
	) name55 (
		_w20_,
		_w69_,
		_w70_,
		_w71_
	);
	LUT4 #(
		.INIT('hea00)
	) name56 (
		\v8_reg/NET0131 ,
		_w64_,
		_w68_,
		_w71_,
		_w72_
	);
	LUT3 #(
		.INIT('h08)
	) name57 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w76_
	);
	LUT3 #(
		.INIT('ha2)
	) name61 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('h0004)
	) name63 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w79_
	);
	LUT3 #(
		.INIT('h0d)
	) name64 (
		_w76_,
		_w77_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w75_,
		_w80_,
		_w81_
	);
	LUT3 #(
		.INIT('h40)
	) name66 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w82_
	);
	LUT4 #(
		.INIT('h4000)
	) name67 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\v2_pad ,
		\v7_reg/NET0131 ,
		_w84_
	);
	LUT3 #(
		.INIT('h02)
	) name69 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		_w85_
	);
	LUT3 #(
		.INIT('he0)
	) name70 (
		_w82_,
		_w83_,
		_w85_,
		_w86_
	);
	LUT4 #(
		.INIT('hef23)
	) name71 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		_w50_,
		_w87_,
		_w88_
	);
	LUT3 #(
		.INIT('h08)
	) name73 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w89_
	);
	LUT3 #(
		.INIT('ha8)
	) name74 (
		_w45_,
		_w73_,
		_w89_,
		_w90_
	);
	LUT3 #(
		.INIT('h01)
	) name75 (
		_w88_,
		_w90_,
		_w86_,
		_w91_
	);
	LUT4 #(
		.INIT('he400)
	) name76 (
		\v7_reg/NET0131 ,
		_w72_,
		_w81_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		CLR_pad,
		_w92_,
		_w93_
	);
	LUT4 #(
		.INIT('h0100)
	) name78 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w94_
	);
	LUT4 #(
		.INIT('h0800)
	) name79 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w95_
	);
	LUT3 #(
		.INIT('h54)
	) name80 (
		\v1_pad ,
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w97_
	);
	LUT4 #(
		.INIT('h1000)
	) name82 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v8_reg/NET0131 ,
		_w98_
	);
	LUT4 #(
		.INIT('h0100)
	) name83 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w99_
	);
	LUT3 #(
		.INIT('h23)
	) name84 (
		\v8_reg/NET0131 ,
		_w98_,
		_w99_,
		_w100_
	);
	LUT3 #(
		.INIT('h45)
	) name85 (
		\v10_reg/NET0131 ,
		_w96_,
		_w100_,
		_w101_
	);
	LUT4 #(
		.INIT('h0006)
	) name86 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w66_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w104_
	);
	LUT3 #(
		.INIT('h70)
	) name89 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w105_
	);
	LUT4 #(
		.INIT('h0777)
	) name90 (
		_w19_,
		_w54_,
		_w104_,
		_w105_,
		_w106_
	);
	LUT3 #(
		.INIT('h20)
	) name91 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w107_
	);
	LUT4 #(
		.INIT('h2000)
	) name92 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w108_
	);
	LUT3 #(
		.INIT('h20)
	) name93 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w109_
	);
	LUT3 #(
		.INIT('h13)
	) name94 (
		_w17_,
		_w108_,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('h40)
	) name95 (
		_w103_,
		_w106_,
		_w110_,
		_w111_
	);
	LUT3 #(
		.INIT('h40)
	) name96 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w112_
	);
	LUT3 #(
		.INIT('h07)
	) name97 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w113_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name98 (
		\v10_reg/NET0131 ,
		_w94_,
		_w112_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w115_
	);
	LUT4 #(
		.INIT('h0002)
	) name100 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w116_
	);
	LUT4 #(
		.INIT('h4000)
	) name101 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w117_
	);
	LUT3 #(
		.INIT('h54)
	) name102 (
		_w18_,
		_w116_,
		_w117_,
		_w118_
	);
	LUT3 #(
		.INIT('h0d)
	) name103 (
		\v2_pad ,
		_w114_,
		_w118_,
		_w119_
	);
	LUT4 #(
		.INIT('h4555)
	) name104 (
		\v7_reg/NET0131 ,
		_w101_,
		_w111_,
		_w119_,
		_w120_
	);
	LUT4 #(
		.INIT('he000)
	) name105 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w121_
	);
	LUT4 #(
		.INIT('h007f)
	) name106 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w122_
	);
	LUT3 #(
		.INIT('hc4)
	) name107 (
		\v12_reg/NET0131 ,
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w124_
	);
	LUT4 #(
		.INIT('h0001)
	) name109 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w62_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w128_
	);
	LUT3 #(
		.INIT('hc4)
	) name113 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w129_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name114 (
		_w70_,
		_w127_,
		_w128_,
		_w129_,
		_w130_
	);
	LUT3 #(
		.INIT('h10)
	) name115 (
		_w123_,
		_w126_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h8a)
	) name116 (
		CLR_pad,
		_w120_,
		_w131_,
		_w132_
	);
	LUT4 #(
		.INIT('h0400)
	) name117 (
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w133_
	);
	LUT4 #(
		.INIT('h4240)
	) name118 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w134_
	);
	LUT3 #(
		.INIT('h54)
	) name119 (
		\v10_reg/NET0131 ,
		_w133_,
		_w134_,
		_w135_
	);
	LUT3 #(
		.INIT('h02)
	) name120 (
		\v12_reg/NET0131 ,
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w136_
	);
	LUT4 #(
		.INIT('h7773)
	) name121 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\v11_reg/NET0131 ,
		_w137_,
		_w138_
	);
	LUT4 #(
		.INIT('hfa77)
	) name123 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		_w115_,
		_w139_,
		_w140_
	);
	LUT4 #(
		.INIT('h2220)
	) name125 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w141_
	);
	LUT3 #(
		.INIT('h51)
	) name126 (
		\v7_reg/NET0131 ,
		_w76_,
		_w141_,
		_w142_
	);
	LUT3 #(
		.INIT('h10)
	) name127 (
		_w140_,
		_w138_,
		_w142_,
		_w143_
	);
	LUT3 #(
		.INIT('h40)
	) name128 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w144_
	);
	LUT4 #(
		.INIT('h5450)
	) name129 (
		\v2_pad ,
		_w18_,
		_w47_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w146_
	);
	LUT3 #(
		.INIT('h01)
	) name131 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w146_,
		_w147_,
		_w148_
	);
	LUT3 #(
		.INIT('h20)
	) name133 (
		\v0_pad ,
		\v1_pad ,
		\v6_pad ,
		_w149_
	);
	LUT4 #(
		.INIT('h8000)
	) name134 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w150_
	);
	LUT4 #(
		.INIT('h6200)
	) name135 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w151_
	);
	LUT3 #(
		.INIT('h0b)
	) name136 (
		_w149_,
		_w150_,
		_w151_,
		_w152_
	);
	LUT3 #(
		.INIT('h10)
	) name137 (
		_w145_,
		_w148_,
		_w152_,
		_w153_
	);
	LUT3 #(
		.INIT('h32)
	) name138 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w154_
	);
	LUT3 #(
		.INIT('hc8)
	) name139 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w155_
	);
	LUT4 #(
		.INIT('h0527)
	) name140 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w154_,
		_w156_,
		_w157_
	);
	LUT3 #(
		.INIT('h08)
	) name142 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w158_
	);
	LUT3 #(
		.INIT('h2a)
	) name143 (
		\v7_reg/NET0131 ,
		_w21_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		_w157_,
		_w159_,
		_w160_
	);
	LUT4 #(
		.INIT('h5540)
	) name145 (
		_w135_,
		_w143_,
		_w153_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		CLR_pad,
		_w161_,
		_w162_
	);
	LUT3 #(
		.INIT('h08)
	) name147 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w163_
	);
	LUT3 #(
		.INIT('h32)
	) name148 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w164_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name149 (
		\v11_reg/NET0131 ,
		_w84_,
		_w163_,
		_w164_,
		_w165_
	);
	LUT3 #(
		.INIT('he8)
	) name150 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT3 #(
		.INIT('ha8)
	) name153 (
		\v8_reg/NET0131 ,
		_w165_,
		_w168_,
		_w169_
	);
	LUT4 #(
		.INIT('hdf00)
	) name154 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w171_
	);
	LUT3 #(
		.INIT('h53)
	) name156 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w172_
	);
	LUT3 #(
		.INIT('h02)
	) name157 (
		_w171_,
		_w170_,
		_w172_,
		_w173_
	);
	LUT4 #(
		.INIT('h0804)
	) name158 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w175_
	);
	LUT4 #(
		.INIT('h54fc)
	) name160 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w176_
	);
	LUT4 #(
		.INIT('h8088)
	) name161 (
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w177_
	);
	LUT3 #(
		.INIT('h45)
	) name162 (
		_w174_,
		_w176_,
		_w177_,
		_w178_
	);
	LUT3 #(
		.INIT('h45)
	) name163 (
		\v12_reg/NET0131 ,
		_w173_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('he)
	) name164 (
		_w169_,
		_w179_,
		_w180_
	);
	LUT3 #(
		.INIT('h80)
	) name165 (
		_w19_,
		_w54_,
		_w124_,
		_w181_
	);
	LUT4 #(
		.INIT('hf070)
	) name166 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w182_
	);
	LUT3 #(
		.INIT('h04)
	) name167 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w183_
	);
	LUT4 #(
		.INIT('haa08)
	) name168 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w182_,
		_w183_,
		_w184_
	);
	LUT4 #(
		.INIT('h33f8)
	) name169 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w185_
	);
	LUT4 #(
		.INIT('hc080)
	) name170 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w186_
	);
	LUT4 #(
		.INIT('h3302)
	) name171 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w185_,
		_w186_,
		_w187_
	);
	LUT4 #(
		.INIT('heeec)
	) name172 (
		\v2_pad ,
		_w181_,
		_w184_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\v4_pad ,
		\v5_pad ,
		_w189_
	);
	LUT4 #(
		.INIT('h00ba)
	) name174 (
		\v10_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w190_
	);
	LUT3 #(
		.INIT('h04)
	) name175 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w191_
	);
	LUT4 #(
		.INIT('h00ab)
	) name176 (
		\v12_reg/NET0131 ,
		_w155_,
		_w190_,
		_w191_,
		_w192_
	);
	LUT3 #(
		.INIT('h20)
	) name177 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w193_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		_w170_,
		_w193_,
		_w194_
	);
	LUT4 #(
		.INIT('h3323)
	) name179 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w195_
	);
	LUT3 #(
		.INIT('he0)
	) name180 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w196_
	);
	LUT4 #(
		.INIT('h10f0)
	) name181 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w197_
	);
	LUT3 #(
		.INIT('h04)
	) name182 (
		_w26_,
		_w197_,
		_w195_,
		_w198_
	);
	LUT4 #(
		.INIT('hff54)
	) name183 (
		\v7_reg/NET0131 ,
		_w192_,
		_w194_,
		_w198_,
		_w199_
	);
	LUT4 #(
		.INIT('h2000)
	) name184 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w201_
	);
	LUT4 #(
		.INIT('h0004)
	) name186 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v7_reg/NET0131 ,
		_w202_
	);
	LUT4 #(
		.INIT('hf400)
	) name187 (
		_w66_,
		_w74_,
		_w200_,
		_w202_,
		_w203_
	);
	LUT4 #(
		.INIT('h8000)
	) name188 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w204_
	);
	LUT3 #(
		.INIT('h40)
	) name189 (
		\v7_reg/NET0131 ,
		_w34_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w206_
	);
	LUT4 #(
		.INIT('h8088)
	) name191 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v1_pad ,
		\v6_pad ,
		_w207_
	);
	LUT3 #(
		.INIT('ha8)
	) name192 (
		\v3_pad ,
		_w206_,
		_w207_,
		_w208_
	);
	LUT4 #(
		.INIT('h0020)
	) name193 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w209_
	);
	LUT4 #(
		.INIT('hcd00)
	) name194 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT4 #(
		.INIT('h0004)
	) name196 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w212_
	);
	LUT4 #(
		.INIT('h0d00)
	) name197 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w213_
	);
	LUT4 #(
		.INIT('haa80)
	) name198 (
		\v11_reg/NET0131 ,
		_w65_,
		_w212_,
		_w213_,
		_w214_
	);
	LUT4 #(
		.INIT('h0200)
	) name199 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w215_
	);
	LUT3 #(
		.INIT('h54)
	) name200 (
		\v8_reg/NET0131 ,
		_w99_,
		_w215_,
		_w216_
	);
	LUT4 #(
		.INIT('h1011)
	) name201 (
		_w214_,
		_w216_,
		_w208_,
		_w211_,
		_w217_
	);
	LUT4 #(
		.INIT('h7faa)
	) name202 (
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		_w218_
	);
	LUT4 #(
		.INIT('h0080)
	) name203 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w219_
	);
	LUT4 #(
		.INIT('h5504)
	) name204 (
		\v2_pad ,
		_w53_,
		_w218_,
		_w219_,
		_w220_
	);
	LUT4 #(
		.INIT('hc080)
	) name205 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w221_
	);
	LUT3 #(
		.INIT('h10)
	) name206 (
		_w46_,
		_w196_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w220_,
		_w222_,
		_w223_
	);
	LUT4 #(
		.INIT('h02aa)
	) name208 (
		CLR_pad,
		\v7_reg/NET0131 ,
		_w217_,
		_w223_,
		_w224_
	);
	LUT4 #(
		.INIT('h8a88)
	) name209 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		\v9_reg/NET0131 ,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w149_,
		_w204_,
		_w227_
	);
	LUT4 #(
		.INIT('h7000)
	) name212 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w228_
	);
	LUT3 #(
		.INIT('h32)
	) name213 (
		\v10_reg/NET0131 ,
		_w99_,
		_w228_,
		_w229_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name214 (
		\v8_reg/NET0131 ,
		_w226_,
		_w227_,
		_w229_,
		_w230_
	);
	LUT4 #(
		.INIT('h8bbb)
	) name215 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w231_
	);
	LUT4 #(
		.INIT('haf8c)
	) name216 (
		\v10_reg/NET0131 ,
		\v3_pad ,
		_w19_,
		_w231_,
		_w232_
	);
	LUT3 #(
		.INIT('h0b)
	) name217 (
		\v11_reg/NET0131 ,
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w233_
	);
	LUT3 #(
		.INIT('h04)
	) name218 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		_w233_,
		_w234_,
		_w235_
	);
	LUT3 #(
		.INIT('h8a)
	) name220 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w236_
	);
	LUT4 #(
		.INIT('h3020)
	) name221 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w237_
	);
	LUT4 #(
		.INIT('h7077)
	) name222 (
		_w27_,
		_w25_,
		_w236_,
		_w237_,
		_w238_
	);
	LUT4 #(
		.INIT('h0e00)
	) name223 (
		\v11_reg/NET0131 ,
		_w232_,
		_w235_,
		_w238_,
		_w239_
	);
	LUT4 #(
		.INIT('h2000)
	) name224 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w240_
	);
	LUT4 #(
		.INIT('h006f)
	) name225 (
		\v10_reg/NET0131 ,
		_w25_,
		_w50_,
		_w240_,
		_w241_
	);
	LUT4 #(
		.INIT('hba00)
	) name226 (
		\v7_reg/NET0131 ,
		_w230_,
		_w239_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		CLR_pad,
		_w242_,
		_w243_
	);
	LUT3 #(
		.INIT('h40)
	) name228 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v6_pad ,
		_w244_
	);
	LUT4 #(
		.INIT('h8ddd)
	) name229 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v3_pad ,
		\v6_pad ,
		_w245_
	);
	LUT4 #(
		.INIT('hef45)
	) name230 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w172_,
		_w245_,
		_w246_
	);
	LUT4 #(
		.INIT('h80c0)
	) name231 (
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		\v8_reg/NET0131 ,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		\v12_reg/NET0131 ,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w79_,
		_w197_,
		_w249_
	);
	LUT4 #(
		.INIT('h45ff)
	) name234 (
		\v7_reg/NET0131 ,
		_w246_,
		_w248_,
		_w249_,
		_w250_
	);
	LUT3 #(
		.INIT('h40)
	) name235 (
		\v10_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w251_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name236 (
		\v12_reg/NET0131 ,
		_w32_,
		_w107_,
		_w251_,
		_w252_
	);
	LUT4 #(
		.INIT('h5051)
	) name237 (
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w43_,
		_w252_,
		_w253_
	);
	LUT4 #(
		.INIT('h0004)
	) name238 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w254_
	);
	LUT4 #(
		.INIT('hcf57)
	) name239 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w255_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name240 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w128_,
		_w255_,
		_w256_
	);
	LUT4 #(
		.INIT('hff54)
	) name241 (
		\v8_reg/NET0131 ,
		_w253_,
		_w254_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('h54fc)
	) name242 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w258_
	);
	LUT4 #(
		.INIT('h3031)
	) name243 (
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w21_,
		_w258_,
		_w259_
	);
	LUT3 #(
		.INIT('h20)
	) name244 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w260_
	);
	LUT4 #(
		.INIT('h2000)
	) name245 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w261_
	);
	LUT3 #(
		.INIT('ha8)
	) name246 (
		\v10_reg/NET0131 ,
		_w259_,
		_w261_,
		_w262_
	);
	LUT4 #(
		.INIT('hfdea)
	) name247 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w263_
	);
	LUT4 #(
		.INIT('h0a02)
	) name248 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w79_,
		_w263_,
		_w264_
	);
	LUT3 #(
		.INIT('hb0)
	) name249 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w265_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name250 (
		_w18_,
		_w74_,
		_w200_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		\v2_pad ,
		_w186_,
		_w267_
	);
	LUT4 #(
		.INIT('hfc04)
	) name252 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w268_
	);
	LUT3 #(
		.INIT('h06)
	) name253 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w269_
	);
	LUT3 #(
		.INIT('h45)
	) name254 (
		\v7_reg/NET0131 ,
		_w268_,
		_w269_,
		_w270_
	);
	LUT4 #(
		.INIT('hab00)
	) name255 (
		\v12_reg/NET0131 ,
		_w266_,
		_w267_,
		_w270_,
		_w271_
	);
	LUT3 #(
		.INIT('hab)
	) name256 (
		_w262_,
		_w264_,
		_w271_,
		_w272_
	);
	LUT4 #(
		.INIT('h004f)
	) name257 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		\v8_reg/NET0131 ,
		_w273_,
		_w274_
	);
	LUT3 #(
		.INIT('h15)
	) name259 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w276_
	);
	LUT4 #(
		.INIT('hddd0)
	) name261 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w277_
	);
	LUT3 #(
		.INIT('h40)
	) name262 (
		_w276_,
		_w275_,
		_w277_,
		_w278_
	);
	LUT4 #(
		.INIT('h3715)
	) name263 (
		\v8_reg/NET0131 ,
		_w128_,
		_w129_,
		_w196_,
		_w279_
	);
	LUT4 #(
		.INIT('h45ff)
	) name264 (
		\v7_reg/NET0131 ,
		_w274_,
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w281_
	);
	LUT4 #(
		.INIT('h135f)
	) name266 (
		_w53_,
		_w89_,
		_w244_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		_w33_,
		_w282_,
		_w283_
	);
	LUT3 #(
		.INIT('h40)
	) name268 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w284_
	);
	LUT3 #(
		.INIT('ha8)
	) name269 (
		\v11_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w285_
	);
	LUT3 #(
		.INIT('he0)
	) name270 (
		_w212_,
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w35_,
		_w251_,
		_w287_
	);
	LUT3 #(
		.INIT('ha8)
	) name272 (
		_w201_,
		_w286_,
		_w287_,
		_w288_
	);
	LUT3 #(
		.INIT('h80)
	) name273 (
		_w33_,
		_w89_,
		_w281_,
		_w289_
	);
	LUT3 #(
		.INIT('h20)
	) name274 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		_w290_
	);
	LUT4 #(
		.INIT('h135f)
	) name275 (
		_w78_,
		_w104_,
		_w136_,
		_w290_,
		_w291_
	);
	LUT3 #(
		.INIT('h04)
	) name276 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		\v7_reg/NET0131 ,
		_w292_
	);
	LUT3 #(
		.INIT('hba)
	) name277 (
		_w289_,
		_w291_,
		_w292_,
		_w293_
	);
	LUT3 #(
		.INIT('h80)
	) name278 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w294_
	);
	LUT3 #(
		.INIT('h01)
	) name279 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w295_
	);
	LUT4 #(
		.INIT('hf800)
	) name280 (
		_w18_,
		_w35_,
		_w294_,
		_w295_,
		_w296_
	);
	LUT3 #(
		.INIT('h80)
	) name281 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w59_,
		_w297_,
		_w298_
	);
	LUT4 #(
		.INIT('h0100)
	) name283 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w299_
	);
	LUT3 #(
		.INIT('h20)
	) name284 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w301_
	);
	LUT3 #(
		.INIT('he0)
	) name286 (
		_w299_,
		_w300_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('he)
	) name287 (
		_w298_,
		_w302_,
		_w303_
	);
	LUT4 #(
		.INIT('h1000)
	) name288 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v6_pad ,
		_w304_
	);
	LUT4 #(
		.INIT('h0080)
	) name289 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w305_
	);
	LUT4 #(
		.INIT('h8000)
	) name290 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w306_
	);
	LUT4 #(
		.INIT('h00ab)
	) name291 (
		\v9_reg/NET0131 ,
		_w304_,
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		_w124_,
		_w307_,
		_w308_
	);
	LUT4 #(
		.INIT('h9f9e)
	) name293 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v5_pad ,
		_w309_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		_w74_,
		_w309_,
		_w310_
	);
	LUT3 #(
		.INIT('h80)
	) name295 (
		_w97_,
		_w104_,
		_w290_,
		_w311_
	);
	LUT3 #(
		.INIT('h54)
	) name296 (
		\v7_reg/NET0131 ,
		_w310_,
		_w311_,
		_w312_
	);
	LUT3 #(
		.INIT('h90)
	) name297 (
		\v10_reg/NET0131 ,
		_w104_,
		_w128_,
		_w313_
	);
	LUT4 #(
		.INIT('hee5f)
	) name298 (
		\v12_reg/NET0131 ,
		\v5_pad ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w314_
	);
	LUT4 #(
		.INIT('h2300)
	) name299 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT4 #(
		.INIT('h1000)
	) name301 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w317_
	);
	LUT3 #(
		.INIT('h08)
	) name302 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v5_pad ,
		_w318_
	);
	LUT3 #(
		.INIT('h01)
	) name303 (
		\v0_pad ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w319_
	);
	LUT4 #(
		.INIT('hec00)
	) name304 (
		_w124_,
		_w317_,
		_w318_,
		_w319_,
		_w320_
	);
	LUT4 #(
		.INIT('h0057)
	) name305 (
		\v11_reg/NET0131 ,
		_w313_,
		_w316_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('hb)
	) name306 (
		_w312_,
		_w321_,
		_w322_
	);
	LUT3 #(
		.INIT('hc9)
	) name307 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w323_
	);
	LUT4 #(
		.INIT('hcf45)
	) name308 (
		_w50_,
		_w76_,
		_w260_,
		_w323_,
		_w324_
	);
	LUT4 #(
		.INIT('h0200)
	) name309 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w325_
	);
	LUT4 #(
		.INIT('h0042)
	) name310 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w326_
	);
	LUT3 #(
		.INIT('h54)
	) name311 (
		\v9_reg/NET0131 ,
		_w325_,
		_w326_,
		_w327_
	);
	LUT3 #(
		.INIT('h45)
	) name312 (
		\v12_reg/NET0131 ,
		\v4_pad ,
		\v5_pad ,
		_w328_
	);
	LUT3 #(
		.INIT('he0)
	) name313 (
		_w200_,
		_w212_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('h7772)
	) name314 (
		\v7_reg/NET0131 ,
		_w324_,
		_w327_,
		_w329_,
		_w330_
	);
	LUT3 #(
		.INIT('hc8)
	) name315 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w331_
	);
	LUT4 #(
		.INIT('h00fd)
	) name316 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w332_
	);
	LUT3 #(
		.INIT('h45)
	) name317 (
		\v8_reg/NET0131 ,
		_w331_,
		_w332_,
		_w333_
	);
	LUT3 #(
		.INIT('h02)
	) name318 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w334_
	);
	LUT4 #(
		.INIT('h3302)
	) name319 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w335_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w334_,
		_w335_,
		_w336_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name321 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w337_
	);
	LUT4 #(
		.INIT('h0054)
	) name322 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w338_
	);
	LUT4 #(
		.INIT('h020f)
	) name323 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w339_
	);
	LUT4 #(
		.INIT('h0e00)
	) name324 (
		_w189_,
		_w337_,
		_w338_,
		_w339_,
		_w340_
	);
	LUT3 #(
		.INIT('he0)
	) name325 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w341_
	);
	LUT4 #(
		.INIT('h2a00)
	) name326 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w342_
	);
	LUT4 #(
		.INIT('h2022)
	) name327 (
		\v7_reg/NET0131 ,
		_w79_,
		_w341_,
		_w342_,
		_w343_
	);
	LUT4 #(
		.INIT('h00ef)
	) name328 (
		_w333_,
		_w336_,
		_w340_,
		_w343_,
		_w344_
	);
	LUT4 #(
		.INIT('h5040)
	) name329 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w345_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		_w175_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('he)
	) name331 (
		_w344_,
		_w346_,
		_w347_
	);
	LUT4 #(
		.INIT('h1f77)
	) name332 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w348_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		\v9_reg/NET0131 ,
		_w348_,
		_w349_
	);
	LUT3 #(
		.INIT('h04)
	) name334 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w350_
	);
	LUT3 #(
		.INIT('h08)
	) name335 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w351_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w352_
	);
	LUT3 #(
		.INIT('he0)
	) name337 (
		_w350_,
		_w351_,
		_w352_,
		_w353_
	);
	LUT3 #(
		.INIT('h54)
	) name338 (
		\v12_reg/NET0131 ,
		_w349_,
		_w353_,
		_w354_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1759/_1_  = _w58_ ;
	assign \g1762/_1_  = _w93_ ;
	assign \g1764/_1_  = _w132_ ;
	assign \g1765/_0_  = _w162_ ;
	assign \g1786/_2_  = _w180_ ;
	assign \g1791/_3_  = _w188_ ;
	assign \g1808/_3_  = _w199_ ;
	assign \g1822/_2_  = _w203_ ;
	assign \g1929/_3_  = _w205_ ;
	assign \g2713/_1_  = _w224_ ;
	assign \g2744/_0_  = _w243_ ;
	assign \v13_D_11_pad  = _w250_ ;
	assign \v13_D_12_pad  = _w257_ ;
	assign \v13_D_13_pad  = _w272_ ;
	assign \v13_D_14_pad  = _w280_ ;
	assign \v13_D_16_pad  = _w283_ ;
	assign \v13_D_18_pad  = _w288_ ;
	assign \v13_D_19_pad  = _w293_ ;
	assign \v13_D_21_pad  = _w296_ ;
	assign \v13_D_22_pad  = _w303_ ;
	assign \v13_D_23_pad  = _w308_ ;
	assign \v13_D_24_pad  = _w322_ ;
	assign \v13_D_7_pad  = _w330_ ;
	assign \v13_D_8_pad  = _w347_ ;
	assign \v13_D_9_pad  = _w354_ ;
endmodule;