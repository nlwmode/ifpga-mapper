module top (\101(0)_pad , \104(1)_pad , \107(2)_pad , \110(3)_pad , \113(4)_pad , \116(5)_pad , \119(6)_pad , \122(7)_pad , \125(8)_pad , \128(9)_pad , \131(10)_pad , \134(11)_pad , \137(12)_pad , \140(13)_pad , \143(14)_pad , \146(15)_pad , \210(16)_pad , \214(17)_pad , \217(18)_pad , \221(19)_pad , \224(20)_pad , \227(21)_pad , \234(22)_pad , \237(23)_pad , \469(24)_pad , \472(25)_pad , \475(26)_pad , \478(27)_pad , \898(28)_pad , \900(29)_pad , \902(30)_pad , \952(31)_pad , \953(32)_pad , \12(862)_pad , \15(861)_pad , \18(860)_pad , \21(859)_pad , \24(858)_pad , \27(857)_pad , \3(865)_pad , \30(856)_pad , \33(855)_pad , \36(854)_pad , \39(853)_pad , \42(852)_pad , \45(851)_pad , \48(850)_pad , \51(899)_pad , \54(900)_pad , \57(912)_pad , \6(864)_pad , \60(901)_pad , \63(902)_pad , \66(903)_pad , \69(908)_pad , \72(909)_pad , \75(866)_pad , \9(863)_pad );
	input \101(0)_pad  ;
	input \104(1)_pad  ;
	input \107(2)_pad  ;
	input \110(3)_pad  ;
	input \113(4)_pad  ;
	input \116(5)_pad  ;
	input \119(6)_pad  ;
	input \122(7)_pad  ;
	input \125(8)_pad  ;
	input \128(9)_pad  ;
	input \131(10)_pad  ;
	input \134(11)_pad  ;
	input \137(12)_pad  ;
	input \140(13)_pad  ;
	input \143(14)_pad  ;
	input \146(15)_pad  ;
	input \210(16)_pad  ;
	input \214(17)_pad  ;
	input \217(18)_pad  ;
	input \221(19)_pad  ;
	input \224(20)_pad  ;
	input \227(21)_pad  ;
	input \234(22)_pad  ;
	input \237(23)_pad  ;
	input \469(24)_pad  ;
	input \472(25)_pad  ;
	input \475(26)_pad  ;
	input \478(27)_pad  ;
	input \898(28)_pad  ;
	input \900(29)_pad  ;
	input \902(30)_pad  ;
	input \952(31)_pad  ;
	input \953(32)_pad  ;
	output \12(862)_pad  ;
	output \15(861)_pad  ;
	output \18(860)_pad  ;
	output \21(859)_pad  ;
	output \24(858)_pad  ;
	output \27(857)_pad  ;
	output \3(865)_pad  ;
	output \30(856)_pad  ;
	output \33(855)_pad  ;
	output \36(854)_pad  ;
	output \39(853)_pad  ;
	output \42(852)_pad  ;
	output \45(851)_pad  ;
	output \48(850)_pad  ;
	output \51(899)_pad  ;
	output \54(900)_pad  ;
	output \57(912)_pad  ;
	output \6(864)_pad  ;
	output \60(901)_pad  ;
	output \63(902)_pad  ;
	output \66(903)_pad  ;
	output \69(908)_pad  ;
	output \72(909)_pad  ;
	output \75(866)_pad  ;
	output \9(863)_pad  ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\101(0)_pad ,
		\119(6)_pad ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\101(0)_pad ,
		\119(6)_pad ,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w34_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\113(4)_pad ,
		\116(5)_pad ,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\113(4)_pad ,
		\116(5)_pad ,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w37_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w36_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w36_,
		_w39_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\237(23)_pad ,
		\953(32)_pad ,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\210(16)_pad ,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\143(14)_pad ,
		\146(15)_pad ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\143(14)_pad ,
		\146(15)_pad ,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\128(9)_pad ,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\128(9)_pad ,
		_w47_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\131(10)_pad ,
		\134(11)_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\131(10)_pad ,
		\134(11)_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\137(12)_pad ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\137(12)_pad ,
		_w53_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w50_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w50_,
		_w56_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w57_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		_w44_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w44_,
		_w59_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w42_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w42_,
		_w62_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w63_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\902(30)_pad ,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\472(25)_pad ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\472(25)_pad ,
		_w66_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\110(3)_pad ,
		\137(12)_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\110(3)_pad ,
		\137(12)_pad ,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\234(22)_pad ,
		\953(32)_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\221(19)_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\125(8)_pad ,
		\140(13)_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\125(8)_pad ,
		\140(13)_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\146(15)_pad ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\146(15)_pad ,
		_w77_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		_w74_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w74_,
		_w80_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w81_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\119(6)_pad ,
		\128(9)_pad ,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\119(6)_pad ,
		\128(9)_pad ,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		_w83_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w83_,
		_w86_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w87_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w72_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w72_,
		_w89_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w90_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\902(30)_pad ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\234(22)_pad ,
		\902(30)_pad ,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\217(18)_pad ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		_w93_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w93_,
		_w95_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		_w69_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\131(10)_pad ,
		\143(14)_pad ,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\131(10)_pad ,
		\143(14)_pad ,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\122(7)_pad ,
		_w80_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\122(7)_pad ,
		_w80_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w102_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w102_,
		_w105_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\214(17)_pad ,
		_w43_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\104(1)_pad ,
		\113(4)_pad ,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\104(1)_pad ,
		\113(4)_pad ,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		_w109_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w109_,
		_w112_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w113_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w108_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w108_,
		_w115_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		\902(30)_pad ,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\475(26)_pad ,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		\475(26)_pad ,
		_w119_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\217(18)_pad ,
		_w73_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\134(11)_pad ,
		\143(14)_pad ,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\134(11)_pad ,
		\143(14)_pad ,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w124_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		_w123_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w123_,
		_w126_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w127_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\116(5)_pad ,
		\122(7)_pad ,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\116(5)_pad ,
		\122(7)_pad ,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\107(2)_pad ,
		\128(9)_pad ,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\107(2)_pad ,
		\128(9)_pad ,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w132_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w132_,
		_w135_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w136_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w129_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w129_,
		_w138_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w139_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\902(30)_pad ,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\478(27)_pad ,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\478(27)_pad ,
		_w142_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		_w122_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\234(22)_pad ,
		\237(23)_pad ,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\902(30)_pad ,
		\953(32)_pad ,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w147_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		\898(28)_pad ,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\952(31)_pad ,
		\953(32)_pad ,
		_w151_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w147_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w150_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		_w146_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\227(21)_pad ,
		\953(32)_pad ,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w59_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w59_,
		_w155_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\104(1)_pad ,
		\107(2)_pad ,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\104(1)_pad ,
		\107(2)_pad ,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		\110(3)_pad ,
		\140(13)_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\110(3)_pad ,
		\140(13)_pad ,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\101(0)_pad ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		\101(0)_pad ,
		_w164_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w165_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		_w161_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w161_,
		_w167_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w158_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w158_,
		_w170_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w171_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\902(30)_pad ,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\469(24)_pad ,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\469(24)_pad ,
		_w174_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w175_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\221(19)_pad ,
		_w94_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		\237(23)_pad ,
		\902(30)_pad ,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\210(16)_pad ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\110(3)_pad ,
		\122(7)_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		\110(3)_pad ,
		\122(7)_pad ,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		_w161_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w161_,
		_w184_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w42_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w42_,
		_w187_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name157 (
		\224(20)_pad ,
		\953(32)_pad ,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\125(8)_pad ,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		\125(8)_pad ,
		_w191_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w192_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		_w50_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w50_,
		_w194_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w190_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w190_,
		_w197_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w198_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		\902(30)_pad ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		_w181_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name169 (
		_w181_,
		_w201_,
		_w203_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w202_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		\214(17)_pad ,
		_w180_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w179_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w99_,
		_w154_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w207_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\110(3)_pad ,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		\110(3)_pad ,
		_w209_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w122_,
		_w145_,
		_w213_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		_w153_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w69_,
		_w98_,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w177_,
		_w178_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w206_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w215_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w214_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		\113(4)_pad ,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		\113(4)_pad ,
		_w219_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w220_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w122_,
		_w145_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w153_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w218_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		\116(5)_pad ,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		\116(5)_pad ,
		_w225_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w69_,
		_w98_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w154_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w217_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h2)
	) name198 (
		\119(6)_pad ,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		\119(6)_pad ,
		_w231_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w122_,
		_w145_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w69_,
		_w98_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		_w153_,
		_w235_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w217_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		\122(7)_pad ,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		\122(7)_pad ,
		_w239_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		\900(29)_pad ,
		_w149_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w152_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		_w213_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w99_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w217_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		\125(8)_pad ,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		\125(8)_pad ,
		_w247_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w248_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w207_,
		_w215_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w154_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		\101(0)_pad ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\101(0)_pad ,
		_w252_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		_w223_,
		_w244_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w207_,
		_w229_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		\128(9)_pad ,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		\128(9)_pad ,
		_w258_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w259_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		_w204_,
		_w205_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w179_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w215_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w245_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		\131(10)_pad ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		\131(10)_pad ,
		_w265_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w256_,
		_w264_,
		_w269_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\134(11)_pad ,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		\134(11)_pad ,
		_w269_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w270_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		_w146_,
		_w244_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w229_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w263_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\137(12)_pad ,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		\137(12)_pad ,
		_w275_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w276_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w246_,
		_w263_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\140(13)_pad ,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		\140(13)_pad ,
		_w279_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w280_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		_w235_,
		_w244_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w251_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\143(14)_pad ,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		\143(14)_pad ,
		_w284_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w285_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w245_,
		_w257_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		\146(15)_pad ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		\146(15)_pad ,
		_w288_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		\952(31)_pad ,
		\953(32)_pad ,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w247_,
		_w258_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w265_,
		_w269_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w275_,
		_w279_,
		_w295_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w284_,
		_w288_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		_w293_,
		_w294_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w207_,
		_w236_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w224_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w214_,
		_w300_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w209_,
		_w219_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w225_,
		_w231_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w239_,
		_w252_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w301_,
		_w302_,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w303_,
		_w304_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w307_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w299_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\902(30)_pad ,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\210(16)_pad ,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w200_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w200_,
		_w312_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w292_,
		_w313_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\469(24)_pad ,
		_w311_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w173_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		_w173_,
		_w317_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w292_,
		_w318_,
		_w320_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		_w319_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\472(25)_pad ,
		_w311_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w65_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		_w65_,
		_w322_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w292_,
		_w323_,
		_w325_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		\104(1)_pad ,
		_w302_,
		_w327_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		\104(1)_pad ,
		_w302_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\475(26)_pad ,
		_w311_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w118_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		_w118_,
		_w330_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w292_,
		_w331_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w332_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		\478(27)_pad ,
		_w311_,
		_w335_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w141_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		_w141_,
		_w335_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w292_,
		_w336_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w337_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\217(18)_pad ,
		_w311_,
		_w340_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w92_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		_w92_,
		_w340_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w292_,
		_w341_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		\898(28)_pad ,
		\953(32)_pad ,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		\953(32)_pad ,
		_w309_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		\224(20)_pad ,
		\953(32)_pad ,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w190_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w190_,
		_w348_,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w345_,
		_w349_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w350_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		\900(29)_pad ,
		\953(32)_pad ,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		\227(21)_pad ,
		\953(32)_pad ,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\953(32)_pad ,
		_w299_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		_w59_,
		_w77_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w59_,
		_w77_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w357_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w356_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w356_,
		_w359_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w353_,
		_w360_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w361_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w146_,
		_w262_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w216_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w236_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		_w177_,
		_w178_,
		_w367_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w216_,
		_w262_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w217_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name337 (
		_w146_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		_w146_,
		_w205_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w205_,
		_w213_,
		_w373_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		_w223_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w204_,
		_w216_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w372_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		_w374_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		_w236_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		_w371_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w236_,
		_w365_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		_w152_,
		_w229_,
		_w381_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		_w380_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w379_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		_w310_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\952(31)_pad ,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		\953(32)_pad ,
		_w366_,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w385_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\107(2)_pad ,
		_w301_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		\107(2)_pad ,
		_w301_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w388_,
		_w389_,
		_w390_
	);
	assign \12(862)_pad  = _w212_ ;
	assign \15(861)_pad  = _w222_ ;
	assign \18(860)_pad  = _w228_ ;
	assign \21(859)_pad  = _w234_ ;
	assign \24(858)_pad  = _w242_ ;
	assign \27(857)_pad  = _w250_ ;
	assign \3(865)_pad  = _w255_ ;
	assign \30(856)_pad  = _w261_ ;
	assign \33(855)_pad  = _w268_ ;
	assign \36(854)_pad  = _w272_ ;
	assign \39(853)_pad  = _w278_ ;
	assign \42(852)_pad  = _w282_ ;
	assign \45(851)_pad  = _w287_ ;
	assign \48(850)_pad  = _w291_ ;
	assign \51(899)_pad  = _w316_ ;
	assign \54(900)_pad  = _w321_ ;
	assign \57(912)_pad  = _w326_ ;
	assign \6(864)_pad  = _w329_ ;
	assign \60(901)_pad  = _w334_ ;
	assign \63(902)_pad  = _w339_ ;
	assign \66(903)_pad  = _w344_ ;
	assign \69(908)_pad  = _w352_ ;
	assign \72(909)_pad  = _w363_ ;
	assign \75(866)_pad  = _w387_ ;
	assign \9(863)_pad  = _w390_ ;
endmodule;