module top( \100(38)_pad  , \103(39)_pad  , \106(40)_pad  , \109(41)_pad  , \11(2)_pad  , \112(42)_pad  , \113(43)_pad  , \114(44)_pad  , \115(45)_pad  , \116(46)_pad  , \117(47)_pad  , \118(48)_pad  , \119(49)_pad  , \120(50)_pad  , \121(51)_pad  , \122(52)_pad  , \123(53)_pad  , \126(54)_pad  , \127(55)_pad  , \128(56)_pad  , \129(57)_pad  , \130(58)_pad  , \131(59)_pad  , \132(60)_pad  , \135(61)_pad  , \136(62)_pad  , \14(3)_pad  , \140(64)_pad  , \144(354)_pad  , \145(66)_pad  , \146(67)_pad  , \149(68)_pad  , \1497(156)_pad  , \152(69)_pad  , \155(70)_pad  , \158(71)_pad  , \161(72)_pad  , \164(73)_pad  , \167(74)_pad  , \1689(157)_pad  , \1690(158)_pad  , \1691(159)_pad  , \1694(160)_pad  , \17(4)_pad  , \170(75)_pad  , \173(76)_pad  , \176(77)_pad  , \179(78)_pad  , \182(79)_pad  , \185(80)_pad  , \188(81)_pad  , \191(82)_pad  , \194(83)_pad  , \197(84)_pad  , \20(5)_pad  , \200(85)_pad  , \203(86)_pad  , \206(87)_pad  , \209(88)_pad  , \210(89)_pad  , \217(90)_pad  , \2174(161)_pad  , \218(91)_pad  , \225(92)_pad  , \226(93)_pad  , \23(6)_pad  , \233(94)_pad  , \234(95)_pad  , \2358(162)_pad  , \24(7)_pad  , \241(96)_pad  , \242(97)_pad  , \245(98)_pad  , \248(99)_pad  , \25(8)_pad  , \251(100)_pad  , \254(101)_pad  , \257(102)_pad  , \26(9)_pad  , \264(103)_pad  , \265(104)_pad  , \27(10)_pad  , \272(105)_pad  , \273(106)_pad  , \280(107)_pad  , \281(108)_pad  , \2824(163)_pad  , \288(109)_pad  , \289(110)_pad  , \292(111)_pad  , \298(299)_pad  , \302(114)_pad  , \307(115)_pad  , \308(116)_pad  , \31(11)_pad  , \315(117)_pad  , \316(118)_pad  , \323(119)_pad  , \324(120)_pad  , \331(121)_pad  , \332(122)_pad  , \335(123)_pad  , \338(124)_pad  , \34(12)_pad  , \341(125)_pad  , \348(126)_pad  , \351(127)_pad  , \3546(165)_pad  , \3548(166)_pad  , \3550(167)_pad  , \3552(168)_pad  , \358(128)_pad  , \361(129)_pad  , \366(130)_pad  , \369(131)_pad  , \37(13)_pad  , \3717(169)_pad  , \372(132)_pad  , \3724(170)_pad  , \373(133)_pad  , \374(134)_pad  , \386(135)_pad  , \389(136)_pad  , \4(1)_pad  , \40(14)_pad  , \400(137)_pad  , \4087(171)_pad  , \4088(172)_pad  , \4089(173)_pad  , \4090(174)_pad  , \4091(175)_pad  , \4092(176)_pad  , \411(138)_pad  , \4115(177)_pad  , \422(139)_pad  , \43(15)_pad  , \435(140)_pad  , \446(141)_pad  , \457(142)_pad  , \46(16)_pad  , \468(143)_pad  , \479(144)_pad  , \49(17)_pad  , \490(145)_pad  , \503(146)_pad  , \514(147)_pad  , \52(18)_pad  , \523(148)_pad  , \53(19)_pad  , \534(149)_pad  , \54(20)_pad  , \545(150)_pad  , \552(152)_pad  , \556(153)_pad  , \559(154)_pad  , \562(155)_pad  , \61(21)_pad  , \64(22)_pad  , \67(23)_pad  , \70(24)_pad  , \73(25)_pad  , \76(26)_pad  , \79(27)_pad  , \80(28)_pad  , \81(29)_pad  , \82(30)_pad  , \83(31)_pad  , \86(32)_pad  , \87(33)_pad  , \88(34)_pad  , \889(734)_pad  , \892(408)_pad  , \91(35)_pad  , \926(624)_pad  , \94(36)_pad  , \97(37)_pad  , \973(202)_pad  , \993(850)_pad  , \1000(2168)_pad  , \1002(1920)_pad  , \1004(1977)_pad  , \588(1696)_pad  , \593(733)_pad  , \598(1623)_pad  , \599(269)_pad  , \600(259)_pad  , \601(220)_pad  , \604(223)_pad  , \606(407)_pad  , \611(275)_pad  , \612(263)_pad  , \615(1750)_pad  , \618(1925)_pad  , \621(1893)_pad  , \626(1752)_pad  , \632(1692)_pad  , \634(665)_pad  , \636(1280)_pad  , \639(1275)_pad  , \642(2222)_pad  , \645(2271)_pad  , \648(2295)_pad  , \651(2314)_pad  , \654(2315)_pad  , \656(621)_pad  , \658(2483)_pad  , \661(2178)_pad  , \664(2223)_pad  , \667(2224)_pad  , \670(2225)_pad  , \673(1276)_pad  , \676(2229)_pad  , \679(2272)_pad  , \682(2296)_pad  , \685(2316)_pad  , \688(2317)_pad  , \690(2484)_pad  , \693(2179)_pad  , \696(2226)_pad  , \699(2227)_pad  , \702(2228)_pad  , \704(1281)_pad  , \707(1277)_pad  , \712(2297)_pad  , \715(1278)_pad  , \722(2131)_pad  , \727(2298)_pad  , \732(2300)_pad  , \737(2279)_pad  , \742(2238)_pad  , \747(2187)_pad  , \752(2189)_pad  , \757(2190)_pad  , \762(2184)_pad  , \767(2479)_pad  , \772(2299)_pad  , \777(2278)_pad  , \782(2239)_pad  , \787(2186)_pad  , \792(2188)_pad  , \797(2191)_pad  , \802(2183)_pad  , \807(2480)_pad  , \809(655)_pad  , \810(356)_pad  , \813(2260)_pad  , \815(627)_pad  , \820(1283)_pad  , \822(1933)_pad  , \824(2274)_pad  , \826(2275)_pad  , \828(2233)_pad  , \830(2182)_pad  , \832(2133)_pad  , \834(2123)_pad  , \836(2128)_pad  , \838(2064)_pad  , \843(2455)_pad  , \845(845)_pad  , \847(465)_pad  , \848(330)_pad  , \849(219)_pad  , \850(217)_pad  , \851(218)_pad  , \854(2268)_pad  , \859(2132)_pad  , \861(2070)_pad  , \863(2276)_pad  , \865(2277)_pad  , \867(2237)_pad  , \869(2181)_pad  , \871(2127)_pad  , \873(2124)_pad  , \875(2125)_pad  , \877(2126)_pad  , \882(2456)_pad  , \998(2163)_pad  , \u2023_syn_3  , \u2095_syn_3  , \u2109_syn_3  , \u2318_syn_3  , \u3086_syn_3  );
  input \100(38)_pad  ;
  input \103(39)_pad  ;
  input \106(40)_pad  ;
  input \109(41)_pad  ;
  input \11(2)_pad  ;
  input \112(42)_pad  ;
  input \113(43)_pad  ;
  input \114(44)_pad  ;
  input \115(45)_pad  ;
  input \116(46)_pad  ;
  input \117(47)_pad  ;
  input \118(48)_pad  ;
  input \119(49)_pad  ;
  input \120(50)_pad  ;
  input \121(51)_pad  ;
  input \122(52)_pad  ;
  input \123(53)_pad  ;
  input \126(54)_pad  ;
  input \127(55)_pad  ;
  input \128(56)_pad  ;
  input \129(57)_pad  ;
  input \130(58)_pad  ;
  input \131(59)_pad  ;
  input \132(60)_pad  ;
  input \135(61)_pad  ;
  input \136(62)_pad  ;
  input \14(3)_pad  ;
  input \140(64)_pad  ;
  input \144(354)_pad  ;
  input \145(66)_pad  ;
  input \146(67)_pad  ;
  input \149(68)_pad  ;
  input \1497(156)_pad  ;
  input \152(69)_pad  ;
  input \155(70)_pad  ;
  input \158(71)_pad  ;
  input \161(72)_pad  ;
  input \164(73)_pad  ;
  input \167(74)_pad  ;
  input \1689(157)_pad  ;
  input \1690(158)_pad  ;
  input \1691(159)_pad  ;
  input \1694(160)_pad  ;
  input \17(4)_pad  ;
  input \170(75)_pad  ;
  input \173(76)_pad  ;
  input \176(77)_pad  ;
  input \179(78)_pad  ;
  input \182(79)_pad  ;
  input \185(80)_pad  ;
  input \188(81)_pad  ;
  input \191(82)_pad  ;
  input \194(83)_pad  ;
  input \197(84)_pad  ;
  input \20(5)_pad  ;
  input \200(85)_pad  ;
  input \203(86)_pad  ;
  input \206(87)_pad  ;
  input \209(88)_pad  ;
  input \210(89)_pad  ;
  input \217(90)_pad  ;
  input \2174(161)_pad  ;
  input \218(91)_pad  ;
  input \225(92)_pad  ;
  input \226(93)_pad  ;
  input \23(6)_pad  ;
  input \233(94)_pad  ;
  input \234(95)_pad  ;
  input \2358(162)_pad  ;
  input \24(7)_pad  ;
  input \241(96)_pad  ;
  input \242(97)_pad  ;
  input \245(98)_pad  ;
  input \248(99)_pad  ;
  input \25(8)_pad  ;
  input \251(100)_pad  ;
  input \254(101)_pad  ;
  input \257(102)_pad  ;
  input \26(9)_pad  ;
  input \264(103)_pad  ;
  input \265(104)_pad  ;
  input \27(10)_pad  ;
  input \272(105)_pad  ;
  input \273(106)_pad  ;
  input \280(107)_pad  ;
  input \281(108)_pad  ;
  input \2824(163)_pad  ;
  input \288(109)_pad  ;
  input \289(110)_pad  ;
  input \292(111)_pad  ;
  input \298(299)_pad  ;
  input \302(114)_pad  ;
  input \307(115)_pad  ;
  input \308(116)_pad  ;
  input \31(11)_pad  ;
  input \315(117)_pad  ;
  input \316(118)_pad  ;
  input \323(119)_pad  ;
  input \324(120)_pad  ;
  input \331(121)_pad  ;
  input \332(122)_pad  ;
  input \335(123)_pad  ;
  input \338(124)_pad  ;
  input \34(12)_pad  ;
  input \341(125)_pad  ;
  input \348(126)_pad  ;
  input \351(127)_pad  ;
  input \3546(165)_pad  ;
  input \3548(166)_pad  ;
  input \3550(167)_pad  ;
  input \3552(168)_pad  ;
  input \358(128)_pad  ;
  input \361(129)_pad  ;
  input \366(130)_pad  ;
  input \369(131)_pad  ;
  input \37(13)_pad  ;
  input \3717(169)_pad  ;
  input \372(132)_pad  ;
  input \3724(170)_pad  ;
  input \373(133)_pad  ;
  input \374(134)_pad  ;
  input \386(135)_pad  ;
  input \389(136)_pad  ;
  input \4(1)_pad  ;
  input \40(14)_pad  ;
  input \400(137)_pad  ;
  input \4087(171)_pad  ;
  input \4088(172)_pad  ;
  input \4089(173)_pad  ;
  input \4090(174)_pad  ;
  input \4091(175)_pad  ;
  input \4092(176)_pad  ;
  input \411(138)_pad  ;
  input \4115(177)_pad  ;
  input \422(139)_pad  ;
  input \43(15)_pad  ;
  input \435(140)_pad  ;
  input \446(141)_pad  ;
  input \457(142)_pad  ;
  input \46(16)_pad  ;
  input \468(143)_pad  ;
  input \479(144)_pad  ;
  input \49(17)_pad  ;
  input \490(145)_pad  ;
  input \503(146)_pad  ;
  input \514(147)_pad  ;
  input \52(18)_pad  ;
  input \523(148)_pad  ;
  input \53(19)_pad  ;
  input \534(149)_pad  ;
  input \54(20)_pad  ;
  input \545(150)_pad  ;
  input \552(152)_pad  ;
  input \556(153)_pad  ;
  input \559(154)_pad  ;
  input \562(155)_pad  ;
  input \61(21)_pad  ;
  input \64(22)_pad  ;
  input \67(23)_pad  ;
  input \70(24)_pad  ;
  input \73(25)_pad  ;
  input \76(26)_pad  ;
  input \79(27)_pad  ;
  input \80(28)_pad  ;
  input \81(29)_pad  ;
  input \82(30)_pad  ;
  input \83(31)_pad  ;
  input \86(32)_pad  ;
  input \87(33)_pad  ;
  input \88(34)_pad  ;
  input \889(734)_pad  ;
  input \892(408)_pad  ;
  input \91(35)_pad  ;
  input \926(624)_pad  ;
  input \94(36)_pad  ;
  input \97(37)_pad  ;
  input \973(202)_pad  ;
  input \993(850)_pad  ;
  output \1000(2168)_pad  ;
  output \1002(1920)_pad  ;
  output \1004(1977)_pad  ;
  output \588(1696)_pad  ;
  output \593(733)_pad  ;
  output \598(1623)_pad  ;
  output \599(269)_pad  ;
  output \600(259)_pad  ;
  output \601(220)_pad  ;
  output \604(223)_pad  ;
  output \606(407)_pad  ;
  output \611(275)_pad  ;
  output \612(263)_pad  ;
  output \615(1750)_pad  ;
  output \618(1925)_pad  ;
  output \621(1893)_pad  ;
  output \626(1752)_pad  ;
  output \632(1692)_pad  ;
  output \634(665)_pad  ;
  output \636(1280)_pad  ;
  output \639(1275)_pad  ;
  output \642(2222)_pad  ;
  output \645(2271)_pad  ;
  output \648(2295)_pad  ;
  output \651(2314)_pad  ;
  output \654(2315)_pad  ;
  output \656(621)_pad  ;
  output \658(2483)_pad  ;
  output \661(2178)_pad  ;
  output \664(2223)_pad  ;
  output \667(2224)_pad  ;
  output \670(2225)_pad  ;
  output \673(1276)_pad  ;
  output \676(2229)_pad  ;
  output \679(2272)_pad  ;
  output \682(2296)_pad  ;
  output \685(2316)_pad  ;
  output \688(2317)_pad  ;
  output \690(2484)_pad  ;
  output \693(2179)_pad  ;
  output \696(2226)_pad  ;
  output \699(2227)_pad  ;
  output \702(2228)_pad  ;
  output \704(1281)_pad  ;
  output \707(1277)_pad  ;
  output \712(2297)_pad  ;
  output \715(1278)_pad  ;
  output \722(2131)_pad  ;
  output \727(2298)_pad  ;
  output \732(2300)_pad  ;
  output \737(2279)_pad  ;
  output \742(2238)_pad  ;
  output \747(2187)_pad  ;
  output \752(2189)_pad  ;
  output \757(2190)_pad  ;
  output \762(2184)_pad  ;
  output \767(2479)_pad  ;
  output \772(2299)_pad  ;
  output \777(2278)_pad  ;
  output \782(2239)_pad  ;
  output \787(2186)_pad  ;
  output \792(2188)_pad  ;
  output \797(2191)_pad  ;
  output \802(2183)_pad  ;
  output \807(2480)_pad  ;
  output \809(655)_pad  ;
  output \810(356)_pad  ;
  output \813(2260)_pad  ;
  output \815(627)_pad  ;
  output \820(1283)_pad  ;
  output \822(1933)_pad  ;
  output \824(2274)_pad  ;
  output \826(2275)_pad  ;
  output \828(2233)_pad  ;
  output \830(2182)_pad  ;
  output \832(2133)_pad  ;
  output \834(2123)_pad  ;
  output \836(2128)_pad  ;
  output \838(2064)_pad  ;
  output \843(2455)_pad  ;
  output \845(845)_pad  ;
  output \847(465)_pad  ;
  output \848(330)_pad  ;
  output \849(219)_pad  ;
  output \850(217)_pad  ;
  output \851(218)_pad  ;
  output \854(2268)_pad  ;
  output \859(2132)_pad  ;
  output \861(2070)_pad  ;
  output \863(2276)_pad  ;
  output \865(2277)_pad  ;
  output \867(2237)_pad  ;
  output \869(2181)_pad  ;
  output \871(2127)_pad  ;
  output \873(2124)_pad  ;
  output \875(2125)_pad  ;
  output \877(2126)_pad  ;
  output \882(2456)_pad  ;
  output \998(2163)_pad  ;
  output \u2023_syn_3  ;
  output \u2095_syn_3  ;
  output \u2109_syn_3  ;
  output \u2318_syn_3  ;
  output \u3086_syn_3  ;
  wire n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 ;
  assign n179 = \233(94)_pad  & \335(123)_pad  ;
  assign n180 = \226(93)_pad  & ~\335(123)_pad  ;
  assign n181 = ~n179 & ~n180 ;
  assign n182 = \264(103)_pad  & \335(123)_pad  ;
  assign n183 = \257(102)_pad  & ~\335(123)_pad  ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = \280(107)_pad  & \335(123)_pad  ;
  assign n186 = \273(106)_pad  & ~\335(123)_pad  ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = ~n184 & ~n187 ;
  assign n189 = n184 & n187 ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = n181 & ~n190 ;
  assign n192 = ~n181 & n190 ;
  assign n193 = ~n191 & ~n192 ;
  assign n194 = \241(96)_pad  & \335(123)_pad  ;
  assign n195 = \234(95)_pad  & ~\335(123)_pad  ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = \288(109)_pad  & \335(123)_pad  ;
  assign n198 = \281(108)_pad  & ~\335(123)_pad  ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = n196 & ~n199 ;
  assign n201 = ~n196 & n199 ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = \272(105)_pad  & \335(123)_pad  ;
  assign n204 = \265(104)_pad  & ~\335(123)_pad  ;
  assign n205 = ~n203 & ~n204 ;
  assign n206 = \217(90)_pad  & \335(123)_pad  ;
  assign n207 = \210(89)_pad  & ~\335(123)_pad  ;
  assign n208 = ~n206 & ~n207 ;
  assign n209 = ~n205 & ~n208 ;
  assign n210 = n205 & n208 ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = ~\292(111)_pad  & \335(123)_pad  ;
  assign n213 = ~\289(110)_pad  & ~\335(123)_pad  ;
  assign n214 = ~n212 & ~n213 ;
  assign n215 = n211 & ~n214 ;
  assign n216 = ~n211 & n214 ;
  assign n217 = ~n215 & ~n216 ;
  assign n218 = n202 & n217 ;
  assign n219 = ~n202 & ~n217 ;
  assign n220 = ~n218 & ~n219 ;
  assign n221 = \225(92)_pad  & \335(123)_pad  ;
  assign n222 = \218(91)_pad  & ~\335(123)_pad  ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = \209(88)_pad  & \335(123)_pad  ;
  assign n225 = \206(87)_pad  & ~\335(123)_pad  ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = n223 & ~n226 ;
  assign n228 = ~n223 & n226 ;
  assign n229 = ~n227 & ~n228 ;
  assign n230 = n220 & ~n229 ;
  assign n231 = ~n220 & n229 ;
  assign n232 = ~n230 & ~n231 ;
  assign n233 = n193 & n232 ;
  assign n234 = ~n193 & ~n232 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = \316(118)_pad  & ~\369(131)_pad  ;
  assign n237 = ~\316(118)_pad  & \369(131)_pad  ;
  assign n238 = ~n236 & ~n237 ;
  assign n239 = ~\324(120)_pad  & ~\341(125)_pad  ;
  assign n240 = \324(120)_pad  & \341(125)_pad  ;
  assign n241 = ~n239 & ~n240 ;
  assign n242 = n238 & ~n241 ;
  assign n243 = ~n238 & n241 ;
  assign n244 = ~n242 & ~n243 ;
  assign n245 = ~\308(116)_pad  & ~\361(129)_pad  ;
  assign n246 = \308(116)_pad  & \361(129)_pad  ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = \298(299)_pad  & n247 ;
  assign n249 = ~\298(299)_pad  & ~n247 ;
  assign n250 = ~n248 & ~n249 ;
  assign n251 = \302(114)_pad  & ~\351(127)_pad  ;
  assign n252 = ~\302(114)_pad  & \351(127)_pad  ;
  assign n253 = ~n251 & ~n252 ;
  assign n254 = n250 & ~n253 ;
  assign n255 = ~n250 & n253 ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = n244 & n256 ;
  assign n258 = ~n244 & ~n256 ;
  assign n259 = ~n257 & ~n258 ;
  assign n260 = \218(91)_pad  & ~\281(108)_pad  ;
  assign n261 = ~\218(91)_pad  & \281(108)_pad  ;
  assign n262 = ~n260 & ~n261 ;
  assign n263 = ~\206(87)_pad  & ~\289(110)_pad  ;
  assign n264 = \206(87)_pad  & \289(110)_pad  ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = n262 & ~n265 ;
  assign n267 = ~n262 & n265 ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = ~\257(102)_pad  & ~\265(104)_pad  ;
  assign n270 = \257(102)_pad  & \265(104)_pad  ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = \210(89)_pad  & ~\273(106)_pad  ;
  assign n273 = ~\210(89)_pad  & \273(106)_pad  ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = n271 & n274 ;
  assign n276 = ~n271 & ~n274 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = \226(93)_pad  & ~\234(95)_pad  ;
  assign n279 = ~\226(93)_pad  & \234(95)_pad  ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = n277 & ~n280 ;
  assign n282 = ~n277 & n280 ;
  assign n283 = ~n281 & ~n282 ;
  assign n284 = n268 & n283 ;
  assign n285 = ~n268 & ~n283 ;
  assign n286 = ~n284 & ~n285 ;
  assign n294 = \374(134)_pad  & ~n199 ;
  assign n295 = ~\374(134)_pad  & n199 ;
  assign n296 = ~n294 & ~n295 ;
  assign n297 = \411(138)_pad  & ~n187 ;
  assign n298 = ~\411(138)_pad  & n187 ;
  assign n299 = ~n297 & ~n298 ;
  assign n300 = \400(137)_pad  & ~n205 ;
  assign n301 = ~\400(137)_pad  & n205 ;
  assign n302 = ~n300 & ~n301 ;
  assign n303 = n299 & n302 ;
  assign n304 = n296 & n303 ;
  assign n305 = \435(140)_pad  & ~n196 ;
  assign n306 = ~\435(140)_pad  & n196 ;
  assign n307 = ~n305 & ~n306 ;
  assign n308 = \389(136)_pad  & ~n184 ;
  assign n309 = ~\389(136)_pad  & n184 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = n307 & n310 ;
  assign n312 = n304 & n311 ;
  assign n287 = \422(139)_pad  & ~n181 ;
  assign n288 = \468(143)_pad  & ~n223 ;
  assign n289 = ~\468(143)_pad  & n223 ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = ~\422(139)_pad  & n181 ;
  assign n292 = n290 & ~n291 ;
  assign n293 = ~n287 & n292 ;
  assign n313 = \446(141)_pad  & ~n226 ;
  assign n314 = ~\446(141)_pad  & n226 ;
  assign n315 = ~n313 & ~n314 ;
  assign n316 = \457(142)_pad  & ~n208 ;
  assign n317 = ~\457(142)_pad  & n208 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = n315 & n318 ;
  assign n320 = n293 & n319 ;
  assign n321 = n312 & n320 ;
  assign n323 = ~\248(99)_pad  & \316(118)_pad  ;
  assign n322 = ~\251(100)_pad  & ~\316(118)_pad  ;
  assign n324 = \490(145)_pad  & ~n322 ;
  assign n325 = ~n323 & n324 ;
  assign n327 = \242(97)_pad  & \316(118)_pad  ;
  assign n326 = \254(101)_pad  & ~\316(118)_pad  ;
  assign n328 = ~\490(145)_pad  & ~n326 ;
  assign n329 = ~n327 & n328 ;
  assign n330 = ~n325 & ~n329 ;
  assign n332 = ~\248(99)_pad  & \308(116)_pad  ;
  assign n331 = ~\251(100)_pad  & ~\308(116)_pad  ;
  assign n333 = \479(144)_pad  & ~n331 ;
  assign n334 = ~n332 & n333 ;
  assign n336 = \242(97)_pad  & \308(116)_pad  ;
  assign n335 = \254(101)_pad  & ~\308(116)_pad  ;
  assign n337 = ~\479(144)_pad  & ~n335 ;
  assign n338 = ~n336 & n337 ;
  assign n339 = ~n334 & ~n338 ;
  assign n340 = ~n330 & ~n339 ;
  assign n345 = \341(125)_pad  & \3552(168)_pad  ;
  assign n344 = ~\341(125)_pad  & \3550(167)_pad  ;
  assign n346 = \523(148)_pad  & ~n344 ;
  assign n347 = ~n345 & n346 ;
  assign n349 = \341(125)_pad  & ~\3546(165)_pad  ;
  assign n348 = ~\341(125)_pad  & ~\3548(166)_pad  ;
  assign n350 = ~\523(148)_pad  & ~n348 ;
  assign n351 = ~n349 & n350 ;
  assign n352 = ~n347 & ~n351 ;
  assign n371 = \254(101)_pad  & ~\298(299)_pad  ;
  assign n372 = \242(97)_pad  & \298(299)_pad  ;
  assign n373 = ~n371 & ~n372 ;
  assign n374 = \251(100)_pad  & ~\302(114)_pad  ;
  assign n375 = \248(99)_pad  & \302(114)_pad  ;
  assign n376 = ~n374 & ~n375 ;
  assign n377 = n373 & ~n376 ;
  assign n341 = \251(100)_pad  & ~\361(129)_pad  ;
  assign n342 = \248(99)_pad  & \361(129)_pad  ;
  assign n343 = ~n341 & ~n342 ;
  assign n378 = ~\3552(168)_pad  & \514(147)_pad  ;
  assign n379 = \3546(165)_pad  & ~\514(147)_pad  ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n343 & ~n380 ;
  assign n382 = n377 & n381 ;
  assign n383 = ~n352 & n382 ;
  assign n354 = \324(120)_pad  & \3552(168)_pad  ;
  assign n353 = ~\324(120)_pad  & \3550(167)_pad  ;
  assign n355 = \503(146)_pad  & ~n353 ;
  assign n356 = ~n354 & n355 ;
  assign n358 = \324(120)_pad  & ~\3546(165)_pad  ;
  assign n357 = ~\324(120)_pad  & ~\3548(166)_pad  ;
  assign n359 = ~\503(146)_pad  & ~n357 ;
  assign n360 = ~n358 & n359 ;
  assign n361 = ~n356 & ~n360 ;
  assign n363 = \351(127)_pad  & \3552(168)_pad  ;
  assign n362 = ~\351(127)_pad  & \3550(167)_pad  ;
  assign n364 = \534(149)_pad  & ~n362 ;
  assign n365 = ~n363 & n364 ;
  assign n367 = \351(127)_pad  & ~\3546(165)_pad  ;
  assign n366 = ~\351(127)_pad  & ~\3548(166)_pad  ;
  assign n368 = ~\534(149)_pad  & ~n366 ;
  assign n369 = ~n367 & n368 ;
  assign n370 = ~n365 & ~n369 ;
  assign n384 = ~n361 & ~n370 ;
  assign n385 = n383 & n384 ;
  assign n386 = n340 & n385 ;
  assign n387 = \552(152)_pad  & \562(155)_pad  ;
  assign n388 = \332(122)_pad  & ~\338(124)_pad  ;
  assign n389 = ~\514(147)_pad  & n388 ;
  assign n390 = \514(147)_pad  & ~n388 ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = \332(122)_pad  & \348(126)_pad  ;
  assign n393 = ~\332(122)_pad  & \341(125)_pad  ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = \523(148)_pad  & ~n394 ;
  assign n396 = ~\523(148)_pad  & n394 ;
  assign n397 = ~n395 & ~n396 ;
  assign n398 = \332(122)_pad  & \358(128)_pad  ;
  assign n399 = ~\332(122)_pad  & \351(127)_pad  ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = \534(149)_pad  & ~n400 ;
  assign n402 = ~\534(149)_pad  & n400 ;
  assign n403 = ~n401 & ~n402 ;
  assign n404 = n397 & n403 ;
  assign n405 = \332(122)_pad  & \366(130)_pad  ;
  assign n406 = ~\332(122)_pad  & \361(129)_pad  ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = n404 & n407 ;
  assign n409 = n391 & n408 ;
  assign n410 = ~\324(120)_pad  & ~\332(122)_pad  ;
  assign n411 = ~\331(121)_pad  & \332(122)_pad  ;
  assign n412 = ~n410 & ~n411 ;
  assign n413 = \503(146)_pad  & n412 ;
  assign n414 = ~\503(146)_pad  & ~n412 ;
  assign n415 = ~n413 & ~n414 ;
  assign n416 = n409 & n415 ;
  assign n417 = \332(122)_pad  & \889(734)_pad  ;
  assign n418 = \298(299)_pad  & ~\332(122)_pad  ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = \307(115)_pad  & \332(122)_pad  ;
  assign n421 = \302(114)_pad  & ~\332(122)_pad  ;
  assign n422 = ~n420 & ~n421 ;
  assign n423 = n419 & n422 ;
  assign n424 = \315(117)_pad  & \332(122)_pad  ;
  assign n425 = \308(116)_pad  & ~\332(122)_pad  ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = \479(144)_pad  & ~n426 ;
  assign n428 = ~\479(144)_pad  & n426 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = \323(119)_pad  & \332(122)_pad  ;
  assign n431 = \316(118)_pad  & ~\332(122)_pad  ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = \490(145)_pad  & ~n432 ;
  assign n434 = ~\490(145)_pad  & n432 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = n429 & n435 ;
  assign n437 = n423 & n436 ;
  assign n438 = n416 & n437 ;
  assign n441 = ~n402 & ~n407 ;
  assign n442 = ~n395 & ~n401 ;
  assign n443 = ~n441 & n442 ;
  assign n444 = ~n396 & ~n443 ;
  assign n445 = ~n390 & ~n444 ;
  assign n446 = ~n389 & ~n445 ;
  assign n447 = ~n413 & ~n446 ;
  assign n448 = ~n414 & ~n447 ;
  assign n449 = n437 & n448 ;
  assign n439 = n429 & n433 ;
  assign n440 = ~n427 & ~n439 ;
  assign n450 = n423 & n440 ;
  assign n451 = ~n449 & n450 ;
  assign n452 = n287 & n290 ;
  assign n453 = ~n288 & ~n452 ;
  assign n454 = ~n316 & n453 ;
  assign n455 = n294 & ~n298 ;
  assign n456 = ~n297 & ~n300 ;
  assign n457 = ~n455 & n456 ;
  assign n458 = ~n301 & ~n457 ;
  assign n459 = ~n309 & n458 ;
  assign n460 = ~n308 & ~n459 ;
  assign n461 = ~n305 & n460 ;
  assign n462 = ~n306 & ~n461 ;
  assign n463 = n293 & n462 ;
  assign n464 = n454 & ~n463 ;
  assign n465 = ~n314 & ~n317 ;
  assign n466 = ~n464 & n465 ;
  assign n467 = ~n313 & ~n466 ;
  assign n468 = \373(133)_pad  & \993(850)_pad  ;
  assign n471 = \2358(162)_pad  & ~\87(33)_pad  ;
  assign n469 = \27(10)_pad  & \31(11)_pad  ;
  assign n470 = ~\2358(162)_pad  & ~\86(32)_pad  ;
  assign n472 = n469 & ~n470 ;
  assign n473 = ~n471 & n472 ;
  assign n475 = \2358(162)_pad  & \25(8)_pad  ;
  assign n474 = ~\2358(162)_pad  & \24(7)_pad  ;
  assign n476 = n469 & ~n474 ;
  assign n477 = ~n475 & n476 ;
  assign n478 = \144(354)_pad  & ~n477 ;
  assign n508 = ~\1689(157)_pad  & ~\1690(158)_pad  ;
  assign n491 = \4091(175)_pad  & ~\4092(176)_pad  ;
  assign n510 = \54(20)_pad  & n408 ;
  assign n511 = n391 & n510 ;
  assign n512 = ~n446 & ~n511 ;
  assign n513 = n415 & ~n512 ;
  assign n514 = ~n415 & n512 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = n491 & n515 ;
  assign n480 = ~\4091(175)_pad  & ~\4092(176)_pad  ;
  assign n509 = n361 & n480 ;
  assign n499 = ~\4091(175)_pad  & \4092(176)_pad  ;
  assign n517 = \52(18)_pad  & n499 ;
  assign n518 = ~n509 & ~n517 ;
  assign n519 = ~n516 & n518 ;
  assign n520 = n508 & ~n519 ;
  assign n479 = \1689(157)_pad  & ~\1690(158)_pad  ;
  assign n492 = \4(1)_pad  & n304 ;
  assign n493 = n310 & n492 ;
  assign n494 = n460 & ~n493 ;
  assign n495 = n307 & n494 ;
  assign n496 = ~n307 & ~n494 ;
  assign n497 = ~n495 & ~n496 ;
  assign n498 = n491 & ~n497 ;
  assign n482 = \234(95)_pad  & \3552(168)_pad  ;
  assign n481 = ~\234(95)_pad  & \3550(167)_pad  ;
  assign n483 = \435(140)_pad  & ~n481 ;
  assign n484 = ~n482 & n483 ;
  assign n486 = \234(95)_pad  & ~\3546(165)_pad  ;
  assign n485 = ~\234(95)_pad  & ~\3548(166)_pad  ;
  assign n487 = ~\435(140)_pad  & ~n485 ;
  assign n488 = ~n486 & n487 ;
  assign n489 = ~n484 & ~n488 ;
  assign n490 = n480 & n489 ;
  assign n500 = \122(52)_pad  & n499 ;
  assign n501 = ~n490 & ~n500 ;
  assign n502 = ~n498 & n501 ;
  assign n503 = n479 & ~n502 ;
  assign n504 = \1689(157)_pad  & \1690(158)_pad  ;
  assign n505 = \170(75)_pad  & n504 ;
  assign n506 = ~\1689(157)_pad  & \1690(158)_pad  ;
  assign n507 = \200(85)_pad  & n506 ;
  assign n521 = ~n505 & ~n507 ;
  assign n522 = ~n503 & n521 ;
  assign n523 = ~n520 & n522 ;
  assign n524 = \926(624)_pad  & ~n523 ;
  assign n549 = ~n413 & ~n513 ;
  assign n550 = ~n435 & ~n549 ;
  assign n551 = n435 & n549 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = n491 & ~n552 ;
  assign n548 = n330 & n480 ;
  assign n554 = \112(42)_pad  & n499 ;
  assign n555 = ~n548 & ~n554 ;
  assign n556 = ~n553 & n555 ;
  assign n557 = n508 & ~n556 ;
  assign n535 = ~n287 & ~n291 ;
  assign n536 = n461 & ~n493 ;
  assign n537 = ~n306 & ~n536 ;
  assign n538 = ~n535 & n537 ;
  assign n539 = n535 & ~n537 ;
  assign n540 = ~n538 & ~n539 ;
  assign n541 = n491 & ~n540 ;
  assign n526 = \226(93)_pad  & \3552(168)_pad  ;
  assign n525 = ~\226(93)_pad  & \3550(167)_pad  ;
  assign n527 = \422(139)_pad  & ~n525 ;
  assign n528 = ~n526 & n527 ;
  assign n530 = \226(93)_pad  & ~\3546(165)_pad  ;
  assign n529 = ~\226(93)_pad  & ~\3548(166)_pad  ;
  assign n531 = ~\422(139)_pad  & ~n529 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = ~n528 & ~n532 ;
  assign n534 = n480 & n533 ;
  assign n542 = \113(43)_pad  & n499 ;
  assign n543 = ~n534 & ~n542 ;
  assign n544 = ~n541 & n543 ;
  assign n545 = n479 & ~n544 ;
  assign n546 = \173(76)_pad  & n504 ;
  assign n547 = \203(86)_pad  & n506 ;
  assign n558 = ~n546 & ~n547 ;
  assign n559 = ~n545 & n558 ;
  assign n560 = ~n557 & n559 ;
  assign n561 = \926(624)_pad  & ~n560 ;
  assign n590 = ~n429 & n551 ;
  assign n586 = n429 & ~n434 ;
  assign n587 = ~n429 & n434 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = ~n551 & ~n588 ;
  assign n591 = n491 & ~n589 ;
  assign n592 = ~n590 & n591 ;
  assign n584 = n339 & n480 ;
  assign n585 = \116(46)_pad  & n499 ;
  assign n593 = ~n584 & ~n585 ;
  assign n594 = ~n592 & n593 ;
  assign n595 = n508 & ~n594 ;
  assign n573 = ~n290 & n291 ;
  assign n574 = ~n292 & ~n573 ;
  assign n576 = n539 & n574 ;
  assign n575 = ~n539 & ~n574 ;
  assign n577 = n491 & ~n575 ;
  assign n578 = ~n576 & n577 ;
  assign n563 = \218(91)_pad  & \3552(168)_pad  ;
  assign n562 = ~\218(91)_pad  & \3550(167)_pad  ;
  assign n564 = \468(143)_pad  & ~n562 ;
  assign n565 = ~n563 & n564 ;
  assign n567 = \218(91)_pad  & ~\3546(165)_pad  ;
  assign n566 = ~\218(91)_pad  & ~\3548(166)_pad  ;
  assign n568 = ~\468(143)_pad  & ~n566 ;
  assign n569 = ~n567 & n568 ;
  assign n570 = ~n565 & ~n569 ;
  assign n571 = n480 & n570 ;
  assign n572 = \53(19)_pad  & n499 ;
  assign n579 = ~n571 & ~n572 ;
  assign n580 = ~n578 & n579 ;
  assign n581 = n479 & ~n580 ;
  assign n582 = \167(74)_pad  & n504 ;
  assign n583 = \197(84)_pad  & n506 ;
  assign n596 = ~n582 & ~n583 ;
  assign n597 = ~n581 & n596 ;
  assign n598 = ~n595 & n597 ;
  assign n599 = \926(624)_pad  & ~n598 ;
  assign n624 = n436 & ~n549 ;
  assign n625 = n440 & ~n624 ;
  assign n626 = ~n422 & ~n625 ;
  assign n627 = n422 & n625 ;
  assign n628 = ~n626 & ~n627 ;
  assign n629 = n491 & ~n628 ;
  assign n623 = n376 & n480 ;
  assign n630 = \121(51)_pad  & n499 ;
  assign n631 = ~n623 & ~n630 ;
  assign n632 = ~n629 & n631 ;
  assign n633 = n508 & ~n632 ;
  assign n610 = n453 & ~n537 ;
  assign n611 = ~n288 & ~n292 ;
  assign n612 = ~n610 & ~n611 ;
  assign n613 = n318 & n612 ;
  assign n614 = ~n318 & ~n612 ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = n491 & n615 ;
  assign n601 = \210(89)_pad  & \3552(168)_pad  ;
  assign n600 = ~\210(89)_pad  & \3550(167)_pad  ;
  assign n602 = \457(142)_pad  & ~n600 ;
  assign n603 = ~n601 & n602 ;
  assign n605 = \210(89)_pad  & ~\3546(165)_pad  ;
  assign n604 = ~\210(89)_pad  & ~\3548(166)_pad  ;
  assign n606 = ~\457(142)_pad  & ~n604 ;
  assign n607 = ~n605 & n606 ;
  assign n608 = ~n603 & ~n607 ;
  assign n609 = n480 & n608 ;
  assign n617 = \114(44)_pad  & n499 ;
  assign n618 = ~n609 & ~n617 ;
  assign n619 = ~n616 & n618 ;
  assign n620 = n479 & ~n619 ;
  assign n621 = \164(73)_pad  & n504 ;
  assign n622 = \194(83)_pad  & n506 ;
  assign n634 = ~n621 & ~n622 ;
  assign n635 = ~n620 & n634 ;
  assign n636 = ~n633 & n635 ;
  assign n637 = \926(624)_pad  & ~n636 ;
  assign n664 = ~n419 & n627 ;
  assign n665 = n419 & ~n627 ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = n491 & n666 ;
  assign n662 = ~n373 & n480 ;
  assign n663 = \123(53)_pad  & n499 ;
  assign n668 = ~n662 & ~n663 ;
  assign n669 = ~n667 & n668 ;
  assign n670 = n508 & ~n669 ;
  assign n648 = ~n293 & n454 ;
  assign n649 = ~n317 & ~n648 ;
  assign n650 = n454 & ~n537 ;
  assign n651 = n649 & ~n650 ;
  assign n652 = n315 & n651 ;
  assign n653 = ~n315 & ~n651 ;
  assign n654 = ~n652 & ~n653 ;
  assign n655 = n491 & n654 ;
  assign n639 = \206(87)_pad  & ~\248(99)_pad  ;
  assign n638 = ~\206(87)_pad  & ~\251(100)_pad  ;
  assign n640 = \446(141)_pad  & ~n638 ;
  assign n641 = ~n639 & n640 ;
  assign n643 = \206(87)_pad  & \242(97)_pad  ;
  assign n642 = ~\206(87)_pad  & \254(101)_pad  ;
  assign n644 = ~\446(141)_pad  & ~n642 ;
  assign n645 = ~n643 & n644 ;
  assign n646 = ~n641 & ~n645 ;
  assign n647 = n480 & n646 ;
  assign n656 = \115(45)_pad  & n499 ;
  assign n657 = ~n647 & ~n656 ;
  assign n658 = ~n655 & n657 ;
  assign n659 = n479 & ~n658 ;
  assign n660 = \161(72)_pad  & n504 ;
  assign n661 = \191(82)_pad  & n506 ;
  assign n671 = ~n660 & ~n661 ;
  assign n672 = ~n659 & n671 ;
  assign n673 = ~n670 & n672 ;
  assign n674 = \926(624)_pad  & ~n673 ;
  assign n675 = \140(64)_pad  & n469 ;
  assign n676 = \4092(176)_pad  & \97(37)_pad  ;
  assign n677 = ~n307 & ~n310 ;
  assign n678 = ~n311 & ~n677 ;
  assign n679 = ~n294 & ~n297 ;
  assign n680 = ~n455 & ~n679 ;
  assign n681 = ~n308 & ~n458 ;
  assign n682 = ~n459 & ~n681 ;
  assign n683 = n680 & ~n682 ;
  assign n684 = ~n680 & n682 ;
  assign n685 = ~n683 & ~n684 ;
  assign n686 = ~n296 & ~n685 ;
  assign n687 = ~n304 & ~n458 ;
  assign n688 = ~n309 & ~n687 ;
  assign n689 = ~n308 & n687 ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = n295 & ~n297 ;
  assign n692 = ~n295 & ~n298 ;
  assign n693 = ~n691 & ~n692 ;
  assign n695 = ~n690 & n693 ;
  assign n694 = n690 & ~n693 ;
  assign n696 = n296 & ~n694 ;
  assign n697 = ~n695 & n696 ;
  assign n698 = ~n686 & ~n697 ;
  assign n699 = \1497(156)_pad  & ~n698 ;
  assign n700 = n296 & n685 ;
  assign n701 = ~\1497(156)_pad  & ~n686 ;
  assign n702 = ~n700 & n701 ;
  assign n703 = ~n699 & ~n702 ;
  assign n704 = n678 & ~n703 ;
  assign n705 = ~n678 & n703 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n299 & ~n302 ;
  assign n708 = ~n303 & ~n707 ;
  assign n709 = \1497(156)_pad  & n312 ;
  assign n710 = ~n462 & ~n709 ;
  assign n711 = ~n317 & ~n453 ;
  assign n712 = ~n454 & ~n711 ;
  assign n713 = ~n315 & n712 ;
  assign n714 = ~n315 & ~n318 ;
  assign n715 = ~n319 & ~n714 ;
  assign n716 = ~n712 & n715 ;
  assign n717 = ~n713 & ~n716 ;
  assign n718 = ~n574 & ~n717 ;
  assign n719 = n574 & n717 ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = n710 & ~n720 ;
  assign n722 = ~n287 & ~n290 ;
  assign n723 = ~n452 & ~n722 ;
  assign n724 = n715 & n723 ;
  assign n725 = ~n715 & ~n723 ;
  assign n726 = ~n724 & ~n725 ;
  assign n727 = ~n611 & ~n649 ;
  assign n728 = ~n293 & n316 ;
  assign n729 = n453 & n728 ;
  assign n730 = ~n727 & ~n729 ;
  assign n732 = n726 & n730 ;
  assign n731 = ~n726 & ~n730 ;
  assign n733 = ~n710 & ~n731 ;
  assign n734 = ~n732 & n733 ;
  assign n735 = ~n721 & ~n734 ;
  assign n736 = n708 & ~n735 ;
  assign n737 = ~n708 & n735 ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = ~n706 & n738 ;
  assign n740 = n706 & ~n738 ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = \4091(175)_pad  & n741 ;
  assign n744 = \234(95)_pad  & ~\248(99)_pad  ;
  assign n743 = ~\234(95)_pad  & ~\251(100)_pad  ;
  assign n745 = \435(140)_pad  & ~n743 ;
  assign n746 = ~n744 & n745 ;
  assign n748 = \234(95)_pad  & \242(97)_pad  ;
  assign n747 = ~\234(95)_pad  & \254(101)_pad  ;
  assign n749 = ~\435(140)_pad  & ~n747 ;
  assign n750 = ~n748 & n749 ;
  assign n751 = ~n746 & ~n750 ;
  assign n753 = \226(93)_pad  & ~\248(99)_pad  ;
  assign n752 = ~\226(93)_pad  & ~\251(100)_pad  ;
  assign n754 = \422(139)_pad  & ~n752 ;
  assign n755 = ~n753 & n754 ;
  assign n757 = \226(93)_pad  & \242(97)_pad  ;
  assign n756 = ~\226(93)_pad  & \254(101)_pad  ;
  assign n758 = ~\422(139)_pad  & ~n756 ;
  assign n759 = ~n757 & n758 ;
  assign n760 = ~n755 & ~n759 ;
  assign n761 = n751 & ~n760 ;
  assign n762 = ~n751 & n760 ;
  assign n763 = ~n761 & ~n762 ;
  assign n765 = \210(89)_pad  & ~\248(99)_pad  ;
  assign n764 = ~\210(89)_pad  & ~\251(100)_pad  ;
  assign n766 = \457(142)_pad  & ~n764 ;
  assign n767 = ~n765 & n766 ;
  assign n769 = \210(89)_pad  & \242(97)_pad  ;
  assign n768 = ~\210(89)_pad  & \254(101)_pad  ;
  assign n770 = ~\457(142)_pad  & ~n768 ;
  assign n771 = ~n769 & n770 ;
  assign n772 = ~n767 & ~n771 ;
  assign n773 = ~n646 & n772 ;
  assign n774 = n646 & ~n772 ;
  assign n775 = ~n773 & ~n774 ;
  assign n777 = \218(91)_pad  & ~\248(99)_pad  ;
  assign n776 = ~\218(91)_pad  & ~\251(100)_pad  ;
  assign n778 = \468(143)_pad  & ~n776 ;
  assign n779 = ~n777 & n778 ;
  assign n781 = \218(91)_pad  & \242(97)_pad  ;
  assign n780 = ~\218(91)_pad  & \254(101)_pad  ;
  assign n782 = ~\468(143)_pad  & ~n780 ;
  assign n783 = ~n781 & n782 ;
  assign n784 = ~n779 & ~n783 ;
  assign n785 = n775 & ~n784 ;
  assign n786 = ~n775 & n784 ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = n763 & n787 ;
  assign n789 = ~n763 & ~n787 ;
  assign n790 = ~n788 & ~n789 ;
  assign n792 = ~\248(99)_pad  & \257(102)_pad  ;
  assign n791 = ~\251(100)_pad  & ~\257(102)_pad  ;
  assign n793 = \389(136)_pad  & ~n791 ;
  assign n794 = ~n792 & n793 ;
  assign n796 = \242(97)_pad  & \257(102)_pad  ;
  assign n795 = \254(101)_pad  & ~\257(102)_pad  ;
  assign n797 = ~\389(136)_pad  & ~n795 ;
  assign n798 = ~n796 & n797 ;
  assign n799 = ~n794 & ~n798 ;
  assign n801 = ~\248(99)_pad  & \281(108)_pad  ;
  assign n800 = ~\251(100)_pad  & ~\281(108)_pad  ;
  assign n802 = \374(134)_pad  & ~n800 ;
  assign n803 = ~n801 & n802 ;
  assign n805 = \242(97)_pad  & \281(108)_pad  ;
  assign n804 = \254(101)_pad  & ~\281(108)_pad  ;
  assign n806 = ~\374(134)_pad  & ~n804 ;
  assign n807 = ~n805 & n806 ;
  assign n808 = ~n803 & ~n807 ;
  assign n810 = ~\248(99)_pad  & \273(106)_pad  ;
  assign n809 = ~\251(100)_pad  & ~\273(106)_pad  ;
  assign n811 = \411(138)_pad  & ~n809 ;
  assign n812 = ~n810 & n811 ;
  assign n814 = \242(97)_pad  & \273(106)_pad  ;
  assign n813 = \254(101)_pad  & ~\273(106)_pad  ;
  assign n815 = ~\411(138)_pad  & ~n813 ;
  assign n816 = ~n814 & n815 ;
  assign n817 = ~n812 & ~n816 ;
  assign n818 = ~n808 & n817 ;
  assign n819 = n808 & ~n817 ;
  assign n820 = ~n818 & ~n819 ;
  assign n822 = ~\248(99)_pad  & \265(104)_pad  ;
  assign n821 = ~\251(100)_pad  & ~\265(104)_pad  ;
  assign n823 = \400(137)_pad  & ~n821 ;
  assign n824 = ~n822 & n823 ;
  assign n826 = \242(97)_pad  & \265(104)_pad  ;
  assign n825 = \254(101)_pad  & ~\265(104)_pad  ;
  assign n827 = ~\400(137)_pad  & ~n825 ;
  assign n828 = ~n826 & n827 ;
  assign n829 = ~n824 & ~n828 ;
  assign n830 = n820 & ~n829 ;
  assign n831 = ~n820 & n829 ;
  assign n832 = ~n830 & ~n831 ;
  assign n833 = n799 & n832 ;
  assign n834 = ~n799 & ~n832 ;
  assign n835 = ~n833 & ~n834 ;
  assign n837 = ~n790 & n835 ;
  assign n836 = n790 & ~n835 ;
  assign n838 = ~\4091(175)_pad  & ~n836 ;
  assign n839 = ~n837 & n838 ;
  assign n840 = ~\4092(176)_pad  & ~n839 ;
  assign n841 = ~n742 & n840 ;
  assign n842 = ~n676 & ~n841 ;
  assign n843 = n479 & ~n842 ;
  assign n844 = \4092(176)_pad  & \94(36)_pad  ;
  assign n845 = ~n397 & ~n403 ;
  assign n846 = ~n404 & ~n845 ;
  assign n847 = n391 & ~n415 ;
  assign n848 = ~n391 & n415 ;
  assign n849 = ~n847 & ~n848 ;
  assign n850 = n846 & n849 ;
  assign n851 = ~n846 & ~n849 ;
  assign n852 = ~n850 & ~n851 ;
  assign n853 = ~n395 & n402 ;
  assign n854 = ~n396 & ~n402 ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = ~n409 & ~n855 ;
  assign n857 = ~n446 & ~n856 ;
  assign n858 = n446 & ~n855 ;
  assign n859 = ~n857 & ~n858 ;
  assign n860 = ~n407 & ~n859 ;
  assign n861 = n407 & n859 ;
  assign n862 = ~n860 & ~n861 ;
  assign n863 = \2174(161)_pad  & ~n862 ;
  assign n864 = ~n389 & n444 ;
  assign n865 = ~n445 & ~n864 ;
  assign n867 = n401 & n865 ;
  assign n866 = ~n401 & ~n865 ;
  assign n868 = n407 & ~n866 ;
  assign n869 = ~n867 & n868 ;
  assign n870 = ~\2174(161)_pad  & ~n860 ;
  assign n871 = ~n869 & n870 ;
  assign n872 = ~n863 & ~n871 ;
  assign n873 = \2174(161)_pad  & n416 ;
  assign n874 = ~n448 & ~n873 ;
  assign n875 = ~n422 & ~n440 ;
  assign n876 = n419 & ~n875 ;
  assign n877 = ~n419 & n875 ;
  assign n878 = ~n876 & ~n877 ;
  assign n879 = n588 & ~n878 ;
  assign n880 = ~n588 & n878 ;
  assign n881 = ~n879 & ~n880 ;
  assign n882 = n874 & ~n881 ;
  assign n883 = ~n429 & ~n433 ;
  assign n884 = ~n439 & ~n883 ;
  assign n885 = ~n427 & ~n586 ;
  assign n886 = ~n422 & ~n885 ;
  assign n887 = n419 & ~n886 ;
  assign n888 = ~n419 & n886 ;
  assign n889 = ~n887 & ~n888 ;
  assign n890 = n884 & n889 ;
  assign n891 = ~n884 & ~n889 ;
  assign n892 = ~n890 & ~n891 ;
  assign n893 = ~n874 & ~n892 ;
  assign n894 = ~n882 & ~n893 ;
  assign n895 = n872 & ~n894 ;
  assign n896 = ~n872 & n894 ;
  assign n897 = ~n895 & ~n896 ;
  assign n898 = n852 & n897 ;
  assign n899 = ~n852 & ~n897 ;
  assign n900 = ~n898 & ~n899 ;
  assign n901 = \4091(175)_pad  & n900 ;
  assign n902 = ~\248(99)_pad  & \514(147)_pad  ;
  assign n903 = \242(97)_pad  & ~\514(147)_pad  ;
  assign n904 = ~n902 & ~n903 ;
  assign n905 = ~n373 & n376 ;
  assign n906 = ~n377 & ~n905 ;
  assign n907 = n330 & n339 ;
  assign n908 = ~n340 & ~n907 ;
  assign n909 = n906 & ~n908 ;
  assign n910 = ~n906 & n908 ;
  assign n911 = ~n909 & ~n910 ;
  assign n912 = n904 & n911 ;
  assign n913 = ~n904 & ~n911 ;
  assign n914 = ~n912 & ~n913 ;
  assign n916 = ~\248(99)_pad  & \324(120)_pad  ;
  assign n915 = ~\251(100)_pad  & ~\324(120)_pad  ;
  assign n917 = \503(146)_pad  & ~n915 ;
  assign n918 = ~n916 & n917 ;
  assign n920 = \242(97)_pad  & \324(120)_pad  ;
  assign n919 = \254(101)_pad  & ~\324(120)_pad  ;
  assign n921 = ~\503(146)_pad  & ~n919 ;
  assign n922 = ~n920 & n921 ;
  assign n923 = ~n918 & ~n922 ;
  assign n924 = n343 & ~n923 ;
  assign n925 = ~n343 & n923 ;
  assign n926 = ~n924 & ~n925 ;
  assign n928 = ~\248(99)_pad  & \341(125)_pad  ;
  assign n927 = ~\251(100)_pad  & ~\341(125)_pad  ;
  assign n929 = \523(148)_pad  & ~n927 ;
  assign n930 = ~n928 & n929 ;
  assign n932 = \242(97)_pad  & \341(125)_pad  ;
  assign n931 = \254(101)_pad  & ~\341(125)_pad  ;
  assign n933 = ~\523(148)_pad  & ~n931 ;
  assign n934 = ~n932 & n933 ;
  assign n935 = ~n930 & ~n934 ;
  assign n937 = ~\248(99)_pad  & \351(127)_pad  ;
  assign n936 = ~\251(100)_pad  & ~\351(127)_pad  ;
  assign n938 = \534(149)_pad  & ~n936 ;
  assign n939 = ~n937 & n938 ;
  assign n941 = \242(97)_pad  & \351(127)_pad  ;
  assign n940 = \254(101)_pad  & ~\351(127)_pad  ;
  assign n942 = ~\534(149)_pad  & ~n940 ;
  assign n943 = ~n941 & n942 ;
  assign n944 = ~n939 & ~n943 ;
  assign n945 = n935 & ~n944 ;
  assign n946 = ~n935 & n944 ;
  assign n947 = ~n945 & ~n946 ;
  assign n948 = n926 & n947 ;
  assign n949 = ~n926 & ~n947 ;
  assign n950 = ~n948 & ~n949 ;
  assign n952 = n914 & n950 ;
  assign n951 = ~n914 & ~n950 ;
  assign n953 = ~\4091(175)_pad  & ~n951 ;
  assign n954 = ~n952 & n953 ;
  assign n955 = ~\4092(176)_pad  & ~n954 ;
  assign n956 = ~n901 & n955 ;
  assign n957 = ~n844 & ~n956 ;
  assign n958 = n508 & ~n957 ;
  assign n959 = \179(78)_pad  & n504 ;
  assign n960 = \176(77)_pad  & n506 ;
  assign n961 = ~n959 & ~n960 ;
  assign n962 = ~n958 & n961 ;
  assign n963 = ~n843 & n962 ;
  assign n964 = \926(624)_pad  & ~n963 ;
  assign n986 = \4(1)_pad  & n296 ;
  assign n987 = ~\4(1)_pad  & ~n296 ;
  assign n988 = ~n986 & ~n987 ;
  assign n989 = n491 & n988 ;
  assign n977 = \281(108)_pad  & \3552(168)_pad  ;
  assign n976 = ~\281(108)_pad  & \3550(167)_pad  ;
  assign n978 = \374(134)_pad  & ~n976 ;
  assign n979 = ~n977 & n978 ;
  assign n981 = \281(108)_pad  & ~\3546(165)_pad  ;
  assign n980 = ~\281(108)_pad  & ~\3548(166)_pad  ;
  assign n982 = ~\374(134)_pad  & ~n980 ;
  assign n983 = ~n981 & n982 ;
  assign n984 = ~n979 & ~n983 ;
  assign n985 = n480 & n984 ;
  assign n990 = \117(47)_pad  & n499 ;
  assign n991 = ~n985 & ~n990 ;
  assign n992 = ~n989 & n991 ;
  assign n993 = n479 & ~n992 ;
  assign n966 = \54(20)_pad  & ~n407 ;
  assign n967 = ~\54(20)_pad  & n407 ;
  assign n968 = ~n966 & ~n967 ;
  assign n969 = n491 & ~n968 ;
  assign n965 = n343 & n480 ;
  assign n970 = \131(59)_pad  & n499 ;
  assign n971 = ~n965 & ~n970 ;
  assign n972 = ~n969 & n971 ;
  assign n973 = n508 & ~n972 ;
  assign n974 = \185(80)_pad  & n504 ;
  assign n975 = \182(79)_pad  & n506 ;
  assign n994 = ~n974 & ~n975 ;
  assign n995 = ~n973 & n994 ;
  assign n996 = ~n993 & n995 ;
  assign n997 = \926(624)_pad  & ~n996 ;
  assign n1020 = \4(1)_pad  & ~n295 ;
  assign n1021 = ~n294 & ~n1020 ;
  assign n1022 = n299 & ~n1021 ;
  assign n1023 = ~n299 & n1021 ;
  assign n1024 = ~n1022 & ~n1023 ;
  assign n1025 = n491 & n1024 ;
  assign n1011 = \273(106)_pad  & \3552(168)_pad  ;
  assign n1010 = ~\273(106)_pad  & \3550(167)_pad  ;
  assign n1012 = \411(138)_pad  & ~n1010 ;
  assign n1013 = ~n1011 & n1012 ;
  assign n1015 = \273(106)_pad  & ~\3546(165)_pad  ;
  assign n1014 = ~\273(106)_pad  & ~\3548(166)_pad  ;
  assign n1016 = ~\411(138)_pad  & ~n1014 ;
  assign n1017 = ~n1015 & n1016 ;
  assign n1018 = ~n1013 & ~n1017 ;
  assign n1019 = n480 & n1018 ;
  assign n1026 = \126(54)_pad  & n499 ;
  assign n1027 = ~n1019 & ~n1026 ;
  assign n1028 = ~n1025 & n1027 ;
  assign n1029 = n479 & ~n1028 ;
  assign n1001 = ~n402 & ~n967 ;
  assign n1002 = ~n401 & n1001 ;
  assign n1000 = ~n403 & n967 ;
  assign n1003 = n491 & ~n1000 ;
  assign n1004 = ~n1002 & n1003 ;
  assign n998 = n370 & n480 ;
  assign n999 = \129(57)_pad  & n499 ;
  assign n1005 = ~n998 & ~n999 ;
  assign n1006 = ~n1004 & n1005 ;
  assign n1007 = n508 & ~n1006 ;
  assign n1008 = \158(71)_pad  & n504 ;
  assign n1009 = \188(81)_pad  & n506 ;
  assign n1030 = ~n1008 & ~n1009 ;
  assign n1031 = ~n1007 & n1030 ;
  assign n1032 = ~n1029 & n1031 ;
  assign n1033 = \926(624)_pad  & ~n1032 ;
  assign n1056 = ~n298 & ~n1021 ;
  assign n1057 = ~n297 & ~n1056 ;
  assign n1058 = n302 & ~n1057 ;
  assign n1059 = ~n302 & n1057 ;
  assign n1060 = ~n1058 & ~n1059 ;
  assign n1061 = n491 & n1060 ;
  assign n1047 = \265(104)_pad  & \3552(168)_pad  ;
  assign n1046 = ~\265(104)_pad  & \3550(167)_pad  ;
  assign n1048 = \400(137)_pad  & ~n1046 ;
  assign n1049 = ~n1047 & n1048 ;
  assign n1051 = \265(104)_pad  & ~\3546(165)_pad  ;
  assign n1050 = ~\265(104)_pad  & ~\3548(166)_pad  ;
  assign n1052 = ~\400(137)_pad  & ~n1050 ;
  assign n1053 = ~n1051 & n1052 ;
  assign n1054 = ~n1049 & ~n1053 ;
  assign n1055 = n480 & n1054 ;
  assign n1062 = \127(55)_pad  & n499 ;
  assign n1063 = ~n1055 & ~n1062 ;
  assign n1064 = ~n1061 & n1063 ;
  assign n1065 = n479 & ~n1064 ;
  assign n1035 = ~n401 & ~n1001 ;
  assign n1036 = n397 & n1035 ;
  assign n1037 = ~n397 & ~n1035 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = n491 & ~n1038 ;
  assign n1034 = n352 & n480 ;
  assign n1040 = \119(49)_pad  & n499 ;
  assign n1041 = ~n1034 & ~n1040 ;
  assign n1042 = ~n1039 & n1041 ;
  assign n1043 = n508 & ~n1042 ;
  assign n1044 = \152(69)_pad  & n504 ;
  assign n1045 = \155(70)_pad  & n506 ;
  assign n1066 = ~n1044 & ~n1045 ;
  assign n1067 = ~n1043 & n1066 ;
  assign n1068 = ~n1065 & n1067 ;
  assign n1069 = \926(624)_pad  & ~n1068 ;
  assign n1092 = ~n458 & ~n492 ;
  assign n1093 = n310 & n1092 ;
  assign n1094 = ~n310 & ~n1092 ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = n491 & ~n1095 ;
  assign n1083 = \257(102)_pad  & \3552(168)_pad  ;
  assign n1082 = ~\257(102)_pad  & \3550(167)_pad  ;
  assign n1084 = \389(136)_pad  & ~n1082 ;
  assign n1085 = ~n1083 & n1084 ;
  assign n1087 = \257(102)_pad  & ~\3546(165)_pad  ;
  assign n1086 = ~\257(102)_pad  & ~\3548(166)_pad  ;
  assign n1088 = ~\389(136)_pad  & ~n1086 ;
  assign n1089 = ~n1087 & n1088 ;
  assign n1090 = ~n1085 & ~n1089 ;
  assign n1091 = n480 & n1090 ;
  assign n1097 = \128(56)_pad  & n499 ;
  assign n1098 = ~n1091 & ~n1097 ;
  assign n1099 = ~n1096 & n1098 ;
  assign n1100 = n479 & ~n1099 ;
  assign n1071 = ~n444 & ~n510 ;
  assign n1072 = n391 & n1071 ;
  assign n1073 = ~n391 & ~n1071 ;
  assign n1074 = ~n1072 & ~n1073 ;
  assign n1075 = n491 & ~n1074 ;
  assign n1070 = n380 & n480 ;
  assign n1076 = \130(58)_pad  & n499 ;
  assign n1077 = ~n1070 & ~n1076 ;
  assign n1078 = ~n1075 & n1077 ;
  assign n1079 = n508 & ~n1078 ;
  assign n1080 = \146(67)_pad  & n504 ;
  assign n1081 = \149(68)_pad  & n506 ;
  assign n1101 = ~n1080 & ~n1081 ;
  assign n1102 = ~n1079 & n1101 ;
  assign n1103 = ~n1100 & n1102 ;
  assign n1104 = \926(624)_pad  & ~n1103 ;
  assign n1106 = \2358(162)_pad  & \81(29)_pad  ;
  assign n1105 = ~\2358(162)_pad  & \26(9)_pad  ;
  assign n1107 = n469 & ~n1105 ;
  assign n1108 = ~n1106 & n1107 ;
  assign n1109 = \144(354)_pad  & ~n1108 ;
  assign n1116 = ~\1691(159)_pad  & ~\1694(160)_pad  ;
  assign n1117 = ~n519 & n1116 ;
  assign n1110 = \1691(159)_pad  & ~\1694(160)_pad  ;
  assign n1111 = ~n502 & n1110 ;
  assign n1112 = \1691(159)_pad  & \1694(160)_pad  ;
  assign n1113 = \170(75)_pad  & n1112 ;
  assign n1114 = ~\1691(159)_pad  & \1694(160)_pad  ;
  assign n1115 = \200(85)_pad  & n1114 ;
  assign n1118 = ~n1113 & ~n1115 ;
  assign n1119 = ~n1111 & n1118 ;
  assign n1120 = ~n1117 & n1119 ;
  assign n1121 = \926(624)_pad  & ~n1120 ;
  assign n1125 = ~n556 & n1116 ;
  assign n1122 = ~n544 & n1110 ;
  assign n1123 = \173(76)_pad  & n1112 ;
  assign n1124 = \203(86)_pad  & n1114 ;
  assign n1126 = ~n1123 & ~n1124 ;
  assign n1127 = ~n1122 & n1126 ;
  assign n1128 = ~n1125 & n1127 ;
  assign n1129 = \926(624)_pad  & ~n1128 ;
  assign n1133 = ~n594 & n1116 ;
  assign n1130 = ~n580 & n1110 ;
  assign n1131 = \167(74)_pad  & n1112 ;
  assign n1132 = \197(84)_pad  & n1114 ;
  assign n1134 = ~n1131 & ~n1132 ;
  assign n1135 = ~n1130 & n1134 ;
  assign n1136 = ~n1133 & n1135 ;
  assign n1137 = \926(624)_pad  & ~n1136 ;
  assign n1141 = ~n632 & n1116 ;
  assign n1138 = ~n619 & n1110 ;
  assign n1139 = \164(73)_pad  & n1112 ;
  assign n1140 = \194(83)_pad  & n1114 ;
  assign n1142 = ~n1139 & ~n1140 ;
  assign n1143 = ~n1138 & n1142 ;
  assign n1144 = ~n1141 & n1143 ;
  assign n1145 = \926(624)_pad  & ~n1144 ;
  assign n1149 = ~n669 & n1116 ;
  assign n1146 = ~n658 & n1110 ;
  assign n1147 = \161(72)_pad  & n1112 ;
  assign n1148 = \191(82)_pad  & n1114 ;
  assign n1150 = ~n1147 & ~n1148 ;
  assign n1151 = ~n1146 & n1150 ;
  assign n1152 = ~n1149 & n1151 ;
  assign n1153 = \926(624)_pad  & ~n1152 ;
  assign n1154 = ~n842 & n1110 ;
  assign n1155 = ~n957 & n1116 ;
  assign n1156 = \179(78)_pad  & n1112 ;
  assign n1157 = \176(77)_pad  & n1114 ;
  assign n1158 = ~n1156 & ~n1157 ;
  assign n1159 = ~n1155 & n1158 ;
  assign n1160 = ~n1154 & n1159 ;
  assign n1161 = \926(624)_pad  & ~n1160 ;
  assign n1165 = ~n992 & n1110 ;
  assign n1162 = ~n972 & n1116 ;
  assign n1163 = \185(80)_pad  & n1112 ;
  assign n1164 = \182(79)_pad  & n1114 ;
  assign n1166 = ~n1163 & ~n1164 ;
  assign n1167 = ~n1162 & n1166 ;
  assign n1168 = ~n1165 & n1167 ;
  assign n1169 = \926(624)_pad  & ~n1168 ;
  assign n1173 = ~n1028 & n1110 ;
  assign n1170 = ~n1006 & n1116 ;
  assign n1171 = \158(71)_pad  & n1112 ;
  assign n1172 = \188(81)_pad  & n1114 ;
  assign n1174 = ~n1171 & ~n1172 ;
  assign n1175 = ~n1170 & n1174 ;
  assign n1176 = ~n1173 & n1175 ;
  assign n1177 = \926(624)_pad  & ~n1176 ;
  assign n1181 = ~n1064 & n1110 ;
  assign n1178 = ~n1042 & n1116 ;
  assign n1179 = \152(69)_pad  & n1112 ;
  assign n1180 = \155(70)_pad  & n1114 ;
  assign n1182 = ~n1179 & ~n1180 ;
  assign n1183 = ~n1178 & n1182 ;
  assign n1184 = ~n1181 & n1183 ;
  assign n1185 = \926(624)_pad  & ~n1184 ;
  assign n1189 = ~n1099 & n1110 ;
  assign n1186 = ~n1078 & n1116 ;
  assign n1187 = \146(67)_pad  & n1112 ;
  assign n1188 = \149(68)_pad  & n1114 ;
  assign n1190 = ~n1187 & ~n1188 ;
  assign n1191 = ~n1186 & n1190 ;
  assign n1192 = ~n1189 & n1191 ;
  assign n1193 = \926(624)_pad  & ~n1192 ;
  assign n1195 = \2358(162)_pad  & ~\34(12)_pad  ;
  assign n1194 = ~\2358(162)_pad  & ~\88(34)_pad  ;
  assign n1196 = n469 & ~n1194 ;
  assign n1197 = ~n1195 & n1196 ;
  assign n1199 = \23(6)_pad  & \2358(162)_pad  ;
  assign n1198 = ~\2358(162)_pad  & \79(27)_pad  ;
  assign n1200 = n469 & ~n1198 ;
  assign n1201 = ~n1199 & n1200 ;
  assign n1202 = \144(354)_pad  & ~n1201 ;
  assign n1209 = ~\4089(173)_pad  & ~\4090(174)_pad  ;
  assign n1210 = ~n669 & n1209 ;
  assign n1203 = \4089(173)_pad  & ~\4090(174)_pad  ;
  assign n1204 = ~n658 & n1203 ;
  assign n1205 = \4089(173)_pad  & \4090(174)_pad  ;
  assign n1206 = \106(40)_pad  & n1205 ;
  assign n1207 = ~\4089(173)_pad  & \4090(174)_pad  ;
  assign n1208 = \109(41)_pad  & n1207 ;
  assign n1211 = ~n1206 & ~n1208 ;
  assign n1212 = ~n1204 & n1211 ;
  assign n1213 = ~n1210 & n1212 ;
  assign n1215 = \2358(162)_pad  & \80(28)_pad  ;
  assign n1214 = ~\2358(162)_pad  & \82(30)_pad  ;
  assign n1216 = n469 & ~n1214 ;
  assign n1217 = ~n1215 & n1216 ;
  assign n1218 = \144(354)_pad  & ~n1217 ;
  assign n1225 = ~\4087(171)_pad  & \4088(172)_pad  ;
  assign n1226 = ~n992 & n1225 ;
  assign n1219 = ~\4087(171)_pad  & ~\4088(172)_pad  ;
  assign n1220 = ~n972 & n1219 ;
  assign n1221 = \4087(171)_pad  & \4088(172)_pad  ;
  assign n1222 = \61(21)_pad  & n1221 ;
  assign n1223 = \4087(171)_pad  & ~\4088(172)_pad  ;
  assign n1224 = \11(2)_pad  & n1223 ;
  assign n1227 = ~n1222 & ~n1224 ;
  assign n1228 = ~n1220 & n1227 ;
  assign n1229 = ~n1226 & n1228 ;
  assign n1233 = ~n669 & n1219 ;
  assign n1230 = ~n658 & n1225 ;
  assign n1231 = \106(40)_pad  & n1221 ;
  assign n1232 = \109(41)_pad  & n1223 ;
  assign n1234 = ~n1231 & ~n1232 ;
  assign n1235 = ~n1230 & n1234 ;
  assign n1236 = ~n1233 & n1235 ;
  assign n1240 = ~n632 & n1219 ;
  assign n1237 = ~n619 & n1225 ;
  assign n1238 = \49(17)_pad  & n1221 ;
  assign n1239 = \46(16)_pad  & n1223 ;
  assign n1241 = ~n1238 & ~n1239 ;
  assign n1242 = ~n1237 & n1241 ;
  assign n1243 = ~n1240 & n1242 ;
  assign n1247 = ~n594 & n1219 ;
  assign n1244 = ~n580 & n1225 ;
  assign n1245 = \103(39)_pad  & n1221 ;
  assign n1246 = \100(38)_pad  & n1223 ;
  assign n1248 = ~n1245 & ~n1246 ;
  assign n1249 = ~n1244 & n1248 ;
  assign n1250 = ~n1247 & n1249 ;
  assign n1254 = ~n556 & n1219 ;
  assign n1251 = ~n544 & n1225 ;
  assign n1252 = \40(14)_pad  & n1221 ;
  assign n1253 = \91(35)_pad  & n1223 ;
  assign n1255 = ~n1252 & ~n1253 ;
  assign n1256 = ~n1251 & n1255 ;
  assign n1257 = ~n1254 & n1256 ;
  assign n1261 = ~n519 & n1219 ;
  assign n1258 = ~n502 & n1225 ;
  assign n1259 = \37(13)_pad  & n1221 ;
  assign n1260 = \43(15)_pad  & n1223 ;
  assign n1262 = ~n1259 & ~n1260 ;
  assign n1263 = ~n1258 & n1262 ;
  assign n1264 = ~n1261 & n1263 ;
  assign n1268 = ~n1099 & n1225 ;
  assign n1265 = ~n1078 & n1219 ;
  assign n1266 = \20(5)_pad  & n1221 ;
  assign n1267 = \76(26)_pad  & n1223 ;
  assign n1269 = ~n1266 & ~n1267 ;
  assign n1270 = ~n1265 & n1269 ;
  assign n1271 = ~n1268 & n1270 ;
  assign n1275 = ~n1064 & n1225 ;
  assign n1272 = ~n1042 & n1219 ;
  assign n1273 = \17(4)_pad  & n1221 ;
  assign n1274 = \73(25)_pad  & n1223 ;
  assign n1276 = ~n1273 & ~n1274 ;
  assign n1277 = ~n1272 & n1276 ;
  assign n1278 = ~n1275 & n1277 ;
  assign n1282 = ~n1028 & n1225 ;
  assign n1279 = ~n1006 & n1219 ;
  assign n1280 = \70(24)_pad  & n1221 ;
  assign n1281 = \67(23)_pad  & n1223 ;
  assign n1283 = ~n1280 & ~n1281 ;
  assign n1284 = ~n1279 & n1283 ;
  assign n1285 = ~n1282 & n1284 ;
  assign n1289 = ~n842 & n1225 ;
  assign n1286 = ~n957 & n1219 ;
  assign n1287 = \64(22)_pad  & n1221 ;
  assign n1288 = \14(3)_pad  & n1223 ;
  assign n1290 = ~n1287 & ~n1288 ;
  assign n1291 = ~n1286 & n1290 ;
  assign n1292 = ~n1289 & n1291 ;
  assign n1296 = ~n632 & n1209 ;
  assign n1293 = ~n619 & n1203 ;
  assign n1294 = \49(17)_pad  & n1205 ;
  assign n1295 = \46(16)_pad  & n1207 ;
  assign n1297 = ~n1294 & ~n1295 ;
  assign n1298 = ~n1293 & n1297 ;
  assign n1299 = ~n1296 & n1298 ;
  assign n1303 = ~n594 & n1209 ;
  assign n1300 = ~n580 & n1203 ;
  assign n1301 = \103(39)_pad  & n1205 ;
  assign n1302 = \100(38)_pad  & n1207 ;
  assign n1304 = ~n1301 & ~n1302 ;
  assign n1305 = ~n1300 & n1304 ;
  assign n1306 = ~n1303 & n1305 ;
  assign n1310 = ~n556 & n1209 ;
  assign n1307 = ~n544 & n1203 ;
  assign n1308 = \40(14)_pad  & n1205 ;
  assign n1309 = \91(35)_pad  & n1207 ;
  assign n1311 = ~n1308 & ~n1309 ;
  assign n1312 = ~n1307 & n1311 ;
  assign n1313 = ~n1310 & n1312 ;
  assign n1317 = ~n519 & n1209 ;
  assign n1314 = ~n502 & n1203 ;
  assign n1315 = \37(13)_pad  & n1205 ;
  assign n1316 = \43(15)_pad  & n1207 ;
  assign n1318 = ~n1315 & ~n1316 ;
  assign n1319 = ~n1314 & n1318 ;
  assign n1320 = ~n1317 & n1319 ;
  assign n1324 = ~n1099 & n1203 ;
  assign n1321 = ~n1078 & n1209 ;
  assign n1322 = \20(5)_pad  & n1205 ;
  assign n1323 = \76(26)_pad  & n1207 ;
  assign n1325 = ~n1322 & ~n1323 ;
  assign n1326 = ~n1321 & n1325 ;
  assign n1327 = ~n1324 & n1326 ;
  assign n1331 = ~n1064 & n1203 ;
  assign n1328 = ~n1042 & n1209 ;
  assign n1329 = \17(4)_pad  & n1205 ;
  assign n1330 = \73(25)_pad  & n1207 ;
  assign n1332 = ~n1329 & ~n1330 ;
  assign n1333 = ~n1328 & n1332 ;
  assign n1334 = ~n1331 & n1333 ;
  assign n1338 = ~n1028 & n1203 ;
  assign n1335 = ~n1006 & n1209 ;
  assign n1336 = \70(24)_pad  & n1205 ;
  assign n1337 = \67(23)_pad  & n1207 ;
  assign n1339 = ~n1336 & ~n1337 ;
  assign n1340 = ~n1335 & n1339 ;
  assign n1341 = ~n1338 & n1340 ;
  assign n1345 = ~n842 & n1203 ;
  assign n1342 = ~n957 & n1209 ;
  assign n1343 = \64(22)_pad  & n1205 ;
  assign n1344 = \14(3)_pad  & n1207 ;
  assign n1346 = ~n1343 & ~n1344 ;
  assign n1347 = ~n1342 & n1346 ;
  assign n1348 = ~n1345 & n1347 ;
  assign n1349 = \144(354)_pad  & \145(66)_pad  ;
  assign n1350 = \132(60)_pad  & ~n627 ;
  assign n1351 = ~\132(60)_pad  & n627 ;
  assign n1352 = ~n1350 & ~n1351 ;
  assign n1353 = \136(62)_pad  & ~\973(202)_pad  ;
  assign n1354 = \83(31)_pad  & n469 ;
  assign n1355 = n491 & n900 ;
  assign n1356 = ~n499 & ~n955 ;
  assign n1357 = \120(50)_pad  & n499 ;
  assign n1358 = ~n1356 & ~n1357 ;
  assign n1359 = ~n1355 & n1358 ;
  assign n1360 = \27(10)_pad  & ~\2824(163)_pad  ;
  assign n1361 = \386(135)_pad  & \556(153)_pad  ;
  assign n1362 = n394 & ~n422 ;
  assign n1363 = ~n394 & n422 ;
  assign n1364 = ~n1362 & ~n1363 ;
  assign n1365 = ~\332(122)_pad  & \369(131)_pad  ;
  assign n1366 = \332(122)_pad  & \372(132)_pad  ;
  assign n1367 = ~n1365 & ~n1366 ;
  assign n1368 = n426 & ~n1367 ;
  assign n1369 = ~n426 & n1367 ;
  assign n1370 = ~n1368 & ~n1369 ;
  assign n1371 = n1364 & ~n1370 ;
  assign n1372 = ~n1364 & n1370 ;
  assign n1373 = ~n1371 & ~n1372 ;
  assign n1374 = ~n407 & ~n419 ;
  assign n1375 = n407 & n419 ;
  assign n1376 = ~n1374 & ~n1375 ;
  assign n1377 = n400 & ~n1376 ;
  assign n1378 = ~n400 & n1376 ;
  assign n1379 = ~n1377 & ~n1378 ;
  assign n1380 = n432 & n1379 ;
  assign n1381 = ~n432 & ~n1379 ;
  assign n1382 = ~n1380 & ~n1381 ;
  assign n1383 = ~n388 & n412 ;
  assign n1384 = ~\331(121)_pad  & n388 ;
  assign n1385 = ~n1383 & ~n1384 ;
  assign n1386 = n1382 & ~n1385 ;
  assign n1387 = ~n1382 & n1385 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = n1373 & n1388 ;
  assign n1390 = ~n1373 & ~n1388 ;
  assign n1391 = ~n1389 & ~n1390 ;
  assign n1392 = \245(98)_pad  & \559(154)_pad  ;
  assign n1393 = n387 & n1392 ;
  assign n1394 = n1361 & n1393 ;
  assign n1395 = n259 & n1394 ;
  assign n1396 = n286 & n1395 ;
  assign n1397 = ~n235 & n1396 ;
  assign n1398 = n1391 & n1397 ;
  assign n1402 = ~n992 & n1203 ;
  assign n1399 = ~n972 & n1209 ;
  assign n1400 = \61(21)_pad  & n1205 ;
  assign n1401 = \11(2)_pad  & n1207 ;
  assign n1403 = ~n1400 & ~n1401 ;
  assign n1404 = ~n1399 & n1403 ;
  assign n1405 = ~n1402 & n1404 ;
  assign n1406 = n491 & n741 ;
  assign n1407 = ~n499 & ~n840 ;
  assign n1408 = \118(48)_pad  & n499 ;
  assign n1409 = ~n1407 & ~n1408 ;
  assign n1410 = ~n1406 & n1409 ;
  assign n1420 = \3724(170)_pad  & n666 ;
  assign n1419 = \123(53)_pad  & ~\3724(170)_pad  ;
  assign n1421 = \3717(169)_pad  & ~n1419 ;
  assign n1422 = ~n1420 & n1421 ;
  assign n1411 = \135(61)_pad  & \4115(177)_pad  ;
  assign n1413 = \132(60)_pad  & ~n419 ;
  assign n1414 = ~\132(60)_pad  & n419 ;
  assign n1415 = ~n1413 & ~n1414 ;
  assign n1416 = \3724(170)_pad  & ~n1415 ;
  assign n1412 = ~\3724(170)_pad  & ~n373 ;
  assign n1417 = ~\3717(169)_pad  & ~n1412 ;
  assign n1418 = ~n1416 & n1417 ;
  assign n1423 = ~n1411 & ~n1418 ;
  assign n1424 = ~n1422 & n1423 ;
  assign n1425 = ~n574 & ~n988 ;
  assign n1426 = ~n1024 & n1425 ;
  assign n1427 = ~n1060 & n1426 ;
  assign n1428 = n1095 & n1427 ;
  assign n1429 = n497 & n1428 ;
  assign n1430 = n540 & n1429 ;
  assign n1431 = ~n615 & n1430 ;
  assign n1432 = ~n654 & n1431 ;
  assign n1433 = n403 & n968 ;
  assign n1434 = ~n588 & n1433 ;
  assign n1435 = n1038 & n1434 ;
  assign n1436 = n1074 & n1435 ;
  assign n1437 = ~n515 & n1436 ;
  assign n1438 = n552 & n1437 ;
  assign n1439 = n628 & n1438 ;
  assign n1440 = ~n666 & n1439 ;
  assign n1444 = ~n1018 & ~n1054 ;
  assign n1445 = ~n1090 & n1444 ;
  assign n1441 = ~n489 & ~n533 ;
  assign n1442 = ~n570 & ~n608 ;
  assign n1443 = ~n646 & ~n984 ;
  assign n1446 = n1442 & n1443 ;
  assign n1447 = n1441 & n1446 ;
  assign n1448 = n1445 & n1447 ;
  assign \1000(2168)_pad  = n235 ;
  assign \1002(1920)_pad  = ~n259 ;
  assign \1004(1977)_pad  = ~n286 ;
  assign \588(1696)_pad  = n321 ;
  assign \593(733)_pad  = ~\889(734)_pad  ;
  assign \598(1623)_pad  = n386 ;
  assign \599(269)_pad  = ~\348(126)_pad  ;
  assign \600(259)_pad  = ~\366(130)_pad  ;
  assign \601(220)_pad  = n387 ;
  assign \604(223)_pad  = ~\545(150)_pad  ;
  assign \606(407)_pad  = ~\892(408)_pad  ;
  assign \611(275)_pad  = ~\338(124)_pad  ;
  assign \612(263)_pad  = ~\358(128)_pad  ;
  assign \615(1750)_pad  = n438 ;
  assign \618(1925)_pad  = ~n451 ;
  assign \621(1893)_pad  = ~n467 ;
  assign \626(1752)_pad  = n438 ;
  assign \632(1692)_pad  = n321 ;
  assign \634(665)_pad  = n468 ;
  assign \636(1280)_pad  = ~n473 ;
  assign \639(1275)_pad  = n478 ;
  assign \642(2222)_pad  = n524 ;
  assign \645(2271)_pad  = n561 ;
  assign \648(2295)_pad  = n599 ;
  assign \651(2314)_pad  = n637 ;
  assign \654(2315)_pad  = n674 ;
  assign \656(621)_pad  = ~n675 ;
  assign \658(2483)_pad  = ~n964 ;
  assign \661(2178)_pad  = n997 ;
  assign \664(2223)_pad  = n1033 ;
  assign \667(2224)_pad  = n1069 ;
  assign \670(2225)_pad  = n1104 ;
  assign \673(1276)_pad  = n1109 ;
  assign \676(2229)_pad  = n1121 ;
  assign \679(2272)_pad  = n1129 ;
  assign \682(2296)_pad  = n1137 ;
  assign \685(2316)_pad  = n1145 ;
  assign \688(2317)_pad  = n1153 ;
  assign \690(2484)_pad  = ~n1161 ;
  assign \693(2179)_pad  = n1169 ;
  assign \696(2226)_pad  = n1177 ;
  assign \699(2227)_pad  = n1185 ;
  assign \702(2228)_pad  = n1193 ;
  assign \704(1281)_pad  = ~n1197 ;
  assign \707(1277)_pad  = n1202 ;
  assign \712(2297)_pad  = ~n1213 ;
  assign \715(1278)_pad  = n1218 ;
  assign \722(2131)_pad  = ~n1229 ;
  assign \727(2298)_pad  = ~n1236 ;
  assign \732(2300)_pad  = ~n1243 ;
  assign \737(2279)_pad  = ~n1250 ;
  assign \742(2238)_pad  = ~n1257 ;
  assign \747(2187)_pad  = ~n1264 ;
  assign \752(2189)_pad  = ~n1271 ;
  assign \757(2190)_pad  = ~n1278 ;
  assign \762(2184)_pad  = ~n1285 ;
  assign \767(2479)_pad  = ~n1292 ;
  assign \772(2299)_pad  = ~n1299 ;
  assign \777(2278)_pad  = ~n1306 ;
  assign \782(2239)_pad  = ~n1313 ;
  assign \787(2186)_pad  = ~n1320 ;
  assign \792(2188)_pad  = ~n1327 ;
  assign \797(2191)_pad  = ~n1334 ;
  assign \802(2183)_pad  = ~n1341 ;
  assign \807(2480)_pad  = ~n1348 ;
  assign \809(655)_pad  = ~n469 ;
  assign \810(356)_pad  = n1349 ;
  assign \813(2260)_pad  = n1352 ;
  assign \815(627)_pad  = n1353 ;
  assign \820(1283)_pad  = ~n1354 ;
  assign \822(1933)_pad  = n972 ;
  assign \824(2274)_pad  = n669 ;
  assign \826(2275)_pad  = n632 ;
  assign \828(2233)_pad  = n594 ;
  assign \830(2182)_pad  = n556 ;
  assign \832(2133)_pad  = n519 ;
  assign \834(2123)_pad  = n1078 ;
  assign \836(2128)_pad  = n1042 ;
  assign \838(2064)_pad  = n1006 ;
  assign \843(2455)_pad  = ~n1359 ;
  assign \845(845)_pad  = ~n1360 ;
  assign \847(465)_pad  = ~n1361 ;
  assign \848(330)_pad  = ~\245(98)_pad  ;
  assign \849(219)_pad  = ~\552(152)_pad  ;
  assign \850(217)_pad  = ~\562(155)_pad  ;
  assign \851(218)_pad  = ~\559(154)_pad  ;
  assign \854(2268)_pad  = n1398 ;
  assign \859(2132)_pad  = ~n1405 ;
  assign \861(2070)_pad  = n992 ;
  assign \863(2276)_pad  = n658 ;
  assign \865(2277)_pad  = n619 ;
  assign \867(2237)_pad  = n580 ;
  assign \869(2181)_pad  = n544 ;
  assign \871(2127)_pad  = n502 ;
  assign \873(2124)_pad  = n1099 ;
  assign \875(2125)_pad  = n1064 ;
  assign \877(2126)_pad  = n1028 ;
  assign \882(2456)_pad  = ~n1410 ;
  assign \998(2163)_pad  = ~n1391 ;
  assign \u2023_syn_3  = n1424 ;
  assign \u2095_syn_3  = n1432 ;
  assign \u2109_syn_3  = n1440 ;
  assign \u2318_syn_3  = ~n666 ;
  assign \u3086_syn_3  = n1448 ;
endmodule
