module top( \C_0_pad  , \C_10_pad  , \C_11_pad  , \C_12_pad  , \C_13_pad  , \C_14_pad  , \C_15_pad  , \C_16_pad  , \C_17_pad  , \C_18_pad  , \C_19_pad  , \C_1_pad  , \C_20_pad  , \C_21_pad  , \C_22_pad  , \C_23_pad  , \C_24_pad  , \C_25_pad  , \C_26_pad  , \C_27_pad  , \C_28_pad  , \C_29_pad  , \C_2_pad  , \C_30_pad  , \C_31_pad  , \C_32_pad  , \C_3_pad  , \C_4_pad  , \C_5_pad  , \C_6_pad  , \C_7_pad  , \C_8_pad  , \C_9_pad  , \P_0_pad  , \X_10_reg/NET0131  , \X_11_reg/NET0131  , \X_12_reg/NET0131  , \X_13_reg/NET0131  , \X_14_reg/NET0131  , \X_15_reg/NET0131  , \X_16_reg/NET0131  , \X_17_reg/NET0131  , \X_18_reg/NET0131  , \X_19_reg/NET0131  , \X_1_reg/NET0131  , \X_20_reg/NET0131  , \X_21_reg/NET0131  , \X_22_reg/NET0131  , \X_23_reg/NET0131  , \X_24_reg/NET0131  , \X_25_reg/NET0131  , \X_26_reg/NET0131  , \X_27_reg/NET0131  , \X_28_reg/NET0131  , \X_29_reg/NET0131  , \X_2_reg/NET0131  , \X_30_reg/P0002  , \X_31_reg/P0002  , \X_32_reg/P0002  , \X_3_reg/NET0131  , \X_4_reg/NET0131  , \X_5_reg/NET0131  , \X_6_reg/NET0131  , \X_7_reg/NET0131  , \X_8_reg/NET0131  , \X_9_reg/NET0131  , \X_30_reg/P0000  , \X_31_reg/P0000  , \X_32_reg/P0000  , Z_pad , \_al_n0  , \_al_n1  , \g1375/_1_  , \g1387/_0_  , \g1398/_0_  , \g1400/_0_  , \g1419/_0_  , \g1433/_0_  , \g1443/_0_  , \g1457/_0_  , \g1458/_0_  , \g1468/_0_  , \g1483/_0_  , \g1486/_0_  , \g1493/_0_  , \g1504/_0_  , \g1505/_0_  , \g1512/_0_  , \g1525/_0_  , \g1535/_0_  , \g1544/_0_  , \g1565/_0_  , \g1871/_0_  , \g1900/_0_  , \g1955/_0_  , \g1961/_0_  , \g1991/_0_  , \g2026/_0_  , \g2040/_0_  , \g2046/_0_  , \g2051/_1_  , \g2098/_0_  , \g21/_0_  , \g2101/_0_  );
  input \C_0_pad  ;
  input \C_10_pad  ;
  input \C_11_pad  ;
  input \C_12_pad  ;
  input \C_13_pad  ;
  input \C_14_pad  ;
  input \C_15_pad  ;
  input \C_16_pad  ;
  input \C_17_pad  ;
  input \C_18_pad  ;
  input \C_19_pad  ;
  input \C_1_pad  ;
  input \C_20_pad  ;
  input \C_21_pad  ;
  input \C_22_pad  ;
  input \C_23_pad  ;
  input \C_24_pad  ;
  input \C_25_pad  ;
  input \C_26_pad  ;
  input \C_27_pad  ;
  input \C_28_pad  ;
  input \C_29_pad  ;
  input \C_2_pad  ;
  input \C_30_pad  ;
  input \C_31_pad  ;
  input \C_32_pad  ;
  input \C_3_pad  ;
  input \C_4_pad  ;
  input \C_5_pad  ;
  input \C_6_pad  ;
  input \C_7_pad  ;
  input \C_8_pad  ;
  input \C_9_pad  ;
  input \P_0_pad  ;
  input \X_10_reg/NET0131  ;
  input \X_11_reg/NET0131  ;
  input \X_12_reg/NET0131  ;
  input \X_13_reg/NET0131  ;
  input \X_14_reg/NET0131  ;
  input \X_15_reg/NET0131  ;
  input \X_16_reg/NET0131  ;
  input \X_17_reg/NET0131  ;
  input \X_18_reg/NET0131  ;
  input \X_19_reg/NET0131  ;
  input \X_1_reg/NET0131  ;
  input \X_20_reg/NET0131  ;
  input \X_21_reg/NET0131  ;
  input \X_22_reg/NET0131  ;
  input \X_23_reg/NET0131  ;
  input \X_24_reg/NET0131  ;
  input \X_25_reg/NET0131  ;
  input \X_26_reg/NET0131  ;
  input \X_27_reg/NET0131  ;
  input \X_28_reg/NET0131  ;
  input \X_29_reg/NET0131  ;
  input \X_2_reg/NET0131  ;
  input \X_30_reg/P0002  ;
  input \X_31_reg/P0002  ;
  input \X_32_reg/P0002  ;
  input \X_3_reg/NET0131  ;
  input \X_4_reg/NET0131  ;
  input \X_5_reg/NET0131  ;
  input \X_6_reg/NET0131  ;
  input \X_7_reg/NET0131  ;
  input \X_8_reg/NET0131  ;
  input \X_9_reg/NET0131  ;
  output \X_30_reg/P0000  ;
  output \X_31_reg/P0000  ;
  output \X_32_reg/P0000  ;
  output Z_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1375/_1_  ;
  output \g1387/_0_  ;
  output \g1398/_0_  ;
  output \g1400/_0_  ;
  output \g1419/_0_  ;
  output \g1433/_0_  ;
  output \g1443/_0_  ;
  output \g1457/_0_  ;
  output \g1458/_0_  ;
  output \g1468/_0_  ;
  output \g1483/_0_  ;
  output \g1486/_0_  ;
  output \g1493/_0_  ;
  output \g1504/_0_  ;
  output \g1505/_0_  ;
  output \g1512/_0_  ;
  output \g1525/_0_  ;
  output \g1535/_0_  ;
  output \g1544/_0_  ;
  output \g1565/_0_  ;
  output \g1871/_0_  ;
  output \g1900/_0_  ;
  output \g1955/_0_  ;
  output \g1961/_0_  ;
  output \g1991/_0_  ;
  output \g2026/_0_  ;
  output \g2040/_0_  ;
  output \g2046/_0_  ;
  output \g2051/_1_  ;
  output \g2098/_0_  ;
  output \g21/_0_  ;
  output \g2101/_0_  ;
  wire n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 ;
  assign n72 = ~\X_7_reg/NET0131  & ~\X_8_reg/NET0131  ;
  assign n73 = ~\X_4_reg/NET0131  & ~\X_5_reg/NET0131  ;
  assign n74 = ~\X_6_reg/NET0131  & n73 ;
  assign n75 = n72 & n74 ;
  assign n93 = ~\X_20_reg/NET0131  & ~\X_2_reg/NET0131  ;
  assign n94 = ~\X_3_reg/NET0131  & n93 ;
  assign n91 = ~\X_17_reg/NET0131  & ~\X_18_reg/NET0131  ;
  assign n92 = ~\X_19_reg/NET0131  & ~\X_1_reg/NET0131  ;
  assign n95 = n91 & n92 ;
  assign n96 = n94 & n95 ;
  assign n67 = ~\X_10_reg/NET0131  & ~\X_9_reg/NET0131  ;
  assign n68 = ~\X_11_reg/NET0131  & ~\X_12_reg/NET0131  ;
  assign n69 = n67 & n68 ;
  assign n88 = ~\X_13_reg/NET0131  & ~\X_14_reg/NET0131  ;
  assign n89 = ~\X_15_reg/NET0131  & ~\X_16_reg/NET0131  ;
  assign n90 = n88 & n89 ;
  assign n97 = n69 & n90 ;
  assign n98 = n96 & n97 ;
  assign n99 = n75 & n98 ;
  assign n100 = ~\C_21_pad  & \X_21_reg/NET0131  ;
  assign n102 = \C_23_pad  & ~\X_22_reg/NET0131  ;
  assign n103 = \X_23_reg/NET0131  & n102 ;
  assign n101 = \C_22_pad  & \X_22_reg/NET0131  ;
  assign n104 = ~\X_21_reg/NET0131  & ~n101 ;
  assign n105 = ~n103 & n104 ;
  assign n106 = ~n100 & ~n105 ;
  assign n107 = n99 & n106 ;
  assign n70 = ~\X_1_reg/NET0131  & ~\X_2_reg/NET0131  ;
  assign n71 = ~\X_3_reg/NET0131  & n70 ;
  assign n76 = n71 & n75 ;
  assign n77 = \C_14_pad  & \X_14_reg/NET0131  ;
  assign n78 = \C_16_pad  & ~\X_14_reg/NET0131  ;
  assign n79 = ~\X_15_reg/NET0131  & \X_16_reg/NET0131  ;
  assign n80 = n78 & n79 ;
  assign n81 = ~n77 & ~n80 ;
  assign n82 = ~\X_13_reg/NET0131  & n69 ;
  assign n83 = ~n81 & n82 ;
  assign n84 = n76 & n83 ;
  assign n85 = ~\X_4_reg/NET0131  & n71 ;
  assign n86 = \C_5_pad  & \X_5_reg/NET0131  ;
  assign n87 = n85 & n86 ;
  assign n108 = ~\C_0_pad  & ~n87 ;
  assign n109 = ~n84 & n108 ;
  assign n110 = ~n107 & n109 ;
  assign n111 = \P_0_pad  & ~n110 ;
  assign n165 = ~\X_21_reg/NET0131  & ~\X_22_reg/NET0131  ;
  assign n166 = n99 & n165 ;
  assign n167 = \C_24_pad  & \P_0_pad  ;
  assign n168 = ~\X_23_reg/NET0131  & \X_24_reg/NET0131  ;
  assign n169 = n167 & n168 ;
  assign n170 = n166 & n169 ;
  assign n129 = \P_0_pad  & n76 ;
  assign n132 = \C_11_pad  & \X_11_reg/NET0131  ;
  assign n133 = \C_12_pad  & ~\X_11_reg/NET0131  ;
  assign n134 = \X_12_reg/NET0131  & n133 ;
  assign n135 = ~n132 & ~n134 ;
  assign n136 = n67 & ~n135 ;
  assign n137 = \C_9_pad  & \X_9_reg/NET0131  ;
  assign n138 = \C_10_pad  & \X_10_reg/NET0131  ;
  assign n139 = ~\X_9_reg/NET0131  & n138 ;
  assign n140 = ~n137 & ~n139 ;
  assign n141 = ~n136 & n140 ;
  assign n142 = n129 & ~n141 ;
  assign n156 = \C_8_pad  & ~\X_7_reg/NET0131  ;
  assign n157 = \X_8_reg/NET0131  & n156 ;
  assign n158 = \C_7_pad  & \X_7_reg/NET0131  ;
  assign n159 = ~\X_6_reg/NET0131  & ~n158 ;
  assign n160 = ~n157 & n159 ;
  assign n155 = ~\C_6_pad  & \X_6_reg/NET0131  ;
  assign n161 = \P_0_pad  & ~\X_5_reg/NET0131  ;
  assign n162 = ~n155 & n161 ;
  assign n163 = n85 & n162 ;
  assign n164 = ~n160 & n163 ;
  assign n143 = \P_0_pad  & ~\X_1_reg/NET0131  ;
  assign n144 = \C_2_pad  & \X_2_reg/NET0131  ;
  assign n145 = \C_4_pad  & ~\X_2_reg/NET0131  ;
  assign n146 = ~\X_3_reg/NET0131  & \X_4_reg/NET0131  ;
  assign n147 = n145 & n146 ;
  assign n148 = ~n144 & ~n147 ;
  assign n149 = n143 & ~n148 ;
  assign n150 = \P_0_pad  & \X_1_reg/NET0131  ;
  assign n151 = \C_1_pad  & n150 ;
  assign n152 = \C_3_pad  & ~\X_2_reg/NET0131  ;
  assign n153 = \X_3_reg/NET0131  & n152 ;
  assign n154 = n143 & n153 ;
  assign n201 = ~n151 & ~n154 ;
  assign n202 = ~n149 & n201 ;
  assign n203 = ~n164 & n202 ;
  assign n204 = ~n142 & n203 ;
  assign n205 = ~n170 & n204 ;
  assign n206 = ~n111 & n205 ;
  assign n112 = \C_17_pad  & \X_17_reg/NET0131  ;
  assign n113 = \C_19_pad  & \X_19_reg/NET0131  ;
  assign n114 = \C_20_pad  & ~\X_19_reg/NET0131  ;
  assign n115 = \X_20_reg/NET0131  & n114 ;
  assign n116 = ~n113 & ~n115 ;
  assign n117 = n91 & ~n116 ;
  assign n118 = ~n112 & ~n117 ;
  assign n119 = n90 & ~n118 ;
  assign n123 = \C_18_pad  & ~\X_17_reg/NET0131  ;
  assign n124 = \X_18_reg/NET0131  & n123 ;
  assign n125 = n90 & n124 ;
  assign n120 = \C_13_pad  & \X_13_reg/NET0131  ;
  assign n121 = \C_15_pad  & \X_15_reg/NET0131  ;
  assign n122 = n88 & n121 ;
  assign n126 = ~n120 & ~n122 ;
  assign n127 = ~n125 & n126 ;
  assign n128 = ~n119 & n127 ;
  assign n130 = n69 & n129 ;
  assign n131 = ~n128 & n130 ;
  assign n171 = \C_25_pad  & \X_25_reg/NET0131  ;
  assign n173 = \C_28_pad  & ~\X_27_reg/NET0131  ;
  assign n174 = \X_28_reg/NET0131  & n173 ;
  assign n175 = \C_27_pad  & \X_27_reg/NET0131  ;
  assign n176 = ~\X_26_reg/NET0131  & ~n175 ;
  assign n177 = ~n174 & n176 ;
  assign n172 = ~\C_26_pad  & \X_26_reg/NET0131  ;
  assign n178 = ~\X_25_reg/NET0131  & ~n172 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = ~n171 & ~n179 ;
  assign n181 = \P_0_pad  & ~n180 ;
  assign n183 = \C_31_pad  & \X_31_reg/P0002  ;
  assign n184 = \C_32_pad  & ~\X_31_reg/P0002  ;
  assign n185 = \X_32_reg/P0002  & n184 ;
  assign n186 = ~n183 & ~n185 ;
  assign n187 = ~\X_30_reg/P0002  & ~n186 ;
  assign n182 = \C_30_pad  & \X_30_reg/P0002  ;
  assign n188 = ~\X_29_reg/NET0131  & ~n182 ;
  assign n189 = ~n187 & n188 ;
  assign n192 = ~\X_26_reg/NET0131  & ~\X_27_reg/NET0131  ;
  assign n193 = ~\X_28_reg/NET0131  & n192 ;
  assign n190 = ~\C_29_pad  & \X_29_reg/NET0131  ;
  assign n191 = \P_0_pad  & ~\X_25_reg/NET0131  ;
  assign n194 = ~n190 & n191 ;
  assign n195 = n193 & n194 ;
  assign n196 = ~n189 & n195 ;
  assign n197 = ~n181 & ~n196 ;
  assign n198 = ~\X_23_reg/NET0131  & ~\X_24_reg/NET0131  ;
  assign n199 = n166 & n198 ;
  assign n200 = ~n197 & n199 ;
  assign n207 = ~n131 & ~n200 ;
  assign n208 = n206 & n207 ;
  assign n209 = \X_7_reg/NET0131  & \X_8_reg/NET0131  ;
  assign n210 = \X_10_reg/NET0131  & \X_9_reg/NET0131  ;
  assign n211 = n209 & n210 ;
  assign n212 = \X_11_reg/NET0131  & \X_12_reg/NET0131  ;
  assign n213 = \X_5_reg/NET0131  & \X_6_reg/NET0131  ;
  assign n214 = n212 & n213 ;
  assign n215 = n211 & n214 ;
  assign n216 = \X_14_reg/NET0131  & \X_15_reg/NET0131  ;
  assign n217 = \X_16_reg/NET0131  & n216 ;
  assign n220 = \X_20_reg/NET0131  & \X_3_reg/NET0131  ;
  assign n221 = \X_4_reg/NET0131  & n220 ;
  assign n218 = \X_17_reg/NET0131  & \X_18_reg/NET0131  ;
  assign n219 = \X_19_reg/NET0131  & \X_1_reg/NET0131  ;
  assign n222 = n218 & n219 ;
  assign n223 = n221 & n222 ;
  assign n224 = n217 & n223 ;
  assign n225 = n215 & n224 ;
  assign n228 = \X_21_reg/NET0131  & \X_22_reg/NET0131  ;
  assign n229 = \X_23_reg/NET0131  & n228 ;
  assign n230 = \X_24_reg/NET0131  & n229 ;
  assign n226 = \P_0_pad  & \X_13_reg/NET0131  ;
  assign n227 = \X_2_reg/NET0131  & n226 ;
  assign n231 = \X_25_reg/NET0131  & n227 ;
  assign n232 = n230 & n231 ;
  assign n233 = n225 & n232 ;
  assign n234 = \X_26_reg/NET0131  & n233 ;
  assign n235 = \X_27_reg/NET0131  & \X_28_reg/NET0131  ;
  assign n236 = n234 & n235 ;
  assign n237 = \X_29_reg/NET0131  & n236 ;
  assign n238 = \X_30_reg/P0002  & n237 ;
  assign n239 = \X_31_reg/P0002  & n238 ;
  assign n240 = ~\X_26_reg/NET0131  & ~n233 ;
  assign n241 = ~n234 & ~n240 ;
  assign n242 = n225 & n227 ;
  assign n243 = \X_21_reg/NET0131  & n242 ;
  assign n244 = ~\X_22_reg/NET0131  & ~n243 ;
  assign n245 = n228 & n242 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = \X_27_reg/NET0131  & n234 ;
  assign n248 = ~\X_27_reg/NET0131  & ~n234 ;
  assign n249 = ~n247 & ~n248 ;
  assign n250 = ~\X_23_reg/NET0131  & ~n245 ;
  assign n251 = n229 & n242 ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = ~\X_21_reg/NET0131  & ~n242 ;
  assign n254 = ~n243 & ~n253 ;
  assign n255 = \X_2_reg/NET0131  & n150 ;
  assign n256 = \X_3_reg/NET0131  & n255 ;
  assign n257 = \X_4_reg/NET0131  & n256 ;
  assign n258 = n215 & n257 ;
  assign n259 = \X_13_reg/NET0131  & n258 ;
  assign n260 = n217 & n259 ;
  assign n261 = n218 & n260 ;
  assign n262 = \X_19_reg/NET0131  & n261 ;
  assign n263 = ~\X_19_reg/NET0131  & ~n261 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = \X_5_reg/NET0131  & n257 ;
  assign n266 = \X_6_reg/NET0131  & n265 ;
  assign n267 = n211 & n266 ;
  assign n268 = \X_11_reg/NET0131  & n267 ;
  assign n269 = ~\X_12_reg/NET0131  & ~n268 ;
  assign n270 = ~n258 & ~n269 ;
  assign n271 = \X_17_reg/NET0131  & n260 ;
  assign n272 = ~\X_17_reg/NET0131  & ~n260 ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = \X_14_reg/NET0131  & n259 ;
  assign n275 = ~\X_15_reg/NET0131  & ~n274 ;
  assign n276 = \X_15_reg/NET0131  & n274 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = ~\X_13_reg/NET0131  & ~n258 ;
  assign n279 = ~n259 & ~n278 ;
  assign n280 = ~\X_6_reg/NET0131  & ~n265 ;
  assign n281 = ~n266 & ~n280 ;
  assign n282 = ~\X_11_reg/NET0131  & ~n267 ;
  assign n283 = ~n268 & ~n282 ;
  assign n284 = ~\X_4_reg/NET0131  & ~n256 ;
  assign n285 = ~n257 & ~n284 ;
  assign n286 = n209 & n266 ;
  assign n287 = \X_9_reg/NET0131  & n286 ;
  assign n288 = ~\X_9_reg/NET0131  & ~n286 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = ~\X_7_reg/NET0131  & n266 ;
  assign n291 = \X_7_reg/NET0131  & ~n266 ;
  assign n292 = ~n290 & ~n291 ;
  assign n293 = ~\X_5_reg/NET0131  & ~n257 ;
  assign n294 = ~n265 & ~n293 ;
  assign n295 = ~\X_3_reg/NET0131  & ~n255 ;
  assign n296 = ~n256 & ~n295 ;
  assign n297 = ~\X_2_reg/NET0131  & ~n150 ;
  assign n298 = ~n255 & ~n297 ;
  assign n299 = ~\P_0_pad  & \X_1_reg/NET0131  ;
  assign n300 = ~n143 & ~n299 ;
  assign n301 = \X_20_reg/NET0131  & ~n262 ;
  assign n302 = ~\X_20_reg/NET0131  & n262 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = ~\X_14_reg/NET0131  & ~n259 ;
  assign n305 = ~n274 & ~n304 ;
  assign n306 = ~\X_18_reg/NET0131  & ~n271 ;
  assign n307 = ~n261 & ~n306 ;
  assign n308 = ~\X_24_reg/NET0131  & ~n251 ;
  assign n309 = n230 & n242 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = ~\X_25_reg/NET0131  & ~n309 ;
  assign n312 = ~n233 & ~n311 ;
  assign n313 = ~\X_29_reg/NET0131  & ~n236 ;
  assign n314 = ~n237 & ~n313 ;
  assign n315 = ~n72 & ~n209 ;
  assign n316 = ~n291 & ~n315 ;
  assign n317 = n291 & n315 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = ~\X_28_reg/NET0131  & ~n247 ;
  assign n320 = ~n236 & ~n319 ;
  assign n321 = ~\X_16_reg/NET0131  & ~n276 ;
  assign n322 = ~n260 & ~n321 ;
  assign n323 = ~\X_10_reg/NET0131  & ~n287 ;
  assign n324 = ~n267 & ~n323 ;
  assign \X_30_reg/P0000  = ~\X_30_reg/P0002  ;
  assign \X_31_reg/P0000  = ~\X_31_reg/P0002  ;
  assign \X_32_reg/P0000  = ~\X_32_reg/P0002  ;
  assign Z_pad = ~n208 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1375/_1_  = n239 ;
  assign \g1387/_0_  = n241 ;
  assign \g1398/_0_  = n246 ;
  assign \g1400/_0_  = n249 ;
  assign \g1419/_0_  = n252 ;
  assign \g1433/_0_  = n254 ;
  assign \g1443/_0_  = n264 ;
  assign \g1457/_0_  = n270 ;
  assign \g1458/_0_  = n273 ;
  assign \g1468/_0_  = n277 ;
  assign \g1483/_0_  = n279 ;
  assign \g1486/_0_  = n281 ;
  assign \g1493/_0_  = n283 ;
  assign \g1504/_0_  = n285 ;
  assign \g1505/_0_  = n289 ;
  assign \g1512/_0_  = ~n292 ;
  assign \g1525/_0_  = n294 ;
  assign \g1535/_0_  = n296 ;
  assign \g1544/_0_  = n298 ;
  assign \g1565/_0_  = ~n300 ;
  assign \g1871/_0_  = ~n303 ;
  assign \g1900/_0_  = n305 ;
  assign \g1955/_0_  = n307 ;
  assign \g1961/_0_  = n310 ;
  assign \g1991/_0_  = n312 ;
  assign \g2026/_0_  = n314 ;
  assign \g2040/_0_  = n318 ;
  assign \g2046/_0_  = n238 ;
  assign \g2051/_1_  = n237 ;
  assign \g2098/_0_  = n320 ;
  assign \g21/_0_  = n322 ;
  assign \g2101/_0_  = n324 ;
endmodule
