module top( \P1_B_reg/NET0131  , \P1_IR_reg[0]/NET0131  , \P1_IR_reg[10]/NET0131  , \P1_IR_reg[11]/NET0131  , \P1_IR_reg[12]/NET0131  , \P1_IR_reg[13]/NET0131  , \P1_IR_reg[14]/NET0131  , \P1_IR_reg[15]/NET0131  , \P1_IR_reg[16]/NET0131  , \P1_IR_reg[17]/NET0131  , \P1_IR_reg[18]/NET0131  , \P1_IR_reg[19]/NET0131  , \P1_IR_reg[1]/NET0131  , \P1_IR_reg[20]/NET0131  , \P1_IR_reg[21]/NET0131  , \P1_IR_reg[22]/NET0131  , \P1_IR_reg[23]/NET0131  , \P1_IR_reg[24]/NET0131  , \P1_IR_reg[25]/NET0131  , \P1_IR_reg[26]/NET0131  , \P1_IR_reg[27]/NET0131  , \P1_IR_reg[28]/NET0131  , \P1_IR_reg[29]/NET0131  , \P1_IR_reg[2]/NET0131  , \P1_IR_reg[30]/NET0131  , \P1_IR_reg[31]/NET0131  , \P1_IR_reg[3]/NET0131  , \P1_IR_reg[4]/NET0131  , \P1_IR_reg[5]/NET0131  , \P1_IR_reg[6]/NET0131  , \P1_IR_reg[7]/NET0131  , \P1_IR_reg[8]/NET0131  , \P1_IR_reg[9]/NET0131  , \P1_addr_reg[0]/NET0131  , \P1_addr_reg[10]/NET0131  , \P1_addr_reg[11]/NET0131  , \P1_addr_reg[12]/NET0131  , \P1_addr_reg[13]/NET0131  , \P1_addr_reg[14]/NET0131  , \P1_addr_reg[15]/NET0131  , \P1_addr_reg[16]/NET0131  , \P1_addr_reg[17]/NET0131  , \P1_addr_reg[18]/NET0131  , \P1_addr_reg[19]/NET0131  , \P1_addr_reg[1]/NET0131  , \P1_addr_reg[2]/NET0131  , \P1_addr_reg[3]/NET0131  , \P1_addr_reg[4]/NET0131  , \P1_addr_reg[5]/NET0131  , \P1_addr_reg[6]/NET0131  , \P1_addr_reg[7]/NET0131  , \P1_addr_reg[8]/NET0131  , \P1_addr_reg[9]/NET0131  , \P1_d_reg[0]/NET0131  , \P1_d_reg[1]/NET0131  , \P1_datao_reg[0]/NET0131  , \P1_datao_reg[10]/NET0131  , \P1_datao_reg[11]/NET0131  , \P1_datao_reg[12]/NET0131  , \P1_datao_reg[13]/NET0131  , \P1_datao_reg[14]/NET0131  , \P1_datao_reg[15]/NET0131  , \P1_datao_reg[16]/NET0131  , \P1_datao_reg[17]/NET0131  , \P1_datao_reg[18]/NET0131  , \P1_datao_reg[19]/NET0131  , \P1_datao_reg[1]/NET0131  , \P1_datao_reg[20]/NET0131  , \P1_datao_reg[21]/NET0131  , \P1_datao_reg[22]/NET0131  , \P1_datao_reg[23]/NET0131  , \P1_datao_reg[24]/NET0131  , \P1_datao_reg[25]/NET0131  , \P1_datao_reg[26]/NET0131  , \P1_datao_reg[27]/NET0131  , \P1_datao_reg[28]/NET0131  , \P1_datao_reg[29]/NET0131  , \P1_datao_reg[2]/NET0131  , \P1_datao_reg[30]/NET0131  , \P1_datao_reg[31]/NET0131  , \P1_datao_reg[3]/NET0131  , \P1_datao_reg[4]/NET0131  , \P1_datao_reg[5]/NET0131  , \P1_datao_reg[6]/NET0131  , \P1_datao_reg[7]/NET0131  , \P1_datao_reg[8]/NET0131  , \P1_datao_reg[9]/NET0131  , \P1_rd_reg/NET0131  , \P1_reg0_reg[0]/NET0131  , \P1_reg0_reg[10]/NET0131  , \P1_reg0_reg[11]/NET0131  , \P1_reg0_reg[12]/NET0131  , \P1_reg0_reg[13]/NET0131  , \P1_reg0_reg[14]/NET0131  , \P1_reg0_reg[15]/NET0131  , \P1_reg0_reg[16]/NET0131  , \P1_reg0_reg[17]/NET0131  , \P1_reg0_reg[18]/NET0131  , \P1_reg0_reg[19]/NET0131  , \P1_reg0_reg[1]/NET0131  , \P1_reg0_reg[20]/NET0131  , \P1_reg0_reg[21]/NET0131  , \P1_reg0_reg[22]/NET0131  , \P1_reg0_reg[23]/NET0131  , \P1_reg0_reg[24]/NET0131  , \P1_reg0_reg[25]/NET0131  , \P1_reg0_reg[26]/NET0131  , \P1_reg0_reg[27]/NET0131  , \P1_reg0_reg[28]/NET0131  , \P1_reg0_reg[29]/NET0131  , \P1_reg0_reg[2]/NET0131  , \P1_reg0_reg[30]/NET0131  , \P1_reg0_reg[31]/NET0131  , \P1_reg0_reg[3]/NET0131  , \P1_reg0_reg[4]/NET0131  , \P1_reg0_reg[5]/NET0131  , \P1_reg0_reg[6]/NET0131  , \P1_reg0_reg[7]/NET0131  , \P1_reg0_reg[8]/NET0131  , \P1_reg0_reg[9]/NET0131  , \P1_reg1_reg[0]/NET0131  , \P1_reg1_reg[10]/NET0131  , \P1_reg1_reg[11]/NET0131  , \P1_reg1_reg[12]/NET0131  , \P1_reg1_reg[13]/NET0131  , \P1_reg1_reg[14]/NET0131  , \P1_reg1_reg[15]/NET0131  , \P1_reg1_reg[16]/NET0131  , \P1_reg1_reg[17]/NET0131  , \P1_reg1_reg[18]/NET0131  , \P1_reg1_reg[19]/NET0131  , \P1_reg1_reg[1]/NET0131  , \P1_reg1_reg[20]/NET0131  , \P1_reg1_reg[21]/NET0131  , \P1_reg1_reg[22]/NET0131  , \P1_reg1_reg[23]/NET0131  , \P1_reg1_reg[24]/NET0131  , \P1_reg1_reg[25]/NET0131  , \P1_reg1_reg[26]/NET0131  , \P1_reg1_reg[27]/NET0131  , \P1_reg1_reg[28]/NET0131  , \P1_reg1_reg[29]/NET0131  , \P1_reg1_reg[2]/NET0131  , \P1_reg1_reg[30]/NET0131  , \P1_reg1_reg[31]/NET0131  , \P1_reg1_reg[3]/NET0131  , \P1_reg1_reg[4]/NET0131  , \P1_reg1_reg[5]/NET0131  , \P1_reg1_reg[6]/NET0131  , \P1_reg1_reg[7]/NET0131  , \P1_reg1_reg[8]/NET0131  , \P1_reg1_reg[9]/NET0131  , \P1_reg2_reg[0]/NET0131  , \P1_reg2_reg[10]/NET0131  , \P1_reg2_reg[11]/NET0131  , \P1_reg2_reg[12]/NET0131  , \P1_reg2_reg[13]/NET0131  , \P1_reg2_reg[14]/NET0131  , \P1_reg2_reg[15]/NET0131  , \P1_reg2_reg[16]/NET0131  , \P1_reg2_reg[17]/NET0131  , \P1_reg2_reg[18]/NET0131  , \P1_reg2_reg[19]/NET0131  , \P1_reg2_reg[1]/NET0131  , \P1_reg2_reg[20]/NET0131  , \P1_reg2_reg[21]/NET0131  , \P1_reg2_reg[22]/NET0131  , \P1_reg2_reg[23]/NET0131  , \P1_reg2_reg[24]/NET0131  , \P1_reg2_reg[25]/NET0131  , \P1_reg2_reg[26]/NET0131  , \P1_reg2_reg[27]/NET0131  , \P1_reg2_reg[28]/NET0131  , \P1_reg2_reg[29]/NET0131  , \P1_reg2_reg[2]/NET0131  , \P1_reg2_reg[30]/NET0131  , \P1_reg2_reg[31]/NET0131  , \P1_reg2_reg[3]/NET0131  , \P1_reg2_reg[4]/NET0131  , \P1_reg2_reg[5]/NET0131  , \P1_reg2_reg[6]/NET0131  , \P1_reg2_reg[7]/NET0131  , \P1_reg2_reg[8]/NET0131  , \P1_reg2_reg[9]/NET0131  , \P1_reg3_reg[0]/NET0131  , \P1_reg3_reg[10]/NET0131  , \P1_reg3_reg[11]/NET0131  , \P1_reg3_reg[12]/NET0131  , \P1_reg3_reg[13]/NET0131  , \P1_reg3_reg[14]/NET0131  , \P1_reg3_reg[15]/NET0131  , \P1_reg3_reg[16]/NET0131  , \P1_reg3_reg[17]/NET0131  , \P1_reg3_reg[18]/NET0131  , \P1_reg3_reg[19]/NET0131  , \P1_reg3_reg[1]/NET0131  , \P1_reg3_reg[20]/NET0131  , \P1_reg3_reg[21]/NET0131  , \P1_reg3_reg[22]/NET0131  , \P1_reg3_reg[23]/NET0131  , \P1_reg3_reg[24]/NET0131  , \P1_reg3_reg[25]/NET0131  , \P1_reg3_reg[26]/NET0131  , \P1_reg3_reg[27]/NET0131  , \P1_reg3_reg[28]/NET0131  , \P1_reg3_reg[2]/NET0131  , \P1_reg3_reg[3]/NET0131  , \P1_reg3_reg[4]/NET0131  , \P1_reg3_reg[5]/NET0131  , \P1_reg3_reg[6]/NET0131  , \P1_reg3_reg[7]/NET0131  , \P1_reg3_reg[8]/NET0131  , \P1_reg3_reg[9]/NET0131  , \P1_state_reg[0]/NET0131  , \P1_wr_reg/NET0131  , \P2_B_reg/NET0131  , \P2_IR_reg[0]/NET0131  , \P2_IR_reg[10]/NET0131  , \P2_IR_reg[11]/NET0131  , \P2_IR_reg[12]/NET0131  , \P2_IR_reg[13]/NET0131  , \P2_IR_reg[14]/NET0131  , \P2_IR_reg[15]/NET0131  , \P2_IR_reg[16]/NET0131  , \P2_IR_reg[17]/NET0131  , \P2_IR_reg[18]/NET0131  , \P2_IR_reg[19]/NET0131  , \P2_IR_reg[1]/NET0131  , \P2_IR_reg[20]/NET0131  , \P2_IR_reg[21]/NET0131  , \P2_IR_reg[22]/NET0131  , \P2_IR_reg[23]/NET0131  , \P2_IR_reg[24]/NET0131  , \P2_IR_reg[25]/NET0131  , \P2_IR_reg[26]/NET0131  , \P2_IR_reg[27]/NET0131  , \P2_IR_reg[28]/NET0131  , \P2_IR_reg[29]/NET0131  , \P2_IR_reg[2]/NET0131  , \P2_IR_reg[30]/NET0131  , \P2_IR_reg[31]/NET0131  , \P2_IR_reg[3]/NET0131  , \P2_IR_reg[4]/NET0131  , \P2_IR_reg[5]/NET0131  , \P2_IR_reg[6]/NET0131  , \P2_IR_reg[7]/NET0131  , \P2_IR_reg[8]/NET0131  , \P2_IR_reg[9]/NET0131  , \P2_addr_reg[0]/NET0131  , \P2_addr_reg[10]/NET0131  , \P2_addr_reg[11]/NET0131  , \P2_addr_reg[12]/NET0131  , \P2_addr_reg[13]/NET0131  , \P2_addr_reg[14]/NET0131  , \P2_addr_reg[15]/NET0131  , \P2_addr_reg[16]/NET0131  , \P2_addr_reg[17]/NET0131  , \P2_addr_reg[18]/NET0131  , \P2_addr_reg[19]/NET0131  , \P2_addr_reg[1]/NET0131  , \P2_addr_reg[2]/NET0131  , \P2_addr_reg[3]/NET0131  , \P2_addr_reg[4]/NET0131  , \P2_addr_reg[5]/NET0131  , \P2_addr_reg[6]/NET0131  , \P2_addr_reg[7]/NET0131  , \P2_addr_reg[8]/NET0131  , \P2_addr_reg[9]/NET0131  , \P2_d_reg[0]/NET0131  , \P2_d_reg[1]/NET0131  , \P2_datao_reg[0]/NET0131  , \P2_datao_reg[10]/NET0131  , \P2_datao_reg[11]/NET0131  , \P2_datao_reg[12]/NET0131  , \P2_datao_reg[13]/NET0131  , \P2_datao_reg[14]/NET0131  , \P2_datao_reg[15]/NET0131  , \P2_datao_reg[16]/NET0131  , \P2_datao_reg[17]/NET0131  , \P2_datao_reg[18]/NET0131  , \P2_datao_reg[19]/NET0131  , \P2_datao_reg[1]/NET0131  , \P2_datao_reg[20]/NET0131  , \P2_datao_reg[21]/NET0131  , \P2_datao_reg[22]/NET0131  , \P2_datao_reg[23]/NET0131  , \P2_datao_reg[24]/NET0131  , \P2_datao_reg[25]/NET0131  , \P2_datao_reg[26]/NET0131  , \P2_datao_reg[27]/NET0131  , \P2_datao_reg[28]/NET0131  , \P2_datao_reg[29]/NET0131  , \P2_datao_reg[2]/NET0131  , \P2_datao_reg[30]/NET0131  , \P2_datao_reg[31]/NET0131  , \P2_datao_reg[3]/NET0131  , \P2_datao_reg[4]/NET0131  , \P2_datao_reg[5]/NET0131  , \P2_datao_reg[6]/NET0131  , \P2_datao_reg[7]/NET0131  , \P2_datao_reg[8]/NET0131  , \P2_datao_reg[9]/NET0131  , \P2_rd_reg/NET0131  , \P2_reg0_reg[0]/NET0131  , \P2_reg0_reg[10]/NET0131  , \P2_reg0_reg[11]/NET0131  , \P2_reg0_reg[12]/NET0131  , \P2_reg0_reg[13]/NET0131  , \P2_reg0_reg[14]/NET0131  , \P2_reg0_reg[15]/NET0131  , \P2_reg0_reg[16]/NET0131  , \P2_reg0_reg[17]/NET0131  , \P2_reg0_reg[18]/NET0131  , \P2_reg0_reg[19]/NET0131  , \P2_reg0_reg[1]/NET0131  , \P2_reg0_reg[20]/NET0131  , \P2_reg0_reg[21]/NET0131  , \P2_reg0_reg[22]/NET0131  , \P2_reg0_reg[23]/NET0131  , \P2_reg0_reg[24]/NET0131  , \P2_reg0_reg[25]/NET0131  , \P2_reg0_reg[26]/NET0131  , \P2_reg0_reg[27]/NET0131  , \P2_reg0_reg[28]/NET0131  , \P2_reg0_reg[29]/NET0131  , \P2_reg0_reg[2]/NET0131  , \P2_reg0_reg[30]/NET0131  , \P2_reg0_reg[31]/NET0131  , \P2_reg0_reg[3]/NET0131  , \P2_reg0_reg[4]/NET0131  , \P2_reg0_reg[5]/NET0131  , \P2_reg0_reg[6]/NET0131  , \P2_reg0_reg[7]/NET0131  , \P2_reg0_reg[8]/NET0131  , \P2_reg0_reg[9]/NET0131  , \P2_reg1_reg[0]/NET0131  , \P2_reg1_reg[10]/NET0131  , \P2_reg1_reg[11]/NET0131  , \P2_reg1_reg[12]/NET0131  , \P2_reg1_reg[13]/NET0131  , \P2_reg1_reg[14]/NET0131  , \P2_reg1_reg[15]/NET0131  , \P2_reg1_reg[16]/NET0131  , \P2_reg1_reg[17]/NET0131  , \P2_reg1_reg[18]/NET0131  , \P2_reg1_reg[19]/NET0131  , \P2_reg1_reg[1]/NET0131  , \P2_reg1_reg[20]/NET0131  , \P2_reg1_reg[21]/NET0131  , \P2_reg1_reg[22]/NET0131  , \P2_reg1_reg[23]/NET0131  , \P2_reg1_reg[24]/NET0131  , \P2_reg1_reg[25]/NET0131  , \P2_reg1_reg[26]/NET0131  , \P2_reg1_reg[27]/NET0131  , \P2_reg1_reg[28]/NET0131  , \P2_reg1_reg[29]/NET0131  , \P2_reg1_reg[2]/NET0131  , \P2_reg1_reg[30]/NET0131  , \P2_reg1_reg[31]/NET0131  , \P2_reg1_reg[3]/NET0131  , \P2_reg1_reg[4]/NET0131  , \P2_reg1_reg[5]/NET0131  , \P2_reg1_reg[6]/NET0131  , \P2_reg1_reg[7]/NET0131  , \P2_reg1_reg[8]/NET0131  , \P2_reg1_reg[9]/NET0131  , \P2_reg2_reg[0]/NET0131  , \P2_reg2_reg[10]/NET0131  , \P2_reg2_reg[11]/NET0131  , \P2_reg2_reg[12]/NET0131  , \P2_reg2_reg[13]/NET0131  , \P2_reg2_reg[14]/NET0131  , \P2_reg2_reg[15]/NET0131  , \P2_reg2_reg[16]/NET0131  , \P2_reg2_reg[17]/NET0131  , \P2_reg2_reg[18]/NET0131  , \P2_reg2_reg[19]/NET0131  , \P2_reg2_reg[1]/NET0131  , \P2_reg2_reg[20]/NET0131  , \P2_reg2_reg[21]/NET0131  , \P2_reg2_reg[22]/NET0131  , \P2_reg2_reg[23]/NET0131  , \P2_reg2_reg[24]/NET0131  , \P2_reg2_reg[25]/NET0131  , \P2_reg2_reg[26]/NET0131  , \P2_reg2_reg[27]/NET0131  , \P2_reg2_reg[28]/NET0131  , \P2_reg2_reg[29]/NET0131  , \P2_reg2_reg[2]/NET0131  , \P2_reg2_reg[30]/NET0131  , \P2_reg2_reg[31]/NET0131  , \P2_reg2_reg[3]/NET0131  , \P2_reg2_reg[4]/NET0131  , \P2_reg2_reg[5]/NET0131  , \P2_reg2_reg[6]/NET0131  , \P2_reg2_reg[7]/NET0131  , \P2_reg2_reg[8]/NET0131  , \P2_reg2_reg[9]/NET0131  , \P2_reg3_reg[0]/NET0131  , \P2_reg3_reg[10]/NET0131  , \P2_reg3_reg[11]/NET0131  , \P2_reg3_reg[12]/NET0131  , \P2_reg3_reg[13]/NET0131  , \P2_reg3_reg[14]/NET0131  , \P2_reg3_reg[15]/NET0131  , \P2_reg3_reg[16]/NET0131  , \P2_reg3_reg[17]/NET0131  , \P2_reg3_reg[18]/NET0131  , \P2_reg3_reg[19]/NET0131  , \P2_reg3_reg[1]/NET0131  , \P2_reg3_reg[20]/NET0131  , \P2_reg3_reg[21]/NET0131  , \P2_reg3_reg[22]/NET0131  , \P2_reg3_reg[23]/NET0131  , \P2_reg3_reg[24]/NET0131  , \P2_reg3_reg[25]/NET0131  , \P2_reg3_reg[26]/NET0131  , \P2_reg3_reg[27]/NET0131  , \P2_reg3_reg[28]/NET0131  , \P2_reg3_reg[2]/NET0131  , \P2_reg3_reg[3]/NET0131  , \P2_reg3_reg[4]/NET0131  , \P2_reg3_reg[5]/NET0131  , \P2_reg3_reg[6]/NET0131  , \P2_reg3_reg[7]/NET0131  , \P2_reg3_reg[8]/NET0131  , \P2_reg3_reg[9]/NET0131  , \P2_wr_reg/NET0131  , \si[0]_pad  , \si[10]_pad  , \si[11]_pad  , \si[12]_pad  , \si[13]_pad  , \si[14]_pad  , \si[15]_pad  , \si[16]_pad  , \si[17]_pad  , \si[18]_pad  , \si[19]_pad  , \si[1]_pad  , \si[20]_pad  , \si[21]_pad  , \si[22]_pad  , \si[23]_pad  , \si[24]_pad  , \si[25]_pad  , \si[26]_pad  , \si[27]_pad  , \si[28]_pad  , \si[29]_pad  , \si[2]_pad  , \si[30]_pad  , \si[31]_pad  , \si[3]_pad  , \si[4]_pad  , \si[5]_pad  , \si[6]_pad  , \si[7]_pad  , \si[8]_pad  , \si[9]_pad  , \P1_state_reg[0]/NET0131_syn_2  , \_al_n0  , \_al_n1  , \g35/_0_  , \g73637/_0_  , \g73647/_0_  , \g73648/_0_  , \g73649/_0_  , \g73650/_0_  , \g73667/_0_  , \g73668/_0_  , \g73669/_0_  , \g73670/_0_  , \g73671/_0_  , \g73672/_0_  , \g73674/_0_  , \g73675/_0_  , \g73709/_0_  , \g73710/_0_  , \g73711/_0_  , \g73716/_0_  , \g73717/_0_  , \g73718/_0_  , \g73719/_0_  , \g73720/_0_  , \g73721/_0_  , \g73722/_0_  , \g73723/_0_  , \g73724/_0_  , \g73765/_0_  , \g73769/_0_  , \g73770/_0_  , \g73771/_0_  , \g73772/_0_  , \g73773/_0_  , \g73774/_0_  , \g73775/_0_  , \g73776/_0_  , \g73777/_0_  , \g73778/_0_  , \g73779/_0_  , \g73780/_0_  , \g73781/_0_  , \g73782/_0_  , \g73783/_0_  , \g73784/_0_  , \g73785/_0_  , \g73786/_0_  , \g73787/_0_  , \g73788/_0_  , \g73789/_0_  , \g73790/_0_  , \g73791/_0_  , \g73792/_0_  , \g73845/_0_  , \g73846/_0_  , \g73847/_0_  , \g73848/_0_  , \g73860/_0_  , \g73863/_0_  , \g73864/_0_  , \g73867/_0_  , \g73870/_0_  , \g73871/_0_  , \g73872/_0_  , \g73873/_0_  , \g73874/_0_  , \g73875/_0_  , \g73876/_0_  , \g73877/_0_  , \g73878/_0_  , \g73879/_0_  , \g73880/_0_  , \g73924/_0_  , \g73925/_0_  , \g73949/_0_  , \g73950/_0_  , \g73953/_0_  , \g73954/_0_  , \g73955/_0_  , \g73956/_0_  , \g73957/_0_  , \g73958/_0_  , \g73960/_0_  , \g73961/_0_  , \g73962/_0_  , \g73963/_0_  , \g73964/_0_  , \g73965/_0_  , \g73966/_0_  , \g73967/_0_  , \g73968/_0_  , \g73969/_0_  , \g73970/_0_  , \g73971/_0_  , \g73972/_0_  , \g73973/_0_  , \g73974/_0_  , \g73975/_0_  , \g73976/_0_  , \g73977/_0_  , \g73978/_0_  , \g73979/_0_  , \g73980/_0_  , \g74062/_0_  , \g74063/_0_  , \g74064/_0_  , \g74065/_0_  , \g74066/_0_  , \g74071/_0_  , \g74072/_0_  , \g74105/_0_  , \g74106/_0_  , \g74107/_0_  , \g74108/_0_  , \g74109/_0_  , \g74110/_0_  , \g74111/_0_  , \g74112/_0_  , \g74113/_0_  , \g74114/_0_  , \g74115/_0_  , \g74167/_0_  , \g74168/_0_  , \g74169/_0_  , \g74170/_0_  , \g74172/_0_  , \g74173/_0_  , \g74174/_0_  , \g74175/_0_  , \g74225/_0_  , \g74226/_0_  , \g74227/_0_  , \g74229/_0_  , \g74230/_0_  , \g74231/_0_  , \g74232/_0_  , \g74233/_0_  , \g74234/_0_  , \g74235/_0_  , \g74236/_0_  , \g74237/_0_  , \g74238/_0_  , \g74239/_0_  , \g74240/_0_  , \g74241/_0_  , \g74242/_0_  , \g74243/_0_  , \g74244/_0_  , \g74245/_0_  , \g74246/_0_  , \g74247/_0_  , \g74248/_0_  , \g74249/_0_  , \g74250/_0_  , \g74251/_0_  , \g74252/_0_  , \g74253/_0_  , \g74254/_0_  , \g74255/_0_  , \g74330/_0_  , \g74331/_0_  , \g74333/_0_  , \g74334/_0_  , \g74335/_0_  , \g74390/_0_  , \g74391/_0_  , \g74405/_0_  , \g74407/_0_  , \g74408/_0_  , \g74409/_0_  , \g74410/_0_  , \g74411/_0_  , \g74412/_0_  , \g74413/_0_  , \g74414/_0_  , \g74415/_0_  , \g74416/_0_  , \g74417/_0_  , \g74418/_0_  , \g74419/_0_  , \g74420/_0_  , \g74421/_0_  , \g74422/_0_  , \g74483/_0_  , \g74485/_0_  , \g74486/_0_  , \g74487/_0_  , \g74576/_0_  , \g74578/_0_  , \g74581/_0_  , \g74582/_0_  , \g74583/_0_  , \g74584/_0_  , \g74585/_0_  , \g74588/_0_  , \g74589/_0_  , \g74590/_0_  , \g74591/_0_  , \g74592/_0_  , \g74595/_0_  , \g74596/_0_  , \g74597/_0_  , \g74598/_0_  , \g74599/_0_  , \g74600/_0_  , \g74601/_0_  , \g74602/_0_  , \g74711/_0_  , \g74835/_0_  , \g74836/_0_  , \g74838/_0_  , \g74840/_0_  , \g74841/_0_  , \g74843/_0_  , \g74844/_0_  , \g74963/_0_  , \g75075/_0_  , \g75078/_0_  , \g75079/_0_  , \g75083/_0_  , \g75084/_0_  , \g75089/_0_  , \g75090/_0_  , \g75091/_0_  , \g75224/_0_  , \g75233/_0_  , \g75234/_0_  , \g75427/_0_  , \g75430/_0_  , \g75434/_0_  , \g75436/_0_  , \g75438/_0_  , \g75844/_0_  , \g75850/_0_  , \g75851/_0_  , \g75860/_0_  , \g75865/_0_  , \g75867/_0_  , \g76076/_0_  , \g76375/_0_  , \g76896/_0_  , \g76901/_0_  , \g76905/_0_  , \g77085/_0_  , \g77892/_0_  , \g77897/_0_  , \g77902/_0_  , \g78635/_0_  , \g78636/_0_  , \g78640/_0_  , \g78642/_0_  , \g78645/_0_  , \g78964/_0_  , \g83163/_3_  , \g83164/_3_  , \g83165/_3_  , \g83166/_3_  , \g83167/_3_  , \g83168/_3_  , \g83644/_0_  , \g83645/_0_  , \g83646/_0_  , \g83647/_0_  , \g83648/_0_  , \g83649/_0_  , \g83650/_0_  , \g83651/_0_  , \g83652/_0_  , \g83653/_0_  , \g83654/_0_  , \g83655/_0_  , \g83656/_0_  , \g83657/_0_  , \g83658/_0_  , \g83659/_0_  , \g83660/_0_  , \g83661/_0_  , \g83662/_0_  , \g83663/_0_  , \g83664/_0_  , \g83665/_0_  , \g83666/_0_  , \g83667/_3_  , \g83668/_0_  , \g83669/_0_  , \g83670/_0_  , \g83671/_0_  , \g83715/_3_  , \g83716/_3_  , \g83717/_3_  , \g83718/_3_  , \g83719/_3_  , \g83720/_3_  , \g83721/_3_  , \g83722/_3_  , \g83723/_3_  , \g83724/_3_  , \g83725/_0_  , \g83726/_3_  , \g83727/_3_  , \g83728/_3_  , \g83729/_3_  , \g83730/_3_  , \g83731/_3_  , \g83732/_3_  , \g83733/_3_  , \g83734/_3_  , \g83735/_0_  , \g83736/_0_  , \g83737/_0_  , \g83738/_3_  , \g83739/_3_  , \g83740/_0_  , \g83741/_3_  , \g83742/_3_  , \g84164/_0_  , \g84181/_0_  , \g85146/_0_  , \g85147/_0_  , \g85148/_0_  , \g85149/_0_  , \g85151/_0_  , \g85152/_0_  , \g85154/_0_  , \g85155/_0_  , \g85156/_0_  , \g85157/_0_  , \g85158/_0_  , \g85159/_0_  , \g85160/_0_  , \g85161/_0_  , \g85162/_0_  , \g85163/_0_  , \g85164/_0_  , \g85165/_0_  , \g85166/_0_  , \g85167/_0_  , \g85168/_0_  , \g85169/_0_  , \g85171/_0_  , \g85173/_0_  , \g85174/_0_  , \g85175/_0_  , \g85176/_0_  , \g85178/_0_  , \g85179/_0_  , \g85180/_0_  , \g85181/_0_  , \g85182/_0_  , \g85183/_0_  , \g85184/_0_  , \g85185/_0_  , \g85186/_0_  , \g85187/_0_  , \g85188/_0_  , \g85189/_0_  , \g85190/_0_  , \g85510/_0_  , \g85711/u3_syn_4  , \g85972/_0_  , \g86107/_0_  , \g86200/u3_syn_4  , \g86477/_0_  , \g86548/_0_  , \g86652/u3_syn_4  , \g86807/u3_syn_4  , \g87581/_0_  , \g88104/_0_  , \g88112/_0_  , \g88136/_0_  , \g88148/_0_  , \g88157/_0_  , \g88171/_0_  , \g88179/_0_  , \g88208/_0_  , \g88217/_0_  , \g88222/_0_  , \g88228/_0_  , \g88236/_0_  , \g88242/_0_  , \g88252_dup/_0_  , \g88253/_2_  , \g88259/_0_  , \g88274/_0_  , \g88286/_0_  , \g88296/_0_  , \g88306/_0_  , \g88319/_0_  , \g88330/_0_  , \g88370/_0_  , \g88375/_0_  , \g88388/_0_  , \g88397/_0_  , \g88404/_0_  , \g88793/_0_  , \g88834/_0_  , \g88905/_0_  , \g88910/_0_  , \g88936_dup/_0_  , \g88953/_0_  , \g88962/_0_  , \g89007/_0_  , \g89018/_0_  , \g89024/_0_  , \g89031/_0_  , \g89066/_0_  , \g89082/_0_  , \g89097/_0_  , \g90677/_1__syn_2  , \g96226/_0_  , \g96236/_0_  , \g96261/_0_  , \g96339/_0_  , \g96380/_1_  , \g96418/_0_  , \g96566/_1_  , \g96574/_0_  , \g96620/_0_  , \g96629/_0_  , \g96735/_0_  , \g96866/_0_  , \g96875/_0_  , \g96910/_0_  , \g96946/_0_  , \g96965/_0_  , \g97098/_0_  , \g97228/_0_  , \g97231/_0_  , \g97242/_0_  , \g97384/_0_  , \g97409/_0_  , \g97506/_0_  , \g97626/_0_  , rd_pad , \so[0]_pad  , \so[10]_pad  , \so[11]_pad  , \so[12]_pad  , \so[13]_pad  , \so[14]_pad  , \so[15]_pad  , \so[16]_pad  , \so[17]_pad  , \so[18]_pad  , \so[19]_pad  , \so[1]_pad  , \so[2]_pad  , \so[3]_pad  , \so[4]_pad  , \so[5]_pad  , \so[6]_pad  , \so[7]_pad  , \so[8]_pad  , \so[9]_pad  , wr_pad );
  input \P1_B_reg/NET0131  ;
  input \P1_IR_reg[0]/NET0131  ;
  input \P1_IR_reg[10]/NET0131  ;
  input \P1_IR_reg[11]/NET0131  ;
  input \P1_IR_reg[12]/NET0131  ;
  input \P1_IR_reg[13]/NET0131  ;
  input \P1_IR_reg[14]/NET0131  ;
  input \P1_IR_reg[15]/NET0131  ;
  input \P1_IR_reg[16]/NET0131  ;
  input \P1_IR_reg[17]/NET0131  ;
  input \P1_IR_reg[18]/NET0131  ;
  input \P1_IR_reg[19]/NET0131  ;
  input \P1_IR_reg[1]/NET0131  ;
  input \P1_IR_reg[20]/NET0131  ;
  input \P1_IR_reg[21]/NET0131  ;
  input \P1_IR_reg[22]/NET0131  ;
  input \P1_IR_reg[23]/NET0131  ;
  input \P1_IR_reg[24]/NET0131  ;
  input \P1_IR_reg[25]/NET0131  ;
  input \P1_IR_reg[26]/NET0131  ;
  input \P1_IR_reg[27]/NET0131  ;
  input \P1_IR_reg[28]/NET0131  ;
  input \P1_IR_reg[29]/NET0131  ;
  input \P1_IR_reg[2]/NET0131  ;
  input \P1_IR_reg[30]/NET0131  ;
  input \P1_IR_reg[31]/NET0131  ;
  input \P1_IR_reg[3]/NET0131  ;
  input \P1_IR_reg[4]/NET0131  ;
  input \P1_IR_reg[5]/NET0131  ;
  input \P1_IR_reg[6]/NET0131  ;
  input \P1_IR_reg[7]/NET0131  ;
  input \P1_IR_reg[8]/NET0131  ;
  input \P1_IR_reg[9]/NET0131  ;
  input \P1_addr_reg[0]/NET0131  ;
  input \P1_addr_reg[10]/NET0131  ;
  input \P1_addr_reg[11]/NET0131  ;
  input \P1_addr_reg[12]/NET0131  ;
  input \P1_addr_reg[13]/NET0131  ;
  input \P1_addr_reg[14]/NET0131  ;
  input \P1_addr_reg[15]/NET0131  ;
  input \P1_addr_reg[16]/NET0131  ;
  input \P1_addr_reg[17]/NET0131  ;
  input \P1_addr_reg[18]/NET0131  ;
  input \P1_addr_reg[19]/NET0131  ;
  input \P1_addr_reg[1]/NET0131  ;
  input \P1_addr_reg[2]/NET0131  ;
  input \P1_addr_reg[3]/NET0131  ;
  input \P1_addr_reg[4]/NET0131  ;
  input \P1_addr_reg[5]/NET0131  ;
  input \P1_addr_reg[6]/NET0131  ;
  input \P1_addr_reg[7]/NET0131  ;
  input \P1_addr_reg[8]/NET0131  ;
  input \P1_addr_reg[9]/NET0131  ;
  input \P1_d_reg[0]/NET0131  ;
  input \P1_d_reg[1]/NET0131  ;
  input \P1_datao_reg[0]/NET0131  ;
  input \P1_datao_reg[10]/NET0131  ;
  input \P1_datao_reg[11]/NET0131  ;
  input \P1_datao_reg[12]/NET0131  ;
  input \P1_datao_reg[13]/NET0131  ;
  input \P1_datao_reg[14]/NET0131  ;
  input \P1_datao_reg[15]/NET0131  ;
  input \P1_datao_reg[16]/NET0131  ;
  input \P1_datao_reg[17]/NET0131  ;
  input \P1_datao_reg[18]/NET0131  ;
  input \P1_datao_reg[19]/NET0131  ;
  input \P1_datao_reg[1]/NET0131  ;
  input \P1_datao_reg[20]/NET0131  ;
  input \P1_datao_reg[21]/NET0131  ;
  input \P1_datao_reg[22]/NET0131  ;
  input \P1_datao_reg[23]/NET0131  ;
  input \P1_datao_reg[24]/NET0131  ;
  input \P1_datao_reg[25]/NET0131  ;
  input \P1_datao_reg[26]/NET0131  ;
  input \P1_datao_reg[27]/NET0131  ;
  input \P1_datao_reg[28]/NET0131  ;
  input \P1_datao_reg[29]/NET0131  ;
  input \P1_datao_reg[2]/NET0131  ;
  input \P1_datao_reg[30]/NET0131  ;
  input \P1_datao_reg[31]/NET0131  ;
  input \P1_datao_reg[3]/NET0131  ;
  input \P1_datao_reg[4]/NET0131  ;
  input \P1_datao_reg[5]/NET0131  ;
  input \P1_datao_reg[6]/NET0131  ;
  input \P1_datao_reg[7]/NET0131  ;
  input \P1_datao_reg[8]/NET0131  ;
  input \P1_datao_reg[9]/NET0131  ;
  input \P1_rd_reg/NET0131  ;
  input \P1_reg0_reg[0]/NET0131  ;
  input \P1_reg0_reg[10]/NET0131  ;
  input \P1_reg0_reg[11]/NET0131  ;
  input \P1_reg0_reg[12]/NET0131  ;
  input \P1_reg0_reg[13]/NET0131  ;
  input \P1_reg0_reg[14]/NET0131  ;
  input \P1_reg0_reg[15]/NET0131  ;
  input \P1_reg0_reg[16]/NET0131  ;
  input \P1_reg0_reg[17]/NET0131  ;
  input \P1_reg0_reg[18]/NET0131  ;
  input \P1_reg0_reg[19]/NET0131  ;
  input \P1_reg0_reg[1]/NET0131  ;
  input \P1_reg0_reg[20]/NET0131  ;
  input \P1_reg0_reg[21]/NET0131  ;
  input \P1_reg0_reg[22]/NET0131  ;
  input \P1_reg0_reg[23]/NET0131  ;
  input \P1_reg0_reg[24]/NET0131  ;
  input \P1_reg0_reg[25]/NET0131  ;
  input \P1_reg0_reg[26]/NET0131  ;
  input \P1_reg0_reg[27]/NET0131  ;
  input \P1_reg0_reg[28]/NET0131  ;
  input \P1_reg0_reg[29]/NET0131  ;
  input \P1_reg0_reg[2]/NET0131  ;
  input \P1_reg0_reg[30]/NET0131  ;
  input \P1_reg0_reg[31]/NET0131  ;
  input \P1_reg0_reg[3]/NET0131  ;
  input \P1_reg0_reg[4]/NET0131  ;
  input \P1_reg0_reg[5]/NET0131  ;
  input \P1_reg0_reg[6]/NET0131  ;
  input \P1_reg0_reg[7]/NET0131  ;
  input \P1_reg0_reg[8]/NET0131  ;
  input \P1_reg0_reg[9]/NET0131  ;
  input \P1_reg1_reg[0]/NET0131  ;
  input \P1_reg1_reg[10]/NET0131  ;
  input \P1_reg1_reg[11]/NET0131  ;
  input \P1_reg1_reg[12]/NET0131  ;
  input \P1_reg1_reg[13]/NET0131  ;
  input \P1_reg1_reg[14]/NET0131  ;
  input \P1_reg1_reg[15]/NET0131  ;
  input \P1_reg1_reg[16]/NET0131  ;
  input \P1_reg1_reg[17]/NET0131  ;
  input \P1_reg1_reg[18]/NET0131  ;
  input \P1_reg1_reg[19]/NET0131  ;
  input \P1_reg1_reg[1]/NET0131  ;
  input \P1_reg1_reg[20]/NET0131  ;
  input \P1_reg1_reg[21]/NET0131  ;
  input \P1_reg1_reg[22]/NET0131  ;
  input \P1_reg1_reg[23]/NET0131  ;
  input \P1_reg1_reg[24]/NET0131  ;
  input \P1_reg1_reg[25]/NET0131  ;
  input \P1_reg1_reg[26]/NET0131  ;
  input \P1_reg1_reg[27]/NET0131  ;
  input \P1_reg1_reg[28]/NET0131  ;
  input \P1_reg1_reg[29]/NET0131  ;
  input \P1_reg1_reg[2]/NET0131  ;
  input \P1_reg1_reg[30]/NET0131  ;
  input \P1_reg1_reg[31]/NET0131  ;
  input \P1_reg1_reg[3]/NET0131  ;
  input \P1_reg1_reg[4]/NET0131  ;
  input \P1_reg1_reg[5]/NET0131  ;
  input \P1_reg1_reg[6]/NET0131  ;
  input \P1_reg1_reg[7]/NET0131  ;
  input \P1_reg1_reg[8]/NET0131  ;
  input \P1_reg1_reg[9]/NET0131  ;
  input \P1_reg2_reg[0]/NET0131  ;
  input \P1_reg2_reg[10]/NET0131  ;
  input \P1_reg2_reg[11]/NET0131  ;
  input \P1_reg2_reg[12]/NET0131  ;
  input \P1_reg2_reg[13]/NET0131  ;
  input \P1_reg2_reg[14]/NET0131  ;
  input \P1_reg2_reg[15]/NET0131  ;
  input \P1_reg2_reg[16]/NET0131  ;
  input \P1_reg2_reg[17]/NET0131  ;
  input \P1_reg2_reg[18]/NET0131  ;
  input \P1_reg2_reg[19]/NET0131  ;
  input \P1_reg2_reg[1]/NET0131  ;
  input \P1_reg2_reg[20]/NET0131  ;
  input \P1_reg2_reg[21]/NET0131  ;
  input \P1_reg2_reg[22]/NET0131  ;
  input \P1_reg2_reg[23]/NET0131  ;
  input \P1_reg2_reg[24]/NET0131  ;
  input \P1_reg2_reg[25]/NET0131  ;
  input \P1_reg2_reg[26]/NET0131  ;
  input \P1_reg2_reg[27]/NET0131  ;
  input \P1_reg2_reg[28]/NET0131  ;
  input \P1_reg2_reg[29]/NET0131  ;
  input \P1_reg2_reg[2]/NET0131  ;
  input \P1_reg2_reg[30]/NET0131  ;
  input \P1_reg2_reg[31]/NET0131  ;
  input \P1_reg2_reg[3]/NET0131  ;
  input \P1_reg2_reg[4]/NET0131  ;
  input \P1_reg2_reg[5]/NET0131  ;
  input \P1_reg2_reg[6]/NET0131  ;
  input \P1_reg2_reg[7]/NET0131  ;
  input \P1_reg2_reg[8]/NET0131  ;
  input \P1_reg2_reg[9]/NET0131  ;
  input \P1_reg3_reg[0]/NET0131  ;
  input \P1_reg3_reg[10]/NET0131  ;
  input \P1_reg3_reg[11]/NET0131  ;
  input \P1_reg3_reg[12]/NET0131  ;
  input \P1_reg3_reg[13]/NET0131  ;
  input \P1_reg3_reg[14]/NET0131  ;
  input \P1_reg3_reg[15]/NET0131  ;
  input \P1_reg3_reg[16]/NET0131  ;
  input \P1_reg3_reg[17]/NET0131  ;
  input \P1_reg3_reg[18]/NET0131  ;
  input \P1_reg3_reg[19]/NET0131  ;
  input \P1_reg3_reg[1]/NET0131  ;
  input \P1_reg3_reg[20]/NET0131  ;
  input \P1_reg3_reg[21]/NET0131  ;
  input \P1_reg3_reg[22]/NET0131  ;
  input \P1_reg3_reg[23]/NET0131  ;
  input \P1_reg3_reg[24]/NET0131  ;
  input \P1_reg3_reg[25]/NET0131  ;
  input \P1_reg3_reg[26]/NET0131  ;
  input \P1_reg3_reg[27]/NET0131  ;
  input \P1_reg3_reg[28]/NET0131  ;
  input \P1_reg3_reg[2]/NET0131  ;
  input \P1_reg3_reg[3]/NET0131  ;
  input \P1_reg3_reg[4]/NET0131  ;
  input \P1_reg3_reg[5]/NET0131  ;
  input \P1_reg3_reg[6]/NET0131  ;
  input \P1_reg3_reg[7]/NET0131  ;
  input \P1_reg3_reg[8]/NET0131  ;
  input \P1_reg3_reg[9]/NET0131  ;
  input \P1_state_reg[0]/NET0131  ;
  input \P1_wr_reg/NET0131  ;
  input \P2_B_reg/NET0131  ;
  input \P2_IR_reg[0]/NET0131  ;
  input \P2_IR_reg[10]/NET0131  ;
  input \P2_IR_reg[11]/NET0131  ;
  input \P2_IR_reg[12]/NET0131  ;
  input \P2_IR_reg[13]/NET0131  ;
  input \P2_IR_reg[14]/NET0131  ;
  input \P2_IR_reg[15]/NET0131  ;
  input \P2_IR_reg[16]/NET0131  ;
  input \P2_IR_reg[17]/NET0131  ;
  input \P2_IR_reg[18]/NET0131  ;
  input \P2_IR_reg[19]/NET0131  ;
  input \P2_IR_reg[1]/NET0131  ;
  input \P2_IR_reg[20]/NET0131  ;
  input \P2_IR_reg[21]/NET0131  ;
  input \P2_IR_reg[22]/NET0131  ;
  input \P2_IR_reg[23]/NET0131  ;
  input \P2_IR_reg[24]/NET0131  ;
  input \P2_IR_reg[25]/NET0131  ;
  input \P2_IR_reg[26]/NET0131  ;
  input \P2_IR_reg[27]/NET0131  ;
  input \P2_IR_reg[28]/NET0131  ;
  input \P2_IR_reg[29]/NET0131  ;
  input \P2_IR_reg[2]/NET0131  ;
  input \P2_IR_reg[30]/NET0131  ;
  input \P2_IR_reg[31]/NET0131  ;
  input \P2_IR_reg[3]/NET0131  ;
  input \P2_IR_reg[4]/NET0131  ;
  input \P2_IR_reg[5]/NET0131  ;
  input \P2_IR_reg[6]/NET0131  ;
  input \P2_IR_reg[7]/NET0131  ;
  input \P2_IR_reg[8]/NET0131  ;
  input \P2_IR_reg[9]/NET0131  ;
  input \P2_addr_reg[0]/NET0131  ;
  input \P2_addr_reg[10]/NET0131  ;
  input \P2_addr_reg[11]/NET0131  ;
  input \P2_addr_reg[12]/NET0131  ;
  input \P2_addr_reg[13]/NET0131  ;
  input \P2_addr_reg[14]/NET0131  ;
  input \P2_addr_reg[15]/NET0131  ;
  input \P2_addr_reg[16]/NET0131  ;
  input \P2_addr_reg[17]/NET0131  ;
  input \P2_addr_reg[18]/NET0131  ;
  input \P2_addr_reg[19]/NET0131  ;
  input \P2_addr_reg[1]/NET0131  ;
  input \P2_addr_reg[2]/NET0131  ;
  input \P2_addr_reg[3]/NET0131  ;
  input \P2_addr_reg[4]/NET0131  ;
  input \P2_addr_reg[5]/NET0131  ;
  input \P2_addr_reg[6]/NET0131  ;
  input \P2_addr_reg[7]/NET0131  ;
  input \P2_addr_reg[8]/NET0131  ;
  input \P2_addr_reg[9]/NET0131  ;
  input \P2_d_reg[0]/NET0131  ;
  input \P2_d_reg[1]/NET0131  ;
  input \P2_datao_reg[0]/NET0131  ;
  input \P2_datao_reg[10]/NET0131  ;
  input \P2_datao_reg[11]/NET0131  ;
  input \P2_datao_reg[12]/NET0131  ;
  input \P2_datao_reg[13]/NET0131  ;
  input \P2_datao_reg[14]/NET0131  ;
  input \P2_datao_reg[15]/NET0131  ;
  input \P2_datao_reg[16]/NET0131  ;
  input \P2_datao_reg[17]/NET0131  ;
  input \P2_datao_reg[18]/NET0131  ;
  input \P2_datao_reg[19]/NET0131  ;
  input \P2_datao_reg[1]/NET0131  ;
  input \P2_datao_reg[20]/NET0131  ;
  input \P2_datao_reg[21]/NET0131  ;
  input \P2_datao_reg[22]/NET0131  ;
  input \P2_datao_reg[23]/NET0131  ;
  input \P2_datao_reg[24]/NET0131  ;
  input \P2_datao_reg[25]/NET0131  ;
  input \P2_datao_reg[26]/NET0131  ;
  input \P2_datao_reg[27]/NET0131  ;
  input \P2_datao_reg[28]/NET0131  ;
  input \P2_datao_reg[29]/NET0131  ;
  input \P2_datao_reg[2]/NET0131  ;
  input \P2_datao_reg[30]/NET0131  ;
  input \P2_datao_reg[31]/NET0131  ;
  input \P2_datao_reg[3]/NET0131  ;
  input \P2_datao_reg[4]/NET0131  ;
  input \P2_datao_reg[5]/NET0131  ;
  input \P2_datao_reg[6]/NET0131  ;
  input \P2_datao_reg[7]/NET0131  ;
  input \P2_datao_reg[8]/NET0131  ;
  input \P2_datao_reg[9]/NET0131  ;
  input \P2_rd_reg/NET0131  ;
  input \P2_reg0_reg[0]/NET0131  ;
  input \P2_reg0_reg[10]/NET0131  ;
  input \P2_reg0_reg[11]/NET0131  ;
  input \P2_reg0_reg[12]/NET0131  ;
  input \P2_reg0_reg[13]/NET0131  ;
  input \P2_reg0_reg[14]/NET0131  ;
  input \P2_reg0_reg[15]/NET0131  ;
  input \P2_reg0_reg[16]/NET0131  ;
  input \P2_reg0_reg[17]/NET0131  ;
  input \P2_reg0_reg[18]/NET0131  ;
  input \P2_reg0_reg[19]/NET0131  ;
  input \P2_reg0_reg[1]/NET0131  ;
  input \P2_reg0_reg[20]/NET0131  ;
  input \P2_reg0_reg[21]/NET0131  ;
  input \P2_reg0_reg[22]/NET0131  ;
  input \P2_reg0_reg[23]/NET0131  ;
  input \P2_reg0_reg[24]/NET0131  ;
  input \P2_reg0_reg[25]/NET0131  ;
  input \P2_reg0_reg[26]/NET0131  ;
  input \P2_reg0_reg[27]/NET0131  ;
  input \P2_reg0_reg[28]/NET0131  ;
  input \P2_reg0_reg[29]/NET0131  ;
  input \P2_reg0_reg[2]/NET0131  ;
  input \P2_reg0_reg[30]/NET0131  ;
  input \P2_reg0_reg[31]/NET0131  ;
  input \P2_reg0_reg[3]/NET0131  ;
  input \P2_reg0_reg[4]/NET0131  ;
  input \P2_reg0_reg[5]/NET0131  ;
  input \P2_reg0_reg[6]/NET0131  ;
  input \P2_reg0_reg[7]/NET0131  ;
  input \P2_reg0_reg[8]/NET0131  ;
  input \P2_reg0_reg[9]/NET0131  ;
  input \P2_reg1_reg[0]/NET0131  ;
  input \P2_reg1_reg[10]/NET0131  ;
  input \P2_reg1_reg[11]/NET0131  ;
  input \P2_reg1_reg[12]/NET0131  ;
  input \P2_reg1_reg[13]/NET0131  ;
  input \P2_reg1_reg[14]/NET0131  ;
  input \P2_reg1_reg[15]/NET0131  ;
  input \P2_reg1_reg[16]/NET0131  ;
  input \P2_reg1_reg[17]/NET0131  ;
  input \P2_reg1_reg[18]/NET0131  ;
  input \P2_reg1_reg[19]/NET0131  ;
  input \P2_reg1_reg[1]/NET0131  ;
  input \P2_reg1_reg[20]/NET0131  ;
  input \P2_reg1_reg[21]/NET0131  ;
  input \P2_reg1_reg[22]/NET0131  ;
  input \P2_reg1_reg[23]/NET0131  ;
  input \P2_reg1_reg[24]/NET0131  ;
  input \P2_reg1_reg[25]/NET0131  ;
  input \P2_reg1_reg[26]/NET0131  ;
  input \P2_reg1_reg[27]/NET0131  ;
  input \P2_reg1_reg[28]/NET0131  ;
  input \P2_reg1_reg[29]/NET0131  ;
  input \P2_reg1_reg[2]/NET0131  ;
  input \P2_reg1_reg[30]/NET0131  ;
  input \P2_reg1_reg[31]/NET0131  ;
  input \P2_reg1_reg[3]/NET0131  ;
  input \P2_reg1_reg[4]/NET0131  ;
  input \P2_reg1_reg[5]/NET0131  ;
  input \P2_reg1_reg[6]/NET0131  ;
  input \P2_reg1_reg[7]/NET0131  ;
  input \P2_reg1_reg[8]/NET0131  ;
  input \P2_reg1_reg[9]/NET0131  ;
  input \P2_reg2_reg[0]/NET0131  ;
  input \P2_reg2_reg[10]/NET0131  ;
  input \P2_reg2_reg[11]/NET0131  ;
  input \P2_reg2_reg[12]/NET0131  ;
  input \P2_reg2_reg[13]/NET0131  ;
  input \P2_reg2_reg[14]/NET0131  ;
  input \P2_reg2_reg[15]/NET0131  ;
  input \P2_reg2_reg[16]/NET0131  ;
  input \P2_reg2_reg[17]/NET0131  ;
  input \P2_reg2_reg[18]/NET0131  ;
  input \P2_reg2_reg[19]/NET0131  ;
  input \P2_reg2_reg[1]/NET0131  ;
  input \P2_reg2_reg[20]/NET0131  ;
  input \P2_reg2_reg[21]/NET0131  ;
  input \P2_reg2_reg[22]/NET0131  ;
  input \P2_reg2_reg[23]/NET0131  ;
  input \P2_reg2_reg[24]/NET0131  ;
  input \P2_reg2_reg[25]/NET0131  ;
  input \P2_reg2_reg[26]/NET0131  ;
  input \P2_reg2_reg[27]/NET0131  ;
  input \P2_reg2_reg[28]/NET0131  ;
  input \P2_reg2_reg[29]/NET0131  ;
  input \P2_reg2_reg[2]/NET0131  ;
  input \P2_reg2_reg[30]/NET0131  ;
  input \P2_reg2_reg[31]/NET0131  ;
  input \P2_reg2_reg[3]/NET0131  ;
  input \P2_reg2_reg[4]/NET0131  ;
  input \P2_reg2_reg[5]/NET0131  ;
  input \P2_reg2_reg[6]/NET0131  ;
  input \P2_reg2_reg[7]/NET0131  ;
  input \P2_reg2_reg[8]/NET0131  ;
  input \P2_reg2_reg[9]/NET0131  ;
  input \P2_reg3_reg[0]/NET0131  ;
  input \P2_reg3_reg[10]/NET0131  ;
  input \P2_reg3_reg[11]/NET0131  ;
  input \P2_reg3_reg[12]/NET0131  ;
  input \P2_reg3_reg[13]/NET0131  ;
  input \P2_reg3_reg[14]/NET0131  ;
  input \P2_reg3_reg[15]/NET0131  ;
  input \P2_reg3_reg[16]/NET0131  ;
  input \P2_reg3_reg[17]/NET0131  ;
  input \P2_reg3_reg[18]/NET0131  ;
  input \P2_reg3_reg[19]/NET0131  ;
  input \P2_reg3_reg[1]/NET0131  ;
  input \P2_reg3_reg[20]/NET0131  ;
  input \P2_reg3_reg[21]/NET0131  ;
  input \P2_reg3_reg[22]/NET0131  ;
  input \P2_reg3_reg[23]/NET0131  ;
  input \P2_reg3_reg[24]/NET0131  ;
  input \P2_reg3_reg[25]/NET0131  ;
  input \P2_reg3_reg[26]/NET0131  ;
  input \P2_reg3_reg[27]/NET0131  ;
  input \P2_reg3_reg[28]/NET0131  ;
  input \P2_reg3_reg[2]/NET0131  ;
  input \P2_reg3_reg[3]/NET0131  ;
  input \P2_reg3_reg[4]/NET0131  ;
  input \P2_reg3_reg[5]/NET0131  ;
  input \P2_reg3_reg[6]/NET0131  ;
  input \P2_reg3_reg[7]/NET0131  ;
  input \P2_reg3_reg[8]/NET0131  ;
  input \P2_reg3_reg[9]/NET0131  ;
  input \P2_wr_reg/NET0131  ;
  input \si[0]_pad  ;
  input \si[10]_pad  ;
  input \si[11]_pad  ;
  input \si[12]_pad  ;
  input \si[13]_pad  ;
  input \si[14]_pad  ;
  input \si[15]_pad  ;
  input \si[16]_pad  ;
  input \si[17]_pad  ;
  input \si[18]_pad  ;
  input \si[19]_pad  ;
  input \si[1]_pad  ;
  input \si[20]_pad  ;
  input \si[21]_pad  ;
  input \si[22]_pad  ;
  input \si[23]_pad  ;
  input \si[24]_pad  ;
  input \si[25]_pad  ;
  input \si[26]_pad  ;
  input \si[27]_pad  ;
  input \si[28]_pad  ;
  input \si[29]_pad  ;
  input \si[2]_pad  ;
  input \si[30]_pad  ;
  input \si[31]_pad  ;
  input \si[3]_pad  ;
  input \si[4]_pad  ;
  input \si[5]_pad  ;
  input \si[6]_pad  ;
  input \si[7]_pad  ;
  input \si[8]_pad  ;
  input \si[9]_pad  ;
  output \P1_state_reg[0]/NET0131_syn_2  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g35/_0_  ;
  output \g73637/_0_  ;
  output \g73647/_0_  ;
  output \g73648/_0_  ;
  output \g73649/_0_  ;
  output \g73650/_0_  ;
  output \g73667/_0_  ;
  output \g73668/_0_  ;
  output \g73669/_0_  ;
  output \g73670/_0_  ;
  output \g73671/_0_  ;
  output \g73672/_0_  ;
  output \g73674/_0_  ;
  output \g73675/_0_  ;
  output \g73709/_0_  ;
  output \g73710/_0_  ;
  output \g73711/_0_  ;
  output \g73716/_0_  ;
  output \g73717/_0_  ;
  output \g73718/_0_  ;
  output \g73719/_0_  ;
  output \g73720/_0_  ;
  output \g73721/_0_  ;
  output \g73722/_0_  ;
  output \g73723/_0_  ;
  output \g73724/_0_  ;
  output \g73765/_0_  ;
  output \g73769/_0_  ;
  output \g73770/_0_  ;
  output \g73771/_0_  ;
  output \g73772/_0_  ;
  output \g73773/_0_  ;
  output \g73774/_0_  ;
  output \g73775/_0_  ;
  output \g73776/_0_  ;
  output \g73777/_0_  ;
  output \g73778/_0_  ;
  output \g73779/_0_  ;
  output \g73780/_0_  ;
  output \g73781/_0_  ;
  output \g73782/_0_  ;
  output \g73783/_0_  ;
  output \g73784/_0_  ;
  output \g73785/_0_  ;
  output \g73786/_0_  ;
  output \g73787/_0_  ;
  output \g73788/_0_  ;
  output \g73789/_0_  ;
  output \g73790/_0_  ;
  output \g73791/_0_  ;
  output \g73792/_0_  ;
  output \g73845/_0_  ;
  output \g73846/_0_  ;
  output \g73847/_0_  ;
  output \g73848/_0_  ;
  output \g73860/_0_  ;
  output \g73863/_0_  ;
  output \g73864/_0_  ;
  output \g73867/_0_  ;
  output \g73870/_0_  ;
  output \g73871/_0_  ;
  output \g73872/_0_  ;
  output \g73873/_0_  ;
  output \g73874/_0_  ;
  output \g73875/_0_  ;
  output \g73876/_0_  ;
  output \g73877/_0_  ;
  output \g73878/_0_  ;
  output \g73879/_0_  ;
  output \g73880/_0_  ;
  output \g73924/_0_  ;
  output \g73925/_0_  ;
  output \g73949/_0_  ;
  output \g73950/_0_  ;
  output \g73953/_0_  ;
  output \g73954/_0_  ;
  output \g73955/_0_  ;
  output \g73956/_0_  ;
  output \g73957/_0_  ;
  output \g73958/_0_  ;
  output \g73960/_0_  ;
  output \g73961/_0_  ;
  output \g73962/_0_  ;
  output \g73963/_0_  ;
  output \g73964/_0_  ;
  output \g73965/_0_  ;
  output \g73966/_0_  ;
  output \g73967/_0_  ;
  output \g73968/_0_  ;
  output \g73969/_0_  ;
  output \g73970/_0_  ;
  output \g73971/_0_  ;
  output \g73972/_0_  ;
  output \g73973/_0_  ;
  output \g73974/_0_  ;
  output \g73975/_0_  ;
  output \g73976/_0_  ;
  output \g73977/_0_  ;
  output \g73978/_0_  ;
  output \g73979/_0_  ;
  output \g73980/_0_  ;
  output \g74062/_0_  ;
  output \g74063/_0_  ;
  output \g74064/_0_  ;
  output \g74065/_0_  ;
  output \g74066/_0_  ;
  output \g74071/_0_  ;
  output \g74072/_0_  ;
  output \g74105/_0_  ;
  output \g74106/_0_  ;
  output \g74107/_0_  ;
  output \g74108/_0_  ;
  output \g74109/_0_  ;
  output \g74110/_0_  ;
  output \g74111/_0_  ;
  output \g74112/_0_  ;
  output \g74113/_0_  ;
  output \g74114/_0_  ;
  output \g74115/_0_  ;
  output \g74167/_0_  ;
  output \g74168/_0_  ;
  output \g74169/_0_  ;
  output \g74170/_0_  ;
  output \g74172/_0_  ;
  output \g74173/_0_  ;
  output \g74174/_0_  ;
  output \g74175/_0_  ;
  output \g74225/_0_  ;
  output \g74226/_0_  ;
  output \g74227/_0_  ;
  output \g74229/_0_  ;
  output \g74230/_0_  ;
  output \g74231/_0_  ;
  output \g74232/_0_  ;
  output \g74233/_0_  ;
  output \g74234/_0_  ;
  output \g74235/_0_  ;
  output \g74236/_0_  ;
  output \g74237/_0_  ;
  output \g74238/_0_  ;
  output \g74239/_0_  ;
  output \g74240/_0_  ;
  output \g74241/_0_  ;
  output \g74242/_0_  ;
  output \g74243/_0_  ;
  output \g74244/_0_  ;
  output \g74245/_0_  ;
  output \g74246/_0_  ;
  output \g74247/_0_  ;
  output \g74248/_0_  ;
  output \g74249/_0_  ;
  output \g74250/_0_  ;
  output \g74251/_0_  ;
  output \g74252/_0_  ;
  output \g74253/_0_  ;
  output \g74254/_0_  ;
  output \g74255/_0_  ;
  output \g74330/_0_  ;
  output \g74331/_0_  ;
  output \g74333/_0_  ;
  output \g74334/_0_  ;
  output \g74335/_0_  ;
  output \g74390/_0_  ;
  output \g74391/_0_  ;
  output \g74405/_0_  ;
  output \g74407/_0_  ;
  output \g74408/_0_  ;
  output \g74409/_0_  ;
  output \g74410/_0_  ;
  output \g74411/_0_  ;
  output \g74412/_0_  ;
  output \g74413/_0_  ;
  output \g74414/_0_  ;
  output \g74415/_0_  ;
  output \g74416/_0_  ;
  output \g74417/_0_  ;
  output \g74418/_0_  ;
  output \g74419/_0_  ;
  output \g74420/_0_  ;
  output \g74421/_0_  ;
  output \g74422/_0_  ;
  output \g74483/_0_  ;
  output \g74485/_0_  ;
  output \g74486/_0_  ;
  output \g74487/_0_  ;
  output \g74576/_0_  ;
  output \g74578/_0_  ;
  output \g74581/_0_  ;
  output \g74582/_0_  ;
  output \g74583/_0_  ;
  output \g74584/_0_  ;
  output \g74585/_0_  ;
  output \g74588/_0_  ;
  output \g74589/_0_  ;
  output \g74590/_0_  ;
  output \g74591/_0_  ;
  output \g74592/_0_  ;
  output \g74595/_0_  ;
  output \g74596/_0_  ;
  output \g74597/_0_  ;
  output \g74598/_0_  ;
  output \g74599/_0_  ;
  output \g74600/_0_  ;
  output \g74601/_0_  ;
  output \g74602/_0_  ;
  output \g74711/_0_  ;
  output \g74835/_0_  ;
  output \g74836/_0_  ;
  output \g74838/_0_  ;
  output \g74840/_0_  ;
  output \g74841/_0_  ;
  output \g74843/_0_  ;
  output \g74844/_0_  ;
  output \g74963/_0_  ;
  output \g75075/_0_  ;
  output \g75078/_0_  ;
  output \g75079/_0_  ;
  output \g75083/_0_  ;
  output \g75084/_0_  ;
  output \g75089/_0_  ;
  output \g75090/_0_  ;
  output \g75091/_0_  ;
  output \g75224/_0_  ;
  output \g75233/_0_  ;
  output \g75234/_0_  ;
  output \g75427/_0_  ;
  output \g75430/_0_  ;
  output \g75434/_0_  ;
  output \g75436/_0_  ;
  output \g75438/_0_  ;
  output \g75844/_0_  ;
  output \g75850/_0_  ;
  output \g75851/_0_  ;
  output \g75860/_0_  ;
  output \g75865/_0_  ;
  output \g75867/_0_  ;
  output \g76076/_0_  ;
  output \g76375/_0_  ;
  output \g76896/_0_  ;
  output \g76901/_0_  ;
  output \g76905/_0_  ;
  output \g77085/_0_  ;
  output \g77892/_0_  ;
  output \g77897/_0_  ;
  output \g77902/_0_  ;
  output \g78635/_0_  ;
  output \g78636/_0_  ;
  output \g78640/_0_  ;
  output \g78642/_0_  ;
  output \g78645/_0_  ;
  output \g78964/_0_  ;
  output \g83163/_3_  ;
  output \g83164/_3_  ;
  output \g83165/_3_  ;
  output \g83166/_3_  ;
  output \g83167/_3_  ;
  output \g83168/_3_  ;
  output \g83644/_0_  ;
  output \g83645/_0_  ;
  output \g83646/_0_  ;
  output \g83647/_0_  ;
  output \g83648/_0_  ;
  output \g83649/_0_  ;
  output \g83650/_0_  ;
  output \g83651/_0_  ;
  output \g83652/_0_  ;
  output \g83653/_0_  ;
  output \g83654/_0_  ;
  output \g83655/_0_  ;
  output \g83656/_0_  ;
  output \g83657/_0_  ;
  output \g83658/_0_  ;
  output \g83659/_0_  ;
  output \g83660/_0_  ;
  output \g83661/_0_  ;
  output \g83662/_0_  ;
  output \g83663/_0_  ;
  output \g83664/_0_  ;
  output \g83665/_0_  ;
  output \g83666/_0_  ;
  output \g83667/_3_  ;
  output \g83668/_0_  ;
  output \g83669/_0_  ;
  output \g83670/_0_  ;
  output \g83671/_0_  ;
  output \g83715/_3_  ;
  output \g83716/_3_  ;
  output \g83717/_3_  ;
  output \g83718/_3_  ;
  output \g83719/_3_  ;
  output \g83720/_3_  ;
  output \g83721/_3_  ;
  output \g83722/_3_  ;
  output \g83723/_3_  ;
  output \g83724/_3_  ;
  output \g83725/_0_  ;
  output \g83726/_3_  ;
  output \g83727/_3_  ;
  output \g83728/_3_  ;
  output \g83729/_3_  ;
  output \g83730/_3_  ;
  output \g83731/_3_  ;
  output \g83732/_3_  ;
  output \g83733/_3_  ;
  output \g83734/_3_  ;
  output \g83735/_0_  ;
  output \g83736/_0_  ;
  output \g83737/_0_  ;
  output \g83738/_3_  ;
  output \g83739/_3_  ;
  output \g83740/_0_  ;
  output \g83741/_3_  ;
  output \g83742/_3_  ;
  output \g84164/_0_  ;
  output \g84181/_0_  ;
  output \g85146/_0_  ;
  output \g85147/_0_  ;
  output \g85148/_0_  ;
  output \g85149/_0_  ;
  output \g85151/_0_  ;
  output \g85152/_0_  ;
  output \g85154/_0_  ;
  output \g85155/_0_  ;
  output \g85156/_0_  ;
  output \g85157/_0_  ;
  output \g85158/_0_  ;
  output \g85159/_0_  ;
  output \g85160/_0_  ;
  output \g85161/_0_  ;
  output \g85162/_0_  ;
  output \g85163/_0_  ;
  output \g85164/_0_  ;
  output \g85165/_0_  ;
  output \g85166/_0_  ;
  output \g85167/_0_  ;
  output \g85168/_0_  ;
  output \g85169/_0_  ;
  output \g85171/_0_  ;
  output \g85173/_0_  ;
  output \g85174/_0_  ;
  output \g85175/_0_  ;
  output \g85176/_0_  ;
  output \g85178/_0_  ;
  output \g85179/_0_  ;
  output \g85180/_0_  ;
  output \g85181/_0_  ;
  output \g85182/_0_  ;
  output \g85183/_0_  ;
  output \g85184/_0_  ;
  output \g85185/_0_  ;
  output \g85186/_0_  ;
  output \g85187/_0_  ;
  output \g85188/_0_  ;
  output \g85189/_0_  ;
  output \g85190/_0_  ;
  output \g85510/_0_  ;
  output \g85711/u3_syn_4  ;
  output \g85972/_0_  ;
  output \g86107/_0_  ;
  output \g86200/u3_syn_4  ;
  output \g86477/_0_  ;
  output \g86548/_0_  ;
  output \g86652/u3_syn_4  ;
  output \g86807/u3_syn_4  ;
  output \g87581/_0_  ;
  output \g88104/_0_  ;
  output \g88112/_0_  ;
  output \g88136/_0_  ;
  output \g88148/_0_  ;
  output \g88157/_0_  ;
  output \g88171/_0_  ;
  output \g88179/_0_  ;
  output \g88208/_0_  ;
  output \g88217/_0_  ;
  output \g88222/_0_  ;
  output \g88228/_0_  ;
  output \g88236/_0_  ;
  output \g88242/_0_  ;
  output \g88252_dup/_0_  ;
  output \g88253/_2_  ;
  output \g88259/_0_  ;
  output \g88274/_0_  ;
  output \g88286/_0_  ;
  output \g88296/_0_  ;
  output \g88306/_0_  ;
  output \g88319/_0_  ;
  output \g88330/_0_  ;
  output \g88370/_0_  ;
  output \g88375/_0_  ;
  output \g88388/_0_  ;
  output \g88397/_0_  ;
  output \g88404/_0_  ;
  output \g88793/_0_  ;
  output \g88834/_0_  ;
  output \g88905/_0_  ;
  output \g88910/_0_  ;
  output \g88936_dup/_0_  ;
  output \g88953/_0_  ;
  output \g88962/_0_  ;
  output \g89007/_0_  ;
  output \g89018/_0_  ;
  output \g89024/_0_  ;
  output \g89031/_0_  ;
  output \g89066/_0_  ;
  output \g89082/_0_  ;
  output \g89097/_0_  ;
  output \g90677/_1__syn_2  ;
  output \g96226/_0_  ;
  output \g96236/_0_  ;
  output \g96261/_0_  ;
  output \g96339/_0_  ;
  output \g96380/_1_  ;
  output \g96418/_0_  ;
  output \g96566/_1_  ;
  output \g96574/_0_  ;
  output \g96620/_0_  ;
  output \g96629/_0_  ;
  output \g96735/_0_  ;
  output \g96866/_0_  ;
  output \g96875/_0_  ;
  output \g96910/_0_  ;
  output \g96946/_0_  ;
  output \g96965/_0_  ;
  output \g97098/_0_  ;
  output \g97228/_0_  ;
  output \g97231/_0_  ;
  output \g97242/_0_  ;
  output \g97384/_0_  ;
  output \g97409/_0_  ;
  output \g97506/_0_  ;
  output \g97626/_0_  ;
  output rd_pad ;
  output \so[0]_pad  ;
  output \so[10]_pad  ;
  output \so[11]_pad  ;
  output \so[12]_pad  ;
  output \so[13]_pad  ;
  output \so[14]_pad  ;
  output \so[15]_pad  ;
  output \so[16]_pad  ;
  output \so[17]_pad  ;
  output \so[18]_pad  ;
  output \so[19]_pad  ;
  output \so[1]_pad  ;
  output \so[2]_pad  ;
  output \so[3]_pad  ;
  output \so[4]_pad  ;
  output \so[5]_pad  ;
  output \so[6]_pad  ;
  output \so[7]_pad  ;
  output \so[8]_pad  ;
  output \so[9]_pad  ;
  output wr_pad ;
  wire n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 ;
  assign n462 = ~\P1_IR_reg[6]/NET0131  & ~\P1_IR_reg[7]/NET0131  ;
  assign n463 = ~\P1_IR_reg[0]/NET0131  & ~\P1_IR_reg[1]/NET0131  ;
  assign n464 = ~\P1_IR_reg[2]/NET0131  & ~\P1_IR_reg[3]/NET0131  ;
  assign n465 = n463 & n464 ;
  assign n466 = ~\P1_IR_reg[4]/NET0131  & ~\P1_IR_reg[5]/NET0131  ;
  assign n467 = n465 & n466 ;
  assign n468 = n462 & n467 ;
  assign n469 = ~\P1_IR_reg[8]/NET0131  & n468 ;
  assign n473 = ~\P1_IR_reg[14]/NET0131  & ~\P1_IR_reg[15]/NET0131  ;
  assign n474 = ~\P1_IR_reg[16]/NET0131  & n473 ;
  assign n470 = ~\P1_IR_reg[10]/NET0131  & ~\P1_IR_reg[11]/NET0131  ;
  assign n471 = ~\P1_IR_reg[12]/NET0131  & ~\P1_IR_reg[13]/NET0131  ;
  assign n472 = n470 & n471 ;
  assign n475 = ~\P1_IR_reg[9]/NET0131  & n472 ;
  assign n476 = n474 & n475 ;
  assign n477 = n469 & n476 ;
  assign n480 = ~\P1_IR_reg[19]/NET0131  & ~\P1_IR_reg[20]/NET0131  ;
  assign n481 = ~\P1_IR_reg[17]/NET0131  & ~\P1_IR_reg[18]/NET0131  ;
  assign n482 = n480 & n481 ;
  assign n478 = ~\P1_IR_reg[22]/NET0131  & ~\P1_IR_reg[23]/NET0131  ;
  assign n479 = ~\P1_IR_reg[21]/NET0131  & n478 ;
  assign n483 = ~\P1_IR_reg[24]/NET0131  & n479 ;
  assign n484 = n482 & n483 ;
  assign n485 = n477 & n484 ;
  assign n486 = \P1_IR_reg[31]/NET0131  & ~n485 ;
  assign n487 = ~\P1_IR_reg[27]/NET0131  & ~\P1_IR_reg[28]/NET0131  ;
  assign n488 = ~\P1_IR_reg[25]/NET0131  & ~\P1_IR_reg[26]/NET0131  ;
  assign n489 = n487 & n488 ;
  assign n490 = \P1_IR_reg[31]/NET0131  & ~n489 ;
  assign n491 = ~n486 & ~n490 ;
  assign n492 = \P1_IR_reg[29]/NET0131  & ~n491 ;
  assign n493 = ~\P1_IR_reg[29]/NET0131  & n491 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = ~\P1_IR_reg[8]/NET0131  & ~\P1_IR_reg[9]/NET0131  ;
  assign n496 = n462 & n495 ;
  assign n497 = n467 & n496 ;
  assign n498 = n472 & n497 ;
  assign n499 = ~\P1_IR_reg[21]/NET0131  & n474 ;
  assign n500 = n482 & n499 ;
  assign n501 = n498 & n500 ;
  assign n502 = ~\P1_IR_reg[24]/NET0131  & ~\P1_IR_reg[25]/NET0131  ;
  assign n503 = n478 & n502 ;
  assign n504 = n501 & n503 ;
  assign n505 = \P1_IR_reg[31]/NET0131  & ~n504 ;
  assign n506 = ~\P1_IR_reg[29]/NET0131  & n487 ;
  assign n507 = ~\P1_IR_reg[26]/NET0131  & n506 ;
  assign n508 = \P1_IR_reg[31]/NET0131  & ~n507 ;
  assign n509 = ~n505 & ~n508 ;
  assign n510 = \P1_IR_reg[30]/NET0131  & ~n509 ;
  assign n511 = ~\P1_IR_reg[30]/NET0131  & n509 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = ~n494 & n512 ;
  assign n514 = \P1_reg2_reg[3]/NET0131  & n513 ;
  assign n515 = n494 & ~n512 ;
  assign n516 = \P1_reg1_reg[3]/NET0131  & n515 ;
  assign n521 = ~n514 & ~n516 ;
  assign n517 = ~n494 & ~n512 ;
  assign n518 = \P1_reg0_reg[3]/NET0131  & n517 ;
  assign n519 = n494 & n512 ;
  assign n520 = ~\P1_reg3_reg[3]/NET0131  & n519 ;
  assign n522 = ~n518 & ~n520 ;
  assign n523 = n521 & n522 ;
  assign n524 = ~\P2_IR_reg[10]/NET0131  & ~\P2_IR_reg[11]/NET0131  ;
  assign n525 = ~\P2_IR_reg[9]/NET0131  & n524 ;
  assign n526 = ~\P2_IR_reg[12]/NET0131  & n525 ;
  assign n527 = ~\P2_IR_reg[7]/NET0131  & ~\P2_IR_reg[8]/NET0131  ;
  assign n528 = ~\P2_IR_reg[0]/NET0131  & ~\P2_IR_reg[1]/NET0131  ;
  assign n529 = ~\P2_IR_reg[2]/NET0131  & n528 ;
  assign n530 = ~\P2_IR_reg[3]/NET0131  & n529 ;
  assign n531 = ~\P2_IR_reg[4]/NET0131  & ~\P2_IR_reg[5]/NET0131  ;
  assign n532 = ~\P2_IR_reg[6]/NET0131  & n531 ;
  assign n533 = n530 & n532 ;
  assign n534 = n527 & n533 ;
  assign n535 = n526 & n534 ;
  assign n536 = \P2_IR_reg[31]/NET0131  & ~n535 ;
  assign n538 = ~\P2_IR_reg[14]/NET0131  & ~\P2_IR_reg[15]/NET0131  ;
  assign n539 = ~\P2_IR_reg[16]/NET0131  & n538 ;
  assign n540 = ~\P2_IR_reg[13]/NET0131  & n539 ;
  assign n541 = ~\P2_IR_reg[17]/NET0131  & ~\P2_IR_reg[18]/NET0131  ;
  assign n542 = ~\P2_IR_reg[19]/NET0131  & ~\P2_IR_reg[20]/NET0131  ;
  assign n543 = n541 & n542 ;
  assign n537 = ~\P2_IR_reg[22]/NET0131  & ~\P2_IR_reg[23]/NET0131  ;
  assign n544 = ~\P2_IR_reg[21]/NET0131  & ~\P2_IR_reg[24]/NET0131  ;
  assign n545 = n537 & n544 ;
  assign n546 = n543 & n545 ;
  assign n547 = n540 & n546 ;
  assign n548 = ~\P2_IR_reg[26]/NET0131  & ~\P2_IR_reg[27]/NET0131  ;
  assign n549 = ~\P2_IR_reg[25]/NET0131  & ~\P2_IR_reg[28]/NET0131  ;
  assign n550 = n548 & n549 ;
  assign n551 = n547 & n550 ;
  assign n552 = \P2_IR_reg[31]/NET0131  & ~n551 ;
  assign n553 = ~n536 & ~n552 ;
  assign n554 = \P2_IR_reg[29]/NET0131  & ~n553 ;
  assign n555 = ~\P2_IR_reg[29]/NET0131  & n553 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = ~\P2_IR_reg[7]/NET0131  & n533 ;
  assign n558 = ~\P2_IR_reg[13]/NET0131  & ~\P2_IR_reg[8]/NET0131  ;
  assign n559 = n526 & n558 ;
  assign n560 = n557 & n559 ;
  assign n561 = \P2_IR_reg[31]/NET0131  & ~n560 ;
  assign n563 = ~\P2_IR_reg[17]/NET0131  & n539 ;
  assign n562 = ~\P2_IR_reg[21]/NET0131  & n542 ;
  assign n564 = ~\P2_IR_reg[18]/NET0131  & n562 ;
  assign n565 = n563 & n564 ;
  assign n566 = ~\P2_IR_reg[24]/NET0131  & ~\P2_IR_reg[25]/NET0131  ;
  assign n567 = n537 & n566 ;
  assign n568 = ~\P2_IR_reg[28]/NET0131  & ~\P2_IR_reg[29]/NET0131  ;
  assign n569 = n548 & n568 ;
  assign n570 = n567 & n569 ;
  assign n571 = n565 & n570 ;
  assign n572 = \P2_IR_reg[31]/NET0131  & ~n571 ;
  assign n573 = ~n561 & ~n572 ;
  assign n574 = \P2_IR_reg[30]/NET0131  & ~n573 ;
  assign n575 = ~\P2_IR_reg[30]/NET0131  & n573 ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = n556 & ~n576 ;
  assign n578 = \P2_reg1_reg[15]/NET0131  & n577 ;
  assign n579 = ~n556 & ~n576 ;
  assign n580 = \P2_reg0_reg[15]/NET0131  & n579 ;
  assign n599 = ~n578 & ~n580 ;
  assign n581 = n556 & n576 ;
  assign n582 = ~\P2_reg3_reg[3]/NET0131  & ~\P2_reg3_reg[4]/NET0131  ;
  assign n583 = ~\P2_reg3_reg[5]/NET0131  & n582 ;
  assign n584 = ~\P2_reg3_reg[6]/NET0131  & n583 ;
  assign n585 = ~\P2_reg3_reg[7]/NET0131  & n584 ;
  assign n586 = ~\P2_reg3_reg[8]/NET0131  & ~\P2_reg3_reg[9]/NET0131  ;
  assign n587 = n585 & n586 ;
  assign n588 = ~\P2_reg3_reg[10]/NET0131  & n587 ;
  assign n589 = ~\P2_reg3_reg[11]/NET0131  & ~\P2_reg3_reg[12]/NET0131  ;
  assign n590 = ~\P2_reg3_reg[13]/NET0131  & ~\P2_reg3_reg[14]/NET0131  ;
  assign n591 = n589 & n590 ;
  assign n592 = n588 & n591 ;
  assign n593 = ~\P2_reg3_reg[15]/NET0131  & n592 ;
  assign n594 = \P2_reg3_reg[15]/NET0131  & ~n592 ;
  assign n595 = ~n593 & ~n594 ;
  assign n596 = n581 & ~n595 ;
  assign n597 = ~n556 & n576 ;
  assign n598 = \P2_reg2_reg[15]/NET0131  & n597 ;
  assign n600 = ~n596 & ~n598 ;
  assign n601 = n599 & n600 ;
  assign n602 = n538 & n559 ;
  assign n603 = n557 & n602 ;
  assign n604 = ~\P2_IR_reg[22]/NET0131  & n562 ;
  assign n605 = ~\P2_IR_reg[16]/NET0131  & n541 ;
  assign n606 = ~\P2_IR_reg[23]/NET0131  & n605 ;
  assign n607 = n604 & n606 ;
  assign n608 = n603 & n607 ;
  assign n609 = \P2_IR_reg[31]/NET0131  & ~n608 ;
  assign n610 = n548 & n566 ;
  assign n611 = \P2_IR_reg[31]/NET0131  & ~n610 ;
  assign n612 = ~n609 & ~n611 ;
  assign n613 = \P2_IR_reg[28]/NET0131  & ~n612 ;
  assign n614 = ~\P2_IR_reg[28]/NET0131  & n612 ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = ~\P2_IR_reg[9]/NET0131  & n527 ;
  assign n617 = ~\P2_IR_reg[10]/NET0131  & n616 ;
  assign n618 = n533 & n617 ;
  assign n619 = ~\P2_IR_reg[11]/NET0131  & ~\P2_IR_reg[12]/NET0131  ;
  assign n620 = ~\P2_IR_reg[13]/NET0131  & ~\P2_IR_reg[14]/NET0131  ;
  assign n621 = n619 & n620 ;
  assign n622 = n618 & n621 ;
  assign n623 = ~\P2_IR_reg[15]/NET0131  & n605 ;
  assign n624 = n622 & n623 ;
  assign n625 = \P2_IR_reg[31]/NET0131  & ~n624 ;
  assign n626 = ~\P2_IR_reg[23]/NET0131  & ~\P2_IR_reg[26]/NET0131  ;
  assign n627 = n566 & n626 ;
  assign n628 = n604 & n627 ;
  assign n629 = \P2_IR_reg[31]/NET0131  & ~n628 ;
  assign n630 = ~n625 & ~n629 ;
  assign n631 = \P2_IR_reg[27]/NET0131  & ~n630 ;
  assign n632 = ~\P2_IR_reg[27]/NET0131  & n630 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = ~n615 & ~n633 ;
  assign n635 = ~\P1_addr_reg[19]/NET0131  & ~\P2_addr_reg[19]/NET0131  ;
  assign n636 = ~\P1_rd_reg/NET0131  & n635 ;
  assign n637 = \P1_addr_reg[19]/NET0131  & \P2_addr_reg[19]/NET0131  ;
  assign n638 = ~\P2_rd_reg/NET0131  & n637 ;
  assign n639 = ~n636 & ~n638 ;
  assign n640 = \P1_datao_reg[15]/NET0131  & ~n639 ;
  assign n654 = ~\P1_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n655 = \P1_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n656 = \P1_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n657 = ~n655 & ~n656 ;
  assign n658 = ~n654 & ~n657 ;
  assign n659 = ~\P1_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n660 = ~\P1_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n661 = \P1_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n662 = ~\P1_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n663 = n661 & ~n662 ;
  assign n664 = \P1_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n665 = \P1_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = ~n663 & n666 ;
  assign n668 = ~n660 & ~n667 ;
  assign n669 = ~n659 & n668 ;
  assign n670 = \P1_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n671 = \P1_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n672 = ~n670 & ~n671 ;
  assign n673 = ~n669 & n672 ;
  assign n674 = ~\P1_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n675 = ~\P1_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = ~n654 & n676 ;
  assign n678 = ~n673 & n677 ;
  assign n679 = ~n658 & ~n678 ;
  assign n646 = ~\P1_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n641 = ~\P1_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n647 = ~\P1_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n648 = ~n641 & ~n647 ;
  assign n649 = ~n646 & n648 ;
  assign n680 = ~\P1_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n681 = n649 & ~n680 ;
  assign n682 = ~n679 & n681 ;
  assign n642 = \P1_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n643 = \P1_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = ~n641 & ~n644 ;
  assign n650 = \P1_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n651 = \P1_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n652 = ~n650 & ~n651 ;
  assign n653 = n649 & ~n652 ;
  assign n683 = ~n645 & ~n653 ;
  assign n684 = ~n682 & n683 ;
  assign n685 = ~\P1_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n686 = ~\P1_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n687 = ~n685 & ~n686 ;
  assign n688 = ~\P1_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n689 = ~\P1_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = n687 & n690 ;
  assign n692 = ~n684 & n691 ;
  assign n693 = \P1_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n694 = \P1_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n695 = ~n693 & ~n694 ;
  assign n696 = ~n688 & ~n695 ;
  assign n697 = \P1_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n698 = \P1_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n699 = ~n697 & ~n698 ;
  assign n700 = ~n685 & n690 ;
  assign n701 = ~n699 & n700 ;
  assign n702 = ~n696 & ~n701 ;
  assign n703 = ~n692 & n702 ;
  assign n704 = ~\P1_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n705 = \P1_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n706 = ~n704 & ~n705 ;
  assign n708 = ~n703 & n706 ;
  assign n707 = n703 & ~n706 ;
  assign n709 = n639 & ~n707 ;
  assign n710 = ~n708 & n709 ;
  assign n711 = ~n640 & ~n710 ;
  assign n712 = ~n634 & ~n711 ;
  assign n713 = \P2_IR_reg[31]/NET0131  & ~n622 ;
  assign n714 = \P2_IR_reg[15]/NET0131  & n713 ;
  assign n715 = ~\P2_IR_reg[15]/NET0131  & ~n713 ;
  assign n716 = ~n714 & ~n715 ;
  assign n717 = n634 & n716 ;
  assign n718 = ~n712 & ~n717 ;
  assign n719 = n601 & ~n718 ;
  assign n720 = \P1_datao_reg[14]/NET0131  & ~n639 ;
  assign n721 = ~n693 & ~n697 ;
  assign n722 = ~n642 & ~n698 ;
  assign n723 = n687 & ~n722 ;
  assign n724 = n721 & ~n723 ;
  assign n725 = ~n689 & ~n724 ;
  assign n726 = ~n663 & ~n664 ;
  assign n727 = ~n660 & ~n726 ;
  assign n728 = ~n665 & ~n671 ;
  assign n729 = ~n727 & n728 ;
  assign n730 = ~n659 & ~n729 ;
  assign n731 = n676 & n730 ;
  assign n732 = ~n655 & ~n670 ;
  assign n733 = ~n675 & ~n732 ;
  assign n734 = ~n731 & ~n733 ;
  assign n735 = ~n646 & ~n680 ;
  assign n736 = ~n647 & n735 ;
  assign n737 = ~n654 & n736 ;
  assign n738 = ~n734 & n737 ;
  assign n739 = ~n643 & ~n650 ;
  assign n740 = ~n647 & ~n739 ;
  assign n741 = ~n651 & ~n656 ;
  assign n742 = n736 & ~n741 ;
  assign n743 = ~n740 & ~n742 ;
  assign n744 = ~n738 & n743 ;
  assign n745 = ~n641 & ~n689 ;
  assign n746 = n687 & n745 ;
  assign n747 = ~n744 & n746 ;
  assign n748 = ~n725 & ~n747 ;
  assign n749 = ~n688 & ~n694 ;
  assign n751 = ~n748 & n749 ;
  assign n750 = n748 & ~n749 ;
  assign n752 = n639 & ~n750 ;
  assign n753 = ~n751 & n752 ;
  assign n754 = ~n720 & ~n753 ;
  assign n755 = ~n634 & ~n754 ;
  assign n756 = ~\P2_IR_reg[14]/NET0131  & ~n561 ;
  assign n757 = \P2_IR_reg[14]/NET0131  & n561 ;
  assign n758 = ~n756 & ~n757 ;
  assign n759 = n634 & n758 ;
  assign n760 = ~n755 & ~n759 ;
  assign n761 = \P2_reg2_reg[14]/NET0131  & n597 ;
  assign n762 = \P2_reg0_reg[14]/NET0131  & n579 ;
  assign n770 = ~n761 & ~n762 ;
  assign n763 = ~\P2_reg3_reg[11]/NET0131  & n588 ;
  assign n764 = ~\P2_reg3_reg[12]/NET0131  & n763 ;
  assign n765 = ~\P2_reg3_reg[13]/NET0131  & n764 ;
  assign n766 = \P2_reg3_reg[14]/NET0131  & ~n765 ;
  assign n767 = ~n592 & ~n766 ;
  assign n768 = n581 & ~n767 ;
  assign n769 = \P2_reg1_reg[14]/NET0131  & n577 ;
  assign n771 = ~n768 & ~n769 ;
  assign n772 = n770 & n771 ;
  assign n773 = ~n760 & n772 ;
  assign n774 = ~n719 & ~n773 ;
  assign n775 = \P2_reg1_reg[13]/NET0131  & n577 ;
  assign n776 = \P2_reg3_reg[13]/NET0131  & ~n764 ;
  assign n777 = ~n765 & ~n776 ;
  assign n778 = n581 & ~n777 ;
  assign n781 = ~n775 & ~n778 ;
  assign n779 = \P2_reg0_reg[13]/NET0131  & n579 ;
  assign n780 = \P2_reg2_reg[13]/NET0131  & n597 ;
  assign n782 = ~n779 & ~n780 ;
  assign n783 = n781 & n782 ;
  assign n784 = \P1_datao_reg[13]/NET0131  & ~n639 ;
  assign n787 = ~n673 & ~n674 ;
  assign n788 = ~n654 & ~n680 ;
  assign n789 = ~n646 & ~n675 ;
  assign n790 = n788 & n789 ;
  assign n791 = n787 & n790 ;
  assign n785 = ~n651 & ~n658 ;
  assign n786 = n735 & ~n785 ;
  assign n792 = ~n650 & ~n786 ;
  assign n793 = ~n791 & n792 ;
  assign n794 = n648 & n687 ;
  assign n795 = ~n793 & n794 ;
  assign n796 = ~n645 & ~n698 ;
  assign n797 = n687 & ~n796 ;
  assign n798 = ~n697 & ~n797 ;
  assign n799 = ~n795 & n798 ;
  assign n800 = ~n689 & ~n693 ;
  assign n802 = ~n799 & n800 ;
  assign n801 = n799 & ~n800 ;
  assign n803 = n639 & ~n801 ;
  assign n804 = ~n802 & n803 ;
  assign n805 = ~n784 & ~n804 ;
  assign n806 = ~n634 & ~n805 ;
  assign n807 = ~\P2_IR_reg[13]/NET0131  & ~n536 ;
  assign n808 = \P2_IR_reg[13]/NET0131  & n536 ;
  assign n809 = ~n807 & ~n808 ;
  assign n810 = n634 & n809 ;
  assign n811 = ~n806 & ~n810 ;
  assign n812 = n783 & ~n811 ;
  assign n813 = ~n783 & n811 ;
  assign n814 = \P2_reg3_reg[12]/NET0131  & ~n763 ;
  assign n815 = ~n764 & ~n814 ;
  assign n816 = n581 & ~n815 ;
  assign n817 = \P2_reg0_reg[12]/NET0131  & n579 ;
  assign n820 = ~n816 & ~n817 ;
  assign n818 = \P2_reg2_reg[12]/NET0131  & n597 ;
  assign n819 = \P2_reg1_reg[12]/NET0131  & n577 ;
  assign n821 = ~n818 & ~n819 ;
  assign n822 = n820 & n821 ;
  assign n823 = \P1_datao_reg[12]/NET0131  & ~n639 ;
  assign n824 = ~n685 & ~n697 ;
  assign n825 = n731 & n788 ;
  assign n826 = ~n656 & ~n733 ;
  assign n827 = n788 & ~n826 ;
  assign n828 = ~n651 & ~n827 ;
  assign n829 = ~n825 & n828 ;
  assign n830 = n649 & ~n686 ;
  assign n831 = ~n829 & n830 ;
  assign n832 = ~n642 & ~n740 ;
  assign n833 = ~n641 & ~n686 ;
  assign n834 = ~n832 & n833 ;
  assign n835 = ~n698 & ~n834 ;
  assign n836 = ~n831 & n835 ;
  assign n838 = ~n824 & n836 ;
  assign n837 = n824 & ~n836 ;
  assign n839 = n639 & ~n837 ;
  assign n840 = ~n838 & n839 ;
  assign n841 = ~n823 & ~n840 ;
  assign n842 = ~n634 & ~n841 ;
  assign n843 = \P2_IR_reg[31]/NET0131  & ~n534 ;
  assign n844 = \P2_IR_reg[31]/NET0131  & ~n525 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = \P2_IR_reg[12]/NET0131  & ~n845 ;
  assign n847 = ~\P2_IR_reg[12]/NET0131  & n845 ;
  assign n848 = ~n846 & ~n847 ;
  assign n849 = n634 & n848 ;
  assign n850 = ~n842 & ~n849 ;
  assign n851 = ~n822 & n850 ;
  assign n852 = ~n813 & ~n851 ;
  assign n853 = ~n812 & ~n852 ;
  assign n854 = n774 & n853 ;
  assign n855 = ~n601 & n718 ;
  assign n856 = n760 & ~n772 ;
  assign n857 = ~n855 & ~n856 ;
  assign n858 = ~n719 & ~n857 ;
  assign n859 = ~n854 & ~n858 ;
  assign n860 = \P2_reg3_reg[11]/NET0131  & ~n588 ;
  assign n861 = ~n763 & ~n860 ;
  assign n862 = n581 & ~n861 ;
  assign n863 = \P2_reg0_reg[11]/NET0131  & n579 ;
  assign n866 = ~n862 & ~n863 ;
  assign n864 = \P2_reg2_reg[11]/NET0131  & n597 ;
  assign n865 = \P2_reg1_reg[11]/NET0131  & n577 ;
  assign n867 = ~n864 & ~n865 ;
  assign n868 = n866 & n867 ;
  assign n869 = \P1_datao_reg[11]/NET0131  & ~n639 ;
  assign n870 = ~n686 & ~n698 ;
  assign n872 = n684 & ~n870 ;
  assign n871 = ~n684 & n870 ;
  assign n873 = n639 & ~n871 ;
  assign n874 = ~n872 & n873 ;
  assign n875 = ~n869 & ~n874 ;
  assign n876 = ~n634 & ~n875 ;
  assign n877 = \P2_IR_reg[31]/NET0131  & ~n618 ;
  assign n878 = \P2_IR_reg[11]/NET0131  & n877 ;
  assign n879 = ~\P2_IR_reg[11]/NET0131  & ~n877 ;
  assign n880 = ~n878 & ~n879 ;
  assign n881 = n634 & n880 ;
  assign n882 = ~n876 & ~n881 ;
  assign n883 = ~n868 & n882 ;
  assign n884 = n868 & ~n882 ;
  assign n885 = \P2_reg1_reg[10]/NET0131  & n577 ;
  assign n886 = \P2_reg2_reg[10]/NET0131  & n597 ;
  assign n891 = ~n885 & ~n886 ;
  assign n887 = \P2_reg3_reg[10]/NET0131  & ~n587 ;
  assign n888 = ~n588 & ~n887 ;
  assign n889 = n581 & ~n888 ;
  assign n890 = \P2_reg0_reg[10]/NET0131  & n579 ;
  assign n892 = ~n889 & ~n890 ;
  assign n893 = n891 & n892 ;
  assign n894 = \P1_datao_reg[10]/NET0131  & ~n639 ;
  assign n895 = ~n641 & ~n642 ;
  assign n897 = n744 & ~n895 ;
  assign n896 = ~n744 & n895 ;
  assign n898 = n639 & ~n896 ;
  assign n899 = ~n897 & n898 ;
  assign n900 = ~n894 & ~n899 ;
  assign n901 = ~n634 & ~n900 ;
  assign n902 = \P2_IR_reg[31]/NET0131  & ~n533 ;
  assign n903 = \P2_IR_reg[31]/NET0131  & ~n616 ;
  assign n904 = ~n902 & ~n903 ;
  assign n905 = \P2_IR_reg[10]/NET0131  & ~n904 ;
  assign n906 = ~\P2_IR_reg[10]/NET0131  & n904 ;
  assign n907 = ~n905 & ~n906 ;
  assign n908 = n634 & n907 ;
  assign n909 = ~n901 & ~n908 ;
  assign n910 = n893 & ~n909 ;
  assign n911 = ~n884 & ~n910 ;
  assign n912 = \P2_reg0_reg[9]/NET0131  & n579 ;
  assign n913 = ~\P2_reg3_reg[8]/NET0131  & n585 ;
  assign n914 = \P2_reg3_reg[9]/NET0131  & ~n913 ;
  assign n915 = ~n587 & ~n914 ;
  assign n916 = n581 & ~n915 ;
  assign n919 = ~n912 & ~n916 ;
  assign n917 = \P2_reg1_reg[9]/NET0131  & n577 ;
  assign n918 = \P2_reg2_reg[9]/NET0131  & n597 ;
  assign n920 = ~n917 & ~n918 ;
  assign n921 = n919 & n920 ;
  assign n922 = \P1_datao_reg[9]/NET0131  & ~n639 ;
  assign n923 = ~n643 & ~n647 ;
  assign n925 = n793 & ~n923 ;
  assign n924 = ~n793 & n923 ;
  assign n926 = n639 & ~n924 ;
  assign n927 = ~n925 & n926 ;
  assign n928 = ~n922 & ~n927 ;
  assign n929 = ~n634 & ~n928 ;
  assign n930 = \P2_IR_reg[9]/NET0131  & ~n843 ;
  assign n931 = ~\P2_IR_reg[9]/NET0131  & n843 ;
  assign n932 = ~n930 & ~n931 ;
  assign n933 = n634 & ~n932 ;
  assign n934 = ~n929 & ~n933 ;
  assign n935 = n921 & ~n934 ;
  assign n936 = \P2_reg2_reg[8]/NET0131  & n597 ;
  assign n937 = \P2_reg0_reg[8]/NET0131  & n579 ;
  assign n942 = ~n936 & ~n937 ;
  assign n938 = \P2_reg3_reg[8]/NET0131  & ~n585 ;
  assign n939 = ~n913 & ~n938 ;
  assign n940 = n581 & ~n939 ;
  assign n941 = \P2_reg1_reg[8]/NET0131  & n577 ;
  assign n943 = ~n940 & ~n941 ;
  assign n944 = n942 & n943 ;
  assign n945 = \P1_datao_reg[8]/NET0131  & ~n639 ;
  assign n946 = ~n646 & ~n650 ;
  assign n948 = n829 & ~n946 ;
  assign n947 = ~n829 & n946 ;
  assign n949 = n639 & ~n947 ;
  assign n950 = ~n948 & n949 ;
  assign n951 = ~n945 & ~n950 ;
  assign n952 = ~n634 & ~n951 ;
  assign n953 = \P2_IR_reg[31]/NET0131  & ~n557 ;
  assign n954 = ~\P2_IR_reg[8]/NET0131  & ~n953 ;
  assign n955 = \P2_IR_reg[8]/NET0131  & n953 ;
  assign n956 = ~n954 & ~n955 ;
  assign n957 = n634 & n956 ;
  assign n958 = ~n952 & ~n957 ;
  assign n959 = n944 & ~n958 ;
  assign n960 = ~n935 & ~n959 ;
  assign n961 = ~n921 & n934 ;
  assign n962 = ~n893 & n909 ;
  assign n963 = ~n961 & ~n962 ;
  assign n964 = ~n960 & n963 ;
  assign n965 = n911 & ~n964 ;
  assign n966 = ~n883 & ~n965 ;
  assign n967 = n822 & ~n850 ;
  assign n968 = ~n812 & ~n967 ;
  assign n969 = ~n813 & ~n856 ;
  assign n970 = ~n968 & n969 ;
  assign n971 = n774 & ~n970 ;
  assign n972 = ~n855 & ~n971 ;
  assign n973 = ~n966 & ~n972 ;
  assign n974 = n859 & ~n973 ;
  assign n978 = \P2_reg0_reg[6]/NET0131  & n579 ;
  assign n979 = \P2_reg2_reg[6]/NET0131  & n597 ;
  assign n984 = ~n978 & ~n979 ;
  assign n980 = \P2_reg3_reg[6]/NET0131  & ~n583 ;
  assign n981 = ~n584 & ~n980 ;
  assign n982 = n581 & ~n981 ;
  assign n983 = \P2_reg1_reg[6]/NET0131  & n577 ;
  assign n985 = ~n982 & ~n983 ;
  assign n986 = n984 & n985 ;
  assign n987 = \P1_datao_reg[6]/NET0131  & ~n639 ;
  assign n988 = ~n654 & ~n656 ;
  assign n990 = n734 & ~n988 ;
  assign n989 = ~n734 & n988 ;
  assign n991 = n639 & ~n989 ;
  assign n992 = ~n990 & n991 ;
  assign n993 = ~n987 & ~n992 ;
  assign n994 = ~n634 & ~n993 ;
  assign n995 = ~\P2_IR_reg[4]/NET0131  & n530 ;
  assign n996 = \P2_IR_reg[31]/NET0131  & ~n995 ;
  assign n997 = \P2_IR_reg[31]/NET0131  & \P2_IR_reg[5]/NET0131  ;
  assign n998 = ~n996 & ~n997 ;
  assign n999 = \P2_IR_reg[6]/NET0131  & ~n998 ;
  assign n1000 = ~\P2_IR_reg[6]/NET0131  & n998 ;
  assign n1001 = ~n999 & ~n1000 ;
  assign n1002 = n634 & n1001 ;
  assign n1003 = ~n994 & ~n1002 ;
  assign n1004 = n986 & ~n1003 ;
  assign n1005 = \P2_reg0_reg[7]/NET0131  & n579 ;
  assign n1006 = \P2_reg3_reg[7]/NET0131  & ~n584 ;
  assign n1007 = ~n585 & ~n1006 ;
  assign n1008 = n581 & ~n1007 ;
  assign n1011 = ~n1005 & ~n1008 ;
  assign n1009 = \P2_reg2_reg[7]/NET0131  & n597 ;
  assign n1010 = \P2_reg1_reg[7]/NET0131  & n577 ;
  assign n1012 = ~n1009 & ~n1010 ;
  assign n1013 = n1011 & n1012 ;
  assign n1014 = \P1_datao_reg[7]/NET0131  & ~n639 ;
  assign n1015 = ~n651 & ~n680 ;
  assign n1017 = n679 & ~n1015 ;
  assign n1016 = ~n679 & n1015 ;
  assign n1018 = n639 & ~n1016 ;
  assign n1019 = ~n1017 & n1018 ;
  assign n1020 = ~n1014 & ~n1019 ;
  assign n1021 = ~n634 & ~n1020 ;
  assign n1022 = ~\P2_IR_reg[7]/NET0131  & ~n902 ;
  assign n1023 = \P2_IR_reg[7]/NET0131  & n902 ;
  assign n1024 = ~n1022 & ~n1023 ;
  assign n1025 = n634 & n1024 ;
  assign n1026 = ~n1021 & ~n1025 ;
  assign n1027 = n1013 & ~n1026 ;
  assign n1028 = ~n1004 & ~n1027 ;
  assign n1029 = \P2_reg3_reg[5]/NET0131  & ~n582 ;
  assign n1030 = ~n583 & ~n1029 ;
  assign n1031 = n581 & ~n1030 ;
  assign n1032 = \P2_reg0_reg[5]/NET0131  & n579 ;
  assign n1035 = ~n1031 & ~n1032 ;
  assign n1033 = \P2_reg1_reg[5]/NET0131  & n577 ;
  assign n1034 = \P2_reg2_reg[5]/NET0131  & n597 ;
  assign n1036 = ~n1033 & ~n1034 ;
  assign n1037 = n1035 & n1036 ;
  assign n1038 = \P1_datao_reg[5]/NET0131  & ~n639 ;
  assign n1039 = ~n655 & ~n675 ;
  assign n1041 = n787 & n1039 ;
  assign n1040 = ~n787 & ~n1039 ;
  assign n1042 = n639 & ~n1040 ;
  assign n1043 = ~n1041 & n1042 ;
  assign n1044 = ~n1038 & ~n1043 ;
  assign n1045 = ~n634 & ~n1044 ;
  assign n1046 = \P2_IR_reg[5]/NET0131  & ~n996 ;
  assign n1047 = ~\P2_IR_reg[5]/NET0131  & n996 ;
  assign n1048 = ~n1046 & ~n1047 ;
  assign n1049 = n634 & ~n1048 ;
  assign n1050 = ~n1045 & ~n1049 ;
  assign n1051 = ~n1037 & n1050 ;
  assign n1052 = ~n986 & n1003 ;
  assign n1053 = ~n1051 & ~n1052 ;
  assign n1054 = \P2_reg3_reg[3]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n1055 = ~n582 & ~n1054 ;
  assign n1056 = n581 & ~n1055 ;
  assign n1057 = \P2_reg0_reg[4]/NET0131  & n579 ;
  assign n1060 = ~n1056 & ~n1057 ;
  assign n1058 = \P2_reg1_reg[4]/NET0131  & n577 ;
  assign n1059 = \P2_reg2_reg[4]/NET0131  & n597 ;
  assign n1061 = ~n1058 & ~n1059 ;
  assign n1062 = n1060 & n1061 ;
  assign n1063 = \P1_datao_reg[4]/NET0131  & ~n639 ;
  assign n1064 = ~n670 & ~n674 ;
  assign n1066 = n730 & n1064 ;
  assign n1065 = ~n730 & ~n1064 ;
  assign n1067 = n639 & ~n1065 ;
  assign n1068 = ~n1066 & n1067 ;
  assign n1069 = ~n1063 & ~n1068 ;
  assign n1070 = ~n634 & ~n1069 ;
  assign n1071 = \P2_IR_reg[31]/NET0131  & ~n530 ;
  assign n1072 = \P2_IR_reg[4]/NET0131  & n1071 ;
  assign n1073 = ~\P2_IR_reg[4]/NET0131  & ~n1071 ;
  assign n1074 = ~n1072 & ~n1073 ;
  assign n1075 = n634 & n1074 ;
  assign n1076 = ~n1070 & ~n1075 ;
  assign n1077 = n1062 & ~n1076 ;
  assign n1078 = n1037 & ~n1050 ;
  assign n1079 = ~n1077 & ~n1078 ;
  assign n1080 = \P2_reg0_reg[3]/NET0131  & n579 ;
  assign n1081 = \P2_reg2_reg[3]/NET0131  & n597 ;
  assign n1084 = ~n1080 & ~n1081 ;
  assign n1082 = ~\P2_reg3_reg[3]/NET0131  & n581 ;
  assign n1083 = \P2_reg1_reg[3]/NET0131  & n577 ;
  assign n1085 = ~n1082 & ~n1083 ;
  assign n1086 = n1084 & n1085 ;
  assign n1087 = \P2_IR_reg[31]/NET0131  & ~n529 ;
  assign n1088 = \P2_IR_reg[3]/NET0131  & n1087 ;
  assign n1089 = ~\P2_IR_reg[3]/NET0131  & ~n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1091 = n634 & n1090 ;
  assign n1092 = ~\P1_datao_reg[3]/NET0131  & ~n639 ;
  assign n1093 = ~n659 & ~n671 ;
  assign n1095 = n668 & ~n1093 ;
  assign n1094 = ~n668 & n1093 ;
  assign n1096 = n639 & ~n1094 ;
  assign n1097 = ~n1095 & n1096 ;
  assign n1098 = ~n1092 & ~n1097 ;
  assign n1099 = ~n634 & n1098 ;
  assign n1100 = ~n1091 & ~n1099 ;
  assign n1101 = ~n1086 & n1100 ;
  assign n1102 = ~n1062 & n1076 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = \P2_reg2_reg[2]/NET0131  & n597 ;
  assign n1105 = \P2_reg0_reg[2]/NET0131  & n579 ;
  assign n1108 = ~n1104 & ~n1105 ;
  assign n1106 = \P2_reg3_reg[2]/NET0131  & n581 ;
  assign n1107 = \P2_reg1_reg[2]/NET0131  & n577 ;
  assign n1109 = ~n1106 & ~n1107 ;
  assign n1110 = n1108 & n1109 ;
  assign n1111 = \P1_datao_reg[2]/NET0131  & ~n639 ;
  assign n1112 = ~n660 & ~n665 ;
  assign n1114 = ~n726 & n1112 ;
  assign n1113 = n726 & ~n1112 ;
  assign n1115 = n639 & ~n1113 ;
  assign n1116 = ~n1114 & n1115 ;
  assign n1117 = ~n1111 & ~n1116 ;
  assign n1118 = ~n634 & ~n1117 ;
  assign n1119 = \P2_IR_reg[31]/NET0131  & ~n528 ;
  assign n1120 = ~\P2_IR_reg[2]/NET0131  & n1119 ;
  assign n1121 = \P2_IR_reg[2]/NET0131  & ~n1119 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = n634 & ~n1122 ;
  assign n1124 = ~n1118 & ~n1123 ;
  assign n1125 = n1110 & ~n1124 ;
  assign n1126 = n1086 & ~n1100 ;
  assign n1127 = ~n1125 & ~n1126 ;
  assign n1128 = \P2_reg1_reg[1]/NET0131  & n577 ;
  assign n1129 = \P2_reg3_reg[1]/NET0131  & n581 ;
  assign n1132 = ~n1128 & ~n1129 ;
  assign n1130 = \P2_reg2_reg[1]/NET0131  & n597 ;
  assign n1131 = \P2_reg0_reg[1]/NET0131  & n579 ;
  assign n1133 = ~n1130 & ~n1131 ;
  assign n1134 = n1132 & n1133 ;
  assign n1135 = \P2_IR_reg[0]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n1136 = ~\P2_IR_reg[1]/NET0131  & n1135 ;
  assign n1137 = \P2_IR_reg[1]/NET0131  & ~n1135 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = n634 & ~n1138 ;
  assign n1140 = ~\P1_datao_reg[1]/NET0131  & ~n639 ;
  assign n1141 = ~n662 & ~n664 ;
  assign n1143 = n661 & ~n1141 ;
  assign n1142 = ~n661 & n1141 ;
  assign n1144 = n639 & ~n1142 ;
  assign n1145 = ~n1143 & n1144 ;
  assign n1146 = ~n1140 & ~n1145 ;
  assign n1147 = ~n634 & n1146 ;
  assign n1148 = ~n1139 & ~n1147 ;
  assign n1151 = n1134 & ~n1148 ;
  assign n1152 = \P2_reg3_reg[0]/NET0131  & n581 ;
  assign n1153 = \P2_reg2_reg[0]/NET0131  & n597 ;
  assign n1156 = ~n1152 & ~n1153 ;
  assign n1154 = \P2_reg1_reg[0]/NET0131  & n577 ;
  assign n1155 = \P2_reg0_reg[0]/NET0131  & n579 ;
  assign n1157 = ~n1154 & ~n1155 ;
  assign n1158 = n1156 & n1157 ;
  assign n1159 = \si[0]_pad  & n639 ;
  assign n1160 = ~\P1_datao_reg[0]/NET0131  & ~n1159 ;
  assign n1161 = \P1_datao_reg[0]/NET0131  & n1159 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = ~n634 & n1162 ;
  assign n1164 = \P2_IR_reg[0]/NET0131  & n634 ;
  assign n1165 = ~n1163 & ~n1164 ;
  assign n1166 = ~n1158 & n1165 ;
  assign n1167 = ~n1151 & n1166 ;
  assign n1149 = ~n1134 & n1148 ;
  assign n1150 = ~n1110 & n1124 ;
  assign n1168 = ~n1149 & ~n1150 ;
  assign n1169 = ~n1167 & n1168 ;
  assign n1170 = n1127 & ~n1169 ;
  assign n1171 = n1103 & ~n1170 ;
  assign n1172 = n1079 & ~n1171 ;
  assign n1173 = n1053 & ~n1172 ;
  assign n1174 = n1028 & ~n1173 ;
  assign n975 = ~n883 & ~n962 ;
  assign n976 = ~n944 & n958 ;
  assign n977 = ~n961 & ~n976 ;
  assign n1175 = ~n1013 & n1026 ;
  assign n1176 = n977 & ~n1175 ;
  assign n1177 = n975 & n1176 ;
  assign n1178 = n852 & n1177 ;
  assign n1179 = n857 & n1178 ;
  assign n1180 = ~n1174 & n1179 ;
  assign n1181 = ~n974 & ~n1180 ;
  assign n1182 = \P2_reg2_reg[17]/NET0131  & n597 ;
  assign n1183 = \P2_reg0_reg[17]/NET0131  & n579 ;
  assign n1191 = ~n1182 & ~n1183 ;
  assign n1184 = ~\P2_reg3_reg[15]/NET0131  & ~\P2_reg3_reg[16]/NET0131  ;
  assign n1185 = n592 & n1184 ;
  assign n1186 = ~\P2_reg3_reg[17]/NET0131  & n1185 ;
  assign n1187 = \P2_reg3_reg[17]/NET0131  & ~n1185 ;
  assign n1188 = ~n1186 & ~n1187 ;
  assign n1189 = n581 & ~n1188 ;
  assign n1190 = \P2_reg1_reg[17]/NET0131  & n577 ;
  assign n1192 = ~n1189 & ~n1190 ;
  assign n1193 = n1191 & n1192 ;
  assign n1194 = \P1_datao_reg[17]/NET0131  & ~n639 ;
  assign n1195 = ~\P1_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n1196 = \P1_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n1197 = ~n1195 & ~n1196 ;
  assign n1198 = ~\P1_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n1199 = ~n704 & ~n1198 ;
  assign n1200 = n690 & n1199 ;
  assign n1201 = n795 & n1200 ;
  assign n1202 = \P1_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n1203 = ~n696 & ~n705 ;
  assign n1204 = n1199 & ~n1203 ;
  assign n1205 = ~n1202 & ~n1204 ;
  assign n1206 = ~n798 & n1200 ;
  assign n1207 = n1205 & ~n1206 ;
  assign n1208 = ~n1201 & n1207 ;
  assign n1210 = ~n1197 & n1208 ;
  assign n1209 = n1197 & ~n1208 ;
  assign n1211 = n639 & ~n1209 ;
  assign n1212 = ~n1210 & n1211 ;
  assign n1213 = ~n1194 & ~n1212 ;
  assign n1214 = ~n634 & ~n1213 ;
  assign n1215 = n535 & n540 ;
  assign n1216 = \P2_IR_reg[31]/NET0131  & ~n1215 ;
  assign n1217 = ~\P2_IR_reg[17]/NET0131  & ~n1216 ;
  assign n1218 = \P2_IR_reg[17]/NET0131  & n1216 ;
  assign n1219 = ~n1217 & ~n1218 ;
  assign n1220 = n634 & n1219 ;
  assign n1221 = ~n1214 & ~n1220 ;
  assign n1222 = ~n1193 & n1221 ;
  assign n1223 = \P2_reg2_reg[16]/NET0131  & n597 ;
  assign n1224 = \P2_reg1_reg[16]/NET0131  & n577 ;
  assign n1229 = ~n1223 & ~n1224 ;
  assign n1225 = \P2_reg3_reg[16]/NET0131  & ~n593 ;
  assign n1226 = ~n1185 & ~n1225 ;
  assign n1227 = n581 & ~n1226 ;
  assign n1228 = \P2_reg0_reg[16]/NET0131  & n579 ;
  assign n1230 = ~n1227 & ~n1228 ;
  assign n1231 = n1229 & n1230 ;
  assign n1232 = \P1_datao_reg[16]/NET0131  & ~n639 ;
  assign n1233 = n690 & ~n704 ;
  assign n1234 = ~n685 & n1233 ;
  assign n1235 = n831 & n1234 ;
  assign n1236 = ~n694 & ~n705 ;
  assign n1237 = ~n704 & ~n1236 ;
  assign n1238 = ~n685 & ~n835 ;
  assign n1239 = n721 & ~n1238 ;
  assign n1240 = n1233 & ~n1239 ;
  assign n1241 = ~n1237 & ~n1240 ;
  assign n1242 = ~n1235 & n1241 ;
  assign n1243 = ~n1198 & ~n1202 ;
  assign n1245 = ~n1242 & n1243 ;
  assign n1244 = n1242 & ~n1243 ;
  assign n1246 = n639 & ~n1244 ;
  assign n1247 = ~n1245 & n1246 ;
  assign n1248 = ~n1232 & ~n1247 ;
  assign n1249 = ~n634 & ~n1248 ;
  assign n1250 = \P2_IR_reg[31]/NET0131  & ~n603 ;
  assign n1251 = ~\P2_IR_reg[16]/NET0131  & ~n1250 ;
  assign n1252 = \P2_IR_reg[16]/NET0131  & n1250 ;
  assign n1253 = ~n1251 & ~n1252 ;
  assign n1254 = n634 & n1253 ;
  assign n1255 = ~n1249 & ~n1254 ;
  assign n1256 = ~n1231 & n1255 ;
  assign n1257 = ~n1222 & ~n1256 ;
  assign n1258 = \P2_reg1_reg[19]/NET0131  & n577 ;
  assign n1259 = \P2_reg2_reg[19]/NET0131  & n597 ;
  assign n1267 = ~n1258 & ~n1259 ;
  assign n1260 = ~\P2_reg3_reg[17]/NET0131  & ~\P2_reg3_reg[18]/NET0131  ;
  assign n1261 = n1185 & n1260 ;
  assign n1262 = \P2_reg3_reg[19]/NET0131  & ~n1261 ;
  assign n1263 = ~\P2_reg3_reg[19]/NET0131  & n1261 ;
  assign n1264 = ~n1262 & ~n1263 ;
  assign n1265 = n581 & ~n1264 ;
  assign n1266 = \P2_reg0_reg[19]/NET0131  & n579 ;
  assign n1268 = ~n1265 & ~n1266 ;
  assign n1269 = n1267 & n1268 ;
  assign n1270 = \P1_datao_reg[19]/NET0131  & ~n639 ;
  assign n1271 = ~\P1_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n1272 = \P1_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = ~\P1_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n1275 = ~n1195 & ~n1274 ;
  assign n1276 = n1199 & n1275 ;
  assign n1277 = n692 & n1276 ;
  assign n1278 = ~n702 & n1276 ;
  assign n1279 = \P1_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n1280 = ~n1275 & ~n1279 ;
  assign n1281 = ~n1196 & ~n1279 ;
  assign n1282 = ~n1274 & ~n1281 ;
  assign n1283 = n705 & ~n1198 ;
  assign n1284 = ~n1202 & ~n1283 ;
  assign n1285 = ~n1282 & n1284 ;
  assign n1286 = ~n1280 & ~n1285 ;
  assign n1287 = ~n1278 & ~n1286 ;
  assign n1288 = ~n1277 & n1287 ;
  assign n1290 = ~n1273 & n1288 ;
  assign n1289 = n1273 & ~n1288 ;
  assign n1291 = n639 & ~n1289 ;
  assign n1292 = ~n1290 & n1291 ;
  assign n1293 = ~n1270 & ~n1292 ;
  assign n1294 = ~n634 & ~n1293 ;
  assign n1295 = \P2_IR_reg[19]/NET0131  & ~n625 ;
  assign n1296 = ~\P2_IR_reg[19]/NET0131  & n625 ;
  assign n1297 = ~n1295 & ~n1296 ;
  assign n1298 = n634 & ~n1297 ;
  assign n1299 = ~n1294 & ~n1298 ;
  assign n1300 = ~n1269 & n1299 ;
  assign n1301 = \P2_reg2_reg[18]/NET0131  & n597 ;
  assign n1302 = \P2_reg0_reg[18]/NET0131  & n579 ;
  assign n1307 = ~n1301 & ~n1302 ;
  assign n1303 = \P2_reg3_reg[18]/NET0131  & ~n1186 ;
  assign n1304 = ~n1261 & ~n1303 ;
  assign n1305 = n581 & ~n1304 ;
  assign n1306 = \P2_reg1_reg[18]/NET0131  & n577 ;
  assign n1308 = ~n1305 & ~n1306 ;
  assign n1309 = n1307 & n1308 ;
  assign n1310 = \P1_datao_reg[18]/NET0131  & ~n639 ;
  assign n1311 = ~n1274 & ~n1279 ;
  assign n1312 = ~n688 & ~n1195 ;
  assign n1313 = n1199 & n1312 ;
  assign n1314 = n747 & n1313 ;
  assign n1315 = ~n1195 & ~n1198 ;
  assign n1316 = ~n1202 & ~n1237 ;
  assign n1317 = n1315 & ~n1316 ;
  assign n1318 = ~n1196 & ~n1317 ;
  assign n1319 = n725 & n1313 ;
  assign n1320 = n1318 & ~n1319 ;
  assign n1321 = ~n1314 & n1320 ;
  assign n1323 = ~n1311 & n1321 ;
  assign n1322 = n1311 & ~n1321 ;
  assign n1324 = n639 & ~n1322 ;
  assign n1325 = ~n1323 & n1324 ;
  assign n1326 = ~n1310 & ~n1325 ;
  assign n1327 = ~n634 & ~n1326 ;
  assign n1328 = \P2_IR_reg[31]/NET0131  & ~n563 ;
  assign n1329 = ~n561 & ~n1328 ;
  assign n1330 = \P2_IR_reg[18]/NET0131  & ~n1329 ;
  assign n1331 = ~\P2_IR_reg[18]/NET0131  & n1329 ;
  assign n1332 = ~n1330 & ~n1331 ;
  assign n1333 = n634 & n1332 ;
  assign n1334 = ~n1327 & ~n1333 ;
  assign n1335 = ~n1309 & n1334 ;
  assign n1336 = ~n1300 & ~n1335 ;
  assign n1337 = n1257 & n1336 ;
  assign n1338 = ~n1181 & n1337 ;
  assign n1339 = n1309 & ~n1334 ;
  assign n1340 = n1269 & ~n1299 ;
  assign n1341 = ~n1339 & ~n1340 ;
  assign n1342 = n1193 & ~n1221 ;
  assign n1343 = n1231 & ~n1255 ;
  assign n1344 = ~n1342 & ~n1343 ;
  assign n1345 = ~n1222 & ~n1335 ;
  assign n1346 = ~n1344 & n1345 ;
  assign n1347 = n1341 & ~n1346 ;
  assign n1348 = ~n1300 & ~n1347 ;
  assign n1349 = ~n1338 & ~n1348 ;
  assign n1350 = \P1_datao_reg[21]/NET0131  & ~n639 ;
  assign n1351 = ~\P1_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n1352 = \P1_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = ~\P1_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n1355 = \P1_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n1356 = ~n1272 & ~n1355 ;
  assign n1357 = ~n1354 & ~n1356 ;
  assign n1358 = ~n1271 & ~n1354 ;
  assign n1359 = n1282 & n1358 ;
  assign n1360 = ~n1357 & ~n1359 ;
  assign n1361 = ~n799 & n1200 ;
  assign n1362 = n1205 & ~n1361 ;
  assign n1363 = n1275 & n1358 ;
  assign n1364 = ~n1362 & n1363 ;
  assign n1365 = n1360 & ~n1364 ;
  assign n1367 = ~n1353 & n1365 ;
  assign n1366 = n1353 & ~n1365 ;
  assign n1368 = n639 & ~n1366 ;
  assign n1369 = ~n1367 & n1368 ;
  assign n1370 = ~n1350 & ~n1369 ;
  assign n1371 = ~n634 & ~n1370 ;
  assign n1375 = ~\P2_reg3_reg[20]/NET0131  & n1263 ;
  assign n1376 = ~\P2_reg3_reg[21]/NET0131  & n1375 ;
  assign n1377 = \P2_reg3_reg[21]/NET0131  & ~n1375 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1379 = n581 & ~n1378 ;
  assign n1374 = \P2_reg2_reg[21]/NET0131  & n597 ;
  assign n1372 = \P2_reg1_reg[21]/NET0131  & n577 ;
  assign n1373 = \P2_reg0_reg[21]/NET0131  & n579 ;
  assign n1380 = ~n1372 & ~n1373 ;
  assign n1381 = ~n1374 & n1380 ;
  assign n1382 = ~n1379 & n1381 ;
  assign n1383 = ~n1371 & ~n1382 ;
  assign n1384 = \P1_datao_reg[20]/NET0131  & ~n639 ;
  assign n1385 = ~n1271 & ~n1274 ;
  assign n1386 = n1315 & n1385 ;
  assign n1387 = ~n1242 & n1386 ;
  assign n1388 = ~n1272 & ~n1279 ;
  assign n1389 = ~n1271 & ~n1388 ;
  assign n1390 = ~n1196 & ~n1202 ;
  assign n1391 = ~n1195 & n1385 ;
  assign n1392 = ~n1390 & n1391 ;
  assign n1393 = ~n1389 & ~n1392 ;
  assign n1394 = ~n1387 & n1393 ;
  assign n1395 = ~n1354 & ~n1355 ;
  assign n1397 = ~n1394 & n1395 ;
  assign n1396 = n1394 & ~n1395 ;
  assign n1398 = n639 & ~n1396 ;
  assign n1399 = ~n1397 & n1398 ;
  assign n1400 = ~n1384 & ~n1399 ;
  assign n1401 = ~n634 & ~n1400 ;
  assign n1405 = \P2_reg3_reg[20]/NET0131  & ~n1263 ;
  assign n1406 = ~n1375 & ~n1405 ;
  assign n1407 = n581 & ~n1406 ;
  assign n1404 = \P2_reg0_reg[20]/NET0131  & n579 ;
  assign n1402 = \P2_reg1_reg[20]/NET0131  & n577 ;
  assign n1403 = \P2_reg2_reg[20]/NET0131  & n597 ;
  assign n1408 = ~n1402 & ~n1403 ;
  assign n1409 = ~n1404 & n1408 ;
  assign n1410 = ~n1407 & n1409 ;
  assign n1411 = ~n1401 & ~n1410 ;
  assign n1412 = ~n1383 & ~n1411 ;
  assign n1413 = \P1_datao_reg[23]/NET0131  & ~n639 ;
  assign n1414 = ~\P1_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n1415 = \P1_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = \P1_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n1418 = ~\P1_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n1419 = ~n1351 & ~n1418 ;
  assign n1420 = ~n1352 & ~n1357 ;
  assign n1421 = n1419 & ~n1420 ;
  assign n1422 = ~n1417 & ~n1421 ;
  assign n1423 = n1358 & n1419 ;
  assign n1424 = n1286 & n1423 ;
  assign n1425 = n1422 & ~n1424 ;
  assign n1426 = n1276 & n1423 ;
  assign n1427 = ~n703 & n1426 ;
  assign n1428 = n1425 & ~n1427 ;
  assign n1430 = ~n1416 & n1428 ;
  assign n1429 = n1416 & ~n1428 ;
  assign n1431 = n639 & ~n1429 ;
  assign n1432 = ~n1430 & n1431 ;
  assign n1433 = ~n1413 & ~n1432 ;
  assign n1434 = ~n634 & ~n1433 ;
  assign n1438 = ~\P2_reg3_reg[22]/NET0131  & n1376 ;
  assign n1439 = \P2_reg3_reg[23]/NET0131  & ~n1438 ;
  assign n1440 = ~\P2_reg3_reg[23]/NET0131  & n1438 ;
  assign n1441 = ~n1439 & ~n1440 ;
  assign n1442 = n581 & ~n1441 ;
  assign n1437 = \P2_reg1_reg[23]/NET0131  & n577 ;
  assign n1435 = \P2_reg0_reg[23]/NET0131  & n579 ;
  assign n1436 = \P2_reg2_reg[23]/NET0131  & n597 ;
  assign n1443 = ~n1435 & ~n1436 ;
  assign n1444 = ~n1437 & n1443 ;
  assign n1445 = ~n1442 & n1444 ;
  assign n1446 = ~n1434 & ~n1445 ;
  assign n1447 = \P1_datao_reg[22]/NET0131  & ~n639 ;
  assign n1448 = ~n1417 & ~n1418 ;
  assign n1449 = ~n1351 & ~n1354 ;
  assign n1450 = n1389 & n1449 ;
  assign n1451 = ~n1352 & ~n1355 ;
  assign n1452 = ~n1351 & ~n1451 ;
  assign n1453 = ~n1450 & ~n1452 ;
  assign n1454 = n1385 & n1449 ;
  assign n1455 = ~n1318 & n1454 ;
  assign n1456 = n1453 & ~n1455 ;
  assign n1457 = n1313 & n1454 ;
  assign n1458 = ~n748 & n1457 ;
  assign n1459 = n1456 & ~n1458 ;
  assign n1461 = ~n1448 & n1459 ;
  assign n1460 = n1448 & ~n1459 ;
  assign n1462 = n639 & ~n1460 ;
  assign n1463 = ~n1461 & n1462 ;
  assign n1464 = ~n1447 & ~n1463 ;
  assign n1465 = ~n634 & ~n1464 ;
  assign n1469 = \P2_reg3_reg[22]/NET0131  & ~n1376 ;
  assign n1470 = ~n1438 & ~n1469 ;
  assign n1471 = n581 & ~n1470 ;
  assign n1468 = \P2_reg2_reg[22]/NET0131  & n597 ;
  assign n1466 = \P2_reg0_reg[22]/NET0131  & n579 ;
  assign n1467 = \P2_reg1_reg[22]/NET0131  & n577 ;
  assign n1472 = ~n1466 & ~n1467 ;
  assign n1473 = ~n1468 & n1472 ;
  assign n1474 = ~n1471 & n1473 ;
  assign n1475 = ~n1465 & ~n1474 ;
  assign n1476 = ~n1446 & ~n1475 ;
  assign n1477 = n1412 & n1476 ;
  assign n1478 = ~n1349 & n1477 ;
  assign n1479 = n1465 & n1474 ;
  assign n1480 = n1434 & n1445 ;
  assign n1481 = ~n1479 & ~n1480 ;
  assign n1482 = n1371 & n1382 ;
  assign n1483 = n1401 & n1410 ;
  assign n1484 = ~n1482 & ~n1483 ;
  assign n1485 = ~n1383 & ~n1475 ;
  assign n1486 = ~n1484 & n1485 ;
  assign n1487 = n1481 & ~n1486 ;
  assign n1488 = ~n1446 & ~n1487 ;
  assign n1489 = ~n1478 & ~n1488 ;
  assign n1490 = \P1_datao_reg[25]/NET0131  & ~n639 ;
  assign n1491 = ~\P1_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n1492 = \P1_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1494 = ~\P1_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n1495 = \P1_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n1496 = ~n1415 & ~n1495 ;
  assign n1497 = ~n1494 & ~n1496 ;
  assign n1498 = ~n1414 & ~n1418 ;
  assign n1499 = ~n1494 & n1498 ;
  assign n1500 = ~n1352 & ~n1417 ;
  assign n1501 = n1499 & ~n1500 ;
  assign n1502 = ~n1497 & ~n1501 ;
  assign n1503 = ~n1351 & n1499 ;
  assign n1504 = ~n1208 & n1363 ;
  assign n1505 = n1360 & ~n1504 ;
  assign n1506 = n1503 & ~n1505 ;
  assign n1507 = n1502 & ~n1506 ;
  assign n1509 = ~n1493 & n1507 ;
  assign n1508 = n1493 & ~n1507 ;
  assign n1510 = n639 & ~n1508 ;
  assign n1511 = ~n1509 & n1510 ;
  assign n1512 = ~n1490 & ~n1511 ;
  assign n1513 = ~n634 & ~n1512 ;
  assign n1517 = ~\P2_reg3_reg[23]/NET0131  & ~\P2_reg3_reg[24]/NET0131  ;
  assign n1518 = n1438 & n1517 ;
  assign n1519 = \P2_reg3_reg[25]/NET0131  & ~n1518 ;
  assign n1520 = ~\P2_reg3_reg[25]/NET0131  & n1518 ;
  assign n1521 = ~n1519 & ~n1520 ;
  assign n1522 = n581 & ~n1521 ;
  assign n1516 = \P2_reg2_reg[25]/NET0131  & n597 ;
  assign n1514 = \P2_reg1_reg[25]/NET0131  & n577 ;
  assign n1515 = \P2_reg0_reg[25]/NET0131  & n579 ;
  assign n1523 = ~n1514 & ~n1515 ;
  assign n1524 = ~n1516 & n1523 ;
  assign n1525 = ~n1522 & n1524 ;
  assign n1526 = ~n1513 & ~n1525 ;
  assign n1527 = \P1_datao_reg[24]/NET0131  & ~n639 ;
  assign n1528 = ~n1494 & ~n1495 ;
  assign n1529 = ~n1417 & ~n1452 ;
  assign n1530 = n1498 & ~n1529 ;
  assign n1531 = ~n1415 & ~n1530 ;
  assign n1532 = n1449 & n1498 ;
  assign n1533 = ~n1394 & n1532 ;
  assign n1534 = n1531 & ~n1533 ;
  assign n1536 = ~n1528 & n1534 ;
  assign n1535 = n1528 & ~n1534 ;
  assign n1537 = n639 & ~n1535 ;
  assign n1538 = ~n1536 & n1537 ;
  assign n1539 = ~n1527 & ~n1538 ;
  assign n1540 = ~n634 & ~n1539 ;
  assign n1544 = \P2_reg3_reg[24]/NET0131  & ~n1440 ;
  assign n1545 = ~n1518 & ~n1544 ;
  assign n1546 = n581 & ~n1545 ;
  assign n1543 = \P2_reg1_reg[24]/NET0131  & n577 ;
  assign n1541 = \P2_reg2_reg[24]/NET0131  & n597 ;
  assign n1542 = \P2_reg0_reg[24]/NET0131  & n579 ;
  assign n1547 = ~n1541 & ~n1542 ;
  assign n1548 = ~n1543 & n1547 ;
  assign n1549 = ~n1546 & n1548 ;
  assign n1550 = ~n1540 & ~n1549 ;
  assign n1551 = ~n1526 & ~n1550 ;
  assign n1552 = \P1_datao_reg[26]/NET0131  & ~n639 ;
  assign n1553 = ~\P1_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n1554 = \P1_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n1555 = ~n1553 & ~n1554 ;
  assign n1556 = ~n1492 & ~n1495 ;
  assign n1557 = ~n1491 & ~n1556 ;
  assign n1558 = ~n1491 & ~n1494 ;
  assign n1559 = ~n1414 & n1558 ;
  assign n1560 = ~n1415 & ~n1417 ;
  assign n1561 = n1559 & ~n1560 ;
  assign n1562 = ~n1557 & ~n1561 ;
  assign n1563 = ~n1321 & n1454 ;
  assign n1564 = n1453 & ~n1563 ;
  assign n1565 = n1498 & n1558 ;
  assign n1566 = ~n1564 & n1565 ;
  assign n1567 = n1562 & ~n1566 ;
  assign n1569 = ~n1555 & n1567 ;
  assign n1568 = n1555 & ~n1567 ;
  assign n1570 = n639 & ~n1568 ;
  assign n1571 = ~n1569 & n1570 ;
  assign n1572 = ~n1552 & ~n1571 ;
  assign n1573 = ~n634 & ~n1572 ;
  assign n1577 = \P2_reg3_reg[26]/NET0131  & ~n1520 ;
  assign n1578 = ~\P2_reg3_reg[21]/NET0131  & ~\P2_reg3_reg[22]/NET0131  ;
  assign n1579 = ~\P2_reg3_reg[25]/NET0131  & ~\P2_reg3_reg[26]/NET0131  ;
  assign n1580 = n1578 & n1579 ;
  assign n1581 = n1517 & n1580 ;
  assign n1582 = n1375 & n1581 ;
  assign n1583 = ~n1577 & ~n1582 ;
  assign n1584 = n581 & ~n1583 ;
  assign n1576 = \P2_reg0_reg[26]/NET0131  & n579 ;
  assign n1574 = \P2_reg2_reg[26]/NET0131  & n597 ;
  assign n1575 = \P2_reg1_reg[26]/NET0131  & n577 ;
  assign n1585 = ~n1574 & ~n1575 ;
  assign n1586 = ~n1576 & n1585 ;
  assign n1587 = ~n1584 & n1586 ;
  assign n1588 = ~n1573 & ~n1587 ;
  assign n1589 = \P1_datao_reg[27]/NET0131  & ~n639 ;
  assign n1590 = ~\P1_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n1591 = \P1_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n1592 = ~n1590 & ~n1591 ;
  assign n1593 = ~n1492 & ~n1554 ;
  assign n1594 = ~n1553 & ~n1593 ;
  assign n1595 = ~n1491 & ~n1553 ;
  assign n1596 = n1497 & n1595 ;
  assign n1597 = ~n1594 & ~n1596 ;
  assign n1598 = ~n1553 & n1559 ;
  assign n1599 = ~n1288 & n1423 ;
  assign n1600 = n1422 & ~n1599 ;
  assign n1601 = n1598 & ~n1600 ;
  assign n1602 = n1597 & ~n1601 ;
  assign n1604 = ~n1592 & n1602 ;
  assign n1603 = n1592 & ~n1602 ;
  assign n1605 = n639 & ~n1603 ;
  assign n1606 = ~n1604 & n1605 ;
  assign n1607 = ~n1589 & ~n1606 ;
  assign n1608 = ~n634 & ~n1607 ;
  assign n1612 = ~\P2_reg3_reg[27]/NET0131  & n1582 ;
  assign n1613 = \P2_reg3_reg[27]/NET0131  & ~n1582 ;
  assign n1614 = ~n1612 & ~n1613 ;
  assign n1615 = n581 & ~n1614 ;
  assign n1611 = \P2_reg0_reg[27]/NET0131  & n579 ;
  assign n1609 = \P2_reg1_reg[27]/NET0131  & n577 ;
  assign n1610 = \P2_reg2_reg[27]/NET0131  & n597 ;
  assign n1616 = ~n1609 & ~n1610 ;
  assign n1617 = ~n1611 & n1616 ;
  assign n1618 = ~n1615 & n1617 ;
  assign n1619 = ~n1608 & ~n1618 ;
  assign n1620 = ~n1588 & ~n1619 ;
  assign n1621 = n1551 & n1620 ;
  assign n1622 = ~n1489 & n1621 ;
  assign n1623 = n1573 & n1587 ;
  assign n1624 = n1608 & n1618 ;
  assign n1625 = ~n1623 & ~n1624 ;
  assign n1626 = n1513 & n1525 ;
  assign n1627 = n1540 & n1549 ;
  assign n1628 = ~n1626 & ~n1627 ;
  assign n1629 = ~n1526 & ~n1588 ;
  assign n1630 = ~n1628 & n1629 ;
  assign n1631 = n1625 & ~n1630 ;
  assign n1632 = ~n1619 & ~n1631 ;
  assign n1633 = ~n1622 & ~n1632 ;
  assign n1634 = \P1_datao_reg[29]/NET0131  & ~n639 ;
  assign n1635 = ~\P1_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n1636 = \P1_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n1637 = ~n1635 & ~n1636 ;
  assign n1638 = ~\P1_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n1642 = ~n1590 & ~n1638 ;
  assign n1646 = n1595 & n1642 ;
  assign n1647 = n1503 & n1646 ;
  assign n1648 = ~n1365 & n1647 ;
  assign n1639 = \P1_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n1640 = ~n1591 & ~n1639 ;
  assign n1641 = ~n1638 & ~n1640 ;
  assign n1643 = ~n1502 & n1595 ;
  assign n1644 = ~n1594 & ~n1643 ;
  assign n1645 = n1642 & ~n1644 ;
  assign n1649 = ~n1641 & ~n1645 ;
  assign n1650 = ~n1648 & n1649 ;
  assign n1652 = ~n1637 & n1650 ;
  assign n1651 = n1637 & ~n1650 ;
  assign n1653 = n639 & ~n1651 ;
  assign n1654 = ~n1652 & n1653 ;
  assign n1655 = ~n1634 & ~n1654 ;
  assign n1656 = ~n634 & ~n1655 ;
  assign n1660 = ~\P2_reg3_reg[27]/NET0131  & ~\P2_reg3_reg[28]/NET0131  ;
  assign n1661 = n1582 & n1660 ;
  assign n1662 = n581 & n1661 ;
  assign n1659 = \P2_reg0_reg[29]/NET0131  & n579 ;
  assign n1657 = \P2_reg2_reg[29]/NET0131  & n597 ;
  assign n1658 = \P2_reg1_reg[29]/NET0131  & n577 ;
  assign n1663 = ~n1657 & ~n1658 ;
  assign n1664 = ~n1659 & n1663 ;
  assign n1665 = ~n1662 & n1664 ;
  assign n1666 = ~n1656 & ~n1665 ;
  assign n1667 = \P1_datao_reg[28]/NET0131  & ~n639 ;
  assign n1668 = ~n1638 & ~n1639 ;
  assign n1669 = ~n1553 & ~n1590 ;
  assign n1670 = n1558 & n1669 ;
  assign n1671 = n1533 & n1670 ;
  assign n1672 = ~n1554 & ~n1591 ;
  assign n1673 = ~n1590 & ~n1672 ;
  assign n1674 = ~n1531 & n1558 ;
  assign n1675 = ~n1557 & ~n1674 ;
  assign n1676 = n1669 & ~n1675 ;
  assign n1677 = ~n1673 & ~n1676 ;
  assign n1678 = ~n1671 & n1677 ;
  assign n1680 = ~n1668 & n1678 ;
  assign n1679 = n1668 & ~n1678 ;
  assign n1681 = n639 & ~n1679 ;
  assign n1682 = ~n1680 & n1681 ;
  assign n1683 = ~n1667 & ~n1682 ;
  assign n1684 = ~n634 & ~n1683 ;
  assign n1688 = \P2_reg3_reg[28]/NET0131  & ~n1612 ;
  assign n1689 = ~n1661 & ~n1688 ;
  assign n1690 = n581 & ~n1689 ;
  assign n1687 = \P2_reg1_reg[28]/NET0131  & n577 ;
  assign n1685 = \P2_reg0_reg[28]/NET0131  & n579 ;
  assign n1686 = \P2_reg2_reg[28]/NET0131  & n597 ;
  assign n1691 = ~n1685 & ~n1686 ;
  assign n1692 = ~n1687 & n1691 ;
  assign n1693 = ~n1690 & n1692 ;
  assign n1694 = ~n1684 & ~n1693 ;
  assign n1695 = ~n1666 & ~n1694 ;
  assign n1698 = \P2_reg1_reg[31]/NET0131  & n577 ;
  assign n1696 = \P2_reg2_reg[31]/NET0131  & n597 ;
  assign n1697 = \P2_reg0_reg[31]/NET0131  & n579 ;
  assign n1699 = ~n1696 & ~n1697 ;
  assign n1700 = ~n1698 & n1699 ;
  assign n1701 = ~n1662 & n1700 ;
  assign n1702 = ~\P1_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n1703 = ~n1635 & ~n1702 ;
  assign n1704 = n1642 & n1703 ;
  assign n1705 = n1598 & n1704 ;
  assign n1706 = n1427 & n1705 ;
  assign n1708 = ~n1425 & n1598 ;
  assign n1709 = n1597 & ~n1708 ;
  assign n1710 = n1704 & ~n1709 ;
  assign n1707 = \P1_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n1711 = ~n1636 & ~n1641 ;
  assign n1712 = n1703 & ~n1711 ;
  assign n1713 = ~n1707 & ~n1712 ;
  assign n1714 = ~n1710 & n1713 ;
  assign n1715 = ~n1706 & n1714 ;
  assign n1717 = ~\si[31]_pad  & n1715 ;
  assign n1716 = \si[31]_pad  & ~n1715 ;
  assign n1718 = n639 & ~n1716 ;
  assign n1719 = ~n1717 & n1718 ;
  assign n1720 = \P1_datao_reg[31]/NET0131  & n1719 ;
  assign n1721 = ~\P1_datao_reg[31]/NET0131  & ~n1719 ;
  assign n1722 = ~n1720 & ~n1721 ;
  assign n1723 = ~n634 & n1722 ;
  assign n1724 = n1701 & n1723 ;
  assign n1725 = \P1_datao_reg[30]/NET0131  & ~n639 ;
  assign n1726 = ~n1702 & ~n1707 ;
  assign n1727 = ~n1635 & ~n1638 ;
  assign n1728 = n1669 & n1727 ;
  assign n1729 = n1565 & n1728 ;
  assign n1730 = n1458 & n1729 ;
  assign n1733 = ~n1456 & n1565 ;
  assign n1734 = n1562 & ~n1733 ;
  assign n1735 = n1728 & ~n1734 ;
  assign n1731 = ~n1639 & ~n1673 ;
  assign n1732 = n1727 & ~n1731 ;
  assign n1736 = ~n1636 & ~n1732 ;
  assign n1737 = ~n1735 & n1736 ;
  assign n1738 = ~n1730 & n1737 ;
  assign n1740 = ~n1726 & n1738 ;
  assign n1739 = n1726 & ~n1738 ;
  assign n1741 = n639 & ~n1739 ;
  assign n1742 = ~n1740 & n1741 ;
  assign n1743 = ~n1725 & ~n1742 ;
  assign n1744 = ~n634 & ~n1743 ;
  assign n1747 = \P2_reg1_reg[30]/NET0131  & n577 ;
  assign n1745 = \P2_reg2_reg[30]/NET0131  & n597 ;
  assign n1746 = \P2_reg0_reg[30]/NET0131  & n579 ;
  assign n1748 = ~n1745 & ~n1746 ;
  assign n1749 = ~n1747 & n1748 ;
  assign n1750 = ~n1662 & n1749 ;
  assign n1751 = ~n1744 & ~n1750 ;
  assign n1752 = ~n1724 & ~n1751 ;
  assign n1753 = n1695 & n1752 ;
  assign n1754 = ~n1633 & n1753 ;
  assign n1755 = ~n1701 & ~n1723 ;
  assign n1756 = n1744 & n1750 ;
  assign n1757 = ~n1755 & ~n1756 ;
  assign n1758 = ~n1724 & ~n1757 ;
  assign n1759 = n1656 & n1665 ;
  assign n1760 = n1684 & n1693 ;
  assign n1761 = ~n1759 & ~n1760 ;
  assign n1762 = ~n1666 & n1752 ;
  assign n1763 = ~n1761 & n1762 ;
  assign n1764 = ~n1758 & ~n1763 ;
  assign n1765 = ~n1754 & n1764 ;
  assign n1766 = ~\P2_B_reg/NET0131  & n1765 ;
  assign n1767 = \P2_IR_reg[31]/NET0131  & ~n543 ;
  assign n1768 = ~n1216 & ~n1767 ;
  assign n1769 = \P2_IR_reg[21]/NET0131  & ~n1768 ;
  assign n1770 = ~\P2_IR_reg[21]/NET0131  & n1768 ;
  assign n1771 = ~n1769 & ~n1770 ;
  assign n1772 = ~\P2_IR_reg[19]/NET0131  & n605 ;
  assign n1773 = \P2_IR_reg[31]/NET0131  & ~n1772 ;
  assign n1774 = ~n1250 & ~n1773 ;
  assign n1775 = \P2_IR_reg[20]/NET0131  & ~n1774 ;
  assign n1776 = ~\P2_IR_reg[20]/NET0131  & n1774 ;
  assign n1777 = ~n1775 & ~n1776 ;
  assign n1778 = ~n1771 & ~n1777 ;
  assign n1779 = n560 & n565 ;
  assign n1780 = \P2_IR_reg[31]/NET0131  & ~n1779 ;
  assign n1781 = ~\P2_IR_reg[22]/NET0131  & ~n1780 ;
  assign n1782 = \P2_IR_reg[22]/NET0131  & n1780 ;
  assign n1783 = ~n1781 & ~n1782 ;
  assign n1784 = \P2_IR_reg[31]/NET0131  & ~n604 ;
  assign n1785 = ~n625 & ~n1784 ;
  assign n1786 = \P2_IR_reg[23]/NET0131  & ~n1785 ;
  assign n1787 = ~\P2_IR_reg[23]/NET0131  & n1785 ;
  assign n1788 = ~n1786 & ~n1787 ;
  assign n1789 = n1783 & n1788 ;
  assign n1790 = n1778 & n1789 ;
  assign n1791 = ~n1766 & n1790 ;
  assign n1792 = ~n1695 & ~n1759 ;
  assign n1793 = ~n1756 & n1792 ;
  assign n1794 = n1752 & ~n1793 ;
  assign n1795 = ~n1755 & ~n1794 ;
  assign n1796 = n1625 & n1628 ;
  assign n1797 = n1481 & n1484 ;
  assign n1820 = ~n1257 & ~n1342 ;
  assign n1821 = n1341 & n1820 ;
  assign n1822 = ~n1336 & ~n1340 ;
  assign n1823 = ~n1821 & ~n1822 ;
  assign n1798 = n1341 & n1344 ;
  assign n1800 = n774 & n968 ;
  assign n1824 = ~n935 & ~n977 ;
  assign n1825 = n911 & n1824 ;
  assign n1826 = ~n884 & ~n975 ;
  assign n1827 = ~n1825 & ~n1826 ;
  assign n1828 = n1800 & ~n1827 ;
  assign n1829 = n859 & ~n1828 ;
  assign n1830 = n1798 & ~n1829 ;
  assign n1831 = n1823 & ~n1830 ;
  assign n1832 = n1797 & ~n1831 ;
  assign n1799 = n1797 & n1798 ;
  assign n1801 = n1158 & ~n1165 ;
  assign n1802 = ~n1149 & n1801 ;
  assign n1803 = ~n1151 & ~n1802 ;
  assign n1804 = n1127 & n1803 ;
  assign n1805 = ~n1101 & ~n1150 ;
  assign n1806 = ~n1126 & ~n1805 ;
  assign n1807 = ~n1804 & ~n1806 ;
  assign n1808 = n1079 & ~n1807 ;
  assign n1809 = ~n1051 & ~n1102 ;
  assign n1810 = ~n1078 & ~n1809 ;
  assign n1811 = ~n1808 & ~n1810 ;
  assign n1812 = n1028 & ~n1811 ;
  assign n1813 = ~n1052 & ~n1175 ;
  assign n1814 = ~n1027 & ~n1813 ;
  assign n1815 = ~n1812 & ~n1814 ;
  assign n1816 = n911 & n960 ;
  assign n1817 = ~n1815 & n1816 ;
  assign n1818 = n1800 & n1817 ;
  assign n1819 = n1799 & n1818 ;
  assign n1833 = ~n1412 & ~n1482 ;
  assign n1834 = n1481 & n1833 ;
  assign n1835 = ~n1476 & ~n1480 ;
  assign n1836 = ~n1834 & ~n1835 ;
  assign n1837 = ~n1819 & n1836 ;
  assign n1838 = ~n1832 & n1837 ;
  assign n1839 = n1796 & ~n1838 ;
  assign n1840 = ~n1551 & ~n1626 ;
  assign n1841 = ~n1623 & n1840 ;
  assign n1842 = n1620 & ~n1841 ;
  assign n1843 = ~n1624 & ~n1842 ;
  assign n1844 = ~n1839 & ~n1843 ;
  assign n1845 = n1757 & n1761 ;
  assign n1846 = ~n1844 & n1845 ;
  assign n1847 = ~n1795 & ~n1846 ;
  assign n1848 = ~\P2_B_reg/NET0131  & n1847 ;
  assign n1849 = ~n1783 & n1788 ;
  assign n1850 = ~n1771 & n1777 ;
  assign n1851 = n1849 & n1850 ;
  assign n1852 = ~n1848 & n1851 ;
  assign n1853 = ~n1783 & ~n1788 ;
  assign n1854 = n1850 & n1853 ;
  assign n1855 = ~n1847 & n1854 ;
  assign n1856 = ~n1818 & n1829 ;
  assign n1857 = n1799 & ~n1856 ;
  assign n1858 = n1797 & ~n1823 ;
  assign n1859 = n1836 & ~n1858 ;
  assign n1860 = ~n1857 & n1859 ;
  assign n1861 = ~n1701 & ~n1750 ;
  assign n1862 = n1744 & ~n1861 ;
  assign n1863 = ~n1755 & ~n1862 ;
  assign n1864 = n1761 & n1863 ;
  assign n1865 = n1796 & n1864 ;
  assign n1866 = ~n1860 & n1865 ;
  assign n1867 = n1843 & n1864 ;
  assign n1868 = n1792 & n1863 ;
  assign n1869 = ~n1701 & ~n1751 ;
  assign n1870 = n1723 & ~n1869 ;
  assign n1871 = ~n1868 & ~n1870 ;
  assign n1872 = ~n1867 & n1871 ;
  assign n1873 = ~n1866 & n1872 ;
  assign n1874 = ~\P2_B_reg/NET0131  & ~n1873 ;
  assign n1875 = n1771 & n1789 ;
  assign n1876 = ~n1777 & n1875 ;
  assign n1877 = ~n1874 & n1876 ;
  assign n1878 = n1777 & n1875 ;
  assign n1879 = ~n1873 & n1878 ;
  assign n1880 = n1849 & ~n1850 ;
  assign n1881 = ~n1878 & ~n1880 ;
  assign n1882 = \P2_B_reg/NET0131  & ~n1881 ;
  assign n1883 = ~n1573 & n1587 ;
  assign n1884 = n1573 & ~n1587 ;
  assign n1885 = ~n1883 & ~n1884 ;
  assign n1886 = ~n1684 & n1693 ;
  assign n1887 = n1684 & ~n1693 ;
  assign n1888 = ~n1886 & ~n1887 ;
  assign n1977 = ~n1885 & ~n1888 ;
  assign n1889 = n1608 & ~n1618 ;
  assign n1890 = ~n1608 & n1618 ;
  assign n1891 = ~n1889 & ~n1890 ;
  assign n1892 = ~n1666 & ~n1759 ;
  assign n1978 = ~n1891 & n1892 ;
  assign n1979 = n1977 & n1978 ;
  assign n1939 = ~n1540 & n1549 ;
  assign n1940 = n1540 & ~n1549 ;
  assign n1941 = ~n1939 & ~n1940 ;
  assign n1936 = ~n1513 & n1525 ;
  assign n1937 = n1513 & ~n1525 ;
  assign n1938 = ~n1936 & ~n1937 ;
  assign n1948 = ~n1300 & ~n1340 ;
  assign n1942 = ~n1465 & n1474 ;
  assign n1943 = n1465 & ~n1474 ;
  assign n1944 = ~n1942 & ~n1943 ;
  assign n1945 = n1434 & ~n1445 ;
  assign n1946 = ~n1434 & n1445 ;
  assign n1947 = ~n1945 & ~n1946 ;
  assign n1967 = ~n1944 & ~n1947 ;
  assign n1968 = n1948 & n1967 ;
  assign n1974 = ~n1938 & n1968 ;
  assign n1975 = ~n1941 & n1974 ;
  assign n1933 = n1371 & ~n1382 ;
  assign n1934 = ~n1371 & n1382 ;
  assign n1935 = ~n1933 & ~n1934 ;
  assign n1971 = ~n1724 & ~n1755 ;
  assign n1972 = ~n1935 & n1971 ;
  assign n1965 = ~n1751 & ~n1756 ;
  assign n1893 = ~n1401 & n1410 ;
  assign n1894 = n1401 & ~n1410 ;
  assign n1895 = ~n1893 & ~n1894 ;
  assign n1896 = n1309 & n1334 ;
  assign n1897 = ~n1309 & ~n1334 ;
  assign n1898 = ~n1896 & ~n1897 ;
  assign n1966 = ~n1895 & ~n1898 ;
  assign n1969 = n1965 & n1966 ;
  assign n1932 = ~n1256 & ~n1343 ;
  assign n1928 = n601 & n718 ;
  assign n1929 = ~n601 & ~n718 ;
  assign n1930 = ~n1928 & ~n1929 ;
  assign n1931 = ~n773 & ~n856 ;
  assign n1962 = ~n1930 & n1931 ;
  assign n1963 = n1932 & n1962 ;
  assign n1913 = ~n812 & ~n813 ;
  assign n1910 = n822 & n850 ;
  assign n1911 = ~n822 & ~n850 ;
  assign n1912 = ~n1910 & ~n1911 ;
  assign n1903 = ~n1027 & ~n1175 ;
  assign n1904 = ~n1149 & ~n1151 ;
  assign n1949 = n1903 & n1904 ;
  assign n1908 = ~n1166 & ~n1801 ;
  assign n1909 = ~n1051 & ~n1078 ;
  assign n1950 = n1908 & n1909 ;
  assign n1954 = n1949 & n1950 ;
  assign n1914 = n944 & n958 ;
  assign n1915 = ~n944 & ~n958 ;
  assign n1916 = ~n1914 & ~n1915 ;
  assign n1927 = ~n935 & ~n961 ;
  assign n1955 = ~n1916 & n1927 ;
  assign n1956 = n1954 & n1955 ;
  assign n1959 = ~n1912 & n1956 ;
  assign n1960 = n1913 & n1959 ;
  assign n1899 = ~n1222 & ~n1342 ;
  assign n1905 = ~n893 & ~n909 ;
  assign n1906 = n893 & n909 ;
  assign n1907 = ~n1905 & ~n1906 ;
  assign n1900 = n868 & n882 ;
  assign n1901 = ~n868 & ~n882 ;
  assign n1902 = ~n1900 & ~n1901 ;
  assign n1917 = ~n1125 & ~n1150 ;
  assign n1918 = n986 & n1003 ;
  assign n1919 = ~n986 & ~n1003 ;
  assign n1920 = ~n1918 & ~n1919 ;
  assign n1951 = n1917 & ~n1920 ;
  assign n1921 = n1062 & n1076 ;
  assign n1922 = ~n1062 & ~n1076 ;
  assign n1923 = ~n1921 & ~n1922 ;
  assign n1924 = n1086 & n1100 ;
  assign n1925 = ~n1086 & ~n1100 ;
  assign n1926 = ~n1924 & ~n1925 ;
  assign n1952 = ~n1923 & ~n1926 ;
  assign n1953 = n1951 & n1952 ;
  assign n1957 = ~n1902 & n1953 ;
  assign n1958 = ~n1907 & n1957 ;
  assign n1961 = n1899 & n1958 ;
  assign n1964 = n1960 & n1961 ;
  assign n1970 = n1963 & n1964 ;
  assign n1973 = n1969 & n1970 ;
  assign n1976 = n1972 & n1973 ;
  assign n1980 = n1975 & n1976 ;
  assign n1981 = n1979 & n1980 ;
  assign n1983 = n1777 & n1981 ;
  assign n1982 = ~n1777 & ~n1981 ;
  assign n1984 = n1771 & ~n1783 ;
  assign n1985 = ~n1982 & n1984 ;
  assign n1986 = ~n1983 & n1985 ;
  assign n2004 = ~n1882 & ~n1986 ;
  assign n2005 = ~n1879 & n2004 ;
  assign n2006 = ~n1877 & n2005 ;
  assign n2007 = ~n1855 & n2006 ;
  assign n1987 = n1778 & ~n1783 ;
  assign n1988 = n1847 & n1987 ;
  assign n1992 = ~n1777 & ~n1873 ;
  assign n1989 = n1783 & ~n1788 ;
  assign n1990 = n1771 & n1989 ;
  assign n1991 = n1777 & n1873 ;
  assign n1993 = n1990 & ~n1991 ;
  assign n1994 = ~n1992 & n1993 ;
  assign n2008 = ~n1988 & ~n1994 ;
  assign n2009 = n2007 & n2008 ;
  assign n2010 = ~n1852 & n2009 ;
  assign n2011 = ~n1791 & n2010 ;
  assign n1995 = ~\P2_B_reg/NET0131  & ~n1765 ;
  assign n1996 = n1789 & n1850 ;
  assign n1997 = ~n1995 & n1996 ;
  assign n1998 = ~n1771 & n1989 ;
  assign n1999 = n1777 & n1998 ;
  assign n2000 = n1765 & ~n1999 ;
  assign n2001 = ~n1777 & n1998 ;
  assign n2002 = ~n1765 & ~n2001 ;
  assign n2003 = ~n2000 & ~n2002 ;
  assign n2012 = ~n1997 & ~n2003 ;
  assign n2013 = n2011 & n2012 ;
  assign n2014 = \P1_state_reg[0]/NET0131  & n1788 ;
  assign n2015 = ~n2013 & n2014 ;
  assign n2016 = \P2_B_reg/NET0131  & ~n2014 ;
  assign n2017 = ~n2015 & ~n2016 ;
  assign n2028 = \P2_IR_reg[31]/NET0131  & ~n567 ;
  assign n2029 = ~n1780 & ~n2028 ;
  assign n2030 = \P2_IR_reg[26]/NET0131  & ~n2029 ;
  assign n2031 = ~\P2_IR_reg[26]/NET0131  & n2029 ;
  assign n2032 = ~n2030 & ~n2031 ;
  assign n2020 = \P2_IR_reg[31]/NET0131  & ~n547 ;
  assign n2021 = ~n536 & ~n2020 ;
  assign n2022 = \P2_IR_reg[25]/NET0131  & ~n2021 ;
  assign n2023 = ~\P2_IR_reg[25]/NET0131  & n2021 ;
  assign n2024 = ~n2022 & ~n2023 ;
  assign n2025 = ~\P2_IR_reg[24]/NET0131  & ~n609 ;
  assign n2026 = \P2_IR_reg[24]/NET0131  & n609 ;
  assign n2027 = ~n2025 & ~n2026 ;
  assign n2033 = n2024 & n2027 ;
  assign n2034 = n2032 & n2033 ;
  assign n2035 = ~n1788 & n2034 ;
  assign n2036 = ~n1614 & n2035 ;
  assign n2037 = ~n1788 & ~n2034 ;
  assign n2038 = ~\P2_B_reg/NET0131  & ~n2024 ;
  assign n2039 = n2032 & ~n2038 ;
  assign n2040 = n2027 & ~n2039 ;
  assign n2041 = \P2_B_reg/NET0131  & ~n2027 ;
  assign n2042 = ~n2024 & n2041 ;
  assign n2043 = ~\P2_d_reg[0]/NET0131  & ~n2042 ;
  assign n2044 = n2032 & ~n2043 ;
  assign n2045 = ~n2040 & ~n2044 ;
  assign n2046 = ~\P2_B_reg/NET0131  & n2027 ;
  assign n2047 = ~n2041 & ~n2046 ;
  assign n2048 = ~n2024 & ~n2047 ;
  assign n2049 = ~\P2_d_reg[1]/NET0131  & n2032 ;
  assign n2050 = ~n2048 & n2049 ;
  assign n2051 = ~n2024 & ~n2032 ;
  assign n2052 = ~n2050 & ~n2051 ;
  assign n2053 = ~n2045 & n2052 ;
  assign n2054 = ~n1614 & ~n2053 ;
  assign n2055 = ~n719 & ~n1343 ;
  assign n2056 = ~n1339 & ~n1342 ;
  assign n2057 = n2055 & n2056 ;
  assign n2058 = ~n1004 & ~n1053 ;
  assign n2059 = ~n1150 & ~n1803 ;
  assign n2060 = n1127 & ~n2059 ;
  assign n2061 = n1103 & ~n2060 ;
  assign n2062 = ~n1004 & n1079 ;
  assign n2063 = ~n2061 & n2062 ;
  assign n2064 = ~n2058 & ~n2063 ;
  assign n2065 = ~n959 & ~n1027 ;
  assign n2066 = ~n910 & ~n935 ;
  assign n2067 = n2065 & n2066 ;
  assign n2068 = ~n2064 & n2067 ;
  assign n2069 = ~n976 & ~n1175 ;
  assign n2070 = ~n959 & ~n2069 ;
  assign n2071 = n2066 & n2070 ;
  assign n2072 = ~n910 & ~n963 ;
  assign n2073 = ~n2071 & ~n2072 ;
  assign n2074 = ~n2068 & n2073 ;
  assign n2075 = ~n773 & ~n812 ;
  assign n2076 = ~n884 & ~n967 ;
  assign n2077 = n2075 & n2076 ;
  assign n2078 = ~n2074 & n2077 ;
  assign n2079 = n2057 & n2078 ;
  assign n2080 = n883 & ~n967 ;
  assign n2081 = ~n851 & ~n2080 ;
  assign n2082 = n2075 & ~n2081 ;
  assign n2083 = ~n773 & ~n969 ;
  assign n2084 = ~n2082 & ~n2083 ;
  assign n2085 = n2057 & ~n2084 ;
  assign n2086 = ~n855 & ~n1256 ;
  assign n2087 = ~n1343 & ~n2086 ;
  assign n2088 = n2056 & n2087 ;
  assign n2089 = ~n1339 & ~n1345 ;
  assign n2090 = ~n2088 & ~n2089 ;
  assign n2091 = ~n2085 & n2090 ;
  assign n2092 = ~n2079 & n2091 ;
  assign n2093 = ~n1340 & ~n1483 ;
  assign n2094 = ~n1479 & ~n1482 ;
  assign n2095 = n2093 & n2094 ;
  assign n2096 = ~n1623 & ~n1626 ;
  assign n2097 = ~n1480 & ~n1627 ;
  assign n2098 = n2096 & n2097 ;
  assign n2099 = n2095 & n2098 ;
  assign n2100 = ~n2092 & n2099 ;
  assign n2104 = n1300 & ~n1483 ;
  assign n2105 = ~n1411 & ~n2104 ;
  assign n2106 = n2094 & ~n2105 ;
  assign n2107 = ~n1479 & ~n1485 ;
  assign n2108 = ~n2106 & ~n2107 ;
  assign n2109 = n2098 & ~n2108 ;
  assign n2101 = n1446 & ~n1627 ;
  assign n2102 = ~n1550 & ~n2101 ;
  assign n2103 = n2096 & ~n2102 ;
  assign n2110 = ~n1623 & ~n1629 ;
  assign n2111 = ~n2103 & ~n2110 ;
  assign n2112 = ~n2109 & n2111 ;
  assign n2113 = ~n2100 & n2112 ;
  assign n2114 = n1891 & ~n2113 ;
  assign n2115 = ~n1891 & n2113 ;
  assign n2116 = ~n2114 & ~n2115 ;
  assign n2117 = n2053 & ~n2116 ;
  assign n2118 = ~n2054 & ~n2117 ;
  assign n2119 = ~n1777 & n1849 ;
  assign n2120 = ~n1998 & ~n2119 ;
  assign n2121 = ~n2118 & ~n2120 ;
  assign n2124 = n2045 & ~n2052 ;
  assign n2125 = ~n1614 & ~n2124 ;
  assign n2231 = ~n1158 & ~n1701 ;
  assign n2232 = ~n1134 & n2231 ;
  assign n2233 = ~n1110 & n2232 ;
  assign n2234 = ~n986 & ~n1037 ;
  assign n2235 = ~n1062 & ~n1086 ;
  assign n2236 = n2234 & n2235 ;
  assign n2237 = n2233 & n2236 ;
  assign n2238 = ~n944 & ~n1013 ;
  assign n2239 = n2237 & n2238 ;
  assign n2240 = ~n822 & ~n868 ;
  assign n2241 = ~n893 & ~n921 ;
  assign n2242 = n2240 & n2241 ;
  assign n2243 = n2239 & n2242 ;
  assign n2244 = ~n783 & n2243 ;
  assign n2245 = ~n601 & ~n772 ;
  assign n2246 = ~n1231 & n2245 ;
  assign n2247 = n2244 & n2246 ;
  assign n2248 = ~n1269 & ~n1410 ;
  assign n2249 = ~n1309 & ~n1382 ;
  assign n2250 = n2248 & n2249 ;
  assign n2251 = ~n1193 & ~n1474 ;
  assign n2252 = ~n1445 & n2251 ;
  assign n2253 = n2250 & n2252 ;
  assign n2254 = ~n1549 & n2253 ;
  assign n2255 = n2247 & n2254 ;
  assign n2256 = ~n1525 & ~n1618 ;
  assign n2257 = ~n1587 & n2256 ;
  assign n2258 = n2255 & n2257 ;
  assign n2260 = n1693 & ~n2258 ;
  assign n2259 = ~n1693 & n2258 ;
  assign n2261 = n615 & ~n633 ;
  assign n2262 = ~n615 & n633 ;
  assign n2263 = ~n2261 & ~n2262 ;
  assign n2264 = ~n2259 & n2263 ;
  assign n2265 = ~n2260 & n2264 ;
  assign n2266 = ~n1587 & ~n2263 ;
  assign n2267 = ~n2265 & ~n2266 ;
  assign n2268 = n2124 & ~n2267 ;
  assign n2269 = ~n2125 & ~n2268 ;
  assign n2270 = n1790 & ~n2269 ;
  assign n2228 = ~n1850 & ~n2053 ;
  assign n2229 = n1853 & ~n2228 ;
  assign n2230 = n1608 & n2229 ;
  assign n2271 = ~n1778 & n1789 ;
  assign n2272 = ~n1850 & n1853 ;
  assign n2273 = ~n2053 & n2272 ;
  assign n2274 = ~n2271 & ~n2273 ;
  assign n2275 = ~n1614 & ~n2274 ;
  assign n2276 = ~n2230 & ~n2275 ;
  assign n2277 = ~n2270 & n2276 ;
  assign n2278 = ~n2121 & n2277 ;
  assign n2122 = n1777 & n1849 ;
  assign n2123 = n1771 & n2122 ;
  assign n2126 = n1193 & n1221 ;
  assign n2127 = ~n1896 & ~n2126 ;
  assign n2128 = n1231 & n1255 ;
  assign n2129 = ~n1928 & ~n2128 ;
  assign n2130 = n2127 & n2129 ;
  assign n2132 = ~n1110 & ~n1124 ;
  assign n2133 = ~n1134 & ~n1148 ;
  assign n2134 = n1134 & n1148 ;
  assign n2135 = ~n1158 & ~n1165 ;
  assign n2136 = ~n2134 & n2135 ;
  assign n2137 = ~n2133 & ~n2136 ;
  assign n2138 = ~n2132 & n2137 ;
  assign n2139 = n1110 & n1124 ;
  assign n2140 = ~n1924 & ~n2139 ;
  assign n2141 = ~n1921 & n2140 ;
  assign n2142 = ~n2138 & n2141 ;
  assign n2143 = ~n1922 & ~n1925 ;
  assign n2144 = ~n1921 & ~n2143 ;
  assign n2145 = ~n2142 & ~n2144 ;
  assign n2131 = n1037 & n1050 ;
  assign n2146 = ~n1918 & ~n2131 ;
  assign n2147 = ~n2145 & n2146 ;
  assign n2148 = ~n1037 & ~n1050 ;
  assign n2149 = ~n1918 & n2148 ;
  assign n2150 = ~n1919 & ~n2149 ;
  assign n2151 = ~n2147 & n2150 ;
  assign n2152 = n921 & n934 ;
  assign n2153 = ~n1906 & ~n2152 ;
  assign n2154 = n1013 & n1026 ;
  assign n2155 = ~n1914 & ~n2154 ;
  assign n2156 = n2153 & n2155 ;
  assign n2157 = ~n2151 & n2156 ;
  assign n2158 = ~n1013 & ~n1026 ;
  assign n2159 = ~n1915 & ~n2158 ;
  assign n2160 = ~n1914 & ~n2159 ;
  assign n2161 = n2153 & n2160 ;
  assign n2162 = ~n921 & ~n934 ;
  assign n2163 = ~n1906 & n2162 ;
  assign n2164 = ~n1905 & ~n2163 ;
  assign n2165 = ~n2161 & n2164 ;
  assign n2166 = ~n2157 & n2165 ;
  assign n2167 = n760 & n772 ;
  assign n2168 = n783 & n811 ;
  assign n2169 = ~n2167 & ~n2168 ;
  assign n2170 = ~n1900 & ~n1910 ;
  assign n2171 = n2169 & n2170 ;
  assign n2172 = ~n2166 & n2171 ;
  assign n2173 = n2130 & n2172 ;
  assign n2174 = n1901 & ~n1910 ;
  assign n2175 = ~n1911 & ~n2174 ;
  assign n2176 = n2169 & ~n2175 ;
  assign n2177 = ~n760 & ~n772 ;
  assign n2178 = ~n783 & ~n811 ;
  assign n2179 = ~n2167 & n2178 ;
  assign n2180 = ~n2177 & ~n2179 ;
  assign n2181 = ~n2176 & n2180 ;
  assign n2182 = n2130 & ~n2181 ;
  assign n2183 = ~n1231 & ~n1255 ;
  assign n2184 = n1929 & ~n2128 ;
  assign n2185 = ~n2183 & ~n2184 ;
  assign n2186 = n2127 & ~n2185 ;
  assign n2187 = ~n1193 & ~n1221 ;
  assign n2188 = ~n1896 & n2187 ;
  assign n2189 = ~n1897 & ~n2188 ;
  assign n2190 = ~n2186 & n2189 ;
  assign n2191 = ~n2182 & n2190 ;
  assign n2192 = ~n2173 & n2191 ;
  assign n2193 = ~n1939 & ~n1946 ;
  assign n2194 = ~n1936 & n2193 ;
  assign n2195 = ~n1934 & ~n1942 ;
  assign n2196 = n1269 & n1299 ;
  assign n2197 = ~n1893 & ~n2196 ;
  assign n2198 = n2195 & n2197 ;
  assign n2199 = ~n1883 & n2198 ;
  assign n2200 = n2194 & n2199 ;
  assign n2201 = ~n2192 & n2200 ;
  assign n2206 = ~n1269 & ~n1299 ;
  assign n2207 = ~n1893 & n2206 ;
  assign n2208 = ~n1894 & ~n2207 ;
  assign n2209 = n2195 & ~n2208 ;
  assign n2210 = n1933 & ~n1942 ;
  assign n2211 = ~n1943 & ~n2210 ;
  assign n2212 = ~n2209 & n2211 ;
  assign n2213 = n2194 & ~n2212 ;
  assign n2202 = ~n1884 & ~n1937 ;
  assign n2203 = ~n1939 & n1945 ;
  assign n2204 = ~n1940 & ~n2203 ;
  assign n2205 = ~n1936 & ~n2204 ;
  assign n2214 = n2202 & ~n2205 ;
  assign n2215 = ~n2213 & n2214 ;
  assign n2216 = ~n1883 & ~n2215 ;
  assign n2217 = ~n2201 & ~n2216 ;
  assign n2218 = n1891 & n2217 ;
  assign n2219 = ~n1891 & ~n2217 ;
  assign n2220 = ~n2218 & ~n2219 ;
  assign n2221 = n2124 & ~n2220 ;
  assign n2222 = ~n2125 & ~n2221 ;
  assign n2223 = n2123 & ~n2222 ;
  assign n2224 = ~n1851 & ~n1990 ;
  assign n2225 = n2053 & ~n2220 ;
  assign n2226 = ~n2054 & ~n2225 ;
  assign n2227 = ~n2224 & ~n2226 ;
  assign n2279 = ~n2223 & ~n2227 ;
  assign n2280 = n2278 & n2279 ;
  assign n2281 = n2037 & ~n2280 ;
  assign n2282 = ~n2036 & ~n2281 ;
  assign n2283 = \P1_state_reg[0]/NET0131  & ~n2282 ;
  assign n2018 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[27]/NET0131  ;
  assign n2019 = ~n1614 & n2014 ;
  assign n2284 = ~n2018 & ~n2019 ;
  assign n2285 = ~n2283 & n2284 ;
  assign n2286 = \P1_state_reg[0]/NET0131  & ~n1788 ;
  assign n2287 = \P2_reg2_reg[28]/NET0131  & ~n2286 ;
  assign n2288 = \P2_reg2_reg[28]/NET0131  & n2035 ;
  assign n2289 = n1788 & n1987 ;
  assign n2290 = ~n1998 & ~n2289 ;
  assign n2291 = n2045 & n2052 ;
  assign n2292 = \P2_reg2_reg[28]/NET0131  & ~n2291 ;
  assign n2293 = ~n1817 & n1827 ;
  assign n2294 = n1798 & n1800 ;
  assign n2295 = ~n2293 & n2294 ;
  assign n2296 = ~n859 & n1798 ;
  assign n2297 = n1823 & ~n2296 ;
  assign n2298 = ~n2295 & n2297 ;
  assign n2299 = n1796 & n1797 ;
  assign n2300 = ~n2298 & n2299 ;
  assign n2301 = n1796 & ~n1836 ;
  assign n2302 = ~n1843 & ~n2301 ;
  assign n2303 = ~n2300 & n2302 ;
  assign n2304 = n1888 & ~n2303 ;
  assign n2305 = ~n1888 & n2303 ;
  assign n2306 = ~n2304 & ~n2305 ;
  assign n2307 = n2291 & ~n2306 ;
  assign n2308 = ~n2292 & ~n2307 ;
  assign n2309 = ~n2290 & ~n2308 ;
  assign n2310 = ~n2045 & ~n2052 ;
  assign n2311 = \P2_reg2_reg[28]/NET0131  & ~n2310 ;
  assign n2396 = ~n1618 & ~n2263 ;
  assign n2397 = n1665 & ~n2259 ;
  assign n2398 = ~n1665 & ~n1693 ;
  assign n2399 = n2258 & n2398 ;
  assign n2400 = n2263 & ~n2399 ;
  assign n2401 = ~n2397 & n2400 ;
  assign n2402 = ~n2396 & ~n2401 ;
  assign n2403 = n2310 & ~n2402 ;
  assign n2404 = ~n2311 & ~n2403 ;
  assign n2405 = n1790 & ~n2404 ;
  assign n2394 = n2272 & n2291 ;
  assign n2395 = n1684 & n2394 ;
  assign n2406 = n2272 & ~n2291 ;
  assign n2407 = ~n2271 & ~n2406 ;
  assign n2408 = \P2_reg2_reg[28]/NET0131  & ~n2407 ;
  assign n2409 = ~n1689 & n1854 ;
  assign n2410 = ~n2408 & ~n2409 ;
  assign n2411 = ~n2395 & n2410 ;
  assign n2412 = ~n2405 & n2411 ;
  assign n2413 = ~n2309 & n2412 ;
  assign n2312 = ~n2306 & n2310 ;
  assign n2313 = ~n2311 & ~n2312 ;
  assign n2314 = n1771 & n2119 ;
  assign n2315 = ~n2313 & n2314 ;
  assign n2316 = ~n1918 & ~n2154 ;
  assign n2317 = ~n2137 & n2140 ;
  assign n2318 = ~n1925 & ~n2132 ;
  assign n2319 = ~n1924 & ~n2318 ;
  assign n2320 = ~n2317 & ~n2319 ;
  assign n2321 = ~n1921 & ~n2131 ;
  assign n2322 = ~n2320 & n2321 ;
  assign n2323 = n1922 & ~n2131 ;
  assign n2324 = ~n2148 & ~n2323 ;
  assign n2325 = ~n2322 & n2324 ;
  assign n2326 = n2316 & ~n2325 ;
  assign n2327 = n1919 & ~n2154 ;
  assign n2328 = ~n2158 & ~n2327 ;
  assign n2329 = ~n2326 & n2328 ;
  assign n2330 = ~n1914 & ~n2152 ;
  assign n2331 = ~n1900 & ~n1906 ;
  assign n2332 = n2330 & n2331 ;
  assign n2333 = ~n2329 & n2332 ;
  assign n2334 = ~n1915 & ~n2162 ;
  assign n2335 = ~n2152 & ~n2334 ;
  assign n2336 = n2331 & n2335 ;
  assign n2337 = ~n1900 & n1905 ;
  assign n2338 = ~n1901 & ~n2337 ;
  assign n2339 = ~n2336 & n2338 ;
  assign n2340 = ~n2333 & n2339 ;
  assign n2341 = ~n1928 & ~n2167 ;
  assign n2342 = ~n1910 & ~n2168 ;
  assign n2343 = n2341 & n2342 ;
  assign n2344 = ~n1896 & ~n2196 ;
  assign n2345 = ~n2126 & ~n2128 ;
  assign n2346 = n2344 & n2345 ;
  assign n2347 = n2343 & n2346 ;
  assign n2348 = ~n2340 & n2347 ;
  assign n2349 = ~n1911 & ~n2178 ;
  assign n2350 = ~n2168 & ~n2349 ;
  assign n2351 = n2341 & n2350 ;
  assign n2352 = ~n1928 & n2177 ;
  assign n2353 = ~n1929 & ~n2352 ;
  assign n2354 = ~n2351 & n2353 ;
  assign n2355 = n2346 & ~n2354 ;
  assign n2356 = ~n2126 & n2183 ;
  assign n2357 = ~n2187 & ~n2356 ;
  assign n2358 = n2344 & ~n2357 ;
  assign n2359 = ~n1897 & ~n2206 ;
  assign n2360 = ~n2196 & ~n2359 ;
  assign n2361 = ~n2358 & ~n2360 ;
  assign n2362 = ~n2355 & n2361 ;
  assign n2363 = ~n2348 & n2362 ;
  assign n2364 = ~n1936 & ~n1939 ;
  assign n2365 = ~n1883 & ~n1890 ;
  assign n2366 = n2364 & n2365 ;
  assign n2367 = ~n1893 & ~n1934 ;
  assign n2368 = ~n1942 & ~n1946 ;
  assign n2369 = n2367 & n2368 ;
  assign n2370 = n2366 & n2369 ;
  assign n2371 = ~n2363 & n2370 ;
  assign n2373 = n1894 & ~n1934 ;
  assign n2374 = ~n1933 & ~n2373 ;
  assign n2375 = n2368 & ~n2374 ;
  assign n2376 = n1943 & ~n1946 ;
  assign n2377 = ~n1945 & ~n2376 ;
  assign n2378 = ~n2375 & n2377 ;
  assign n2379 = n2366 & ~n2378 ;
  assign n2380 = ~n1936 & n1940 ;
  assign n2381 = ~n1937 & ~n2380 ;
  assign n2382 = n2365 & ~n2381 ;
  assign n2372 = n1884 & ~n1890 ;
  assign n2383 = ~n1889 & ~n2372 ;
  assign n2384 = ~n2382 & n2383 ;
  assign n2385 = ~n2379 & n2384 ;
  assign n2386 = ~n2371 & n2385 ;
  assign n2387 = n1888 & n2386 ;
  assign n2388 = ~n1888 & ~n2386 ;
  assign n2389 = ~n2387 & ~n2388 ;
  assign n2390 = n2291 & ~n2389 ;
  assign n2391 = ~n2292 & ~n2390 ;
  assign n2392 = ~n1990 & ~n2122 ;
  assign n2393 = ~n2391 & ~n2392 ;
  assign n2414 = ~n2315 & ~n2393 ;
  assign n2415 = n2413 & n2414 ;
  assign n2416 = n2037 & ~n2415 ;
  assign n2417 = ~n2288 & ~n2416 ;
  assign n2418 = \P1_state_reg[0]/NET0131  & ~n2417 ;
  assign n2419 = ~n2287 & ~n2418 ;
  assign n2422 = ~n1689 & n2035 ;
  assign n2423 = ~n1689 & ~n2053 ;
  assign n2424 = n2053 & ~n2306 ;
  assign n2425 = ~n2423 & ~n2424 ;
  assign n2426 = ~n2120 & ~n2425 ;
  assign n2427 = ~n1689 & ~n2124 ;
  assign n2435 = n2124 & ~n2402 ;
  assign n2436 = ~n2427 & ~n2435 ;
  assign n2437 = n1790 & ~n2436 ;
  assign n2434 = ~n1689 & ~n2274 ;
  assign n2438 = n1684 & n2229 ;
  assign n2439 = ~n2434 & ~n2438 ;
  assign n2440 = ~n2437 & n2439 ;
  assign n2441 = ~n2426 & n2440 ;
  assign n2428 = n2124 & ~n2389 ;
  assign n2429 = ~n2427 & ~n2428 ;
  assign n2430 = n2123 & ~n2429 ;
  assign n2431 = n2053 & ~n2389 ;
  assign n2432 = ~n2423 & ~n2431 ;
  assign n2433 = ~n2224 & ~n2432 ;
  assign n2442 = ~n2430 & ~n2433 ;
  assign n2443 = n2441 & n2442 ;
  assign n2444 = n2037 & ~n2443 ;
  assign n2445 = ~n2422 & ~n2444 ;
  assign n2446 = \P1_state_reg[0]/NET0131  & ~n2445 ;
  assign n2420 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[28]/NET0131  ;
  assign n2421 = ~n1689 & n2014 ;
  assign n2447 = ~n2420 & ~n2421 ;
  assign n2448 = ~n2446 & n2447 ;
  assign n2449 = \P2_reg2_reg[27]/NET0131  & ~n2286 ;
  assign n2450 = \P2_reg2_reg[27]/NET0131  & n2035 ;
  assign n2451 = \P2_reg2_reg[27]/NET0131  & ~n2291 ;
  assign n2452 = ~n2116 & n2291 ;
  assign n2453 = ~n2451 & ~n2452 ;
  assign n2454 = ~n2290 & ~n2453 ;
  assign n2458 = \P2_reg2_reg[27]/NET0131  & ~n2310 ;
  assign n2463 = ~n2267 & n2310 ;
  assign n2464 = ~n2458 & ~n2463 ;
  assign n2465 = n1790 & ~n2464 ;
  assign n2462 = n1608 & n2394 ;
  assign n2466 = \P2_reg2_reg[27]/NET0131  & ~n2407 ;
  assign n2467 = ~n1614 & n1854 ;
  assign n2468 = ~n2466 & ~n2467 ;
  assign n2469 = ~n2462 & n2468 ;
  assign n2470 = ~n2465 & n2469 ;
  assign n2471 = ~n2454 & n2470 ;
  assign n2455 = ~n2220 & n2291 ;
  assign n2456 = ~n2451 & ~n2455 ;
  assign n2457 = ~n2392 & ~n2456 ;
  assign n2459 = ~n2116 & n2310 ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = n2314 & ~n2460 ;
  assign n2472 = ~n2457 & ~n2461 ;
  assign n2473 = n2471 & n2472 ;
  assign n2474 = n2037 & ~n2473 ;
  assign n2475 = ~n2450 & ~n2474 ;
  assign n2476 = \P1_state_reg[0]/NET0131  & ~n2475 ;
  assign n2477 = ~n2449 & ~n2476 ;
  assign n2480 = ~n1545 & n2035 ;
  assign n2481 = ~n1545 & ~n2053 ;
  assign n2510 = ~n1838 & n1941 ;
  assign n2511 = n1838 & ~n1941 ;
  assign n2512 = ~n2510 & ~n2511 ;
  assign n2513 = n2053 & ~n2512 ;
  assign n2514 = ~n2481 & ~n2513 ;
  assign n2515 = ~n2120 & ~n2514 ;
  assign n2497 = ~n1545 & ~n2124 ;
  assign n2484 = ~n2339 & n2343 ;
  assign n2485 = n2354 & ~n2484 ;
  assign n2486 = n2346 & ~n2485 ;
  assign n2487 = n2361 & ~n2486 ;
  assign n2488 = n2369 & ~n2487 ;
  assign n2482 = n2347 & n2369 ;
  assign n2483 = n2333 & n2482 ;
  assign n2489 = n2378 & ~n2483 ;
  assign n2490 = ~n2488 & n2489 ;
  assign n2491 = n1941 & n2490 ;
  assign n2492 = ~n1941 & ~n2490 ;
  assign n2493 = ~n2491 & ~n2492 ;
  assign n2507 = n2124 & ~n2493 ;
  assign n2508 = ~n2497 & ~n2507 ;
  assign n2509 = n2123 & ~n2508 ;
  assign n2494 = n2053 & ~n2493 ;
  assign n2495 = ~n2481 & ~n2494 ;
  assign n2496 = ~n2224 & ~n2495 ;
  assign n2499 = ~n1525 & n2255 ;
  assign n2498 = n1525 & ~n2255 ;
  assign n2500 = n2263 & ~n2498 ;
  assign n2501 = ~n2499 & n2500 ;
  assign n2502 = ~n1445 & ~n2263 ;
  assign n2503 = ~n2501 & ~n2502 ;
  assign n2504 = n2124 & ~n2503 ;
  assign n2505 = ~n2497 & ~n2504 ;
  assign n2506 = n1790 & ~n2505 ;
  assign n2516 = ~n1545 & ~n2274 ;
  assign n2517 = n1540 & n2229 ;
  assign n2518 = ~n2516 & ~n2517 ;
  assign n2519 = ~n2506 & n2518 ;
  assign n2520 = ~n2496 & n2519 ;
  assign n2521 = ~n2509 & n2520 ;
  assign n2522 = ~n2515 & n2521 ;
  assign n2523 = n2037 & ~n2522 ;
  assign n2524 = ~n2480 & ~n2523 ;
  assign n2525 = \P1_state_reg[0]/NET0131  & ~n2524 ;
  assign n2478 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[24]/NET0131  ;
  assign n2479 = ~n1545 & n2014 ;
  assign n2526 = ~n2478 & ~n2479 ;
  assign n2527 = ~n2525 & n2526 ;
  assign n2528 = \P2_reg2_reg[24]/NET0131  & ~n2286 ;
  assign n2529 = \P2_reg2_reg[24]/NET0131  & n2035 ;
  assign n2535 = \P2_reg2_reg[24]/NET0131  & ~n2291 ;
  assign n2536 = n2291 & ~n2512 ;
  assign n2537 = ~n2535 & ~n2536 ;
  assign n2538 = ~n2290 & ~n2537 ;
  assign n2531 = \P2_reg2_reg[24]/NET0131  & ~n2310 ;
  assign n2532 = n2310 & ~n2512 ;
  assign n2533 = ~n2531 & ~n2532 ;
  assign n2534 = n2314 & ~n2533 ;
  assign n2539 = n2291 & ~n2493 ;
  assign n2540 = ~n2535 & ~n2539 ;
  assign n2541 = ~n2392 & ~n2540 ;
  assign n2542 = n2310 & ~n2503 ;
  assign n2543 = ~n2531 & ~n2542 ;
  assign n2544 = n1790 & ~n2543 ;
  assign n2530 = n1540 & n2394 ;
  assign n2545 = \P2_reg2_reg[24]/NET0131  & ~n2407 ;
  assign n2546 = ~n1545 & n1854 ;
  assign n2547 = ~n2545 & ~n2546 ;
  assign n2548 = ~n2530 & n2547 ;
  assign n2549 = ~n2544 & n2548 ;
  assign n2550 = ~n2541 & n2549 ;
  assign n2551 = ~n2534 & n2550 ;
  assign n2552 = ~n2538 & n2551 ;
  assign n2553 = n2037 & ~n2552 ;
  assign n2554 = ~n2529 & ~n2553 ;
  assign n2555 = \P1_state_reg[0]/NET0131  & ~n2554 ;
  assign n2556 = ~n2528 & ~n2555 ;
  assign n2557 = \P2_reg0_reg[29]/NET0131  & ~n2286 ;
  assign n2558 = \P2_reg0_reg[29]/NET0131  & n2035 ;
  assign n2559 = \P2_reg0_reg[29]/NET0131  & ~n2124 ;
  assign n2560 = n2056 & n2093 ;
  assign n2561 = n2055 & n2075 ;
  assign n2562 = n2560 & n2561 ;
  assign n2563 = n2072 & n2076 ;
  assign n2564 = n2081 & ~n2563 ;
  assign n2565 = n2063 & n2065 ;
  assign n2566 = n2058 & n2065 ;
  assign n2567 = ~n2070 & ~n2566 ;
  assign n2568 = ~n2565 & n2567 ;
  assign n2569 = n2066 & n2076 ;
  assign n2570 = ~n2568 & n2569 ;
  assign n2571 = n2564 & ~n2570 ;
  assign n2572 = n2562 & ~n2571 ;
  assign n2573 = n2055 & n2083 ;
  assign n2574 = ~n2087 & ~n2573 ;
  assign n2575 = n2560 & ~n2574 ;
  assign n2576 = n2089 & n2093 ;
  assign n2577 = n2105 & ~n2576 ;
  assign n2578 = ~n2575 & n2577 ;
  assign n2579 = ~n2572 & n2578 ;
  assign n2580 = n2094 & n2097 ;
  assign n2581 = ~n1624 & ~n1760 ;
  assign n2582 = n2096 & n2581 ;
  assign n2583 = n2580 & n2582 ;
  assign n2584 = ~n2579 & n2583 ;
  assign n2586 = n2097 & n2107 ;
  assign n2587 = n2102 & ~n2586 ;
  assign n2588 = n2582 & ~n2587 ;
  assign n2585 = n2110 & n2581 ;
  assign n2589 = n1619 & ~n1760 ;
  assign n2590 = ~n1694 & ~n2589 ;
  assign n2591 = ~n2585 & n2590 ;
  assign n2592 = ~n2588 & n2591 ;
  assign n2593 = ~n2584 & n2592 ;
  assign n2594 = ~n1892 & n2593 ;
  assign n2595 = n1892 & ~n2593 ;
  assign n2596 = ~n2594 & ~n2595 ;
  assign n2597 = n2124 & n2596 ;
  assign n2598 = ~n2559 & ~n2597 ;
  assign n2599 = ~n2120 & ~n2598 ;
  assign n2600 = \P2_reg0_reg[29]/NET0131  & ~n2053 ;
  assign n2601 = ~n1693 & ~n2263 ;
  assign n2602 = n1750 & ~n2399 ;
  assign n2603 = ~n1750 & n2399 ;
  assign n2604 = \P2_B_reg/NET0131  & n633 ;
  assign n2605 = n2263 & ~n2604 ;
  assign n2606 = ~n2603 & n2605 ;
  assign n2607 = ~n2602 & n2606 ;
  assign n2608 = ~n2601 & ~n2607 ;
  assign n2609 = n2053 & ~n2608 ;
  assign n2610 = ~n2600 & ~n2609 ;
  assign n2611 = n1790 & ~n2610 ;
  assign n2612 = ~n1854 & ~n2271 ;
  assign n2613 = ~n2124 & n2272 ;
  assign n2614 = n2612 & ~n2613 ;
  assign n2615 = \P2_reg0_reg[29]/NET0131  & ~n2614 ;
  assign n2616 = n2124 & n2272 ;
  assign n2617 = n1656 & n2616 ;
  assign n2661 = ~n2615 & ~n2617 ;
  assign n2662 = ~n2611 & n2661 ;
  assign n2663 = ~n2599 & n2662 ;
  assign n2618 = n2127 & n2197 ;
  assign n2619 = n2129 & n2169 ;
  assign n2620 = n2618 & n2619 ;
  assign n2621 = ~n2164 & n2170 ;
  assign n2622 = n2175 & ~n2621 ;
  assign n2623 = n2147 & n2155 ;
  assign n2624 = ~n2150 & n2155 ;
  assign n2625 = ~n2160 & ~n2624 ;
  assign n2626 = ~n2623 & n2625 ;
  assign n2627 = n2153 & n2170 ;
  assign n2628 = ~n2626 & n2627 ;
  assign n2629 = n2622 & ~n2628 ;
  assign n2630 = n2620 & ~n2629 ;
  assign n2631 = n2129 & ~n2180 ;
  assign n2632 = n2185 & ~n2631 ;
  assign n2633 = n2618 & ~n2632 ;
  assign n2634 = ~n2189 & n2197 ;
  assign n2635 = n2208 & ~n2634 ;
  assign n2636 = ~n2633 & n2635 ;
  assign n2637 = ~n2630 & n2636 ;
  assign n2638 = n2193 & n2195 ;
  assign n2639 = ~n1886 & ~n1936 ;
  assign n2640 = n2365 & n2639 ;
  assign n2641 = n2638 & n2640 ;
  assign n2642 = ~n2637 & n2641 ;
  assign n2643 = ~n2202 & n2365 ;
  assign n2644 = ~n1889 & ~n2643 ;
  assign n2645 = ~n1886 & ~n2644 ;
  assign n2646 = n2193 & ~n2211 ;
  assign n2647 = n2204 & ~n2646 ;
  assign n2648 = n2640 & ~n2647 ;
  assign n2649 = ~n1887 & ~n2648 ;
  assign n2650 = ~n2645 & n2649 ;
  assign n2651 = ~n2642 & n2650 ;
  assign n2652 = ~n1892 & n2651 ;
  assign n2653 = n1892 & ~n2651 ;
  assign n2654 = ~n2652 & ~n2653 ;
  assign n2655 = n2053 & ~n2654 ;
  assign n2656 = ~n2600 & ~n2655 ;
  assign n2657 = n2123 & ~n2656 ;
  assign n2658 = n2124 & ~n2654 ;
  assign n2659 = ~n2559 & ~n2658 ;
  assign n2660 = ~n2224 & ~n2659 ;
  assign n2664 = ~n2657 & ~n2660 ;
  assign n2665 = n2663 & n2664 ;
  assign n2666 = n2037 & ~n2665 ;
  assign n2667 = ~n2558 & ~n2666 ;
  assign n2668 = \P1_state_reg[0]/NET0131  & ~n2667 ;
  assign n2669 = ~n2557 & ~n2668 ;
  assign n2671 = ~\P1_IR_reg[10]/NET0131  & n497 ;
  assign n2672 = ~\P1_IR_reg[11]/NET0131  & ~\P1_IR_reg[14]/NET0131  ;
  assign n2673 = n471 & n2672 ;
  assign n2674 = n2671 & n2673 ;
  assign n2670 = ~\P1_IR_reg[16]/NET0131  & n481 ;
  assign n2675 = ~\P1_IR_reg[15]/NET0131  & n2670 ;
  assign n2676 = n2674 & n2675 ;
  assign n2677 = ~\P1_IR_reg[21]/NET0131  & ~\P1_IR_reg[22]/NET0131  ;
  assign n2678 = n480 & n2677 ;
  assign n2679 = n2676 & n2678 ;
  assign n2680 = \P1_IR_reg[31]/NET0131  & ~n2679 ;
  assign n2681 = ~\P1_IR_reg[23]/NET0131  & ~n2680 ;
  assign n2682 = \P1_IR_reg[23]/NET0131  & n2680 ;
  assign n2683 = ~n2681 & ~n2682 ;
  assign n2690 = n473 & n498 ;
  assign n2691 = ~\P1_IR_reg[19]/NET0131  & n2670 ;
  assign n2692 = n2690 & n2691 ;
  assign n2693 = ~\P1_IR_reg[20]/NET0131  & n479 ;
  assign n2694 = n2692 & n2693 ;
  assign n2695 = \P1_IR_reg[31]/NET0131  & ~n2694 ;
  assign n2696 = ~\P1_IR_reg[24]/NET0131  & ~n2695 ;
  assign n2697 = \P1_IR_reg[24]/NET0131  & n2695 ;
  assign n2698 = ~n2696 & ~n2697 ;
  assign n2684 = \P1_IR_reg[25]/NET0131  & ~n486 ;
  assign n2685 = ~\P1_IR_reg[25]/NET0131  & n486 ;
  assign n2686 = ~n2684 & ~n2685 ;
  assign n2687 = ~\P1_IR_reg[26]/NET0131  & ~n505 ;
  assign n2688 = \P1_IR_reg[26]/NET0131  & n505 ;
  assign n2689 = ~n2687 & ~n2688 ;
  assign n2699 = ~n2686 & n2689 ;
  assign n2700 = n2698 & n2699 ;
  assign n2701 = ~n2683 & ~n2700 ;
  assign n2702 = n2686 & n2689 ;
  assign n2705 = ~\P1_B_reg/NET0131  & n2698 ;
  assign n2706 = n2702 & n2705 ;
  assign n2707 = ~\P1_d_reg[0]/NET0131  & ~n2706 ;
  assign n2708 = n2689 & ~n2707 ;
  assign n2703 = \P1_B_reg/NET0131  & ~n2698 ;
  assign n2704 = n2702 & n2703 ;
  assign n2709 = ~n2689 & n2698 ;
  assign n2710 = ~n2704 & ~n2709 ;
  assign n2711 = ~n2708 & n2710 ;
  assign n2712 = \P1_d_reg[1]/NET0131  & n2689 ;
  assign n2713 = ~n2686 & ~n2689 ;
  assign n2714 = ~n2712 & ~n2713 ;
  assign n2715 = ~n2704 & n2714 ;
  assign n2716 = ~n2706 & n2715 ;
  assign n2717 = n2711 & ~n2716 ;
  assign n2718 = \P1_reg2_reg[29]/NET0131  & ~n2717 ;
  assign n2719 = ~\P1_IR_reg[24]/NET0131  & n488 ;
  assign n2720 = ~\P1_IR_reg[23]/NET0131  & n2719 ;
  assign n2721 = \P1_IR_reg[31]/NET0131  & ~n2720 ;
  assign n2722 = ~n2680 & ~n2721 ;
  assign n2723 = \P1_IR_reg[27]/NET0131  & ~n2722 ;
  assign n2724 = ~\P1_IR_reg[27]/NET0131  & n2722 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = ~\P1_IR_reg[27]/NET0131  & n2719 ;
  assign n2727 = \P1_IR_reg[31]/NET0131  & ~n2726 ;
  assign n2728 = ~n2695 & ~n2727 ;
  assign n2729 = \P1_IR_reg[28]/NET0131  & ~n2728 ;
  assign n2730 = ~\P1_IR_reg[28]/NET0131  & n2728 ;
  assign n2731 = ~n2729 & ~n2730 ;
  assign n2732 = ~n2725 & ~n2731 ;
  assign n2733 = \P2_datao_reg[28]/NET0131  & n639 ;
  assign n2734 = ~\P2_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n2735 = \P2_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n2736 = ~n2734 & ~n2735 ;
  assign n2737 = ~\P2_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n2738 = ~\P2_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n2739 = ~n2737 & ~n2738 ;
  assign n2740 = ~\P2_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n2741 = \P2_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n2742 = \P2_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n2743 = ~n2741 & ~n2742 ;
  assign n2744 = ~n2740 & ~n2743 ;
  assign n2745 = n2739 & n2744 ;
  assign n2746 = \P2_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n2747 = \P2_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n2748 = ~n2746 & ~n2747 ;
  assign n2749 = ~n2738 & ~n2748 ;
  assign n2750 = ~n2745 & ~n2749 ;
  assign n2751 = ~\P2_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n2752 = ~n2740 & ~n2751 ;
  assign n2753 = n2739 & n2752 ;
  assign n2754 = \P2_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n2755 = ~\P2_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n2756 = ~\P2_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n2757 = ~n2755 & ~n2756 ;
  assign n2758 = ~\P2_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n2759 = ~\P2_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n2760 = ~\P2_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n2761 = \P2_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n2762 = \P2_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n2763 = ~n2761 & ~n2762 ;
  assign n2764 = ~n2760 & ~n2763 ;
  assign n2765 = ~n2759 & n2764 ;
  assign n2766 = \P2_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n2767 = \P2_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n2768 = ~n2766 & ~n2767 ;
  assign n2769 = ~n2765 & n2768 ;
  assign n2770 = ~n2758 & ~n2769 ;
  assign n2771 = n2757 & n2770 ;
  assign n2772 = \P2_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n2773 = \P2_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n2774 = \P2_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n2775 = ~n2773 & ~n2774 ;
  assign n2776 = ~n2756 & ~n2775 ;
  assign n2777 = ~n2772 & ~n2776 ;
  assign n2778 = ~n2771 & n2777 ;
  assign n2779 = ~\P2_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n2780 = ~\P2_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n2781 = ~n2779 & ~n2780 ;
  assign n2782 = ~n2778 & n2781 ;
  assign n2783 = ~n2754 & ~n2782 ;
  assign n2784 = ~\P2_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n2785 = ~\P2_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n2786 = ~n2784 & ~n2785 ;
  assign n2787 = ~\P2_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n2788 = n2786 & ~n2787 ;
  assign n2789 = ~\P2_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n2790 = n2788 & ~n2789 ;
  assign n2791 = ~n2783 & n2790 ;
  assign n2792 = ~\P2_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n2793 = ~\P2_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n2794 = ~n2792 & ~n2793 ;
  assign n2795 = ~\P2_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n2796 = ~\P2_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n2797 = ~n2795 & ~n2796 ;
  assign n2798 = n2794 & n2797 ;
  assign n2799 = n2791 & n2798 ;
  assign n2805 = \P2_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n2806 = \P2_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n2807 = \P2_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n2808 = \P2_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n2809 = ~n2807 & ~n2808 ;
  assign n2810 = ~n2785 & ~n2809 ;
  assign n2811 = ~n2806 & ~n2810 ;
  assign n2812 = ~n2784 & ~n2789 ;
  assign n2813 = ~n2811 & n2812 ;
  assign n2814 = ~n2805 & ~n2813 ;
  assign n2815 = n2798 & ~n2814 ;
  assign n2800 = \P2_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n2801 = \P2_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n2802 = ~n2800 & ~n2801 ;
  assign n2803 = ~n2796 & ~n2802 ;
  assign n2804 = n2794 & n2803 ;
  assign n2816 = \P2_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n2817 = \P2_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n2818 = ~n2816 & ~n2817 ;
  assign n2819 = ~n2792 & ~n2818 ;
  assign n2820 = ~n2804 & ~n2819 ;
  assign n2821 = ~n2815 & n2820 ;
  assign n2822 = ~n2799 & n2821 ;
  assign n2823 = n2753 & ~n2822 ;
  assign n2824 = n2750 & ~n2823 ;
  assign n2825 = ~\P2_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n2831 = ~\P2_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n2832 = ~\P2_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n2833 = ~\P2_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2835 = ~n2831 & n2834 ;
  assign n2826 = ~\P2_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n2827 = ~\P2_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n2828 = ~\P2_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n2829 = ~n2827 & ~n2828 ;
  assign n2830 = ~n2826 & n2829 ;
  assign n2836 = ~\P2_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n2837 = n2830 & ~n2836 ;
  assign n2838 = n2835 & n2837 ;
  assign n2839 = ~n2825 & n2838 ;
  assign n2840 = ~n2824 & n2839 ;
  assign n2844 = \P2_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n2845 = \P2_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n2846 = ~n2844 & ~n2845 ;
  assign n2847 = ~n2826 & ~n2846 ;
  assign n2848 = \P2_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n2849 = \P2_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n2850 = ~n2848 & ~n2849 ;
  assign n2851 = n2830 & ~n2850 ;
  assign n2852 = ~n2847 & ~n2851 ;
  assign n2853 = n2835 & ~n2852 ;
  assign n2841 = \P2_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n2842 = \P2_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n2843 = ~n2841 & ~n2842 ;
  assign n2854 = \P2_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n2855 = \P2_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n2856 = ~n2854 & ~n2855 ;
  assign n2857 = ~n2832 & ~n2856 ;
  assign n2858 = ~n2831 & n2857 ;
  assign n2859 = n2843 & ~n2858 ;
  assign n2860 = ~n2853 & n2859 ;
  assign n2861 = ~n2836 & ~n2860 ;
  assign n2862 = ~n2840 & ~n2861 ;
  assign n2864 = ~n2736 & n2862 ;
  assign n2863 = n2736 & ~n2862 ;
  assign n2865 = ~n639 & ~n2863 ;
  assign n2866 = ~n2864 & n2865 ;
  assign n2867 = ~n2733 & ~n2866 ;
  assign n2868 = ~n2732 & ~n2867 ;
  assign n2872 = \P1_reg3_reg[3]/NET0131  & \P1_reg3_reg[4]/NET0131  ;
  assign n2873 = \P1_reg3_reg[5]/NET0131  & n2872 ;
  assign n2874 = \P1_reg3_reg[6]/NET0131  & n2873 ;
  assign n2875 = \P1_reg3_reg[10]/NET0131  & \P1_reg3_reg[7]/NET0131  ;
  assign n2876 = \P1_reg3_reg[8]/NET0131  & \P1_reg3_reg[9]/NET0131  ;
  assign n2877 = n2875 & n2876 ;
  assign n2878 = n2874 & n2877 ;
  assign n2879 = \P1_reg3_reg[11]/NET0131  & \P1_reg3_reg[12]/NET0131  ;
  assign n2880 = n2878 & n2879 ;
  assign n2881 = \P1_reg3_reg[13]/NET0131  & n2880 ;
  assign n2882 = \P1_reg3_reg[14]/NET0131  & n2881 ;
  assign n2883 = \P1_reg3_reg[16]/NET0131  & \P1_reg3_reg[17]/NET0131  ;
  assign n2884 = \P1_reg3_reg[15]/NET0131  & \P1_reg3_reg[18]/NET0131  ;
  assign n2885 = \P1_reg3_reg[19]/NET0131  & \P1_reg3_reg[20]/NET0131  ;
  assign n2886 = n2884 & n2885 ;
  assign n2887 = n2883 & n2886 ;
  assign n2888 = n2882 & n2887 ;
  assign n2889 = \P1_reg3_reg[21]/NET0131  & \P1_reg3_reg[22]/NET0131  ;
  assign n2890 = n2888 & n2889 ;
  assign n2891 = \P1_reg3_reg[23]/NET0131  & n2890 ;
  assign n2892 = \P1_reg3_reg[24]/NET0131  & n2891 ;
  assign n2893 = \P1_reg3_reg[25]/NET0131  & \P1_reg3_reg[26]/NET0131  ;
  assign n2894 = n2892 & n2893 ;
  assign n2895 = \P1_reg3_reg[27]/NET0131  & n2894 ;
  assign n2896 = ~\P1_reg3_reg[28]/NET0131  & ~n2895 ;
  assign n2897 = \P1_reg3_reg[27]/NET0131  & \P1_reg3_reg[28]/NET0131  ;
  assign n2898 = n2893 & n2897 ;
  assign n2899 = n2892 & n2898 ;
  assign n2900 = ~n2896 & ~n2899 ;
  assign n2901 = n519 & n2900 ;
  assign n2871 = \P1_reg0_reg[28]/NET0131  & n517 ;
  assign n2869 = \P1_reg2_reg[28]/NET0131  & n513 ;
  assign n2870 = \P1_reg1_reg[28]/NET0131  & n515 ;
  assign n2902 = ~n2869 & ~n2870 ;
  assign n2903 = ~n2871 & n2902 ;
  assign n2904 = ~n2901 & n2903 ;
  assign n2905 = ~n2868 & n2904 ;
  assign n2906 = \P2_datao_reg[25]/NET0131  & n639 ;
  assign n2907 = ~n2832 & ~n2854 ;
  assign n2908 = ~n2742 & ~n2746 ;
  assign n2909 = ~n2737 & ~n2908 ;
  assign n2910 = ~n2738 & ~n2825 ;
  assign n2911 = n2909 & n2910 ;
  assign n2912 = ~n2747 & ~n2848 ;
  assign n2913 = ~n2825 & ~n2912 ;
  assign n2914 = ~n2911 & ~n2913 ;
  assign n2915 = ~n2737 & ~n2740 ;
  assign n2916 = n2910 & n2915 ;
  assign n2917 = ~n2770 & ~n2774 ;
  assign n2918 = n2757 & ~n2779 ;
  assign n2919 = ~n2780 & ~n2787 ;
  assign n2920 = n2918 & n2919 ;
  assign n2921 = ~n2917 & n2920 ;
  assign n2922 = ~n2772 & ~n2773 ;
  assign n2923 = ~n2779 & ~n2922 ;
  assign n2924 = ~n2754 & ~n2923 ;
  assign n2925 = n2919 & ~n2924 ;
  assign n2926 = ~n2808 & ~n2925 ;
  assign n2927 = ~n2921 & n2926 ;
  assign n2928 = ~n2789 & ~n2795 ;
  assign n2929 = n2786 & n2928 ;
  assign n2930 = ~n2927 & n2929 ;
  assign n2931 = ~n2751 & ~n2792 ;
  assign n2932 = ~n2793 & n2931 ;
  assign n2933 = ~n2796 & n2932 ;
  assign n2934 = n2930 & n2933 ;
  assign n2935 = ~n2741 & ~n2817 ;
  assign n2936 = ~n2751 & ~n2935 ;
  assign n2937 = ~n2801 & ~n2816 ;
  assign n2938 = n2932 & ~n2937 ;
  assign n2939 = ~n2936 & ~n2938 ;
  assign n2940 = ~n2806 & ~n2807 ;
  assign n2941 = ~n2784 & ~n2940 ;
  assign n2942 = ~n2805 & ~n2941 ;
  assign n2943 = n2928 & ~n2942 ;
  assign n2944 = ~n2800 & ~n2943 ;
  assign n2945 = n2933 & ~n2944 ;
  assign n2946 = n2939 & ~n2945 ;
  assign n2947 = ~n2934 & n2946 ;
  assign n2948 = n2916 & ~n2947 ;
  assign n2949 = n2914 & ~n2948 ;
  assign n2950 = n2830 & ~n2833 ;
  assign n2951 = ~n2949 & n2950 ;
  assign n2952 = ~n2844 & ~n2855 ;
  assign n2953 = ~n2845 & ~n2849 ;
  assign n2954 = ~n2828 & ~n2953 ;
  assign n2955 = ~n2826 & n2954 ;
  assign n2956 = n2952 & ~n2955 ;
  assign n2957 = ~n2833 & ~n2956 ;
  assign n2958 = ~n2951 & ~n2957 ;
  assign n2960 = ~n2907 & n2958 ;
  assign n2959 = n2907 & ~n2958 ;
  assign n2961 = ~n639 & ~n2959 ;
  assign n2962 = ~n2960 & n2961 ;
  assign n2963 = ~n2906 & ~n2962 ;
  assign n2964 = ~n2732 & ~n2963 ;
  assign n2968 = \P1_reg3_reg[25]/NET0131  & n2892 ;
  assign n2969 = ~\P1_reg3_reg[25]/NET0131  & ~n2892 ;
  assign n2970 = ~n2968 & ~n2969 ;
  assign n2971 = n519 & n2970 ;
  assign n2967 = \P1_reg2_reg[25]/NET0131  & n513 ;
  assign n2965 = \P1_reg0_reg[25]/NET0131  & n517 ;
  assign n2966 = \P1_reg1_reg[25]/NET0131  & n515 ;
  assign n2972 = ~n2965 & ~n2966 ;
  assign n2973 = ~n2967 & n2972 ;
  assign n2974 = ~n2971 & n2973 ;
  assign n2975 = ~n2964 & n2974 ;
  assign n2976 = \P2_datao_reg[26]/NET0131  & n639 ;
  assign n2977 = ~n2831 & ~n2841 ;
  assign n2978 = ~n2771 & ~n2776 ;
  assign n2979 = ~n2785 & n2919 ;
  assign n2980 = ~n2779 & n2979 ;
  assign n2981 = ~n2978 & n2980 ;
  assign n2982 = ~n2754 & ~n2772 ;
  assign n2983 = n2979 & ~n2982 ;
  assign n2984 = ~n2810 & ~n2983 ;
  assign n2985 = ~n2981 & n2984 ;
  assign n2986 = n2797 & n2812 ;
  assign n2987 = ~n2985 & n2986 ;
  assign n2988 = ~n2740 & n2932 ;
  assign n2989 = n2987 & n2988 ;
  assign n2990 = ~n2805 & ~n2806 ;
  assign n2991 = ~n2796 & n2928 ;
  assign n2992 = ~n2990 & n2991 ;
  assign n2993 = ~n2803 & ~n2992 ;
  assign n2994 = n2988 & ~n2993 ;
  assign n2995 = n2752 & n2819 ;
  assign n2996 = ~n2744 & ~n2995 ;
  assign n2997 = ~n2994 & n2996 ;
  assign n2998 = ~n2989 & n2997 ;
  assign n2999 = ~n2825 & ~n2827 ;
  assign n3000 = n2739 & n2999 ;
  assign n3001 = ~n2998 & n3000 ;
  assign n3002 = n2749 & ~n2825 ;
  assign n3003 = n2850 & ~n3002 ;
  assign n3004 = ~n2827 & ~n3003 ;
  assign n3005 = ~n3001 & ~n3004 ;
  assign n3006 = ~n2826 & ~n2828 ;
  assign n3007 = n2834 & n3006 ;
  assign n3008 = ~n3005 & n3007 ;
  assign n3009 = n2834 & n2847 ;
  assign n3010 = ~n2857 & ~n3009 ;
  assign n3011 = ~n3008 & n3010 ;
  assign n3013 = ~n2977 & n3011 ;
  assign n3012 = n2977 & ~n3011 ;
  assign n3014 = ~n639 & ~n3012 ;
  assign n3015 = ~n3013 & n3014 ;
  assign n3016 = ~n2976 & ~n3015 ;
  assign n3017 = ~n2732 & ~n3016 ;
  assign n3021 = ~\P1_reg3_reg[26]/NET0131  & ~n2968 ;
  assign n3022 = ~n2894 & ~n3021 ;
  assign n3023 = n519 & n3022 ;
  assign n3020 = \P1_reg0_reg[26]/NET0131  & n517 ;
  assign n3018 = \P1_reg2_reg[26]/NET0131  & n513 ;
  assign n3019 = \P1_reg1_reg[26]/NET0131  & n515 ;
  assign n3024 = ~n3018 & ~n3019 ;
  assign n3025 = ~n3020 & n3024 ;
  assign n3026 = ~n3023 & n3025 ;
  assign n3027 = ~n3017 & n3026 ;
  assign n3028 = \P2_datao_reg[27]/NET0131  & n639 ;
  assign n3029 = ~n2836 & ~n2842 ;
  assign n3030 = ~n2841 & ~n2854 ;
  assign n3031 = ~n2831 & ~n3030 ;
  assign n3032 = n2835 & ~n2952 ;
  assign n3033 = ~n3031 & ~n3032 ;
  assign n3034 = ~n2826 & n2835 ;
  assign n3039 = ~n2917 & n2918 ;
  assign n3040 = ~n2923 & ~n3039 ;
  assign n3041 = n2786 & n2919 ;
  assign n3042 = ~n3040 & n3041 ;
  assign n3037 = ~n2754 & ~n2808 ;
  assign n3038 = n2788 & ~n3037 ;
  assign n3043 = ~n2941 & ~n3038 ;
  assign n3044 = ~n3042 & n3043 ;
  assign n3045 = ~n2793 & n2991 ;
  assign n3046 = ~n3044 & n3045 ;
  assign n3047 = n2829 & n2910 ;
  assign n3048 = n2915 & n2931 ;
  assign n3049 = n3047 & n3048 ;
  assign n3050 = n3046 & n3049 ;
  assign n3035 = n2829 & n2913 ;
  assign n3036 = ~n2954 & ~n3035 ;
  assign n3051 = ~n2800 & ~n2805 ;
  assign n3052 = n2797 & ~n3051 ;
  assign n3053 = n2937 & ~n3052 ;
  assign n3054 = ~n2793 & ~n3053 ;
  assign n3055 = n3048 & n3054 ;
  assign n3056 = n2915 & n2936 ;
  assign n3057 = ~n2909 & ~n3056 ;
  assign n3058 = ~n3055 & n3057 ;
  assign n3059 = n3047 & ~n3058 ;
  assign n3060 = n3036 & ~n3059 ;
  assign n3061 = ~n3050 & n3060 ;
  assign n3062 = n3034 & ~n3061 ;
  assign n3063 = n3033 & ~n3062 ;
  assign n3065 = ~n3029 & n3063 ;
  assign n3064 = n3029 & ~n3063 ;
  assign n3066 = ~n639 & ~n3064 ;
  assign n3067 = ~n3065 & n3066 ;
  assign n3068 = ~n3028 & ~n3067 ;
  assign n3069 = ~n2732 & ~n3068 ;
  assign n3073 = ~\P1_reg3_reg[27]/NET0131  & ~n2894 ;
  assign n3074 = ~n2895 & ~n3073 ;
  assign n3075 = n519 & n3074 ;
  assign n3072 = \P1_reg1_reg[27]/NET0131  & n515 ;
  assign n3070 = \P1_reg0_reg[27]/NET0131  & n517 ;
  assign n3071 = \P1_reg2_reg[27]/NET0131  & n513 ;
  assign n3076 = ~n3070 & ~n3071 ;
  assign n3077 = ~n3072 & n3076 ;
  assign n3078 = ~n3075 & n3077 ;
  assign n3079 = ~n3069 & n3078 ;
  assign n3080 = ~n3027 & ~n3079 ;
  assign n3081 = ~n2975 & n3080 ;
  assign n3082 = \P2_datao_reg[24]/NET0131  & n639 ;
  assign n3083 = ~n2833 & ~n2855 ;
  assign n3084 = n2753 & n2799 ;
  assign n3085 = n2753 & ~n2821 ;
  assign n3086 = n2750 & ~n3085 ;
  assign n3087 = ~n3084 & n3086 ;
  assign n3088 = ~n2825 & n2830 ;
  assign n3089 = ~n3087 & n3088 ;
  assign n3090 = n2852 & ~n3089 ;
  assign n3092 = ~n3083 & n3090 ;
  assign n3091 = n3083 & ~n3090 ;
  assign n3093 = ~n639 & ~n3091 ;
  assign n3094 = ~n3092 & n3093 ;
  assign n3095 = ~n3082 & ~n3094 ;
  assign n3096 = ~n2732 & ~n3095 ;
  assign n3097 = \P1_reg0_reg[24]/NET0131  & n517 ;
  assign n3098 = \P1_reg1_reg[24]/NET0131  & n515 ;
  assign n3103 = ~n3097 & ~n3098 ;
  assign n3099 = \P1_reg2_reg[24]/NET0131  & n513 ;
  assign n3100 = ~\P1_reg3_reg[24]/NET0131  & ~n2891 ;
  assign n3101 = ~n2892 & ~n3100 ;
  assign n3102 = n519 & n3101 ;
  assign n3104 = ~n3099 & ~n3102 ;
  assign n3105 = n3103 & n3104 ;
  assign n3106 = ~n3096 & n3105 ;
  assign n3107 = \P2_datao_reg[23]/NET0131  & n639 ;
  assign n3108 = ~n2826 & ~n2844 ;
  assign n3110 = ~n3046 & ~n3054 ;
  assign n3111 = n3049 & ~n3110 ;
  assign n3109 = n3047 & ~n3057 ;
  assign n3112 = n3036 & ~n3109 ;
  assign n3113 = ~n3111 & n3112 ;
  assign n3115 = ~n3108 & n3113 ;
  assign n3114 = n3108 & ~n3113 ;
  assign n3116 = ~n639 & ~n3114 ;
  assign n3117 = ~n3115 & n3116 ;
  assign n3118 = ~n3107 & ~n3117 ;
  assign n3119 = ~n2732 & ~n3118 ;
  assign n3120 = ~\P1_reg3_reg[23]/NET0131  & ~n2890 ;
  assign n3121 = ~n2891 & ~n3120 ;
  assign n3122 = n519 & n3121 ;
  assign n3123 = \P1_reg1_reg[23]/NET0131  & n515 ;
  assign n3126 = ~n3122 & ~n3123 ;
  assign n3124 = \P1_reg2_reg[23]/NET0131  & n513 ;
  assign n3125 = \P1_reg0_reg[23]/NET0131  & n517 ;
  assign n3127 = ~n3124 & ~n3125 ;
  assign n3128 = n3126 & n3127 ;
  assign n3129 = ~n3119 & n3128 ;
  assign n3130 = ~n3106 & ~n3129 ;
  assign n3131 = \P2_datao_reg[22]/NET0131  & n639 ;
  assign n3132 = ~n2828 & ~n2845 ;
  assign n3133 = ~n2987 & n2993 ;
  assign n3134 = n2988 & ~n3133 ;
  assign n3135 = n2996 & ~n3134 ;
  assign n3136 = n3000 & ~n3135 ;
  assign n3137 = ~n3004 & ~n3136 ;
  assign n3139 = ~n3132 & n3137 ;
  assign n3138 = n3132 & ~n3137 ;
  assign n3140 = ~n639 & ~n3138 ;
  assign n3141 = ~n3139 & n3140 ;
  assign n3142 = ~n3131 & ~n3141 ;
  assign n3143 = ~n2732 & ~n3142 ;
  assign n3144 = \P1_reg0_reg[22]/NET0131  & n517 ;
  assign n3145 = \P1_reg1_reg[22]/NET0131  & n515 ;
  assign n3151 = ~n3144 & ~n3145 ;
  assign n3146 = \P1_reg2_reg[22]/NET0131  & n513 ;
  assign n3147 = \P1_reg3_reg[21]/NET0131  & n2888 ;
  assign n3148 = ~\P1_reg3_reg[22]/NET0131  & ~n3147 ;
  assign n3149 = ~n2890 & ~n3148 ;
  assign n3150 = n519 & n3149 ;
  assign n3152 = ~n3146 & ~n3150 ;
  assign n3153 = n3151 & n3152 ;
  assign n3154 = n3143 & ~n3153 ;
  assign n3155 = ~n3143 & n3153 ;
  assign n3156 = \P2_datao_reg[21]/NET0131  & n639 ;
  assign n3157 = ~n2827 & ~n2849 ;
  assign n3158 = ~n2930 & n2944 ;
  assign n3159 = n2933 & ~n3158 ;
  assign n3160 = n2939 & ~n3159 ;
  assign n3161 = n2916 & ~n3160 ;
  assign n3162 = n2914 & ~n3161 ;
  assign n3164 = ~n3157 & n3162 ;
  assign n3163 = n3157 & ~n3162 ;
  assign n3165 = ~n639 & ~n3163 ;
  assign n3166 = ~n3164 & n3165 ;
  assign n3167 = ~n3156 & ~n3166 ;
  assign n3168 = ~n2732 & ~n3167 ;
  assign n3169 = \P1_reg2_reg[21]/NET0131  & n513 ;
  assign n3170 = \P1_reg1_reg[21]/NET0131  & n515 ;
  assign n3175 = ~n3169 & ~n3170 ;
  assign n3171 = ~\P1_reg3_reg[21]/NET0131  & ~n2888 ;
  assign n3172 = ~n3147 & ~n3171 ;
  assign n3173 = n519 & n3172 ;
  assign n3174 = \P1_reg0_reg[21]/NET0131  & n517 ;
  assign n3176 = ~n3173 & ~n3174 ;
  assign n3177 = n3175 & n3176 ;
  assign n3178 = n3168 & ~n3177 ;
  assign n3179 = ~n3155 & n3178 ;
  assign n3180 = ~n3154 & ~n3179 ;
  assign n3181 = n3130 & ~n3180 ;
  assign n3182 = n3096 & ~n3105 ;
  assign n3183 = n3119 & ~n3128 ;
  assign n3184 = ~n3106 & n3183 ;
  assign n3185 = ~n3182 & ~n3184 ;
  assign n3186 = ~n3181 & n3185 ;
  assign n3187 = n3081 & ~n3186 ;
  assign n3189 = n3017 & ~n3026 ;
  assign n3190 = n2964 & ~n2974 ;
  assign n3191 = ~n3189 & ~n3190 ;
  assign n3192 = n3080 & ~n3191 ;
  assign n3188 = n3069 & ~n3078 ;
  assign n3193 = n2868 & ~n2904 ;
  assign n3194 = ~n3188 & ~n3193 ;
  assign n3195 = ~n3192 & n3194 ;
  assign n3196 = ~n3187 & n3195 ;
  assign n3197 = ~n2905 & ~n3196 ;
  assign n3198 = \P1_IR_reg[31]/NET0131  & ~n2671 ;
  assign n3199 = ~\P1_IR_reg[11]/NET0131  & n3198 ;
  assign n3200 = \P1_IR_reg[11]/NET0131  & ~n3198 ;
  assign n3201 = ~n3199 & ~n3200 ;
  assign n3202 = n2732 & n3201 ;
  assign n3203 = \P2_datao_reg[11]/NET0131  & n639 ;
  assign n3204 = ~n2789 & ~n2805 ;
  assign n3206 = n3044 & ~n3204 ;
  assign n3205 = ~n3044 & n3204 ;
  assign n3207 = ~n639 & ~n3205 ;
  assign n3208 = ~n3206 & n3207 ;
  assign n3209 = ~n3203 & ~n3208 ;
  assign n3210 = ~n2732 & n3209 ;
  assign n3211 = ~n3202 & ~n3210 ;
  assign n3212 = \P1_reg3_reg[11]/NET0131  & n2878 ;
  assign n3213 = ~\P1_reg3_reg[11]/NET0131  & ~n2878 ;
  assign n3214 = ~n3212 & ~n3213 ;
  assign n3215 = n519 & n3214 ;
  assign n3216 = \P1_reg1_reg[11]/NET0131  & n515 ;
  assign n3219 = ~n3215 & ~n3216 ;
  assign n3217 = \P1_reg2_reg[11]/NET0131  & n513 ;
  assign n3218 = \P1_reg0_reg[11]/NET0131  & n517 ;
  assign n3220 = ~n3217 & ~n3218 ;
  assign n3221 = n3219 & n3220 ;
  assign n3222 = ~n3211 & n3221 ;
  assign n3223 = \P1_IR_reg[31]/NET0131  & ~n497 ;
  assign n3224 = \P1_IR_reg[31]/NET0131  & ~n470 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = \P1_IR_reg[12]/NET0131  & ~n3225 ;
  assign n3227 = ~\P1_IR_reg[12]/NET0131  & n3225 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = n2732 & ~n3228 ;
  assign n3230 = \P2_datao_reg[12]/NET0131  & n639 ;
  assign n3231 = ~n2795 & ~n2800 ;
  assign n3232 = ~n2791 & n2814 ;
  assign n3234 = ~n3231 & n3232 ;
  assign n3233 = n3231 & ~n3232 ;
  assign n3235 = ~n639 & ~n3233 ;
  assign n3236 = ~n3234 & n3235 ;
  assign n3237 = ~n3230 & ~n3236 ;
  assign n3238 = ~n2732 & n3237 ;
  assign n3239 = ~n3229 & ~n3238 ;
  assign n3240 = \P1_reg2_reg[12]/NET0131  & n513 ;
  assign n3241 = \P1_reg1_reg[12]/NET0131  & n515 ;
  assign n3246 = ~n3240 & ~n3241 ;
  assign n3242 = \P1_reg0_reg[12]/NET0131  & n517 ;
  assign n3243 = ~\P1_reg3_reg[12]/NET0131  & ~n3212 ;
  assign n3244 = ~n2880 & ~n3243 ;
  assign n3245 = n519 & n3244 ;
  assign n3247 = ~n3242 & ~n3245 ;
  assign n3248 = n3246 & n3247 ;
  assign n3249 = ~n3239 & n3248 ;
  assign n3250 = ~n3222 & ~n3249 ;
  assign n3251 = \P1_IR_reg[10]/NET0131  & ~n3223 ;
  assign n3252 = ~\P1_IR_reg[10]/NET0131  & n3223 ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = n2732 & n3253 ;
  assign n3255 = \P2_datao_reg[10]/NET0131  & n639 ;
  assign n3256 = ~n2784 & ~n2806 ;
  assign n3258 = n2985 & ~n3256 ;
  assign n3257 = ~n2985 & n3256 ;
  assign n3259 = ~n639 & ~n3257 ;
  assign n3260 = ~n3258 & n3259 ;
  assign n3261 = ~n3255 & ~n3260 ;
  assign n3262 = ~n2732 & n3261 ;
  assign n3263 = ~n3254 & ~n3262 ;
  assign n3264 = \P1_reg2_reg[10]/NET0131  & n513 ;
  assign n3265 = \P1_reg1_reg[10]/NET0131  & n515 ;
  assign n3273 = ~n3264 & ~n3265 ;
  assign n3266 = \P1_reg0_reg[10]/NET0131  & n517 ;
  assign n3267 = \P1_reg3_reg[7]/NET0131  & n2874 ;
  assign n3268 = \P1_reg3_reg[8]/NET0131  & n3267 ;
  assign n3269 = \P1_reg3_reg[9]/NET0131  & n3268 ;
  assign n3270 = ~\P1_reg3_reg[10]/NET0131  & ~n3269 ;
  assign n3271 = ~n2878 & ~n3270 ;
  assign n3272 = n519 & n3271 ;
  assign n3274 = ~n3266 & ~n3272 ;
  assign n3275 = n3273 & n3274 ;
  assign n3276 = ~n3263 & n3275 ;
  assign n3277 = n3263 & ~n3275 ;
  assign n3278 = \P1_IR_reg[31]/NET0131  & ~n469 ;
  assign n3279 = \P1_IR_reg[9]/NET0131  & ~n3278 ;
  assign n3280 = ~\P1_IR_reg[9]/NET0131  & n3278 ;
  assign n3281 = ~n3279 & ~n3280 ;
  assign n3282 = n2732 & n3281 ;
  assign n3283 = \P2_datao_reg[9]/NET0131  & n639 ;
  assign n3284 = ~n2785 & ~n2807 ;
  assign n3286 = n2927 & ~n3284 ;
  assign n3285 = ~n2927 & n3284 ;
  assign n3287 = ~n639 & ~n3285 ;
  assign n3288 = ~n3286 & n3287 ;
  assign n3289 = ~n3283 & ~n3288 ;
  assign n3290 = ~n2732 & n3289 ;
  assign n3291 = ~n3282 & ~n3290 ;
  assign n3292 = \P1_reg2_reg[9]/NET0131  & n513 ;
  assign n3293 = \P1_reg1_reg[9]/NET0131  & n515 ;
  assign n3298 = ~n3292 & ~n3293 ;
  assign n3294 = \P1_reg0_reg[9]/NET0131  & n517 ;
  assign n3295 = ~\P1_reg3_reg[9]/NET0131  & ~n3268 ;
  assign n3296 = ~n3269 & ~n3295 ;
  assign n3297 = n519 & n3296 ;
  assign n3299 = ~n3294 & ~n3297 ;
  assign n3300 = n3298 & n3299 ;
  assign n3301 = n3291 & ~n3300 ;
  assign n3302 = ~n3277 & ~n3301 ;
  assign n3303 = ~n3276 & ~n3302 ;
  assign n3304 = n3250 & n3303 ;
  assign n3305 = n3239 & ~n3248 ;
  assign n3306 = n3211 & ~n3221 ;
  assign n3307 = ~n3305 & ~n3306 ;
  assign n3308 = ~n3249 & ~n3307 ;
  assign n3309 = ~n3304 & ~n3308 ;
  assign n3310 = \P1_reg0_reg[4]/NET0131  & n517 ;
  assign n3311 = ~\P1_reg3_reg[3]/NET0131  & ~\P1_reg3_reg[4]/NET0131  ;
  assign n3312 = ~n2872 & ~n3311 ;
  assign n3313 = n519 & n3312 ;
  assign n3316 = ~n3310 & ~n3313 ;
  assign n3314 = \P1_reg2_reg[4]/NET0131  & n513 ;
  assign n3315 = \P1_reg1_reg[4]/NET0131  & n515 ;
  assign n3317 = ~n3314 & ~n3315 ;
  assign n3318 = n3316 & n3317 ;
  assign n3319 = \P2_datao_reg[4]/NET0131  & n639 ;
  assign n3320 = ~n2755 & ~n2774 ;
  assign n3322 = n2770 & n3320 ;
  assign n3321 = ~n2770 & ~n3320 ;
  assign n3323 = ~n639 & ~n3321 ;
  assign n3324 = ~n3322 & n3323 ;
  assign n3325 = ~n3319 & ~n3324 ;
  assign n3326 = ~n2732 & ~n3325 ;
  assign n3327 = \P1_IR_reg[31]/NET0131  & ~n465 ;
  assign n3328 = \P1_IR_reg[4]/NET0131  & ~n3327 ;
  assign n3329 = ~\P1_IR_reg[4]/NET0131  & n3327 ;
  assign n3330 = ~n3328 & ~n3329 ;
  assign n3331 = n2732 & ~n3330 ;
  assign n3332 = ~n3326 & ~n3331 ;
  assign n3333 = n3318 & n3332 ;
  assign n3334 = \P1_reg3_reg[2]/NET0131  & n519 ;
  assign n3335 = \P1_reg1_reg[2]/NET0131  & n515 ;
  assign n3338 = ~n3334 & ~n3335 ;
  assign n3336 = \P1_reg2_reg[2]/NET0131  & n513 ;
  assign n3337 = \P1_reg0_reg[2]/NET0131  & n517 ;
  assign n3339 = ~n3336 & ~n3337 ;
  assign n3340 = n3338 & n3339 ;
  assign n3341 = \P2_datao_reg[2]/NET0131  & n639 ;
  assign n3342 = ~n2759 & ~n2767 ;
  assign n3344 = n2764 & n3342 ;
  assign n3343 = ~n2764 & ~n3342 ;
  assign n3345 = ~n639 & ~n3343 ;
  assign n3346 = ~n3344 & n3345 ;
  assign n3347 = ~n3341 & ~n3346 ;
  assign n3348 = ~n2732 & ~n3347 ;
  assign n3349 = \P1_IR_reg[31]/NET0131  & ~n463 ;
  assign n3350 = ~\P1_IR_reg[2]/NET0131  & ~n3349 ;
  assign n3351 = \P1_IR_reg[2]/NET0131  & n3349 ;
  assign n3352 = ~n3350 & ~n3351 ;
  assign n3353 = n2732 & n3352 ;
  assign n3354 = ~n3348 & ~n3353 ;
  assign n3355 = n3340 & n3354 ;
  assign n3356 = \P2_datao_reg[3]/NET0131  & n639 ;
  assign n3357 = ~n2765 & ~n2767 ;
  assign n3358 = ~n2758 & ~n2766 ;
  assign n3360 = ~n3357 & n3358 ;
  assign n3359 = n3357 & ~n3358 ;
  assign n3361 = ~n639 & ~n3359 ;
  assign n3362 = ~n3360 & n3361 ;
  assign n3363 = ~n3356 & ~n3362 ;
  assign n3364 = ~n2732 & ~n3363 ;
  assign n3365 = \P1_IR_reg[2]/NET0131  & \P1_IR_reg[31]/NET0131  ;
  assign n3366 = ~n3349 & ~n3365 ;
  assign n3367 = \P1_IR_reg[3]/NET0131  & ~n3366 ;
  assign n3368 = ~\P1_IR_reg[3]/NET0131  & n3366 ;
  assign n3369 = ~n3367 & ~n3368 ;
  assign n3370 = n2732 & n3369 ;
  assign n3371 = ~n3364 & ~n3370 ;
  assign n3372 = n523 & n3371 ;
  assign n3373 = ~n3355 & ~n3372 ;
  assign n3374 = ~n3340 & ~n3354 ;
  assign n3375 = \P1_reg3_reg[1]/NET0131  & n519 ;
  assign n3376 = \P1_reg2_reg[1]/NET0131  & n513 ;
  assign n3379 = ~n3375 & ~n3376 ;
  assign n3377 = \P1_reg1_reg[1]/NET0131  & n515 ;
  assign n3378 = \P1_reg0_reg[1]/NET0131  & n517 ;
  assign n3380 = ~n3377 & ~n3378 ;
  assign n3381 = n3379 & n3380 ;
  assign n3382 = \P1_IR_reg[0]/NET0131  & \P1_IR_reg[31]/NET0131  ;
  assign n3383 = ~\P1_IR_reg[1]/NET0131  & ~n3382 ;
  assign n3384 = \P1_IR_reg[1]/NET0131  & n3382 ;
  assign n3385 = ~n3383 & ~n3384 ;
  assign n3386 = n2732 & n3385 ;
  assign n3387 = ~\P2_datao_reg[1]/NET0131  & n639 ;
  assign n3388 = ~n2760 & ~n2761 ;
  assign n3390 = ~n2762 & n3388 ;
  assign n3389 = n2762 & ~n3388 ;
  assign n3391 = ~n639 & ~n3389 ;
  assign n3392 = ~n3390 & n3391 ;
  assign n3393 = ~n3387 & ~n3392 ;
  assign n3394 = ~n2732 & n3393 ;
  assign n3395 = ~n3386 & ~n3394 ;
  assign n3396 = ~n3381 & ~n3395 ;
  assign n3397 = n3381 & n3395 ;
  assign n3398 = \P1_reg1_reg[0]/NET0131  & n515 ;
  assign n3399 = \P1_reg0_reg[0]/NET0131  & n517 ;
  assign n3402 = ~n3398 & ~n3399 ;
  assign n3400 = \P1_reg2_reg[0]/NET0131  & n513 ;
  assign n3401 = \P1_reg3_reg[0]/NET0131  & n519 ;
  assign n3403 = ~n3400 & ~n3401 ;
  assign n3404 = n3402 & n3403 ;
  assign n3405 = \si[0]_pad  & ~n639 ;
  assign n3406 = ~\P2_datao_reg[0]/NET0131  & ~n3405 ;
  assign n3407 = ~n639 & n2762 ;
  assign n3408 = ~n3406 & ~n3407 ;
  assign n3409 = ~n2732 & n3408 ;
  assign n3410 = \P1_IR_reg[0]/NET0131  & n2732 ;
  assign n3411 = ~n3409 & ~n3410 ;
  assign n3412 = ~n3404 & ~n3411 ;
  assign n3413 = ~n3397 & n3412 ;
  assign n3414 = ~n3396 & ~n3413 ;
  assign n3415 = ~n3374 & n3414 ;
  assign n3416 = n3373 & ~n3415 ;
  assign n3417 = ~n3318 & ~n3332 ;
  assign n3418 = ~n523 & ~n3371 ;
  assign n3419 = ~n3417 & ~n3418 ;
  assign n3420 = ~n3416 & n3419 ;
  assign n3421 = ~n3333 & ~n3420 ;
  assign n3422 = \P1_IR_reg[31]/NET0131  & ~n468 ;
  assign n3423 = \P1_IR_reg[8]/NET0131  & n3422 ;
  assign n3424 = ~\P1_IR_reg[8]/NET0131  & ~n3422 ;
  assign n3425 = ~n3423 & ~n3424 ;
  assign n3426 = n2732 & ~n3425 ;
  assign n3427 = \P2_datao_reg[8]/NET0131  & n639 ;
  assign n3428 = ~n2787 & ~n2808 ;
  assign n3430 = n2783 & ~n3428 ;
  assign n3429 = ~n2783 & n3428 ;
  assign n3431 = ~n639 & ~n3429 ;
  assign n3432 = ~n3430 & n3431 ;
  assign n3433 = ~n3427 & ~n3432 ;
  assign n3434 = ~n2732 & n3433 ;
  assign n3435 = ~n3426 & ~n3434 ;
  assign n3436 = \P1_reg1_reg[8]/NET0131  & n515 ;
  assign n3437 = \P1_reg2_reg[8]/NET0131  & n513 ;
  assign n3442 = ~n3436 & ~n3437 ;
  assign n3438 = \P1_reg0_reg[8]/NET0131  & n517 ;
  assign n3439 = ~\P1_reg3_reg[8]/NET0131  & ~n3267 ;
  assign n3440 = ~n3268 & ~n3439 ;
  assign n3441 = n519 & n3440 ;
  assign n3443 = ~n3438 & ~n3441 ;
  assign n3444 = n3442 & n3443 ;
  assign n3445 = ~n3435 & n3444 ;
  assign n3446 = \P1_IR_reg[31]/NET0131  & ~n467 ;
  assign n3447 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[6]/NET0131  ;
  assign n3448 = ~n3446 & ~n3447 ;
  assign n3449 = \P1_IR_reg[7]/NET0131  & ~n3448 ;
  assign n3450 = ~\P1_IR_reg[7]/NET0131  & n3448 ;
  assign n3451 = ~n3449 & ~n3450 ;
  assign n3452 = n2732 & ~n3451 ;
  assign n3453 = \P2_datao_reg[7]/NET0131  & n639 ;
  assign n3454 = ~n2754 & ~n2780 ;
  assign n3456 = n3040 & ~n3454 ;
  assign n3455 = ~n3040 & n3454 ;
  assign n3457 = ~n639 & ~n3455 ;
  assign n3458 = ~n3456 & n3457 ;
  assign n3459 = ~n3453 & ~n3458 ;
  assign n3460 = ~n2732 & n3459 ;
  assign n3461 = ~n3452 & ~n3460 ;
  assign n3462 = ~\P1_reg3_reg[7]/NET0131  & ~n2874 ;
  assign n3463 = ~n3267 & ~n3462 ;
  assign n3464 = n519 & n3463 ;
  assign n3465 = \P1_reg0_reg[7]/NET0131  & n517 ;
  assign n3468 = ~n3464 & ~n3465 ;
  assign n3466 = \P1_reg1_reg[7]/NET0131  & n515 ;
  assign n3467 = \P1_reg2_reg[7]/NET0131  & n513 ;
  assign n3469 = ~n3466 & ~n3467 ;
  assign n3470 = n3468 & n3469 ;
  assign n3471 = ~n3461 & n3470 ;
  assign n3472 = ~n3445 & ~n3471 ;
  assign n3473 = \P2_datao_reg[6]/NET0131  & n639 ;
  assign n3474 = ~n2772 & ~n2779 ;
  assign n3476 = n2978 & ~n3474 ;
  assign n3475 = ~n2978 & n3474 ;
  assign n3477 = ~n639 & ~n3475 ;
  assign n3478 = ~n3476 & n3477 ;
  assign n3479 = ~n3473 & ~n3478 ;
  assign n3480 = ~n2732 & ~n3479 ;
  assign n3481 = ~\P1_IR_reg[6]/NET0131  & ~n3446 ;
  assign n3482 = ~n467 & n3447 ;
  assign n3483 = ~n3481 & ~n3482 ;
  assign n3484 = n2732 & n3483 ;
  assign n3485 = ~n3480 & ~n3484 ;
  assign n3486 = \P1_reg1_reg[6]/NET0131  & n515 ;
  assign n3487 = \P1_reg2_reg[6]/NET0131  & n513 ;
  assign n3492 = ~n3486 & ~n3487 ;
  assign n3488 = \P1_reg0_reg[6]/NET0131  & n517 ;
  assign n3489 = ~\P1_reg3_reg[6]/NET0131  & ~n2873 ;
  assign n3490 = ~n2874 & ~n3489 ;
  assign n3491 = n519 & n3490 ;
  assign n3493 = ~n3488 & ~n3491 ;
  assign n3494 = n3492 & n3493 ;
  assign n3495 = n3485 & n3494 ;
  assign n3496 = \P2_datao_reg[5]/NET0131  & n639 ;
  assign n3497 = ~n2756 & ~n2773 ;
  assign n3498 = ~n2755 & ~n2917 ;
  assign n3500 = n3497 & n3498 ;
  assign n3499 = ~n3497 & ~n3498 ;
  assign n3501 = ~n639 & ~n3499 ;
  assign n3502 = ~n3500 & n3501 ;
  assign n3503 = ~n3496 & ~n3502 ;
  assign n3504 = ~n2732 & ~n3503 ;
  assign n3505 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[4]/NET0131  ;
  assign n3506 = ~n3327 & ~n3505 ;
  assign n3507 = \P1_IR_reg[5]/NET0131  & ~n3506 ;
  assign n3508 = ~\P1_IR_reg[5]/NET0131  & n3506 ;
  assign n3509 = ~n3507 & ~n3508 ;
  assign n3510 = n2732 & n3509 ;
  assign n3511 = ~n3504 & ~n3510 ;
  assign n3512 = \P1_reg1_reg[5]/NET0131  & n515 ;
  assign n3513 = \P1_reg2_reg[5]/NET0131  & n513 ;
  assign n3518 = ~n3512 & ~n3513 ;
  assign n3514 = \P1_reg0_reg[5]/NET0131  & n517 ;
  assign n3515 = ~\P1_reg3_reg[5]/NET0131  & ~n2872 ;
  assign n3516 = ~n2873 & ~n3515 ;
  assign n3517 = n519 & n3516 ;
  assign n3519 = ~n3514 & ~n3517 ;
  assign n3520 = n3518 & n3519 ;
  assign n3521 = n3511 & n3520 ;
  assign n3522 = ~n3495 & ~n3521 ;
  assign n3523 = n3472 & n3522 ;
  assign n3524 = n3421 & n3523 ;
  assign n3525 = ~n3485 & ~n3494 ;
  assign n3526 = ~n3511 & ~n3520 ;
  assign n3527 = ~n3525 & ~n3526 ;
  assign n3528 = ~n3495 & ~n3527 ;
  assign n3529 = n3472 & n3528 ;
  assign n3530 = n3435 & ~n3444 ;
  assign n3531 = n3461 & ~n3470 ;
  assign n3532 = ~n3445 & n3531 ;
  assign n3533 = ~n3530 & ~n3532 ;
  assign n3534 = ~n3529 & n3533 ;
  assign n3535 = ~n3524 & n3534 ;
  assign n3536 = ~n3291 & n3300 ;
  assign n3537 = ~n3276 & ~n3536 ;
  assign n3538 = n3250 & n3537 ;
  assign n3539 = ~n3535 & n3538 ;
  assign n3540 = n3309 & ~n3539 ;
  assign n3541 = \P2_datao_reg[20]/NET0131  & n639 ;
  assign n3542 = ~n2825 & ~n2848 ;
  assign n3544 = n2824 & ~n3542 ;
  assign n3543 = ~n2824 & n3542 ;
  assign n3545 = ~n639 & ~n3543 ;
  assign n3546 = ~n3544 & n3545 ;
  assign n3547 = ~n3541 & ~n3546 ;
  assign n3548 = ~n2732 & ~n3547 ;
  assign n3552 = \P1_reg3_reg[15]/NET0131  & n2882 ;
  assign n3553 = n2883 & n3552 ;
  assign n3554 = \P1_reg3_reg[18]/NET0131  & n3553 ;
  assign n3555 = \P1_reg3_reg[19]/NET0131  & n3554 ;
  assign n3556 = ~\P1_reg3_reg[20]/NET0131  & ~n3555 ;
  assign n3557 = ~n2888 & ~n3556 ;
  assign n3558 = n519 & n3557 ;
  assign n3551 = \P1_reg1_reg[20]/NET0131  & n515 ;
  assign n3549 = \P1_reg2_reg[20]/NET0131  & n513 ;
  assign n3550 = \P1_reg0_reg[20]/NET0131  & n517 ;
  assign n3559 = ~n3549 & ~n3550 ;
  assign n3560 = ~n3551 & n3559 ;
  assign n3561 = ~n3558 & n3560 ;
  assign n3562 = ~n3548 & n3561 ;
  assign n3563 = \P1_IR_reg[31]/NET0131  & ~n2676 ;
  assign n3564 = ~\P1_IR_reg[19]/NET0131  & n3563 ;
  assign n3565 = \P1_IR_reg[19]/NET0131  & ~n3563 ;
  assign n3566 = ~n3564 & ~n3565 ;
  assign n3567 = n2732 & n3566 ;
  assign n3568 = \P2_datao_reg[19]/NET0131  & n639 ;
  assign n3569 = ~n2738 & ~n2747 ;
  assign n3570 = n3048 & ~n3110 ;
  assign n3571 = n3057 & ~n3570 ;
  assign n3573 = ~n3569 & n3571 ;
  assign n3572 = n3569 & ~n3571 ;
  assign n3574 = ~n639 & ~n3572 ;
  assign n3575 = ~n3573 & n3574 ;
  assign n3576 = ~n3568 & ~n3575 ;
  assign n3577 = ~n2732 & n3576 ;
  assign n3578 = ~n3567 & ~n3577 ;
  assign n3579 = ~\P1_reg3_reg[19]/NET0131  & ~n3554 ;
  assign n3580 = ~n3555 & ~n3579 ;
  assign n3581 = n519 & n3580 ;
  assign n3582 = \P1_reg1_reg[19]/NET0131  & n515 ;
  assign n3585 = ~n3581 & ~n3582 ;
  assign n3583 = \P1_reg0_reg[19]/NET0131  & n517 ;
  assign n3584 = \P1_reg2_reg[19]/NET0131  & n513 ;
  assign n3586 = ~n3583 & ~n3584 ;
  assign n3587 = n3585 & n3586 ;
  assign n3588 = ~n3578 & n3587 ;
  assign n3589 = ~n3562 & ~n3588 ;
  assign n3590 = \P1_IR_reg[31]/NET0131  & ~n477 ;
  assign n3591 = \P1_IR_reg[17]/NET0131  & ~n3590 ;
  assign n3592 = ~\P1_IR_reg[17]/NET0131  & n3590 ;
  assign n3593 = ~n3591 & ~n3592 ;
  assign n3594 = n2732 & n3593 ;
  assign n3595 = \P2_datao_reg[17]/NET0131  & n639 ;
  assign n3596 = ~n2740 & ~n2742 ;
  assign n3598 = n3160 & ~n3596 ;
  assign n3597 = ~n3160 & n3596 ;
  assign n3599 = ~n639 & ~n3597 ;
  assign n3600 = ~n3598 & n3599 ;
  assign n3601 = ~n3595 & ~n3600 ;
  assign n3602 = ~n2732 & n3601 ;
  assign n3603 = ~n3594 & ~n3602 ;
  assign n3604 = \P1_reg1_reg[17]/NET0131  & n515 ;
  assign n3605 = \P1_reg2_reg[17]/NET0131  & n513 ;
  assign n3611 = ~n3604 & ~n3605 ;
  assign n3606 = \P1_reg0_reg[17]/NET0131  & n517 ;
  assign n3607 = \P1_reg3_reg[16]/NET0131  & n3552 ;
  assign n3608 = ~\P1_reg3_reg[17]/NET0131  & ~n3607 ;
  assign n3609 = ~n3553 & ~n3608 ;
  assign n3610 = n519 & n3609 ;
  assign n3612 = ~n3606 & ~n3610 ;
  assign n3613 = n3611 & n3612 ;
  assign n3614 = ~n3603 & n3613 ;
  assign n3615 = \P1_IR_reg[31]/NET0131  & ~n498 ;
  assign n3616 = ~\P1_IR_reg[17]/NET0131  & n474 ;
  assign n3617 = \P1_IR_reg[31]/NET0131  & ~n3616 ;
  assign n3618 = ~n3615 & ~n3617 ;
  assign n3619 = \P1_IR_reg[18]/NET0131  & ~n3618 ;
  assign n3620 = ~\P1_IR_reg[18]/NET0131  & n3618 ;
  assign n3621 = ~n3619 & ~n3620 ;
  assign n3622 = n2732 & ~n3621 ;
  assign n3623 = \P2_datao_reg[18]/NET0131  & n639 ;
  assign n3624 = ~n2737 & ~n2746 ;
  assign n3626 = n2998 & ~n3624 ;
  assign n3625 = ~n2998 & n3624 ;
  assign n3627 = ~n639 & ~n3625 ;
  assign n3628 = ~n3626 & n3627 ;
  assign n3629 = ~n3623 & ~n3628 ;
  assign n3630 = ~n2732 & n3629 ;
  assign n3631 = ~n3622 & ~n3630 ;
  assign n3632 = ~\P1_reg3_reg[18]/NET0131  & ~n3553 ;
  assign n3633 = ~n3554 & ~n3632 ;
  assign n3634 = n519 & n3633 ;
  assign n3635 = \P1_reg0_reg[18]/NET0131  & n517 ;
  assign n3638 = ~n3634 & ~n3635 ;
  assign n3636 = \P1_reg1_reg[18]/NET0131  & n515 ;
  assign n3637 = \P1_reg2_reg[18]/NET0131  & n513 ;
  assign n3639 = ~n3636 & ~n3637 ;
  assign n3640 = n3638 & n3639 ;
  assign n3641 = ~n3631 & n3640 ;
  assign n3642 = ~n3614 & ~n3641 ;
  assign n3643 = n3589 & n3642 ;
  assign n3644 = \P1_IR_reg[14]/NET0131  & n3615 ;
  assign n3645 = ~\P1_IR_reg[14]/NET0131  & ~n3615 ;
  assign n3646 = ~n3644 & ~n3645 ;
  assign n3647 = n2732 & ~n3646 ;
  assign n3648 = \P2_datao_reg[14]/NET0131  & n639 ;
  assign n3649 = ~n2793 & ~n2816 ;
  assign n3651 = n3133 & ~n3649 ;
  assign n3650 = ~n3133 & n3649 ;
  assign n3652 = ~n639 & ~n3650 ;
  assign n3653 = ~n3651 & n3652 ;
  assign n3654 = ~n3648 & ~n3653 ;
  assign n3655 = ~n2732 & n3654 ;
  assign n3656 = ~n3647 & ~n3655 ;
  assign n3657 = \P1_reg2_reg[14]/NET0131  & n513 ;
  assign n3658 = ~\P1_reg3_reg[14]/NET0131  & ~n2881 ;
  assign n3659 = ~n2882 & ~n3658 ;
  assign n3660 = n519 & n3659 ;
  assign n3663 = ~n3657 & ~n3660 ;
  assign n3661 = \P1_reg1_reg[14]/NET0131  & n515 ;
  assign n3662 = \P1_reg0_reg[14]/NET0131  & n517 ;
  assign n3664 = ~n3661 & ~n3662 ;
  assign n3665 = n3663 & n3664 ;
  assign n3666 = ~n3656 & n3665 ;
  assign n3667 = ~\P1_IR_reg[12]/NET0131  & ~\P1_IR_reg[9]/NET0131  ;
  assign n3668 = n469 & n3667 ;
  assign n3669 = \P1_IR_reg[31]/NET0131  & ~n3668 ;
  assign n3670 = ~n3224 & ~n3669 ;
  assign n3671 = \P1_IR_reg[13]/NET0131  & ~n3670 ;
  assign n3672 = ~\P1_IR_reg[13]/NET0131  & n3670 ;
  assign n3673 = ~n3671 & ~n3672 ;
  assign n3674 = n2732 & ~n3673 ;
  assign n3675 = \P2_datao_reg[13]/NET0131  & n639 ;
  assign n3676 = ~n2796 & ~n2801 ;
  assign n3678 = n3158 & ~n3676 ;
  assign n3677 = ~n3158 & n3676 ;
  assign n3679 = ~n639 & ~n3677 ;
  assign n3680 = ~n3678 & n3679 ;
  assign n3681 = ~n3675 & ~n3680 ;
  assign n3682 = ~n2732 & n3681 ;
  assign n3683 = ~n3674 & ~n3682 ;
  assign n3684 = \P1_reg0_reg[13]/NET0131  & n517 ;
  assign n3685 = ~\P1_reg3_reg[13]/NET0131  & ~n2880 ;
  assign n3686 = ~n2881 & ~n3685 ;
  assign n3687 = n519 & n3686 ;
  assign n3690 = ~n3684 & ~n3687 ;
  assign n3688 = \P1_reg1_reg[13]/NET0131  & n515 ;
  assign n3689 = \P1_reg2_reg[13]/NET0131  & n513 ;
  assign n3691 = ~n3688 & ~n3689 ;
  assign n3692 = n3690 & n3691 ;
  assign n3693 = ~n3683 & n3692 ;
  assign n3694 = ~n3666 & ~n3693 ;
  assign n3695 = \P1_IR_reg[31]/NET0131  & ~n2690 ;
  assign n3696 = \P1_IR_reg[16]/NET0131  & n3695 ;
  assign n3697 = ~\P1_IR_reg[16]/NET0131  & ~n3695 ;
  assign n3698 = ~n3696 & ~n3697 ;
  assign n3699 = n2732 & ~n3698 ;
  assign n3700 = \P2_datao_reg[16]/NET0131  & n639 ;
  assign n3701 = ~n2741 & ~n2751 ;
  assign n3703 = n2822 & ~n3701 ;
  assign n3702 = ~n2822 & n3701 ;
  assign n3704 = ~n639 & ~n3702 ;
  assign n3705 = ~n3703 & n3704 ;
  assign n3706 = ~n3700 & ~n3705 ;
  assign n3707 = ~n2732 & n3706 ;
  assign n3708 = ~n3699 & ~n3707 ;
  assign n3709 = \P1_reg2_reg[16]/NET0131  & n513 ;
  assign n3710 = \P1_reg1_reg[16]/NET0131  & n515 ;
  assign n3715 = ~n3709 & ~n3710 ;
  assign n3711 = \P1_reg0_reg[16]/NET0131  & n517 ;
  assign n3712 = ~\P1_reg3_reg[16]/NET0131  & ~n3552 ;
  assign n3713 = ~n3607 & ~n3712 ;
  assign n3714 = n519 & n3713 ;
  assign n3716 = ~n3711 & ~n3714 ;
  assign n3717 = n3715 & n3716 ;
  assign n3718 = ~n3708 & n3717 ;
  assign n3719 = \P1_IR_reg[31]/NET0131  & ~n2674 ;
  assign n3720 = \P1_IR_reg[15]/NET0131  & n3719 ;
  assign n3721 = ~\P1_IR_reg[15]/NET0131  & ~n3719 ;
  assign n3722 = ~n3720 & ~n3721 ;
  assign n3723 = n2732 & ~n3722 ;
  assign n3724 = \P2_datao_reg[15]/NET0131  & n639 ;
  assign n3725 = ~n2792 & ~n2817 ;
  assign n3727 = n3110 & ~n3725 ;
  assign n3726 = ~n3110 & n3725 ;
  assign n3728 = ~n639 & ~n3726 ;
  assign n3729 = ~n3727 & n3728 ;
  assign n3730 = ~n3724 & ~n3729 ;
  assign n3731 = ~n2732 & n3730 ;
  assign n3732 = ~n3723 & ~n3731 ;
  assign n3733 = \P1_reg2_reg[15]/NET0131  & n513 ;
  assign n3734 = ~\P1_reg3_reg[15]/NET0131  & ~n2882 ;
  assign n3735 = ~n3552 & ~n3734 ;
  assign n3736 = n519 & n3735 ;
  assign n3739 = ~n3733 & ~n3736 ;
  assign n3737 = \P1_reg0_reg[15]/NET0131  & n517 ;
  assign n3738 = \P1_reg1_reg[15]/NET0131  & n515 ;
  assign n3740 = ~n3737 & ~n3738 ;
  assign n3741 = n3739 & n3740 ;
  assign n3742 = ~n3732 & n3741 ;
  assign n3743 = ~n3718 & ~n3742 ;
  assign n3744 = n3694 & n3743 ;
  assign n3745 = n3643 & n3744 ;
  assign n3746 = ~n3540 & n3745 ;
  assign n3747 = n3656 & ~n3665 ;
  assign n3748 = n3683 & ~n3692 ;
  assign n3749 = ~n3747 & ~n3748 ;
  assign n3750 = ~n3666 & ~n3749 ;
  assign n3751 = n3743 & n3750 ;
  assign n3752 = n3708 & ~n3717 ;
  assign n3753 = n3732 & ~n3741 ;
  assign n3754 = ~n3752 & ~n3753 ;
  assign n3755 = ~n3718 & ~n3754 ;
  assign n3756 = ~n3751 & ~n3755 ;
  assign n3757 = n3643 & ~n3756 ;
  assign n3758 = n3631 & ~n3640 ;
  assign n3759 = n3603 & ~n3613 ;
  assign n3760 = ~n3758 & ~n3759 ;
  assign n3761 = ~n3641 & ~n3760 ;
  assign n3762 = n3589 & n3761 ;
  assign n3763 = n3548 & ~n3561 ;
  assign n3764 = n3578 & ~n3587 ;
  assign n3765 = ~n3562 & n3764 ;
  assign n3766 = ~n3763 & ~n3765 ;
  assign n3767 = ~n3762 & n3766 ;
  assign n3768 = ~n3757 & n3767 ;
  assign n3769 = ~n3746 & n3768 ;
  assign n3770 = ~n3168 & n3177 ;
  assign n3771 = ~n3155 & ~n3770 ;
  assign n3772 = n3130 & n3771 ;
  assign n3773 = ~n2905 & n3772 ;
  assign n3774 = n3081 & n3773 ;
  assign n3775 = ~n3769 & n3774 ;
  assign n3776 = ~n3197 & ~n3775 ;
  assign n3777 = \P2_datao_reg[29]/NET0131  & n639 ;
  assign n3778 = \P2_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n3779 = ~\P2_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n3780 = ~n3778 & ~n3779 ;
  assign n3782 = n2838 & ~n3162 ;
  assign n3781 = ~n2735 & ~n2842 ;
  assign n3783 = n2835 & ~n2956 ;
  assign n3784 = ~n3031 & ~n3783 ;
  assign n3785 = ~n2836 & ~n3784 ;
  assign n3786 = n3781 & ~n3785 ;
  assign n3787 = ~n3782 & n3786 ;
  assign n3788 = ~n2734 & ~n3787 ;
  assign n3790 = n3780 & n3788 ;
  assign n3789 = ~n3780 & ~n3788 ;
  assign n3791 = ~n639 & ~n3789 ;
  assign n3792 = ~n3790 & n3791 ;
  assign n3793 = ~n3777 & ~n3792 ;
  assign n3794 = ~n2732 & ~n3793 ;
  assign n3795 = n519 & n2899 ;
  assign n3796 = \P1_reg1_reg[29]/NET0131  & n515 ;
  assign n3799 = ~n3795 & ~n3796 ;
  assign n3797 = \P1_reg2_reg[29]/NET0131  & n513 ;
  assign n3798 = \P1_reg0_reg[29]/NET0131  & n517 ;
  assign n3800 = ~n3797 & ~n3798 ;
  assign n3801 = n3799 & n3800 ;
  assign n3802 = n3794 & n3801 ;
  assign n3803 = ~n3794 & ~n3801 ;
  assign n3804 = ~n3802 & ~n3803 ;
  assign n3805 = n3776 & ~n3804 ;
  assign n3806 = ~n3776 & n3804 ;
  assign n3807 = ~n3805 & ~n3806 ;
  assign n3808 = n2717 & ~n3807 ;
  assign n3809 = ~n2718 & ~n3808 ;
  assign n3810 = \P1_IR_reg[31]/NET0131  & ~n501 ;
  assign n3811 = ~\P1_IR_reg[22]/NET0131  & ~n3810 ;
  assign n3812 = \P1_IR_reg[22]/NET0131  & n3810 ;
  assign n3813 = ~n3811 & ~n3812 ;
  assign n3814 = n2683 & n3813 ;
  assign n3815 = ~n2683 & ~n3813 ;
  assign n3816 = ~n3814 & ~n3815 ;
  assign n3817 = \P1_IR_reg[31]/NET0131  & ~n482 ;
  assign n3818 = ~n3590 & ~n3817 ;
  assign n3819 = \P1_IR_reg[21]/NET0131  & ~n3818 ;
  assign n3820 = ~\P1_IR_reg[21]/NET0131  & n3818 ;
  assign n3821 = ~n3819 & ~n3820 ;
  assign n3822 = n3813 & n3821 ;
  assign n3823 = \P1_IR_reg[31]/NET0131  & ~n2692 ;
  assign n3824 = ~\P1_IR_reg[20]/NET0131  & n3823 ;
  assign n3825 = \P1_IR_reg[20]/NET0131  & ~n3823 ;
  assign n3826 = ~n3824 & ~n3825 ;
  assign n3827 = n2683 & ~n3826 ;
  assign n3828 = ~n3822 & ~n3827 ;
  assign n3829 = n3816 & n3828 ;
  assign n3830 = ~n3809 & n3829 ;
  assign n3831 = n3211 & n3221 ;
  assign n3832 = n3239 & n3248 ;
  assign n3833 = ~n3831 & ~n3832 ;
  assign n3834 = n3263 & n3275 ;
  assign n3835 = ~n3291 & ~n3300 ;
  assign n3836 = ~n3263 & ~n3275 ;
  assign n3837 = ~n3835 & ~n3836 ;
  assign n3838 = ~n3834 & ~n3837 ;
  assign n3839 = n3833 & n3838 ;
  assign n3840 = ~n3239 & ~n3248 ;
  assign n3841 = ~n3211 & ~n3221 ;
  assign n3842 = ~n3832 & n3841 ;
  assign n3843 = ~n3840 & ~n3842 ;
  assign n3844 = ~n3839 & n3843 ;
  assign n3845 = ~n3318 & n3332 ;
  assign n3846 = ~n523 & n3371 ;
  assign n3847 = ~n3845 & ~n3846 ;
  assign n3848 = n3404 & ~n3411 ;
  assign n3849 = n3381 & ~n3395 ;
  assign n3850 = ~n3848 & ~n3849 ;
  assign n3851 = ~n3381 & n3395 ;
  assign n3852 = ~n3340 & n3354 ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3854 = ~n3850 & n3853 ;
  assign n3855 = n3340 & ~n3354 ;
  assign n3856 = n523 & ~n3371 ;
  assign n3857 = ~n3855 & ~n3856 ;
  assign n3858 = ~n3854 & n3857 ;
  assign n3859 = n3847 & ~n3858 ;
  assign n3860 = ~n3485 & n3494 ;
  assign n3861 = n3318 & ~n3332 ;
  assign n3862 = ~n3511 & n3520 ;
  assign n3863 = ~n3861 & ~n3862 ;
  assign n3864 = ~n3860 & n3863 ;
  assign n3865 = ~n3859 & n3864 ;
  assign n3866 = n3485 & ~n3494 ;
  assign n3867 = n3511 & ~n3520 ;
  assign n3868 = ~n3866 & ~n3867 ;
  assign n3869 = ~n3860 & ~n3868 ;
  assign n3870 = ~n3865 & ~n3869 ;
  assign n3871 = n3435 & n3444 ;
  assign n3872 = n3461 & n3470 ;
  assign n3873 = ~n3871 & ~n3872 ;
  assign n3874 = ~n3870 & n3873 ;
  assign n3875 = ~n3435 & ~n3444 ;
  assign n3876 = ~n3461 & ~n3470 ;
  assign n3877 = ~n3875 & ~n3876 ;
  assign n3878 = ~n3871 & ~n3877 ;
  assign n3879 = ~n3874 & ~n3878 ;
  assign n3880 = n3291 & n3300 ;
  assign n3881 = ~n3834 & ~n3880 ;
  assign n3882 = n3833 & n3881 ;
  assign n3883 = ~n3879 & n3882 ;
  assign n3884 = n3844 & ~n3883 ;
  assign n3885 = n3708 & n3717 ;
  assign n3886 = n3732 & n3741 ;
  assign n3887 = ~n3885 & ~n3886 ;
  assign n3888 = n3656 & n3665 ;
  assign n3889 = ~n3683 & ~n3692 ;
  assign n3890 = ~n3656 & ~n3665 ;
  assign n3891 = ~n3889 & ~n3890 ;
  assign n3892 = ~n3888 & ~n3891 ;
  assign n3893 = n3887 & n3892 ;
  assign n3894 = ~n3708 & ~n3717 ;
  assign n3895 = ~n3732 & ~n3741 ;
  assign n3896 = ~n3894 & ~n3895 ;
  assign n3897 = ~n3885 & ~n3896 ;
  assign n3898 = ~n3893 & ~n3897 ;
  assign n3899 = n3548 & n3561 ;
  assign n3900 = n3578 & n3587 ;
  assign n3901 = ~n3899 & ~n3900 ;
  assign n3902 = n3631 & n3640 ;
  assign n3903 = ~n3631 & ~n3640 ;
  assign n3904 = ~n3603 & ~n3613 ;
  assign n3905 = ~n3903 & ~n3904 ;
  assign n3906 = ~n3902 & ~n3905 ;
  assign n3907 = n3901 & n3906 ;
  assign n3908 = ~n3548 & ~n3561 ;
  assign n3909 = ~n3578 & ~n3587 ;
  assign n3910 = ~n3908 & ~n3909 ;
  assign n3911 = ~n3899 & ~n3910 ;
  assign n3912 = ~n3907 & ~n3911 ;
  assign n3913 = n3898 & n3912 ;
  assign n3914 = n3884 & n3913 ;
  assign n3915 = n3603 & n3613 ;
  assign n3916 = ~n3902 & ~n3915 ;
  assign n3917 = n3901 & n3916 ;
  assign n3918 = n3683 & n3692 ;
  assign n3919 = ~n3888 & ~n3918 ;
  assign n3920 = n3887 & n3919 ;
  assign n3921 = n3898 & ~n3920 ;
  assign n3922 = n3917 & ~n3921 ;
  assign n3923 = n3912 & ~n3922 ;
  assign n3924 = n3069 & n3078 ;
  assign n3925 = n2868 & n2904 ;
  assign n3926 = ~n3924 & ~n3925 ;
  assign n3927 = n2964 & n2974 ;
  assign n3928 = n3017 & n3026 ;
  assign n3929 = ~n3927 & ~n3928 ;
  assign n3930 = n3926 & n3929 ;
  assign n3931 = n3168 & n3177 ;
  assign n3932 = n3143 & n3153 ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = n3119 & n3128 ;
  assign n3935 = n3096 & n3105 ;
  assign n3936 = ~n3934 & ~n3935 ;
  assign n3937 = n3933 & n3936 ;
  assign n3938 = n3930 & n3937 ;
  assign n3939 = ~n3923 & n3938 ;
  assign n3940 = ~n3914 & n3939 ;
  assign n3941 = ~n3143 & ~n3153 ;
  assign n3942 = ~n3168 & ~n3177 ;
  assign n3943 = ~n3941 & ~n3942 ;
  assign n3944 = ~n3932 & ~n3943 ;
  assign n3945 = n3936 & n3944 ;
  assign n3946 = ~n3096 & ~n3105 ;
  assign n3947 = ~n3119 & ~n3128 ;
  assign n3948 = ~n3935 & n3947 ;
  assign n3949 = ~n3946 & ~n3948 ;
  assign n3950 = ~n3945 & n3949 ;
  assign n3951 = n3930 & ~n3950 ;
  assign n3952 = ~n3017 & ~n3026 ;
  assign n3953 = ~n2964 & ~n2974 ;
  assign n3954 = ~n3952 & ~n3953 ;
  assign n3955 = ~n3928 & ~n3954 ;
  assign n3956 = n3926 & n3955 ;
  assign n3957 = ~n2868 & ~n2904 ;
  assign n3958 = ~n3069 & ~n3078 ;
  assign n3959 = ~n3925 & n3958 ;
  assign n3960 = ~n3957 & ~n3959 ;
  assign n3961 = ~n3956 & n3960 ;
  assign n3962 = ~n3951 & n3961 ;
  assign n3963 = ~n3940 & n3962 ;
  assign n3964 = ~n3804 & n3963 ;
  assign n3965 = n3804 & ~n3963 ;
  assign n3966 = ~n3964 & ~n3965 ;
  assign n3967 = n2717 & n3966 ;
  assign n3968 = ~n2718 & ~n3967 ;
  assign n3969 = ~n3814 & ~n3828 ;
  assign n3970 = ~n3968 & n3969 ;
  assign n3971 = n2731 & ~n2904 ;
  assign n3974 = ~n3587 & ~n3640 ;
  assign n3975 = ~n3561 & n3974 ;
  assign n3976 = ~n3177 & ~n3613 ;
  assign n3977 = ~n3717 & n3976 ;
  assign n3978 = n3975 & n3977 ;
  assign n3979 = \P1_reg2_reg[31]/NET0131  & n513 ;
  assign n3982 = ~n3795 & ~n3979 ;
  assign n3980 = \P1_reg1_reg[31]/NET0131  & n515 ;
  assign n3981 = \P1_reg0_reg[31]/NET0131  & n517 ;
  assign n3983 = ~n3980 & ~n3981 ;
  assign n3984 = n3982 & n3983 ;
  assign n3985 = ~n3404 & ~n3984 ;
  assign n3986 = ~n3381 & n3985 ;
  assign n3987 = ~n3340 & n3986 ;
  assign n3988 = ~n523 & n3987 ;
  assign n3989 = ~n3318 & n3988 ;
  assign n3990 = ~n3520 & n3989 ;
  assign n3991 = ~n3300 & ~n3444 ;
  assign n3992 = ~n3470 & ~n3494 ;
  assign n3993 = n3991 & n3992 ;
  assign n3994 = n3990 & n3993 ;
  assign n3995 = ~n3221 & ~n3275 ;
  assign n3996 = ~n3248 & n3995 ;
  assign n3997 = ~n3665 & ~n3692 ;
  assign n3998 = ~n3741 & n3997 ;
  assign n3999 = n3996 & n3998 ;
  assign n4000 = n3994 & n3999 ;
  assign n4001 = n3978 & n4000 ;
  assign n4002 = ~n3105 & ~n3128 ;
  assign n4003 = ~n2974 & n4002 ;
  assign n4004 = ~n3026 & n4003 ;
  assign n4005 = ~n3078 & ~n3153 ;
  assign n4006 = n4004 & n4005 ;
  assign n4007 = ~n2904 & n4006 ;
  assign n4008 = n4001 & n4007 ;
  assign n4009 = ~n3801 & n4008 ;
  assign n4010 = \P1_reg2_reg[30]/NET0131  & n513 ;
  assign n4013 = ~n3795 & ~n4010 ;
  assign n4011 = \P1_reg1_reg[30]/NET0131  & n515 ;
  assign n4012 = \P1_reg0_reg[30]/NET0131  & n517 ;
  assign n4014 = ~n4011 & ~n4012 ;
  assign n4015 = n4013 & n4014 ;
  assign n4017 = n4009 & ~n4015 ;
  assign n3972 = ~\P1_B_reg/NET0131  & ~n2731 ;
  assign n3973 = ~n2732 & ~n3972 ;
  assign n4016 = ~n4009 & n4015 ;
  assign n4018 = ~n3973 & ~n4016 ;
  assign n4019 = ~n4017 & n4018 ;
  assign n4020 = ~n3971 & ~n4019 ;
  assign n4021 = n2717 & ~n4020 ;
  assign n4022 = ~n2718 & ~n4021 ;
  assign n4023 = n2683 & n3826 ;
  assign n4024 = ~n3821 & n4023 ;
  assign n4025 = n3813 & n4024 ;
  assign n4026 = ~n4022 & n4025 ;
  assign n4027 = ~n3813 & n3821 ;
  assign n4028 = ~n2683 & n4027 ;
  assign n4029 = n3794 & n4028 ;
  assign n4030 = n3395 & n3411 ;
  assign n4031 = n3354 & n4030 ;
  assign n4032 = n3371 & n4031 ;
  assign n4033 = n3332 & n4032 ;
  assign n4034 = n3485 & n3511 ;
  assign n4035 = n4033 & n4034 ;
  assign n4036 = ~n3461 & n4035 ;
  assign n4037 = ~n3211 & ~n3239 ;
  assign n4038 = ~n3263 & ~n3291 ;
  assign n4039 = ~n3435 & n4038 ;
  assign n4040 = ~n3683 & n4039 ;
  assign n4041 = n4037 & n4040 ;
  assign n4042 = n4036 & n4041 ;
  assign n4043 = ~n3603 & ~n3656 ;
  assign n4044 = ~n3708 & ~n3732 ;
  assign n4045 = n4043 & n4044 ;
  assign n4046 = n4042 & n4045 ;
  assign n4047 = ~n3548 & ~n3631 ;
  assign n4048 = ~n3578 & n4047 ;
  assign n4049 = n4046 & n4048 ;
  assign n4050 = ~n3143 & ~n3168 ;
  assign n4051 = n4049 & n4050 ;
  assign n4052 = ~n2964 & ~n3119 ;
  assign n4053 = ~n3096 & n4052 ;
  assign n4054 = n4051 & n4053 ;
  assign n4055 = ~n2868 & ~n3069 ;
  assign n4056 = ~n3017 & n4055 ;
  assign n4057 = n4054 & n4056 ;
  assign n4058 = n3794 & ~n4057 ;
  assign n4059 = ~n3794 & n4057 ;
  assign n4060 = ~n4058 & ~n4059 ;
  assign n4061 = n3815 & ~n3821 ;
  assign n4062 = n3826 & n4061 ;
  assign n4063 = n4060 & n4062 ;
  assign n4064 = ~n4029 & ~n4063 ;
  assign n4065 = n2717 & ~n4064 ;
  assign n4066 = ~n3821 & n3826 ;
  assign n4067 = n3814 & ~n4066 ;
  assign n4068 = ~n3821 & ~n3826 ;
  assign n4069 = n3815 & ~n4068 ;
  assign n4070 = ~n2717 & n4069 ;
  assign n4071 = ~n4067 & ~n4070 ;
  assign n4072 = \P1_reg2_reg[29]/NET0131  & ~n4071 ;
  assign n4073 = ~n3826 & n4061 ;
  assign n4074 = n2899 & n4073 ;
  assign n4075 = ~n4072 & ~n4074 ;
  assign n4076 = ~n4065 & n4075 ;
  assign n4077 = ~n4026 & n4076 ;
  assign n4078 = ~n3970 & n4077 ;
  assign n4079 = ~n3830 & n4078 ;
  assign n4080 = n2701 & ~n4079 ;
  assign n4081 = ~n2683 & n2700 ;
  assign n4082 = \P1_reg2_reg[29]/NET0131  & n4081 ;
  assign n4083 = ~n4080 & ~n4082 ;
  assign n4084 = \P1_state_reg[0]/NET0131  & ~n4083 ;
  assign n4085 = \P1_state_reg[0]/NET0131  & ~n2683 ;
  assign n4086 = \P1_reg2_reg[29]/NET0131  & ~n4085 ;
  assign n4087 = ~n4084 & ~n4086 ;
  assign n4088 = \P2_reg1_reg[29]/NET0131  & ~n2286 ;
  assign n4089 = \P2_reg1_reg[29]/NET0131  & n2035 ;
  assign n4090 = \P2_reg1_reg[29]/NET0131  & ~n2310 ;
  assign n4091 = n2310 & n2596 ;
  assign n4092 = ~n4090 & ~n4091 ;
  assign n4093 = ~n2290 & ~n4092 ;
  assign n4094 = \P2_reg1_reg[29]/NET0131  & ~n2291 ;
  assign n4095 = n2291 & ~n2608 ;
  assign n4096 = ~n4094 & ~n4095 ;
  assign n4097 = n1790 & ~n4096 ;
  assign n4098 = n2272 & ~n2310 ;
  assign n4099 = n2612 & ~n4098 ;
  assign n4100 = \P2_reg1_reg[29]/NET0131  & ~n4099 ;
  assign n4101 = n2272 & n2310 ;
  assign n4102 = n1656 & n4101 ;
  assign n4109 = ~n4100 & ~n4102 ;
  assign n4110 = ~n4097 & n4109 ;
  assign n4111 = ~n4093 & n4110 ;
  assign n4103 = n2310 & ~n2654 ;
  assign n4104 = ~n4090 & ~n4103 ;
  assign n4105 = ~n2392 & ~n4104 ;
  assign n4106 = n2291 & n2596 ;
  assign n4107 = ~n4094 & ~n4106 ;
  assign n4108 = n2314 & ~n4107 ;
  assign n4112 = ~n4105 & ~n4108 ;
  assign n4113 = n4111 & n4112 ;
  assign n4114 = n2037 & ~n4113 ;
  assign n4115 = ~n4089 & ~n4114 ;
  assign n4116 = \P1_state_reg[0]/NET0131  & ~n4115 ;
  assign n4117 = ~n4088 & ~n4116 ;
  assign n4118 = \P2_reg2_reg[25]/NET0131  & ~n2286 ;
  assign n4119 = \P2_reg2_reg[25]/NET0131  & n2035 ;
  assign n4120 = \P2_reg2_reg[25]/NET0131  & ~n2291 ;
  assign n4124 = n2562 & n2570 ;
  assign n4121 = n2561 & ~n2564 ;
  assign n4122 = n2574 & ~n4121 ;
  assign n4123 = n2560 & ~n4122 ;
  assign n4125 = n2577 & ~n4123 ;
  assign n4126 = ~n4124 & n4125 ;
  assign n4127 = n2580 & ~n4126 ;
  assign n4128 = n2587 & ~n4127 ;
  assign n4129 = n1938 & ~n4128 ;
  assign n4130 = ~n1938 & n4128 ;
  assign n4131 = ~n4129 & ~n4130 ;
  assign n4132 = n2291 & ~n4131 ;
  assign n4133 = ~n4120 & ~n4132 ;
  assign n4134 = ~n2290 & ~n4133 ;
  assign n4149 = \P2_reg2_reg[25]/NET0131  & ~n2310 ;
  assign n4155 = ~n1587 & n2499 ;
  assign n4154 = n1587 & ~n2499 ;
  assign n4156 = n2263 & ~n4154 ;
  assign n4157 = ~n4155 & n4156 ;
  assign n4158 = ~n1549 & ~n2263 ;
  assign n4159 = ~n4157 & ~n4158 ;
  assign n4160 = n2310 & ~n4159 ;
  assign n4161 = ~n4149 & ~n4160 ;
  assign n4162 = n1790 & ~n4161 ;
  assign n4153 = n1513 & n2394 ;
  assign n4163 = \P2_reg2_reg[25]/NET0131  & ~n2407 ;
  assign n4164 = ~n1521 & n1854 ;
  assign n4165 = ~n4163 & ~n4164 ;
  assign n4166 = ~n4153 & n4165 ;
  assign n4167 = ~n4162 & n4166 ;
  assign n4168 = ~n4134 & n4167 ;
  assign n4136 = n2619 & ~n2622 ;
  assign n4137 = n2632 & ~n4136 ;
  assign n4138 = n2618 & ~n4137 ;
  assign n4135 = n2620 & n2628 ;
  assign n4139 = n2635 & ~n4135 ;
  assign n4140 = ~n4138 & n4139 ;
  assign n4141 = n2638 & ~n4140 ;
  assign n4142 = n2647 & ~n4141 ;
  assign n4143 = n1938 & n4142 ;
  assign n4144 = ~n1938 & ~n4142 ;
  assign n4145 = ~n4143 & ~n4144 ;
  assign n4146 = n2291 & ~n4145 ;
  assign n4147 = ~n4120 & ~n4146 ;
  assign n4148 = ~n2392 & ~n4147 ;
  assign n4150 = n2310 & ~n4131 ;
  assign n4151 = ~n4149 & ~n4150 ;
  assign n4152 = n2314 & ~n4151 ;
  assign n4169 = ~n4148 & ~n4152 ;
  assign n4170 = n4168 & n4169 ;
  assign n4171 = n2037 & ~n4170 ;
  assign n4172 = ~n4119 & ~n4171 ;
  assign n4173 = \P1_state_reg[0]/NET0131  & ~n4172 ;
  assign n4174 = ~n4118 & ~n4173 ;
  assign n4175 = \P2_reg2_reg[29]/NET0131  & ~n2286 ;
  assign n4176 = \P2_reg2_reg[29]/NET0131  & n2035 ;
  assign n4177 = \P2_reg2_reg[29]/NET0131  & ~n2291 ;
  assign n4178 = ~n4106 & ~n4177 ;
  assign n4179 = ~n2290 & ~n4178 ;
  assign n4183 = \P2_reg2_reg[29]/NET0131  & ~n2310 ;
  assign n4186 = n2310 & ~n2608 ;
  assign n4187 = ~n4183 & ~n4186 ;
  assign n4188 = n1790 & ~n4187 ;
  assign n4189 = n1656 & n2394 ;
  assign n4190 = \P2_reg2_reg[29]/NET0131  & ~n2407 ;
  assign n4191 = n1661 & n1854 ;
  assign n4192 = ~n4190 & ~n4191 ;
  assign n4193 = ~n4189 & n4192 ;
  assign n4194 = ~n4188 & n4193 ;
  assign n4195 = ~n4179 & n4194 ;
  assign n4180 = n2291 & ~n2654 ;
  assign n4181 = ~n4177 & ~n4180 ;
  assign n4182 = ~n2392 & ~n4181 ;
  assign n4184 = ~n4091 & ~n4183 ;
  assign n4185 = n2314 & ~n4184 ;
  assign n4196 = ~n4182 & ~n4185 ;
  assign n4197 = n4195 & n4196 ;
  assign n4198 = n2037 & ~n4197 ;
  assign n4199 = ~n4176 & ~n4198 ;
  assign n4200 = \P1_state_reg[0]/NET0131  & ~n4199 ;
  assign n4201 = ~n4175 & ~n4200 ;
  assign n4202 = ~n2711 & n2716 ;
  assign n4203 = \P1_reg1_reg[29]/NET0131  & ~n4202 ;
  assign n4204 = ~n3807 & n4202 ;
  assign n4205 = ~n4203 & ~n4204 ;
  assign n4206 = n3829 & ~n4205 ;
  assign n4207 = n3966 & n4202 ;
  assign n4208 = ~n4203 & ~n4207 ;
  assign n4209 = n3969 & ~n4208 ;
  assign n4210 = ~n4020 & n4202 ;
  assign n4211 = ~n4203 & ~n4210 ;
  assign n4212 = n4025 & ~n4211 ;
  assign n4213 = ~n4064 & n4202 ;
  assign n4214 = ~n4067 & ~n4073 ;
  assign n4215 = n4028 & ~n4202 ;
  assign n4216 = n4214 & ~n4215 ;
  assign n4217 = n4062 & ~n4202 ;
  assign n4218 = n4216 & ~n4217 ;
  assign n4219 = \P1_reg1_reg[29]/NET0131  & ~n4218 ;
  assign n4220 = ~n4213 & ~n4219 ;
  assign n4221 = ~n4212 & n4220 ;
  assign n4222 = ~n4209 & n4221 ;
  assign n4223 = ~n4206 & n4222 ;
  assign n4224 = n2701 & ~n4223 ;
  assign n4225 = \P1_reg1_reg[29]/NET0131  & n4081 ;
  assign n4226 = ~n4224 & ~n4225 ;
  assign n4227 = \P1_state_reg[0]/NET0131  & ~n4226 ;
  assign n4228 = \P1_reg1_reg[29]/NET0131  & ~n4085 ;
  assign n4229 = ~n4227 & ~n4228 ;
  assign n4232 = ~n1304 & n2035 ;
  assign n4235 = ~n1304 & ~n2053 ;
  assign n4236 = n2316 & n2330 ;
  assign n4237 = ~n2325 & n4236 ;
  assign n4238 = ~n2328 & n2330 ;
  assign n4239 = ~n2335 & ~n4238 ;
  assign n4240 = ~n4237 & n4239 ;
  assign n4241 = n2331 & n2342 ;
  assign n4242 = ~n4240 & n4241 ;
  assign n4243 = ~n2338 & n2342 ;
  assign n4244 = ~n2350 & ~n4243 ;
  assign n4245 = ~n4242 & n4244 ;
  assign n4246 = n2341 & n2345 ;
  assign n4247 = ~n4245 & n4246 ;
  assign n4248 = n2345 & ~n2353 ;
  assign n4249 = n2357 & ~n4248 ;
  assign n4250 = ~n4247 & n4249 ;
  assign n4251 = n1898 & ~n4250 ;
  assign n4252 = ~n1898 & n4250 ;
  assign n4253 = ~n4251 & ~n4252 ;
  assign n4254 = n2053 & n4253 ;
  assign n4255 = ~n4235 & ~n4254 ;
  assign n4256 = ~n2224 & ~n4255 ;
  assign n4233 = ~n1334 & n2229 ;
  assign n4234 = ~n1304 & ~n2274 ;
  assign n4293 = ~n4233 & ~n4234 ;
  assign n4294 = ~n4256 & n4293 ;
  assign n4272 = n858 & n1344 ;
  assign n4273 = ~n1820 & ~n4272 ;
  assign n4274 = n774 & n1344 ;
  assign n4275 = n968 & n1826 ;
  assign n4276 = ~n853 & ~n4275 ;
  assign n4277 = n960 & n1814 ;
  assign n4278 = ~n1824 & ~n4277 ;
  assign n4279 = n960 & n1028 ;
  assign n4280 = ~n1811 & n4279 ;
  assign n4281 = n4278 & ~n4280 ;
  assign n4282 = n911 & n968 ;
  assign n4283 = ~n4281 & n4282 ;
  assign n4284 = n4276 & ~n4283 ;
  assign n4285 = n4274 & ~n4284 ;
  assign n4286 = n4273 & ~n4285 ;
  assign n4287 = n1898 & ~n4286 ;
  assign n4288 = ~n1898 & n4286 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4290 = n2053 & ~n4289 ;
  assign n4291 = ~n4235 & ~n4290 ;
  assign n4292 = ~n2120 & ~n4291 ;
  assign n4257 = ~n1304 & ~n2124 ;
  assign n4258 = n2124 & n4253 ;
  assign n4259 = ~n4257 & ~n4258 ;
  assign n4260 = n2123 & ~n4259 ;
  assign n4261 = ~n1193 & n2247 ;
  assign n4262 = ~n1309 & n4261 ;
  assign n4264 = ~n1269 & n4262 ;
  assign n4263 = n1269 & ~n4262 ;
  assign n4265 = n2263 & ~n4263 ;
  assign n4266 = ~n4264 & n4265 ;
  assign n4267 = ~n1193 & ~n2263 ;
  assign n4268 = ~n4266 & ~n4267 ;
  assign n4269 = n2124 & ~n4268 ;
  assign n4270 = ~n4257 & ~n4269 ;
  assign n4271 = n1790 & ~n4270 ;
  assign n4295 = ~n4260 & ~n4271 ;
  assign n4296 = ~n4292 & n4295 ;
  assign n4297 = n4294 & n4296 ;
  assign n4298 = n2037 & ~n4297 ;
  assign n4299 = ~n4232 & ~n4298 ;
  assign n4300 = \P1_state_reg[0]/NET0131  & ~n4299 ;
  assign n4230 = ~n1304 & n2014 ;
  assign n4231 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[18]/NET0131  ;
  assign n4301 = ~n4230 & ~n4231 ;
  assign n4302 = ~n4300 & n4301 ;
  assign n4305 = ~n1264 & n2035 ;
  assign n4308 = ~n1264 & ~n2053 ;
  assign n4309 = n1948 & ~n2192 ;
  assign n4310 = ~n1948 & n2192 ;
  assign n4311 = ~n4309 & ~n4310 ;
  assign n4312 = n2053 & ~n4311 ;
  assign n4313 = ~n4308 & ~n4312 ;
  assign n4314 = ~n2224 & ~n4313 ;
  assign n4306 = ~n1264 & ~n2274 ;
  assign n4307 = ~n1299 & n2229 ;
  assign n4334 = ~n4306 & ~n4307 ;
  assign n4335 = ~n4314 & n4334 ;
  assign n4328 = n1948 & ~n2092 ;
  assign n4329 = ~n1948 & n2092 ;
  assign n4330 = ~n4328 & ~n4329 ;
  assign n4331 = n2053 & n4330 ;
  assign n4332 = ~n4308 & ~n4331 ;
  assign n4333 = ~n2120 & ~n4332 ;
  assign n4315 = ~n1264 & ~n2124 ;
  assign n4316 = ~n1309 & ~n2263 ;
  assign n4317 = n1410 & ~n4264 ;
  assign n4318 = n2248 & n4262 ;
  assign n4319 = n2263 & ~n4318 ;
  assign n4320 = ~n4317 & n4319 ;
  assign n4321 = ~n4316 & ~n4320 ;
  assign n4322 = n2124 & ~n4321 ;
  assign n4323 = ~n4315 & ~n4322 ;
  assign n4324 = n1790 & ~n4323 ;
  assign n4325 = n2124 & ~n4311 ;
  assign n4326 = ~n4315 & ~n4325 ;
  assign n4327 = n2123 & ~n4326 ;
  assign n4336 = ~n4324 & ~n4327 ;
  assign n4337 = ~n4333 & n4336 ;
  assign n4338 = n4335 & n4337 ;
  assign n4339 = n2037 & ~n4338 ;
  assign n4340 = ~n4305 & ~n4339 ;
  assign n4341 = \P1_state_reg[0]/NET0131  & ~n4340 ;
  assign n4303 = ~n1264 & n2014 ;
  assign n4304 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[19]/NET0131  ;
  assign n4342 = ~n4303 & ~n4304 ;
  assign n4343 = ~n4341 & n4342 ;
  assign n4346 = ~n1188 & n2035 ;
  assign n4348 = ~n1188 & ~n2053 ;
  assign n4349 = n2619 & ~n2629 ;
  assign n4350 = n2632 & ~n4349 ;
  assign n4351 = n1899 & n4350 ;
  assign n4352 = ~n1899 & ~n4350 ;
  assign n4353 = ~n4351 & ~n4352 ;
  assign n4354 = n2053 & n4353 ;
  assign n4355 = ~n4348 & ~n4354 ;
  assign n4356 = ~n2224 & ~n4355 ;
  assign n4357 = ~n1188 & ~n2124 ;
  assign n4369 = n1309 & ~n4261 ;
  assign n4370 = n2263 & ~n4262 ;
  assign n4371 = ~n4369 & n4370 ;
  assign n4372 = ~n1231 & ~n2263 ;
  assign n4373 = ~n4371 & ~n4372 ;
  assign n4374 = n2124 & ~n4373 ;
  assign n4375 = ~n4357 & ~n4374 ;
  assign n4376 = n1790 & ~n4375 ;
  assign n4347 = ~n1188 & ~n2274 ;
  assign n4377 = ~n1221 & n2229 ;
  assign n4378 = ~n4347 & ~n4377 ;
  assign n4379 = ~n4376 & n4378 ;
  assign n4380 = ~n4356 & n4379 ;
  assign n4358 = n2124 & n4353 ;
  assign n4359 = ~n4357 & ~n4358 ;
  assign n4360 = n2123 & ~n4359 ;
  assign n4361 = n2561 & ~n2571 ;
  assign n4362 = n2574 & ~n4361 ;
  assign n4363 = n1899 & n4362 ;
  assign n4364 = ~n1899 & ~n4362 ;
  assign n4365 = ~n4363 & ~n4364 ;
  assign n4366 = n2053 & ~n4365 ;
  assign n4367 = ~n4348 & ~n4366 ;
  assign n4368 = ~n2120 & ~n4367 ;
  assign n4381 = ~n4360 & ~n4368 ;
  assign n4382 = n4380 & n4381 ;
  assign n4383 = n2037 & ~n4382 ;
  assign n4384 = ~n4346 & ~n4383 ;
  assign n4385 = \P1_state_reg[0]/NET0131  & ~n4384 ;
  assign n4344 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[17]/NET0131  ;
  assign n4345 = ~n1188 & n2014 ;
  assign n4386 = ~n4344 & ~n4345 ;
  assign n4387 = ~n4385 & n4386 ;
  assign n4390 = ~n1470 & n2035 ;
  assign n4403 = ~n1470 & ~n2124 ;
  assign n4392 = n2360 & n2367 ;
  assign n4393 = n2374 & ~n4392 ;
  assign n4394 = n2344 & n2367 ;
  assign n4395 = ~n4250 & n4394 ;
  assign n4396 = n4393 & ~n4395 ;
  assign n4397 = n1944 & n4396 ;
  assign n4398 = ~n1944 & ~n4396 ;
  assign n4399 = ~n4397 & ~n4398 ;
  assign n4404 = n2124 & ~n4399 ;
  assign n4405 = ~n4403 & ~n4404 ;
  assign n4406 = n2123 & ~n4405 ;
  assign n4391 = ~n1470 & ~n2053 ;
  assign n4400 = n2053 & ~n4399 ;
  assign n4401 = ~n4391 & ~n4400 ;
  assign n4402 = ~n2224 & ~n4401 ;
  assign n4408 = n2250 & n4261 ;
  assign n4409 = ~n1474 & n4408 ;
  assign n4411 = n1445 & ~n4409 ;
  assign n4410 = ~n1445 & n4409 ;
  assign n4412 = n2263 & ~n4410 ;
  assign n4413 = ~n4411 & n4412 ;
  assign n4414 = ~n1382 & ~n2263 ;
  assign n4415 = ~n4413 & ~n4414 ;
  assign n4416 = n2124 & ~n4415 ;
  assign n4417 = ~n4403 & ~n4416 ;
  assign n4418 = n1790 & ~n4417 ;
  assign n4419 = n1484 & n1822 ;
  assign n4420 = ~n1833 & ~n4419 ;
  assign n4421 = n1341 & n1484 ;
  assign n4425 = n4274 & n4282 ;
  assign n4426 = n4280 & n4425 ;
  assign n4422 = ~n4278 & n4282 ;
  assign n4423 = n4276 & ~n4422 ;
  assign n4424 = n4274 & ~n4423 ;
  assign n4427 = n4273 & ~n4424 ;
  assign n4428 = ~n4426 & n4427 ;
  assign n4429 = n4421 & ~n4428 ;
  assign n4430 = n4420 & ~n4429 ;
  assign n4431 = n1944 & ~n4430 ;
  assign n4432 = ~n1944 & n4430 ;
  assign n4433 = ~n4431 & ~n4432 ;
  assign n4434 = n2053 & ~n4433 ;
  assign n4435 = ~n4391 & ~n4434 ;
  assign n4436 = ~n2120 & ~n4435 ;
  assign n4407 = ~n1470 & ~n2274 ;
  assign n4437 = n1465 & n2229 ;
  assign n4438 = ~n4407 & ~n4437 ;
  assign n4439 = ~n4436 & n4438 ;
  assign n4440 = ~n4418 & n4439 ;
  assign n4441 = ~n4402 & n4440 ;
  assign n4442 = ~n4406 & n4441 ;
  assign n4443 = n2037 & ~n4442 ;
  assign n4444 = ~n4390 & ~n4443 ;
  assign n4445 = \P1_state_reg[0]/NET0131  & ~n4444 ;
  assign n4388 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[22]/NET0131  ;
  assign n4389 = ~n1470 & n2014 ;
  assign n4446 = ~n4388 & ~n4389 ;
  assign n4447 = ~n4445 & n4446 ;
  assign n4448 = n3074 & n4081 ;
  assign n4449 = ~n2711 & ~n2716 ;
  assign n4450 = n3074 & ~n4449 ;
  assign n4451 = ~n3079 & ~n3188 ;
  assign n4452 = ~n3766 & n3771 ;
  assign n4453 = n3180 & ~n4452 ;
  assign n4454 = ~n2975 & n3130 ;
  assign n4455 = ~n4453 & n4454 ;
  assign n4456 = ~n2975 & ~n3185 ;
  assign n4457 = n3191 & ~n4456 ;
  assign n4458 = ~n4455 & n4457 ;
  assign n4459 = ~n3027 & ~n4458 ;
  assign n4460 = n3421 & n3522 ;
  assign n4461 = ~n3528 & ~n4460 ;
  assign n4462 = n3472 & n3537 ;
  assign n4463 = ~n4461 & n4462 ;
  assign n4464 = ~n3533 & n3537 ;
  assign n4465 = ~n3303 & ~n4464 ;
  assign n4466 = ~n4463 & n4465 ;
  assign n4467 = n3250 & n3694 ;
  assign n4468 = n3642 & n3743 ;
  assign n4469 = n4467 & n4468 ;
  assign n4470 = ~n4466 & n4469 ;
  assign n4471 = n3308 & n3694 ;
  assign n4472 = ~n3750 & ~n4471 ;
  assign n4473 = n4468 & ~n4472 ;
  assign n4474 = n3642 & n3755 ;
  assign n4475 = ~n3761 & ~n4474 ;
  assign n4476 = ~n4473 & n4475 ;
  assign n4477 = ~n4470 & n4476 ;
  assign n4478 = n3589 & n3771 ;
  assign n4479 = ~n3027 & n4454 ;
  assign n4480 = n4478 & n4479 ;
  assign n4481 = ~n4477 & n4480 ;
  assign n4482 = ~n4459 & ~n4481 ;
  assign n4483 = n4451 & n4482 ;
  assign n4484 = ~n4451 & ~n4482 ;
  assign n4485 = ~n4483 & ~n4484 ;
  assign n4486 = n4449 & ~n4485 ;
  assign n4487 = ~n4450 & ~n4486 ;
  assign n4488 = n3829 & ~n4487 ;
  assign n4489 = n3874 & n3881 ;
  assign n4490 = n3878 & n3881 ;
  assign n4491 = ~n3838 & ~n4490 ;
  assign n4492 = ~n4489 & n4491 ;
  assign n4493 = n3833 & n3919 ;
  assign n4494 = n3887 & n3916 ;
  assign n4495 = n4493 & n4494 ;
  assign n4496 = ~n4492 & n4495 ;
  assign n4497 = ~n3843 & n3919 ;
  assign n4498 = ~n3892 & ~n4497 ;
  assign n4499 = n4494 & ~n4498 ;
  assign n4500 = n3897 & n3916 ;
  assign n4501 = ~n3906 & ~n4500 ;
  assign n4502 = ~n4499 & n4501 ;
  assign n4503 = ~n4496 & n4502 ;
  assign n4504 = n3901 & n3933 ;
  assign n4505 = n3929 & n3936 ;
  assign n4506 = n4504 & n4505 ;
  assign n4507 = ~n4503 & n4506 ;
  assign n4508 = n3911 & n3933 ;
  assign n4509 = ~n3944 & ~n4508 ;
  assign n4510 = n4505 & ~n4509 ;
  assign n4511 = n3929 & ~n3949 ;
  assign n4512 = ~n3955 & ~n4511 ;
  assign n4513 = ~n4510 & n4512 ;
  assign n4514 = ~n4507 & n4513 ;
  assign n4515 = n4451 & ~n4514 ;
  assign n4516 = ~n4451 & n4514 ;
  assign n4517 = ~n4515 & ~n4516 ;
  assign n4518 = n4449 & ~n4517 ;
  assign n4519 = ~n4450 & ~n4518 ;
  assign n4520 = n3969 & ~n4519 ;
  assign n4530 = n2731 & ~n3026 ;
  assign n4531 = n4001 & n4006 ;
  assign n4532 = n2904 & ~n4531 ;
  assign n4533 = ~n2731 & ~n4008 ;
  assign n4534 = ~n4532 & n4533 ;
  assign n4535 = ~n4530 & ~n4534 ;
  assign n4536 = n4449 & ~n4535 ;
  assign n4537 = ~n4450 & ~n4536 ;
  assign n4538 = n4025 & ~n4537 ;
  assign n4524 = ~n3017 & n4054 ;
  assign n4525 = n3069 & ~n4524 ;
  assign n4526 = ~n3069 & n4524 ;
  assign n4527 = ~n4525 & ~n4526 ;
  assign n4528 = n4062 & n4527 ;
  assign n4529 = n4449 & n4528 ;
  assign n4521 = n4028 & n4449 ;
  assign n4522 = ~n4073 & ~n4521 ;
  assign n4523 = n3069 & ~n4522 ;
  assign n4539 = n4028 & ~n4449 ;
  assign n4540 = ~n4067 & ~n4539 ;
  assign n4541 = n4062 & ~n4449 ;
  assign n4542 = n4540 & ~n4541 ;
  assign n4543 = n3074 & ~n4542 ;
  assign n4544 = ~n4523 & ~n4543 ;
  assign n4545 = ~n4529 & n4544 ;
  assign n4546 = ~n4538 & n4545 ;
  assign n4547 = ~n4520 & n4546 ;
  assign n4548 = ~n4488 & n4547 ;
  assign n4549 = n2701 & ~n4548 ;
  assign n4550 = ~n4448 & ~n4549 ;
  assign n4551 = \P1_state_reg[0]/NET0131  & ~n4550 ;
  assign n4552 = \P1_state_reg[0]/NET0131  & n2683 ;
  assign n4553 = n3074 & n4552 ;
  assign n4554 = \P1_reg3_reg[27]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4555 = ~n4553 & ~n4554 ;
  assign n4556 = ~n4551 & n4555 ;
  assign n4557 = \P2_reg2_reg[22]/NET0131  & ~n2286 ;
  assign n4558 = \P2_reg2_reg[22]/NET0131  & n2035 ;
  assign n4559 = \P2_reg2_reg[22]/NET0131  & ~n2291 ;
  assign n4560 = n2291 & ~n4399 ;
  assign n4561 = ~n4559 & ~n4560 ;
  assign n4562 = ~n2392 & ~n4561 ;
  assign n4563 = \P2_reg2_reg[22]/NET0131  & ~n2310 ;
  assign n4564 = n2310 & ~n4415 ;
  assign n4565 = ~n4563 & ~n4564 ;
  assign n4566 = n1790 & ~n4565 ;
  assign n4572 = n2310 & ~n4433 ;
  assign n4573 = ~n4563 & ~n4572 ;
  assign n4574 = n2314 & ~n4573 ;
  assign n4567 = n2291 & ~n4433 ;
  assign n4568 = ~n4559 & ~n4567 ;
  assign n4569 = ~n2290 & ~n4568 ;
  assign n4570 = n1465 & n2272 ;
  assign n4571 = n2291 & n4570 ;
  assign n4575 = ~n1470 & n1854 ;
  assign n4576 = \P2_reg2_reg[22]/NET0131  & ~n2407 ;
  assign n4577 = ~n4575 & ~n4576 ;
  assign n4578 = ~n4571 & n4577 ;
  assign n4579 = ~n4569 & n4578 ;
  assign n4580 = ~n4574 & n4579 ;
  assign n4581 = ~n4566 & n4580 ;
  assign n4582 = ~n4562 & n4581 ;
  assign n4583 = n2037 & ~n4582 ;
  assign n4584 = ~n4558 & ~n4583 ;
  assign n4585 = \P1_state_reg[0]/NET0131  & ~n4584 ;
  assign n4586 = ~n4557 & ~n4585 ;
  assign n4587 = \P2_reg0_reg[27]/NET0131  & ~n2286 ;
  assign n4588 = \P2_reg0_reg[27]/NET0131  & n2035 ;
  assign n4589 = \P2_reg0_reg[27]/NET0131  & ~n2124 ;
  assign n4590 = ~n2116 & n2124 ;
  assign n4591 = ~n4589 & ~n4590 ;
  assign n4592 = ~n2120 & ~n4591 ;
  assign n4593 = \P2_reg0_reg[27]/NET0131  & ~n2053 ;
  assign n4599 = n2053 & ~n2267 ;
  assign n4600 = ~n4593 & ~n4599 ;
  assign n4601 = n1790 & ~n4600 ;
  assign n4598 = n1608 & n2616 ;
  assign n4602 = \P2_reg0_reg[27]/NET0131  & ~n2614 ;
  assign n4603 = ~n4598 & ~n4602 ;
  assign n4604 = ~n4601 & n4603 ;
  assign n4605 = ~n4592 & n4604 ;
  assign n4594 = ~n2225 & ~n4593 ;
  assign n4595 = n2123 & ~n4594 ;
  assign n4596 = ~n2221 & ~n4589 ;
  assign n4597 = ~n2224 & ~n4596 ;
  assign n4606 = ~n4595 & ~n4597 ;
  assign n4607 = n4605 & n4606 ;
  assign n4608 = n2037 & ~n4607 ;
  assign n4609 = ~n4588 & ~n4608 ;
  assign n4610 = \P1_state_reg[0]/NET0131  & ~n4609 ;
  assign n4611 = ~n4587 & ~n4610 ;
  assign n4612 = \P2_reg0_reg[28]/NET0131  & ~n2286 ;
  assign n4613 = \P2_reg0_reg[28]/NET0131  & n2035 ;
  assign n4614 = \P2_reg0_reg[28]/NET0131  & ~n2124 ;
  assign n4615 = n2124 & ~n2306 ;
  assign n4616 = ~n4614 & ~n4615 ;
  assign n4617 = ~n2120 & ~n4616 ;
  assign n4620 = \P2_reg0_reg[28]/NET0131  & ~n2053 ;
  assign n4625 = n2053 & ~n2402 ;
  assign n4626 = ~n4620 & ~n4625 ;
  assign n4627 = n1790 & ~n4626 ;
  assign n4623 = n1684 & n2272 ;
  assign n4624 = n2124 & n4623 ;
  assign n4628 = \P2_reg0_reg[28]/NET0131  & ~n2614 ;
  assign n4629 = ~n4624 & ~n4628 ;
  assign n4630 = ~n4627 & n4629 ;
  assign n4631 = ~n4617 & n4630 ;
  assign n4618 = ~n2428 & ~n4614 ;
  assign n4619 = ~n2224 & ~n4618 ;
  assign n4621 = ~n2431 & ~n4620 ;
  assign n4622 = n2123 & ~n4621 ;
  assign n4632 = ~n4619 & ~n4622 ;
  assign n4633 = n4631 & n4632 ;
  assign n4634 = n2037 & ~n4633 ;
  assign n4635 = ~n4613 & ~n4634 ;
  assign n4636 = \P1_state_reg[0]/NET0131  & ~n4635 ;
  assign n4637 = ~n4612 & ~n4636 ;
  assign n4638 = \P1_reg2_reg[28]/NET0131  & ~n4085 ;
  assign n4639 = \P1_reg2_reg[28]/NET0131  & n4081 ;
  assign n4640 = \P1_reg2_reg[28]/NET0131  & ~n2717 ;
  assign n4641 = ~n3471 & ~n3495 ;
  assign n4642 = n3373 & ~n3414 ;
  assign n4643 = ~n3372 & n3374 ;
  assign n4644 = ~n3418 & ~n4643 ;
  assign n4645 = ~n4642 & n4644 ;
  assign n4646 = ~n3333 & ~n3521 ;
  assign n4647 = ~n4645 & n4646 ;
  assign n4648 = ~n3417 & ~n3526 ;
  assign n4649 = ~n3521 & ~n4648 ;
  assign n4650 = ~n4647 & ~n4649 ;
  assign n4651 = n4641 & ~n4650 ;
  assign n4652 = ~n3525 & ~n3531 ;
  assign n4653 = ~n3471 & ~n4652 ;
  assign n4654 = ~n4651 & ~n4653 ;
  assign n4655 = ~n3445 & ~n3536 ;
  assign n4656 = ~n3222 & ~n3276 ;
  assign n4657 = n4655 & n4656 ;
  assign n4658 = ~n4654 & n4657 ;
  assign n4659 = n3530 & ~n3536 ;
  assign n4660 = ~n3301 & ~n4659 ;
  assign n4661 = n4656 & ~n4660 ;
  assign n4662 = ~n3222 & n3277 ;
  assign n4663 = ~n3306 & ~n4662 ;
  assign n4664 = ~n4661 & n4663 ;
  assign n4665 = ~n4658 & n4664 ;
  assign n4666 = ~n3666 & ~n3742 ;
  assign n4667 = ~n3249 & ~n3693 ;
  assign n4668 = n4666 & n4667 ;
  assign n4669 = ~n3614 & ~n3718 ;
  assign n4670 = ~n3588 & ~n3641 ;
  assign n4671 = n4669 & n4670 ;
  assign n4672 = n4668 & n4671 ;
  assign n4673 = ~n4665 & n4672 ;
  assign n4674 = ~n3305 & ~n3748 ;
  assign n4675 = ~n3693 & ~n4674 ;
  assign n4676 = n4666 & n4675 ;
  assign n4677 = ~n3747 & ~n3753 ;
  assign n4678 = ~n3742 & ~n4677 ;
  assign n4679 = ~n4676 & ~n4678 ;
  assign n4680 = n4671 & ~n4679 ;
  assign n4681 = ~n3614 & n3752 ;
  assign n4682 = ~n3759 & ~n4681 ;
  assign n4683 = n4670 & ~n4682 ;
  assign n4684 = ~n3758 & ~n3764 ;
  assign n4685 = ~n3588 & ~n4684 ;
  assign n4686 = ~n4683 & ~n4685 ;
  assign n4687 = ~n4680 & n4686 ;
  assign n4688 = ~n4673 & n4687 ;
  assign n4689 = ~n3562 & ~n3770 ;
  assign n4690 = ~n3129 & ~n3155 ;
  assign n4691 = n4689 & n4690 ;
  assign n4692 = n3081 & ~n3106 ;
  assign n4693 = n4691 & n4692 ;
  assign n4694 = ~n4688 & n4693 ;
  assign n4696 = n3763 & ~n3770 ;
  assign n4697 = ~n3178 & ~n4696 ;
  assign n4698 = n4690 & ~n4697 ;
  assign n4699 = ~n3129 & n3154 ;
  assign n4700 = ~n3183 & ~n4699 ;
  assign n4701 = ~n4698 & n4700 ;
  assign n4702 = n4692 & ~n4701 ;
  assign n4703 = ~n3182 & ~n3190 ;
  assign n4704 = n3081 & ~n4703 ;
  assign n4695 = ~n3079 & n3189 ;
  assign n4705 = ~n3188 & ~n4695 ;
  assign n4706 = ~n4704 & n4705 ;
  assign n4707 = ~n4702 & n4706 ;
  assign n4708 = ~n4694 & n4707 ;
  assign n4709 = ~n2905 & ~n3193 ;
  assign n4710 = n4708 & n4709 ;
  assign n4711 = ~n4708 & ~n4709 ;
  assign n4712 = ~n4710 & ~n4711 ;
  assign n4713 = n2717 & ~n4712 ;
  assign n4714 = ~n4640 & ~n4713 ;
  assign n4715 = n3829 & ~n4714 ;
  assign n4716 = ~n3885 & ~n3915 ;
  assign n4717 = ~n3900 & ~n3902 ;
  assign n4718 = n4716 & n4717 ;
  assign n4725 = ~n3850 & ~n3851 ;
  assign n4726 = n3857 & ~n4725 ;
  assign n4727 = ~n3846 & ~n3852 ;
  assign n4728 = ~n3856 & ~n4727 ;
  assign n4729 = ~n4726 & ~n4728 ;
  assign n4719 = ~n3860 & ~n3872 ;
  assign n4730 = n3863 & n4719 ;
  assign n4731 = ~n4729 & n4730 ;
  assign n4720 = ~n3845 & ~n3867 ;
  assign n4721 = ~n3862 & ~n4720 ;
  assign n4722 = n4719 & n4721 ;
  assign n4723 = n3866 & ~n3872 ;
  assign n4724 = ~n3876 & ~n4723 ;
  assign n4732 = ~n4722 & n4724 ;
  assign n4733 = ~n4731 & n4732 ;
  assign n4734 = ~n3871 & ~n3880 ;
  assign n4735 = ~n3831 & ~n3834 ;
  assign n4736 = n4734 & n4735 ;
  assign n4737 = ~n4733 & n4736 ;
  assign n4738 = ~n3835 & ~n3875 ;
  assign n4739 = ~n3880 & ~n4738 ;
  assign n4740 = n4735 & n4739 ;
  assign n4741 = ~n3836 & ~n3841 ;
  assign n4742 = ~n3831 & ~n4741 ;
  assign n4743 = ~n4740 & ~n4742 ;
  assign n4744 = ~n4737 & n4743 ;
  assign n4745 = ~n3886 & ~n3888 ;
  assign n4746 = ~n3832 & ~n3918 ;
  assign n4747 = n4745 & n4746 ;
  assign n4748 = ~n4744 & n4747 ;
  assign n4749 = n4718 & n4748 ;
  assign n4750 = ~n3840 & ~n3889 ;
  assign n4751 = ~n3918 & ~n4750 ;
  assign n4752 = n4745 & n4751 ;
  assign n4753 = ~n3890 & ~n3895 ;
  assign n4754 = ~n3886 & ~n4753 ;
  assign n4755 = ~n4752 & ~n4754 ;
  assign n4756 = n4718 & ~n4755 ;
  assign n4757 = ~n3894 & ~n3904 ;
  assign n4758 = ~n3915 & ~n4757 ;
  assign n4759 = n4717 & n4758 ;
  assign n4760 = ~n3903 & ~n3909 ;
  assign n4761 = ~n3900 & ~n4760 ;
  assign n4762 = ~n4759 & ~n4761 ;
  assign n4763 = ~n4756 & n4762 ;
  assign n4764 = ~n4749 & n4763 ;
  assign n4765 = ~n3899 & ~n3931 ;
  assign n4766 = ~n3932 & ~n3934 ;
  assign n4767 = n4765 & n4766 ;
  assign n4768 = ~n3927 & ~n3935 ;
  assign n4769 = ~n3924 & ~n3928 ;
  assign n4770 = n4768 & n4769 ;
  assign n4771 = n4767 & n4770 ;
  assign n4772 = ~n4764 & n4771 ;
  assign n4773 = n3908 & ~n3931 ;
  assign n4774 = ~n3942 & ~n4773 ;
  assign n4775 = n4766 & ~n4774 ;
  assign n4776 = ~n3941 & ~n3947 ;
  assign n4777 = ~n3934 & ~n4776 ;
  assign n4778 = ~n4775 & ~n4777 ;
  assign n4779 = n4770 & ~n4778 ;
  assign n4780 = ~n3952 & ~n3958 ;
  assign n4781 = ~n3946 & ~n3953 ;
  assign n4782 = ~n3927 & ~n4781 ;
  assign n4783 = ~n3928 & n4782 ;
  assign n4784 = n4780 & ~n4783 ;
  assign n4785 = ~n3924 & ~n4784 ;
  assign n4786 = ~n4779 & ~n4785 ;
  assign n4787 = ~n4772 & n4786 ;
  assign n4788 = n4709 & ~n4787 ;
  assign n4789 = ~n4709 & n4787 ;
  assign n4790 = ~n4788 & ~n4789 ;
  assign n4791 = n2717 & ~n4790 ;
  assign n4792 = ~n4640 & ~n4791 ;
  assign n4793 = n3969 & ~n4792 ;
  assign n4794 = n2868 & n4028 ;
  assign n4795 = n2868 & ~n4526 ;
  assign n4796 = ~n4057 & ~n4795 ;
  assign n4797 = n4062 & n4796 ;
  assign n4798 = ~n4794 & ~n4797 ;
  assign n4799 = n2717 & ~n4798 ;
  assign n4800 = n3801 & ~n4008 ;
  assign n4801 = ~n4009 & ~n4800 ;
  assign n4802 = ~n2731 & ~n4801 ;
  assign n4803 = n2731 & n3078 ;
  assign n4804 = ~n4802 & ~n4803 ;
  assign n4805 = n2717 & n4804 ;
  assign n4806 = ~n4640 & ~n4805 ;
  assign n4807 = n4025 & ~n4806 ;
  assign n4808 = \P1_reg2_reg[28]/NET0131  & ~n4071 ;
  assign n4809 = n2900 & n4073 ;
  assign n4810 = ~n4808 & ~n4809 ;
  assign n4811 = ~n4807 & n4810 ;
  assign n4812 = ~n4799 & n4811 ;
  assign n4813 = ~n4793 & n4812 ;
  assign n4814 = ~n4715 & n4813 ;
  assign n4815 = n2701 & ~n4814 ;
  assign n4816 = ~n4639 & ~n4815 ;
  assign n4817 = \P1_state_reg[0]/NET0131  & ~n4816 ;
  assign n4818 = ~n4638 & ~n4817 ;
  assign n4819 = \P2_reg1_reg[27]/NET0131  & ~n2286 ;
  assign n4820 = \P2_reg1_reg[27]/NET0131  & n2035 ;
  assign n4821 = \P2_reg1_reg[27]/NET0131  & ~n2310 ;
  assign n4822 = ~n2459 & ~n4821 ;
  assign n4823 = ~n2290 & ~n4822 ;
  assign n4827 = \P2_reg1_reg[27]/NET0131  & ~n2291 ;
  assign n4831 = ~n2267 & n2291 ;
  assign n4832 = ~n4827 & ~n4831 ;
  assign n4833 = n1790 & ~n4832 ;
  assign n4830 = n1608 & n4101 ;
  assign n4834 = \P2_reg1_reg[27]/NET0131  & ~n4099 ;
  assign n4835 = ~n4830 & ~n4834 ;
  assign n4836 = ~n4833 & n4835 ;
  assign n4837 = ~n4823 & n4836 ;
  assign n4824 = ~n2220 & n2310 ;
  assign n4825 = ~n4821 & ~n4824 ;
  assign n4826 = ~n2392 & ~n4825 ;
  assign n4828 = ~n2452 & ~n4827 ;
  assign n4829 = n2314 & ~n4828 ;
  assign n4838 = ~n4826 & ~n4829 ;
  assign n4839 = n4837 & n4838 ;
  assign n4840 = n2037 & ~n4839 ;
  assign n4841 = ~n4820 & ~n4840 ;
  assign n4842 = \P1_state_reg[0]/NET0131  & ~n4841 ;
  assign n4843 = ~n4819 & ~n4842 ;
  assign n4844 = \P2_reg1_reg[28]/NET0131  & ~n2286 ;
  assign n4845 = \P2_reg1_reg[28]/NET0131  & n2035 ;
  assign n4846 = \P2_reg1_reg[28]/NET0131  & ~n2310 ;
  assign n4847 = ~n2312 & ~n4846 ;
  assign n4848 = ~n2290 & ~n4847 ;
  assign n4852 = \P2_reg1_reg[28]/NET0131  & ~n2291 ;
  assign n4856 = n2291 & ~n2402 ;
  assign n4857 = ~n4852 & ~n4856 ;
  assign n4858 = n1790 & ~n4857 ;
  assign n4855 = n2310 & n4623 ;
  assign n4859 = \P2_reg1_reg[28]/NET0131  & ~n4099 ;
  assign n4860 = ~n4855 & ~n4859 ;
  assign n4861 = ~n4858 & n4860 ;
  assign n4862 = ~n4848 & n4861 ;
  assign n4849 = n2310 & ~n2389 ;
  assign n4850 = ~n4846 & ~n4849 ;
  assign n4851 = ~n2392 & ~n4850 ;
  assign n4853 = ~n2307 & ~n4852 ;
  assign n4854 = n2314 & ~n4853 ;
  assign n4863 = ~n4851 & ~n4854 ;
  assign n4864 = n4862 & n4863 ;
  assign n4865 = n2037 & ~n4864 ;
  assign n4866 = ~n4845 & ~n4865 ;
  assign n4867 = \P1_state_reg[0]/NET0131  & ~n4866 ;
  assign n4868 = ~n4844 & ~n4867 ;
  assign n4869 = n2711 & n2716 ;
  assign n4870 = \P1_reg0_reg[29]/NET0131  & ~n4869 ;
  assign n4871 = ~n3807 & n4869 ;
  assign n4872 = ~n4870 & ~n4871 ;
  assign n4873 = n3829 & ~n4872 ;
  assign n4874 = n3966 & n4869 ;
  assign n4875 = ~n4870 & ~n4874 ;
  assign n4876 = n3969 & ~n4875 ;
  assign n4877 = ~n4020 & n4869 ;
  assign n4878 = ~n4870 & ~n4877 ;
  assign n4879 = n4025 & ~n4878 ;
  assign n4880 = n4060 & n4869 ;
  assign n4881 = ~n4870 & ~n4880 ;
  assign n4882 = n4062 & ~n4881 ;
  assign n4883 = \P1_reg0_reg[29]/NET0131  & ~n4214 ;
  assign n4884 = n3794 & n4869 ;
  assign n4885 = ~n4870 & ~n4884 ;
  assign n4886 = n4028 & ~n4885 ;
  assign n4887 = ~n4883 & ~n4886 ;
  assign n4888 = ~n4882 & n4887 ;
  assign n4889 = ~n4879 & n4888 ;
  assign n4890 = ~n4876 & n4889 ;
  assign n4891 = ~n4873 & n4890 ;
  assign n4892 = n2701 & ~n4891 ;
  assign n4893 = \P1_reg0_reg[29]/NET0131  & n4081 ;
  assign n4894 = ~n4892 & ~n4893 ;
  assign n4895 = \P1_state_reg[0]/NET0131  & ~n4894 ;
  assign n4896 = \P1_reg0_reg[29]/NET0131  & ~n4085 ;
  assign n4897 = ~n4895 & ~n4896 ;
  assign n4898 = \P2_reg2_reg[20]/NET0131  & ~n2286 ;
  assign n4899 = \P2_reg2_reg[20]/NET0131  & n2035 ;
  assign n4900 = \P2_reg2_reg[20]/NET0131  & ~n2310 ;
  assign n4901 = ~n1269 & ~n2263 ;
  assign n4902 = n1382 & ~n4318 ;
  assign n4903 = n2263 & ~n4408 ;
  assign n4904 = ~n4902 & n4903 ;
  assign n4905 = ~n4901 & ~n4904 ;
  assign n4906 = n2310 & ~n4905 ;
  assign n4907 = ~n4900 & ~n4906 ;
  assign n4908 = n1790 & ~n4907 ;
  assign n4927 = n1401 & n2394 ;
  assign n4925 = ~n1406 & n1854 ;
  assign n4926 = \P2_reg2_reg[20]/NET0131  & ~n2407 ;
  assign n4928 = ~n4925 & ~n4926 ;
  assign n4929 = ~n4927 & n4928 ;
  assign n4930 = ~n4908 & n4929 ;
  assign n4909 = \P2_reg2_reg[20]/NET0131  & ~n2291 ;
  assign n4916 = n1895 & ~n2298 ;
  assign n4917 = ~n1895 & n2298 ;
  assign n4918 = ~n4916 & ~n4917 ;
  assign n4922 = n2291 & ~n4918 ;
  assign n4923 = ~n4909 & ~n4922 ;
  assign n4924 = ~n2290 & ~n4923 ;
  assign n4910 = n1895 & n2363 ;
  assign n4911 = ~n1895 & ~n2363 ;
  assign n4912 = ~n4910 & ~n4911 ;
  assign n4913 = n2291 & ~n4912 ;
  assign n4914 = ~n4909 & ~n4913 ;
  assign n4915 = ~n2392 & ~n4914 ;
  assign n4919 = n2310 & ~n4918 ;
  assign n4920 = ~n4900 & ~n4919 ;
  assign n4921 = n2314 & ~n4920 ;
  assign n4931 = ~n4915 & ~n4921 ;
  assign n4932 = ~n4924 & n4931 ;
  assign n4933 = n4930 & n4932 ;
  assign n4934 = n2037 & ~n4933 ;
  assign n4935 = ~n4899 & ~n4934 ;
  assign n4936 = \P1_state_reg[0]/NET0131  & ~n4935 ;
  assign n4937 = ~n4898 & ~n4936 ;
  assign n4940 = n3022 & n4081 ;
  assign n4941 = n3022 & ~n4449 ;
  assign n4942 = n3994 & n3996 ;
  assign n4943 = ~n3692 & n4942 ;
  assign n4944 = ~n3665 & n4943 ;
  assign n4945 = ~n3153 & ~n3741 ;
  assign n4946 = n3978 & n4945 ;
  assign n4947 = n4944 & n4946 ;
  assign n4948 = n4004 & n4947 ;
  assign n4949 = n3078 & ~n4948 ;
  assign n4950 = ~n3078 & n4948 ;
  assign n4951 = ~n4949 & ~n4950 ;
  assign n4952 = ~n2731 & ~n4951 ;
  assign n4953 = n2731 & n2974 ;
  assign n4954 = ~n4952 & ~n4953 ;
  assign n4955 = n4449 & n4954 ;
  assign n4956 = ~n4941 & ~n4955 ;
  assign n4957 = n4025 & ~n4956 ;
  assign n5029 = n3017 & ~n4054 ;
  assign n5030 = ~n4524 & ~n5029 ;
  assign n5031 = n4449 & n5030 ;
  assign n5032 = ~n4941 & ~n5031 ;
  assign n5033 = n4062 & ~n5032 ;
  assign n5028 = n3017 & ~n4522 ;
  assign n5034 = n3022 & ~n4540 ;
  assign n5035 = ~n5028 & ~n5034 ;
  assign n5036 = ~n5033 & n5035 ;
  assign n5037 = ~n4957 & n5036 ;
  assign n4958 = ~n3027 & ~n3189 ;
  assign n4959 = n4716 & n4745 ;
  assign n4960 = n3863 & ~n4729 ;
  assign n4961 = ~n4721 & ~n4960 ;
  assign n4962 = n4719 & n4734 ;
  assign n4963 = ~n4961 & n4962 ;
  assign n4964 = ~n4724 & n4734 ;
  assign n4965 = ~n4739 & ~n4964 ;
  assign n4966 = ~n4963 & n4965 ;
  assign n4967 = n4735 & n4746 ;
  assign n4968 = ~n4966 & n4967 ;
  assign n4969 = n4959 & n4968 ;
  assign n4970 = n4742 & n4746 ;
  assign n4971 = ~n4751 & ~n4970 ;
  assign n4972 = n4959 & ~n4971 ;
  assign n4973 = n4716 & n4754 ;
  assign n4974 = ~n4758 & ~n4973 ;
  assign n4975 = ~n4972 & n4974 ;
  assign n4976 = ~n4969 & n4975 ;
  assign n4977 = n4766 & n4768 ;
  assign n4978 = n4717 & n4765 ;
  assign n4979 = n4977 & n4978 ;
  assign n4980 = ~n4976 & n4979 ;
  assign n4981 = n4761 & n4765 ;
  assign n4982 = n4774 & ~n4981 ;
  assign n4983 = n4977 & ~n4982 ;
  assign n4984 = n4768 & n4777 ;
  assign n4985 = ~n4782 & ~n4984 ;
  assign n4986 = ~n4983 & n4985 ;
  assign n4987 = ~n4980 & n4986 ;
  assign n4988 = n4958 & ~n4987 ;
  assign n4989 = ~n4958 & n4987 ;
  assign n4990 = ~n4988 & ~n4989 ;
  assign n4991 = n4449 & ~n4990 ;
  assign n4992 = ~n4941 & ~n4991 ;
  assign n4993 = n3969 & ~n4992 ;
  assign n4994 = n4666 & n4669 ;
  assign n4995 = n4641 & n4655 ;
  assign n4996 = ~n4650 & n4995 ;
  assign n4997 = n4653 & n4655 ;
  assign n4998 = n4660 & ~n4997 ;
  assign n4999 = ~n4996 & n4998 ;
  assign n5000 = n4656 & n4667 ;
  assign n5001 = ~n4999 & n5000 ;
  assign n5002 = n4994 & n5001 ;
  assign n5003 = ~n4663 & n4667 ;
  assign n5004 = ~n4675 & ~n5003 ;
  assign n5005 = n4994 & ~n5004 ;
  assign n5006 = n4669 & n4678 ;
  assign n5007 = n4682 & ~n5006 ;
  assign n5008 = ~n5005 & n5007 ;
  assign n5009 = ~n5002 & n5008 ;
  assign n5010 = n4670 & n4689 ;
  assign n5011 = ~n3155 & n4454 ;
  assign n5012 = n5010 & n5011 ;
  assign n5013 = ~n5009 & n5012 ;
  assign n5014 = n4685 & n4689 ;
  assign n5015 = n4697 & ~n5014 ;
  assign n5016 = n5011 & ~n5015 ;
  assign n5017 = ~n3106 & ~n4700 ;
  assign n5018 = n4703 & ~n5017 ;
  assign n5019 = ~n2975 & ~n5018 ;
  assign n5020 = ~n5016 & ~n5019 ;
  assign n5021 = ~n5013 & n5020 ;
  assign n5022 = n4958 & n5021 ;
  assign n5023 = ~n4958 & ~n5021 ;
  assign n5024 = ~n5022 & ~n5023 ;
  assign n5025 = n4449 & ~n5024 ;
  assign n5026 = ~n4941 & ~n5025 ;
  assign n5027 = n3829 & ~n5026 ;
  assign n5038 = ~n4993 & ~n5027 ;
  assign n5039 = n5037 & n5038 ;
  assign n5040 = n2701 & ~n5039 ;
  assign n5041 = ~n4940 & ~n5040 ;
  assign n5042 = \P1_state_reg[0]/NET0131  & ~n5041 ;
  assign n4938 = \P1_reg3_reg[26]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4939 = n3022 & n4552 ;
  assign n5043 = ~n4938 & ~n4939 ;
  assign n5044 = ~n5042 & n5043 ;
  assign n5045 = \P1_reg2_reg[24]/NET0131  & ~n2717 ;
  assign n5046 = ~n3106 & ~n3182 ;
  assign n5047 = ~n4748 & n4755 ;
  assign n5048 = n4718 & ~n5047 ;
  assign n5049 = n4762 & ~n5048 ;
  assign n5050 = n4767 & ~n5049 ;
  assign n5051 = n4778 & ~n5050 ;
  assign n5052 = n5046 & ~n5051 ;
  assign n5053 = ~n5046 & n5051 ;
  assign n5054 = ~n5052 & ~n5053 ;
  assign n5055 = n2717 & ~n5054 ;
  assign n5056 = ~n5045 & ~n5055 ;
  assign n5057 = n3969 & ~n5056 ;
  assign n5058 = n4658 & n4672 ;
  assign n5059 = ~n4664 & n4668 ;
  assign n5060 = n4679 & ~n5059 ;
  assign n5061 = n4671 & ~n5060 ;
  assign n5062 = n4686 & ~n5061 ;
  assign n5063 = ~n5058 & n5062 ;
  assign n5064 = n4691 & ~n5063 ;
  assign n5065 = n4701 & ~n5064 ;
  assign n5066 = n5046 & n5065 ;
  assign n5067 = ~n5046 & ~n5065 ;
  assign n5068 = ~n5066 & ~n5067 ;
  assign n5069 = n2717 & ~n5068 ;
  assign n5070 = ~n5045 & ~n5069 ;
  assign n5071 = n3829 & ~n5070 ;
  assign n5072 = ~n3128 & ~n3153 ;
  assign n5073 = n4001 & n5072 ;
  assign n5074 = ~n3105 & n5073 ;
  assign n5075 = n2974 & ~n5074 ;
  assign n5076 = ~n2974 & n5074 ;
  assign n5077 = ~n5075 & ~n5076 ;
  assign n5078 = ~n2731 & ~n5077 ;
  assign n5079 = n2731 & n3128 ;
  assign n5080 = ~n5078 & ~n5079 ;
  assign n5081 = n2717 & n5080 ;
  assign n5082 = ~n5045 & ~n5081 ;
  assign n5083 = n4025 & ~n5082 ;
  assign n5085 = n3096 & n4028 ;
  assign n5086 = ~n3119 & n4051 ;
  assign n5087 = n3096 & ~n5086 ;
  assign n5088 = ~n3096 & n5086 ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5090 = n4062 & n5089 ;
  assign n5091 = ~n5085 & ~n5090 ;
  assign n5092 = n2717 & ~n5091 ;
  assign n5084 = \P1_reg2_reg[24]/NET0131  & ~n4071 ;
  assign n5093 = n3101 & n4073 ;
  assign n5094 = ~n5084 & ~n5093 ;
  assign n5095 = ~n5092 & n5094 ;
  assign n5096 = ~n5083 & n5095 ;
  assign n5097 = ~n5071 & n5096 ;
  assign n5098 = ~n5057 & n5097 ;
  assign n5099 = n2701 & ~n5098 ;
  assign n5100 = \P1_reg2_reg[24]/NET0131  & n4081 ;
  assign n5101 = ~n5099 & ~n5100 ;
  assign n5102 = \P1_state_reg[0]/NET0131  & ~n5101 ;
  assign n5103 = \P1_reg2_reg[24]/NET0131  & ~n4085 ;
  assign n5104 = ~n5102 & ~n5103 ;
  assign n5105 = \P1_reg2_reg[25]/NET0131  & ~n4085 ;
  assign n5106 = \P1_reg2_reg[25]/NET0131  & n4081 ;
  assign n5107 = \P1_reg2_reg[25]/NET0131  & ~n2717 ;
  assign n5108 = ~n3026 & ~n5076 ;
  assign n5109 = n3026 & n5076 ;
  assign n5110 = ~n5108 & ~n5109 ;
  assign n5111 = ~n2731 & ~n5110 ;
  assign n5112 = n2731 & ~n3105 ;
  assign n5113 = ~n5111 & ~n5112 ;
  assign n5114 = n2717 & ~n5113 ;
  assign n5115 = ~n5107 & ~n5114 ;
  assign n5116 = n4025 & ~n5115 ;
  assign n5150 = n2964 & ~n5088 ;
  assign n5151 = ~n4054 & ~n5150 ;
  assign n5152 = n2717 & n5151 ;
  assign n5153 = ~n5107 & ~n5152 ;
  assign n5154 = n4062 & ~n5153 ;
  assign n5156 = n2964 & n4028 ;
  assign n5157 = n2717 & n5156 ;
  assign n5147 = ~n2717 & n4028 ;
  assign n5148 = ~n4067 & ~n5147 ;
  assign n5149 = \P1_reg2_reg[25]/NET0131  & ~n5148 ;
  assign n5155 = n2970 & n4073 ;
  assign n5158 = ~n5149 & ~n5155 ;
  assign n5159 = ~n5157 & n5158 ;
  assign n5160 = ~n5154 & n5159 ;
  assign n5161 = ~n5116 & n5160 ;
  assign n5117 = ~n2975 & ~n3190 ;
  assign n5118 = n3539 & n3745 ;
  assign n5119 = ~n3309 & n3744 ;
  assign n5120 = n3756 & ~n5119 ;
  assign n5121 = n3643 & ~n5120 ;
  assign n5122 = n3767 & ~n5121 ;
  assign n5123 = ~n5118 & n5122 ;
  assign n5124 = n3772 & ~n5123 ;
  assign n5125 = n3186 & ~n5124 ;
  assign n5126 = n5117 & n5125 ;
  assign n5127 = ~n5117 & ~n5125 ;
  assign n5128 = ~n5126 & ~n5127 ;
  assign n5129 = n2717 & ~n5128 ;
  assign n5130 = ~n5107 & ~n5129 ;
  assign n5131 = n3829 & ~n5130 ;
  assign n5132 = n3917 & n3920 ;
  assign n5133 = n3883 & n5132 ;
  assign n5134 = ~n3844 & n3920 ;
  assign n5135 = n3898 & ~n5134 ;
  assign n5136 = n3917 & ~n5135 ;
  assign n5137 = n3912 & ~n5136 ;
  assign n5138 = ~n5133 & n5137 ;
  assign n5139 = n3937 & ~n5138 ;
  assign n5140 = n3950 & ~n5139 ;
  assign n5141 = n5117 & ~n5140 ;
  assign n5142 = ~n5117 & n5140 ;
  assign n5143 = ~n5141 & ~n5142 ;
  assign n5144 = n2717 & ~n5143 ;
  assign n5145 = ~n5107 & ~n5144 ;
  assign n5146 = n3969 & ~n5145 ;
  assign n5162 = ~n5131 & ~n5146 ;
  assign n5163 = n5161 & n5162 ;
  assign n5164 = n2701 & ~n5163 ;
  assign n5165 = ~n5106 & ~n5164 ;
  assign n5166 = \P1_state_reg[0]/NET0131  & ~n5165 ;
  assign n5167 = ~n5105 & ~n5166 ;
  assign n5168 = \P2_reg2_reg[17]/NET0131  & ~n2286 ;
  assign n5169 = \P2_reg2_reg[17]/NET0131  & n2035 ;
  assign n5174 = \P2_reg2_reg[17]/NET0131  & ~n2291 ;
  assign n5175 = n2291 & n4353 ;
  assign n5176 = ~n5174 & ~n5175 ;
  assign n5177 = ~n2392 & ~n5176 ;
  assign n5170 = \P2_reg2_reg[17]/NET0131  & ~n2310 ;
  assign n5171 = n2310 & ~n4373 ;
  assign n5172 = ~n5170 & ~n5171 ;
  assign n5173 = n1790 & ~n5172 ;
  assign n5184 = ~n1221 & n2272 ;
  assign n5185 = n2291 & n5184 ;
  assign n5186 = \P2_reg2_reg[17]/NET0131  & ~n2407 ;
  assign n5187 = ~n1188 & n1854 ;
  assign n5188 = ~n5186 & ~n5187 ;
  assign n5189 = ~n5185 & n5188 ;
  assign n5190 = ~n5173 & n5189 ;
  assign n5191 = ~n5177 & n5190 ;
  assign n5178 = n2310 & ~n4365 ;
  assign n5179 = ~n5170 & ~n5178 ;
  assign n5180 = n2314 & ~n5179 ;
  assign n5181 = n2291 & ~n4365 ;
  assign n5182 = ~n5174 & ~n5181 ;
  assign n5183 = ~n2290 & ~n5182 ;
  assign n5192 = ~n5180 & ~n5183 ;
  assign n5193 = n5191 & n5192 ;
  assign n5194 = n2037 & ~n5193 ;
  assign n5195 = ~n5169 & ~n5194 ;
  assign n5196 = \P1_state_reg[0]/NET0131  & ~n5195 ;
  assign n5197 = ~n5168 & ~n5196 ;
  assign n5198 = \P2_reg2_reg[18]/NET0131  & ~n2286 ;
  assign n5199 = \P2_reg2_reg[18]/NET0131  & n2035 ;
  assign n5200 = \P2_reg2_reg[18]/NET0131  & ~n2310 ;
  assign n5201 = n2310 & ~n4268 ;
  assign n5202 = ~n5200 & ~n5201 ;
  assign n5203 = n1790 & ~n5202 ;
  assign n5214 = ~n1334 & n2272 ;
  assign n5215 = n2291 & n5214 ;
  assign n5216 = ~n1304 & n1854 ;
  assign n5217 = \P2_reg2_reg[18]/NET0131  & ~n2407 ;
  assign n5218 = ~n5216 & ~n5217 ;
  assign n5219 = ~n5215 & n5218 ;
  assign n5220 = ~n5203 & n5219 ;
  assign n5211 = n2310 & ~n4289 ;
  assign n5212 = ~n5200 & ~n5211 ;
  assign n5213 = n2314 & ~n5212 ;
  assign n5204 = \P2_reg2_reg[18]/NET0131  & ~n2291 ;
  assign n5205 = n2291 & n4253 ;
  assign n5206 = ~n5204 & ~n5205 ;
  assign n5207 = ~n2392 & ~n5206 ;
  assign n5208 = n2291 & ~n4289 ;
  assign n5209 = ~n5204 & ~n5208 ;
  assign n5210 = ~n2290 & ~n5209 ;
  assign n5221 = ~n5207 & ~n5210 ;
  assign n5222 = ~n5213 & n5221 ;
  assign n5223 = n5220 & n5222 ;
  assign n5224 = n2037 & ~n5223 ;
  assign n5225 = ~n5199 & ~n5224 ;
  assign n5226 = \P1_state_reg[0]/NET0131  & ~n5225 ;
  assign n5227 = ~n5198 & ~n5226 ;
  assign n5228 = \P2_reg2_reg[19]/NET0131  & ~n2286 ;
  assign n5229 = \P2_reg2_reg[19]/NET0131  & n2035 ;
  assign n5230 = \P2_reg2_reg[19]/NET0131  & ~n2310 ;
  assign n5231 = n2310 & ~n4321 ;
  assign n5232 = ~n5230 & ~n5231 ;
  assign n5233 = n1790 & ~n5232 ;
  assign n5244 = ~n1299 & n2272 ;
  assign n5245 = n2291 & n5244 ;
  assign n5246 = ~n1264 & n1854 ;
  assign n5247 = \P2_reg2_reg[19]/NET0131  & ~n2407 ;
  assign n5248 = ~n5246 & ~n5247 ;
  assign n5249 = ~n5245 & n5248 ;
  assign n5250 = ~n5233 & n5249 ;
  assign n5237 = \P2_reg2_reg[19]/NET0131  & ~n2291 ;
  assign n5241 = n2291 & ~n4311 ;
  assign n5242 = ~n5237 & ~n5241 ;
  assign n5243 = ~n2392 & ~n5242 ;
  assign n5234 = n2310 & n4330 ;
  assign n5235 = ~n5230 & ~n5234 ;
  assign n5236 = n2314 & ~n5235 ;
  assign n5238 = n2291 & n4330 ;
  assign n5239 = ~n5237 & ~n5238 ;
  assign n5240 = ~n2290 & ~n5239 ;
  assign n5251 = ~n5236 & ~n5240 ;
  assign n5252 = ~n5243 & n5251 ;
  assign n5253 = n5250 & n5252 ;
  assign n5254 = n2037 & ~n5253 ;
  assign n5255 = ~n5229 & ~n5254 ;
  assign n5256 = \P1_state_reg[0]/NET0131  & ~n5255 ;
  assign n5257 = ~n5228 & ~n5256 ;
  assign n5260 = ~n1406 & n2035 ;
  assign n5262 = ~n1406 & ~n2124 ;
  assign n5263 = n2124 & ~n4912 ;
  assign n5264 = ~n5262 & ~n5263 ;
  assign n5265 = n2123 & ~n5264 ;
  assign n5261 = n1401 & n2229 ;
  assign n5276 = ~n1406 & ~n2274 ;
  assign n5277 = ~n5261 & ~n5276 ;
  assign n5278 = ~n5265 & n5277 ;
  assign n5273 = n2124 & ~n4905 ;
  assign n5274 = ~n5262 & ~n5273 ;
  assign n5275 = n1790 & ~n5274 ;
  assign n5266 = ~n1406 & ~n2053 ;
  assign n5267 = n2053 & ~n4912 ;
  assign n5268 = ~n5266 & ~n5267 ;
  assign n5269 = ~n2224 & ~n5268 ;
  assign n5270 = n2053 & ~n4918 ;
  assign n5271 = ~n5266 & ~n5270 ;
  assign n5272 = ~n2120 & ~n5271 ;
  assign n5279 = ~n5269 & ~n5272 ;
  assign n5280 = ~n5275 & n5279 ;
  assign n5281 = n5278 & n5280 ;
  assign n5282 = n2037 & ~n5281 ;
  assign n5283 = ~n5260 & ~n5282 ;
  assign n5284 = \P1_state_reg[0]/NET0131  & ~n5283 ;
  assign n5258 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[20]/NET0131  ;
  assign n5259 = ~n1406 & n2014 ;
  assign n5285 = ~n5258 & ~n5259 ;
  assign n5286 = ~n5284 & n5285 ;
  assign n5287 = \P1_B_reg/NET0131  & ~n4552 ;
  assign n5288 = \P1_B_reg/NET0131  & n2683 ;
  assign n5297 = n3891 & ~n4746 ;
  assign n5298 = n4745 & ~n5297 ;
  assign n5299 = ~n3895 & ~n5298 ;
  assign n5300 = n3837 & ~n4734 ;
  assign n5301 = n4735 & ~n5300 ;
  assign n5302 = ~n3841 & ~n5301 ;
  assign n5303 = ~n5299 & ~n5302 ;
  assign n5304 = n4755 & ~n5303 ;
  assign n5305 = ~n3404 & n3411 ;
  assign n5306 = ~n3849 & n5305 ;
  assign n5307 = n3853 & ~n5306 ;
  assign n5308 = n3857 & ~n5307 ;
  assign n5309 = n3847 & ~n5308 ;
  assign n5310 = n3863 & ~n5309 ;
  assign n5311 = n3868 & ~n5310 ;
  assign n5312 = n4719 & ~n5311 ;
  assign n5313 = ~n3876 & n4738 ;
  assign n5314 = n4741 & n5313 ;
  assign n5315 = n4750 & n5314 ;
  assign n5316 = n4753 & n5315 ;
  assign n5317 = ~n5312 & n5316 ;
  assign n5318 = ~n5304 & ~n5317 ;
  assign n5294 = n3910 & ~n3942 ;
  assign n5295 = n4776 & n5294 ;
  assign n5319 = ~n3903 & n4757 ;
  assign n5320 = n5295 & n5319 ;
  assign n5321 = ~n5318 & n5320 ;
  assign n5289 = n3943 & ~n4765 ;
  assign n5290 = n4766 & ~n5289 ;
  assign n5291 = ~n3947 & ~n5290 ;
  assign n5292 = n3905 & ~n4716 ;
  assign n5293 = n4717 & ~n5292 ;
  assign n5296 = ~n5293 & n5295 ;
  assign n5322 = ~n5291 & ~n5296 ;
  assign n5323 = ~n5321 & n5322 ;
  assign n5324 = n4780 & n4781 ;
  assign n5325 = ~n5323 & n5324 ;
  assign n5326 = n3954 & ~n4768 ;
  assign n5327 = n4769 & ~n5326 ;
  assign n5328 = ~n3958 & ~n5327 ;
  assign n5329 = ~n5325 & ~n5328 ;
  assign n5330 = ~n3803 & ~n3957 ;
  assign n5332 = ~\P2_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n5333 = ~n2734 & ~n3779 ;
  assign n5334 = ~n2836 & n5333 ;
  assign n5335 = ~n5332 & n5334 ;
  assign n5336 = n3034 & n5335 ;
  assign n5337 = ~n3113 & n5336 ;
  assign n5338 = ~n3033 & n5335 ;
  assign n5331 = \P2_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n5339 = ~n3781 & n5333 ;
  assign n5340 = ~n3778 & ~n5339 ;
  assign n5341 = ~n5332 & ~n5340 ;
  assign n5342 = ~n5331 & ~n5341 ;
  assign n5343 = ~n5338 & n5342 ;
  assign n5344 = ~n5337 & n5343 ;
  assign n5346 = ~\si[31]_pad  & n5344 ;
  assign n5345 = \si[31]_pad  & ~n5344 ;
  assign n5347 = ~n639 & ~n5345 ;
  assign n5348 = ~n5346 & n5347 ;
  assign n5349 = \P2_datao_reg[31]/NET0131  & n5348 ;
  assign n5350 = ~\P2_datao_reg[31]/NET0131  & ~n5348 ;
  assign n5351 = ~n5349 & ~n5350 ;
  assign n5352 = ~n2732 & n5351 ;
  assign n5353 = n3984 & n5352 ;
  assign n5354 = \P2_datao_reg[30]/NET0131  & n639 ;
  assign n5355 = ~n5331 & ~n5332 ;
  assign n5357 = ~n2831 & n5334 ;
  assign n5360 = n3007 & n5357 ;
  assign n5361 = ~n3137 & n5360 ;
  assign n5358 = ~n3010 & n5357 ;
  assign n5359 = ~n2843 & n5334 ;
  assign n5356 = n2735 & ~n3779 ;
  assign n5362 = ~n3778 & ~n5356 ;
  assign n5363 = ~n5359 & n5362 ;
  assign n5364 = ~n5358 & n5363 ;
  assign n5365 = ~n5361 & n5364 ;
  assign n5367 = ~n5355 & n5365 ;
  assign n5366 = n5355 & ~n5365 ;
  assign n5368 = ~n639 & ~n5366 ;
  assign n5369 = ~n5367 & n5368 ;
  assign n5370 = ~n5354 & ~n5369 ;
  assign n5371 = ~n2732 & ~n5370 ;
  assign n5372 = ~n4015 & ~n5371 ;
  assign n5373 = ~n5353 & ~n5372 ;
  assign n5374 = n5330 & n5373 ;
  assign n5375 = ~n5329 & n5374 ;
  assign n5376 = ~n3984 & ~n5352 ;
  assign n5377 = n4015 & n5371 ;
  assign n5378 = ~n5376 & ~n5377 ;
  assign n5379 = ~n3802 & ~n3925 ;
  assign n5380 = ~n3803 & ~n5372 ;
  assign n5381 = ~n5379 & n5380 ;
  assign n5382 = n5378 & ~n5381 ;
  assign n5383 = ~n5353 & ~n5382 ;
  assign n5384 = ~n5375 & ~n5383 ;
  assign n5385 = ~n5288 & ~n5384 ;
  assign n5386 = n4068 & ~n5385 ;
  assign n5387 = ~n5288 & n5384 ;
  assign n5388 = n4066 & ~n5387 ;
  assign n5389 = ~n5386 & ~n5388 ;
  assign n5390 = n3813 & ~n5389 ;
  assign n5391 = n5378 & n5379 ;
  assign n5392 = ~n4762 & n4767 ;
  assign n5393 = n4778 & ~n5392 ;
  assign n5394 = n4770 & ~n5393 ;
  assign n5395 = ~n4785 & ~n5394 ;
  assign n5396 = n5391 & ~n5395 ;
  assign n5397 = ~n3802 & ~n5330 ;
  assign n5398 = ~n5377 & n5397 ;
  assign n5399 = n5373 & ~n5398 ;
  assign n5400 = ~n5376 & ~n5399 ;
  assign n5401 = n4771 & n5391 ;
  assign n5402 = n5048 & n5401 ;
  assign n5403 = ~n5400 & ~n5402 ;
  assign n5404 = ~n5396 & n5403 ;
  assign n5405 = n4068 & ~n5404 ;
  assign n5406 = ~n5288 & ~n5405 ;
  assign n5407 = ~n3813 & ~n5406 ;
  assign n5408 = ~n3813 & n4066 ;
  assign n5409 = n5404 & n5408 ;
  assign n5461 = n3804 & n5373 ;
  assign n5462 = n5378 & n5461 ;
  assign n5433 = ~n3178 & ~n3770 ;
  assign n5417 = ~n3129 & ~n3183 ;
  assign n5432 = ~n3562 & ~n3763 ;
  assign n5451 = ~n5417 & ~n5432 ;
  assign n5452 = ~n5433 & n5451 ;
  assign n5458 = ~n4709 & n5452 ;
  assign n5459 = ~n4958 & n5458 ;
  assign n5412 = ~n3900 & ~n3909 ;
  assign n5410 = ~n3154 & ~n3155 ;
  assign n5455 = ~n5117 & ~n5410 ;
  assign n5456 = n5412 & n5455 ;
  assign n5425 = ~n3718 & ~n3752 ;
  assign n5418 = ~n3742 & ~n3753 ;
  assign n5423 = ~n3614 & ~n3759 ;
  assign n5448 = ~n5418 & ~n5423 ;
  assign n5449 = ~n5425 & n5448 ;
  assign n5419 = ~n3249 & ~n3305 ;
  assign n5413 = ~n3666 & ~n3747 ;
  assign n5420 = ~n3445 & ~n3530 ;
  assign n5414 = ~n3276 & ~n3277 ;
  assign n5415 = ~n3848 & ~n5305 ;
  assign n5416 = ~n3845 & ~n3861 ;
  assign n5434 = n5415 & n5416 ;
  assign n5440 = ~n5414 & n5434 ;
  assign n5441 = ~n5420 & n5440 ;
  assign n5445 = ~n5413 & n5441 ;
  assign n5446 = ~n5419 & n5445 ;
  assign n5411 = ~n3641 & ~n3758 ;
  assign n5431 = ~n3495 & ~n3525 ;
  assign n5428 = ~n3471 & ~n3531 ;
  assign n5429 = ~n3852 & ~n3855 ;
  assign n5437 = ~n5428 & n5429 ;
  assign n5438 = ~n5431 & n5437 ;
  assign n5421 = ~n3835 & ~n3880 ;
  assign n5422 = ~n3521 & ~n3526 ;
  assign n5435 = n5421 & ~n5422 ;
  assign n5426 = ~n3372 & ~n3418 ;
  assign n5427 = ~n3849 & ~n3851 ;
  assign n5436 = ~n5426 & n5427 ;
  assign n5439 = n5435 & n5436 ;
  assign n5442 = n5438 & n5439 ;
  assign n5424 = ~n3831 & ~n3841 ;
  assign n5430 = ~n3693 & ~n3748 ;
  assign n5443 = n5424 & ~n5430 ;
  assign n5444 = n5442 & n5443 ;
  assign n5447 = ~n5411 & n5444 ;
  assign n5450 = n5446 & n5447 ;
  assign n5453 = n5449 & n5450 ;
  assign n5454 = ~n4451 & ~n5046 ;
  assign n5457 = n5453 & n5454 ;
  assign n5460 = n5456 & n5457 ;
  assign n5463 = n5459 & n5460 ;
  assign n5464 = n5462 & n5463 ;
  assign n5466 = ~n3826 & n5464 ;
  assign n5465 = n3826 & ~n5464 ;
  assign n5467 = n4027 & ~n5465 ;
  assign n5468 = ~n5466 & n5467 ;
  assign n5488 = ~n5409 & ~n5468 ;
  assign n5489 = ~n5407 & n5488 ;
  assign n5469 = ~n3984 & ~n4015 ;
  assign n5470 = n5371 & ~n5469 ;
  assign n5471 = ~n5376 & ~n5470 ;
  assign n5473 = n5379 & n5471 ;
  assign n5477 = n4770 & n5473 ;
  assign n5478 = ~n5051 & n5477 ;
  assign n5474 = n4785 & n5473 ;
  assign n5472 = n5397 & n5471 ;
  assign n5475 = ~n3984 & ~n5372 ;
  assign n5476 = n5352 & ~n5475 ;
  assign n5479 = ~n5472 & ~n5476 ;
  assign n5480 = ~n5474 & n5479 ;
  assign n5481 = ~n5478 & n5480 ;
  assign n5482 = ~\P1_B_reg/NET0131  & n5481 ;
  assign n5483 = n3822 & n3827 ;
  assign n5484 = ~n5482 & n5483 ;
  assign n5485 = ~\P1_B_reg/NET0131  & ~n5481 ;
  assign n5486 = n3822 & n4023 ;
  assign n5487 = ~n5485 & n5486 ;
  assign n5490 = ~n5484 & ~n5487 ;
  assign n5491 = n5489 & n5490 ;
  assign n5492 = ~n5390 & n5491 ;
  assign n5493 = n4552 & ~n5492 ;
  assign n5494 = ~n5287 & ~n5493 ;
  assign n5495 = n2900 & n4081 ;
  assign n5496 = n2900 & ~n4449 ;
  assign n5497 = n4449 & ~n4712 ;
  assign n5498 = ~n5496 & ~n5497 ;
  assign n5499 = n3829 & ~n5498 ;
  assign n5500 = n4449 & ~n4790 ;
  assign n5501 = ~n5496 & ~n5500 ;
  assign n5502 = n3969 & ~n5501 ;
  assign n5506 = n4449 & n4797 ;
  assign n5503 = n4449 & n4804 ;
  assign n5504 = ~n5496 & ~n5503 ;
  assign n5505 = n4025 & ~n5504 ;
  assign n5507 = n2868 & ~n4522 ;
  assign n5508 = n2900 & ~n4542 ;
  assign n5509 = ~n5507 & ~n5508 ;
  assign n5510 = ~n5505 & n5509 ;
  assign n5511 = ~n5506 & n5510 ;
  assign n5512 = ~n5502 & n5511 ;
  assign n5513 = ~n5499 & n5512 ;
  assign n5514 = n2701 & ~n5513 ;
  assign n5515 = ~n5495 & ~n5514 ;
  assign n5516 = \P1_state_reg[0]/NET0131  & ~n5515 ;
  assign n5517 = \P1_reg3_reg[28]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5518 = n2900 & n4552 ;
  assign n5519 = ~n5517 & ~n5518 ;
  assign n5520 = ~n5516 & n5519 ;
  assign n5523 = ~n1521 & n2035 ;
  assign n5524 = ~n1521 & ~n2053 ;
  assign n5525 = n2053 & ~n4131 ;
  assign n5526 = ~n5524 & ~n5525 ;
  assign n5527 = ~n2120 & ~n5526 ;
  assign n5531 = ~n1521 & ~n2124 ;
  assign n5536 = n2124 & ~n4159 ;
  assign n5537 = ~n5531 & ~n5536 ;
  assign n5538 = n1790 & ~n5537 ;
  assign n5535 = n1513 & n2229 ;
  assign n5539 = ~n1521 & ~n2274 ;
  assign n5540 = ~n5535 & ~n5539 ;
  assign n5541 = ~n5538 & n5540 ;
  assign n5542 = ~n5527 & n5541 ;
  assign n5528 = n2053 & ~n4145 ;
  assign n5529 = ~n5524 & ~n5528 ;
  assign n5530 = ~n2224 & ~n5529 ;
  assign n5532 = n2124 & ~n4145 ;
  assign n5533 = ~n5531 & ~n5532 ;
  assign n5534 = n2123 & ~n5533 ;
  assign n5543 = ~n5530 & ~n5534 ;
  assign n5544 = n5542 & n5543 ;
  assign n5545 = n2037 & ~n5544 ;
  assign n5546 = ~n5523 & ~n5545 ;
  assign n5547 = \P1_state_reg[0]/NET0131  & ~n5546 ;
  assign n5521 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[25]/NET0131  ;
  assign n5522 = ~n1521 & n2014 ;
  assign n5548 = ~n5521 & ~n5522 ;
  assign n5549 = ~n5547 & n5548 ;
  assign n5550 = ~n1583 & n2035 ;
  assign n5551 = ~n1583 & ~n2124 ;
  assign n5552 = ~n1942 & n2194 ;
  assign n5553 = n4394 & n5552 ;
  assign n5554 = ~n4250 & n5553 ;
  assign n5556 = ~n4393 & n5552 ;
  assign n5555 = n2364 & ~n2377 ;
  assign n5557 = n2381 & ~n5555 ;
  assign n5558 = ~n5556 & n5557 ;
  assign n5559 = ~n5554 & n5558 ;
  assign n5560 = n1885 & n5559 ;
  assign n5561 = ~n1885 & ~n5559 ;
  assign n5562 = ~n5560 & ~n5561 ;
  assign n5563 = n2124 & ~n5562 ;
  assign n5564 = ~n5551 & ~n5563 ;
  assign n5565 = n2123 & ~n5564 ;
  assign n5566 = ~n1525 & ~n2263 ;
  assign n5567 = n1618 & ~n4155 ;
  assign n5568 = ~n2258 & n2263 ;
  assign n5569 = ~n5567 & n5568 ;
  assign n5570 = ~n5566 & ~n5569 ;
  assign n5571 = n2124 & ~n5570 ;
  assign n5572 = ~n5551 & ~n5571 ;
  assign n5573 = n1790 & ~n5572 ;
  assign n5574 = n1573 & n2229 ;
  assign n5575 = ~n1583 & ~n2274 ;
  assign n5594 = ~n5574 & ~n5575 ;
  assign n5595 = ~n5573 & n5594 ;
  assign n5596 = ~n5565 & n5595 ;
  assign n5576 = ~n1583 & ~n2053 ;
  assign n5577 = n2053 & ~n5562 ;
  assign n5578 = ~n5576 & ~n5577 ;
  assign n5579 = ~n2224 & ~n5578 ;
  assign n5580 = n1481 & n1628 ;
  assign n5581 = n4421 & n5580 ;
  assign n5582 = ~n4286 & n5581 ;
  assign n5584 = ~n4420 & n5580 ;
  assign n5583 = n1628 & n1835 ;
  assign n5585 = ~n1840 & ~n5583 ;
  assign n5586 = ~n5584 & n5585 ;
  assign n5587 = ~n5582 & n5586 ;
  assign n5588 = n1885 & ~n5587 ;
  assign n5589 = ~n1885 & n5587 ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5591 = n2053 & ~n5590 ;
  assign n5592 = ~n5576 & ~n5591 ;
  assign n5593 = ~n2120 & ~n5592 ;
  assign n5597 = ~n5579 & ~n5593 ;
  assign n5598 = n5596 & n5597 ;
  assign n5599 = n2037 & ~n5598 ;
  assign n5600 = ~n5550 & ~n5599 ;
  assign n5601 = \P1_state_reg[0]/NET0131  & ~n5600 ;
  assign n5602 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[26]/NET0131  ;
  assign n5603 = ~n1583 & n2014 ;
  assign n5604 = ~n5602 & ~n5603 ;
  assign n5605 = ~n5601 & n5604 ;
  assign n5606 = \P2_reg2_reg[21]/NET0131  & ~n2286 ;
  assign n5607 = \P2_reg2_reg[21]/NET0131  & n2035 ;
  assign n5608 = \P2_reg2_reg[21]/NET0131  & ~n2291 ;
  assign n5609 = n1935 & n2637 ;
  assign n5610 = ~n1935 & ~n2637 ;
  assign n5611 = ~n5609 & ~n5610 ;
  assign n5612 = n2291 & ~n5611 ;
  assign n5613 = ~n5608 & ~n5612 ;
  assign n5614 = ~n2392 & ~n5613 ;
  assign n5633 = n1371 & n2272 ;
  assign n5634 = n2291 & n5633 ;
  assign n5635 = ~n1378 & n1854 ;
  assign n5636 = \P2_reg2_reg[21]/NET0131  & ~n2407 ;
  assign n5637 = ~n5635 & ~n5636 ;
  assign n5638 = ~n5634 & n5637 ;
  assign n5639 = ~n5614 & n5638 ;
  assign n5621 = \P2_reg2_reg[21]/NET0131  & ~n2310 ;
  assign n5625 = n1474 & ~n4408 ;
  assign n5626 = n2263 & ~n4409 ;
  assign n5627 = ~n5625 & n5626 ;
  assign n5628 = ~n1410 & ~n2263 ;
  assign n5629 = ~n5627 & ~n5628 ;
  assign n5630 = n2310 & ~n5629 ;
  assign n5631 = ~n5621 & ~n5630 ;
  assign n5632 = n1790 & ~n5631 ;
  assign n5615 = n1935 & ~n2579 ;
  assign n5616 = ~n1935 & n2579 ;
  assign n5617 = ~n5615 & ~n5616 ;
  assign n5618 = n2291 & ~n5617 ;
  assign n5619 = ~n5608 & ~n5618 ;
  assign n5620 = ~n2290 & ~n5619 ;
  assign n5622 = n2310 & ~n5617 ;
  assign n5623 = ~n5621 & ~n5622 ;
  assign n5624 = n2314 & ~n5623 ;
  assign n5640 = ~n5620 & ~n5624 ;
  assign n5641 = ~n5632 & n5640 ;
  assign n5642 = n5639 & n5641 ;
  assign n5643 = n2037 & ~n5642 ;
  assign n5644 = ~n5607 & ~n5643 ;
  assign n5645 = \P1_state_reg[0]/NET0131  & ~n5644 ;
  assign n5646 = ~n5606 & ~n5645 ;
  assign n5647 = \P2_reg0_reg[24]/NET0131  & ~n2286 ;
  assign n5648 = \P2_reg0_reg[24]/NET0131  & n2035 ;
  assign n5649 = \P2_reg0_reg[24]/NET0131  & ~n2124 ;
  assign n5658 = n2124 & ~n2512 ;
  assign n5659 = ~n5649 & ~n5658 ;
  assign n5660 = ~n2120 & ~n5659 ;
  assign n5652 = \P2_reg0_reg[24]/NET0131  & ~n2053 ;
  assign n5656 = ~n2494 & ~n5652 ;
  assign n5657 = n2123 & ~n5656 ;
  assign n5650 = ~n2507 & ~n5649 ;
  assign n5651 = ~n2224 & ~n5650 ;
  assign n5653 = n2053 & ~n2503 ;
  assign n5654 = ~n5652 & ~n5653 ;
  assign n5655 = n1790 & ~n5654 ;
  assign n5661 = \P2_reg0_reg[24]/NET0131  & ~n2614 ;
  assign n5662 = n1540 & n2272 ;
  assign n5663 = n2124 & n5662 ;
  assign n5664 = ~n5661 & ~n5663 ;
  assign n5665 = ~n5655 & n5664 ;
  assign n5666 = ~n5651 & n5665 ;
  assign n5667 = ~n5657 & n5666 ;
  assign n5668 = ~n5660 & n5667 ;
  assign n5669 = n2037 & ~n5668 ;
  assign n5670 = ~n5648 & ~n5669 ;
  assign n5671 = \P1_state_reg[0]/NET0131  & ~n5670 ;
  assign n5672 = ~n5647 & ~n5671 ;
  assign n5673 = \P2_reg0_reg[25]/NET0131  & ~n2286 ;
  assign n5674 = \P2_reg0_reg[25]/NET0131  & n2035 ;
  assign n5675 = \P2_reg0_reg[25]/NET0131  & ~n2124 ;
  assign n5676 = n2124 & ~n4131 ;
  assign n5677 = ~n5675 & ~n5676 ;
  assign n5678 = ~n2120 & ~n5677 ;
  assign n5681 = \P2_reg0_reg[25]/NET0131  & ~n2053 ;
  assign n5686 = n2053 & ~n4159 ;
  assign n5687 = ~n5681 & ~n5686 ;
  assign n5688 = n1790 & ~n5687 ;
  assign n5684 = n1513 & n2272 ;
  assign n5685 = n2124 & n5684 ;
  assign n5689 = \P2_reg0_reg[25]/NET0131  & ~n2614 ;
  assign n5690 = ~n5685 & ~n5689 ;
  assign n5691 = ~n5688 & n5690 ;
  assign n5692 = ~n5678 & n5691 ;
  assign n5679 = ~n5532 & ~n5675 ;
  assign n5680 = ~n2224 & ~n5679 ;
  assign n5682 = ~n5528 & ~n5681 ;
  assign n5683 = n2123 & ~n5682 ;
  assign n5693 = ~n5680 & ~n5683 ;
  assign n5694 = n5692 & n5693 ;
  assign n5695 = n2037 & ~n5694 ;
  assign n5696 = ~n5674 & ~n5695 ;
  assign n5697 = \P1_state_reg[0]/NET0131  & ~n5696 ;
  assign n5698 = ~n5673 & ~n5697 ;
  assign n5699 = \P2_reg0_reg[26]/NET0131  & ~n2286 ;
  assign n5700 = \P2_reg0_reg[26]/NET0131  & n2035 ;
  assign n5701 = \P2_reg0_reg[26]/NET0131  & ~n2124 ;
  assign n5702 = n2124 & ~n5590 ;
  assign n5703 = ~n5701 & ~n5702 ;
  assign n5704 = ~n2120 & ~n5703 ;
  assign n5705 = \P2_reg0_reg[26]/NET0131  & ~n2053 ;
  assign n5706 = n2053 & ~n5570 ;
  assign n5707 = ~n5705 & ~n5706 ;
  assign n5708 = n1790 & ~n5707 ;
  assign n5709 = n1573 & n2616 ;
  assign n5710 = \P2_reg0_reg[26]/NET0131  & ~n2614 ;
  assign n5715 = ~n5709 & ~n5710 ;
  assign n5716 = ~n5708 & n5715 ;
  assign n5717 = ~n5704 & n5716 ;
  assign n5711 = ~n5577 & ~n5705 ;
  assign n5712 = n2123 & ~n5711 ;
  assign n5713 = ~n5563 & ~n5701 ;
  assign n5714 = ~n2224 & ~n5713 ;
  assign n5718 = ~n5712 & ~n5714 ;
  assign n5719 = n5717 & n5718 ;
  assign n5720 = n2037 & ~n5719 ;
  assign n5721 = ~n5700 & ~n5720 ;
  assign n5722 = \P1_state_reg[0]/NET0131  & ~n5721 ;
  assign n5723 = ~n5699 & ~n5722 ;
  assign n5724 = \P1_reg2_reg[27]/NET0131  & n4081 ;
  assign n5725 = \P1_reg2_reg[27]/NET0131  & ~n2717 ;
  assign n5726 = n2717 & ~n4485 ;
  assign n5727 = ~n5725 & ~n5726 ;
  assign n5728 = n3829 & ~n5727 ;
  assign n5729 = n2717 & ~n4517 ;
  assign n5730 = ~n5725 & ~n5729 ;
  assign n5731 = n3969 & ~n5730 ;
  assign n5733 = n3069 & n4028 ;
  assign n5734 = ~n4528 & ~n5733 ;
  assign n5735 = n2717 & ~n5734 ;
  assign n5736 = n2717 & ~n4535 ;
  assign n5737 = ~n5725 & ~n5736 ;
  assign n5738 = n4025 & ~n5737 ;
  assign n5732 = \P1_reg2_reg[27]/NET0131  & ~n4071 ;
  assign n5739 = n3074 & n4073 ;
  assign n5740 = ~n5732 & ~n5739 ;
  assign n5741 = ~n5738 & n5740 ;
  assign n5742 = ~n5735 & n5741 ;
  assign n5743 = ~n5731 & n5742 ;
  assign n5744 = ~n5728 & n5743 ;
  assign n5745 = n2701 & ~n5744 ;
  assign n5746 = ~n5724 & ~n5745 ;
  assign n5747 = \P1_state_reg[0]/NET0131  & ~n5746 ;
  assign n5748 = \P1_reg2_reg[27]/NET0131  & ~n4085 ;
  assign n5749 = ~n5747 & ~n5748 ;
  assign n5750 = \P2_reg1_reg[24]/NET0131  & ~n2286 ;
  assign n5751 = \P2_reg1_reg[24]/NET0131  & n2035 ;
  assign n5756 = \P2_reg1_reg[24]/NET0131  & ~n2291 ;
  assign n5757 = ~n2536 & ~n5756 ;
  assign n5758 = n2314 & ~n5757 ;
  assign n5753 = \P2_reg1_reg[24]/NET0131  & ~n2310 ;
  assign n5754 = ~n2532 & ~n5753 ;
  assign n5755 = ~n2290 & ~n5754 ;
  assign n5759 = n2310 & ~n2493 ;
  assign n5760 = ~n5753 & ~n5759 ;
  assign n5761 = ~n2392 & ~n5760 ;
  assign n5762 = n2291 & ~n2503 ;
  assign n5763 = ~n5756 & ~n5762 ;
  assign n5764 = n1790 & ~n5763 ;
  assign n5752 = n2310 & n5662 ;
  assign n5765 = \P2_reg1_reg[24]/NET0131  & ~n4099 ;
  assign n5766 = ~n5752 & ~n5765 ;
  assign n5767 = ~n5764 & n5766 ;
  assign n5768 = ~n5761 & n5767 ;
  assign n5769 = ~n5755 & n5768 ;
  assign n5770 = ~n5758 & n5769 ;
  assign n5771 = n2037 & ~n5770 ;
  assign n5772 = ~n5751 & ~n5771 ;
  assign n5773 = \P1_state_reg[0]/NET0131  & ~n5772 ;
  assign n5774 = ~n5750 & ~n5773 ;
  assign n5775 = \P2_reg1_reg[26]/NET0131  & ~n2286 ;
  assign n5776 = \P2_reg1_reg[26]/NET0131  & n2035 ;
  assign n5777 = \P2_reg1_reg[26]/NET0131  & ~n2310 ;
  assign n5778 = n2310 & ~n5590 ;
  assign n5779 = ~n5777 & ~n5778 ;
  assign n5780 = ~n2290 & ~n5779 ;
  assign n5781 = \P2_reg1_reg[26]/NET0131  & ~n2291 ;
  assign n5782 = n2291 & ~n5570 ;
  assign n5783 = ~n5781 & ~n5782 ;
  assign n5784 = n1790 & ~n5783 ;
  assign n5785 = n1573 & n4101 ;
  assign n5786 = \P2_reg1_reg[26]/NET0131  & ~n4099 ;
  assign n5793 = ~n5785 & ~n5786 ;
  assign n5794 = ~n5784 & n5793 ;
  assign n5795 = ~n5780 & n5794 ;
  assign n5787 = n2291 & ~n5590 ;
  assign n5788 = ~n5781 & ~n5787 ;
  assign n5789 = n2314 & ~n5788 ;
  assign n5790 = n2310 & ~n5562 ;
  assign n5791 = ~n5777 & ~n5790 ;
  assign n5792 = ~n2392 & ~n5791 ;
  assign n5796 = ~n5789 & ~n5792 ;
  assign n5797 = n5795 & n5796 ;
  assign n5798 = n2037 & ~n5797 ;
  assign n5799 = ~n5776 & ~n5798 ;
  assign n5800 = \P1_state_reg[0]/NET0131  & ~n5799 ;
  assign n5801 = ~n5775 & ~n5800 ;
  assign n5802 = \P2_reg1_reg[25]/NET0131  & ~n2286 ;
  assign n5803 = \P2_reg1_reg[25]/NET0131  & n2035 ;
  assign n5804 = \P2_reg1_reg[25]/NET0131  & ~n2310 ;
  assign n5805 = ~n4150 & ~n5804 ;
  assign n5806 = ~n2290 & ~n5805 ;
  assign n5810 = \P2_reg1_reg[25]/NET0131  & ~n2291 ;
  assign n5814 = n2291 & ~n4159 ;
  assign n5815 = ~n5810 & ~n5814 ;
  assign n5816 = n1790 & ~n5815 ;
  assign n5813 = n2310 & n5684 ;
  assign n5817 = \P2_reg1_reg[25]/NET0131  & ~n4099 ;
  assign n5818 = ~n5813 & ~n5817 ;
  assign n5819 = ~n5816 & n5818 ;
  assign n5820 = ~n5806 & n5819 ;
  assign n5807 = n2310 & ~n4145 ;
  assign n5808 = ~n5804 & ~n5807 ;
  assign n5809 = ~n2392 & ~n5808 ;
  assign n5811 = ~n4132 & ~n5810 ;
  assign n5812 = n2314 & ~n5811 ;
  assign n5821 = ~n5809 & ~n5812 ;
  assign n5822 = n5820 & n5821 ;
  assign n5823 = n2037 & ~n5822 ;
  assign n5824 = ~n5803 & ~n5823 ;
  assign n5825 = \P1_state_reg[0]/NET0131  & ~n5824 ;
  assign n5826 = ~n5802 & ~n5825 ;
  assign n5827 = \P1_reg0_reg[26]/NET0131  & ~n4085 ;
  assign n5828 = \P1_reg0_reg[26]/NET0131  & n4081 ;
  assign n5829 = \P1_reg0_reg[26]/NET0131  & ~n4869 ;
  assign n5830 = n4869 & n4954 ;
  assign n5831 = ~n5829 & ~n5830 ;
  assign n5832 = n4025 & ~n5831 ;
  assign n5839 = n3017 & n4028 ;
  assign n5840 = n4062 & n5030 ;
  assign n5841 = ~n5839 & ~n5840 ;
  assign n5842 = n4869 & ~n5841 ;
  assign n5843 = n4069 & ~n4869 ;
  assign n5844 = n4214 & ~n5843 ;
  assign n5845 = \P1_reg0_reg[26]/NET0131  & ~n5844 ;
  assign n5846 = ~n5842 & ~n5845 ;
  assign n5847 = ~n5832 & n5846 ;
  assign n5833 = n4869 & ~n5024 ;
  assign n5834 = ~n5829 & ~n5833 ;
  assign n5835 = n3829 & ~n5834 ;
  assign n5836 = n4869 & ~n4990 ;
  assign n5837 = ~n5829 & ~n5836 ;
  assign n5838 = n3969 & ~n5837 ;
  assign n5848 = ~n5835 & ~n5838 ;
  assign n5849 = n5847 & n5848 ;
  assign n5850 = n2701 & ~n5849 ;
  assign n5851 = ~n5828 & ~n5850 ;
  assign n5852 = \P1_state_reg[0]/NET0131  & ~n5851 ;
  assign n5853 = ~n5827 & ~n5852 ;
  assign n5854 = \P1_reg0_reg[27]/NET0131  & n4081 ;
  assign n5855 = \P1_reg0_reg[27]/NET0131  & ~n4869 ;
  assign n5856 = ~n4485 & n4869 ;
  assign n5857 = ~n5855 & ~n5856 ;
  assign n5858 = n3829 & ~n5857 ;
  assign n5859 = ~n4517 & n4869 ;
  assign n5860 = ~n5855 & ~n5859 ;
  assign n5861 = n3969 & ~n5860 ;
  assign n5862 = n4869 & ~n5734 ;
  assign n5863 = n4028 & ~n4869 ;
  assign n5864 = n4214 & ~n5863 ;
  assign n5865 = n4062 & ~n4869 ;
  assign n5866 = n5864 & ~n5865 ;
  assign n5867 = \P1_reg0_reg[27]/NET0131  & ~n5866 ;
  assign n5868 = ~n4535 & n4869 ;
  assign n5869 = ~n5855 & ~n5868 ;
  assign n5870 = n4025 & ~n5869 ;
  assign n5871 = ~n5867 & ~n5870 ;
  assign n5872 = ~n5862 & n5871 ;
  assign n5873 = ~n5861 & n5872 ;
  assign n5874 = ~n5858 & n5873 ;
  assign n5875 = n2701 & ~n5874 ;
  assign n5876 = ~n5854 & ~n5875 ;
  assign n5877 = \P1_state_reg[0]/NET0131  & ~n5876 ;
  assign n5878 = \P1_reg0_reg[27]/NET0131  & ~n4085 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = \P1_reg0_reg[28]/NET0131  & ~n4085 ;
  assign n5881 = \P1_reg0_reg[28]/NET0131  & n4081 ;
  assign n5882 = \P1_reg0_reg[28]/NET0131  & ~n4869 ;
  assign n5883 = ~n4712 & n4869 ;
  assign n5884 = ~n5882 & ~n5883 ;
  assign n5885 = n3829 & ~n5884 ;
  assign n5886 = ~n4790 & n4869 ;
  assign n5887 = ~n5882 & ~n5886 ;
  assign n5888 = n3969 & ~n5887 ;
  assign n5889 = ~n4798 & n4869 ;
  assign n5890 = \P1_reg0_reg[28]/NET0131  & ~n5866 ;
  assign n5891 = n4804 & n4869 ;
  assign n5892 = ~n5882 & ~n5891 ;
  assign n5893 = n4025 & ~n5892 ;
  assign n5894 = ~n5890 & ~n5893 ;
  assign n5895 = ~n5889 & n5894 ;
  assign n5896 = ~n5888 & n5895 ;
  assign n5897 = ~n5885 & n5896 ;
  assign n5898 = n2701 & ~n5897 ;
  assign n5899 = ~n5881 & ~n5898 ;
  assign n5900 = \P1_state_reg[0]/NET0131  & ~n5899 ;
  assign n5901 = ~n5880 & ~n5900 ;
  assign n5902 = \P1_reg1_reg[27]/NET0131  & ~n4085 ;
  assign n5903 = \P1_reg1_reg[27]/NET0131  & ~n4202 ;
  assign n5904 = n4202 & ~n4485 ;
  assign n5905 = ~n5903 & ~n5904 ;
  assign n5906 = n3829 & ~n5905 ;
  assign n5907 = n4202 & ~n4517 ;
  assign n5908 = ~n5903 & ~n5907 ;
  assign n5909 = n3969 & ~n5908 ;
  assign n5911 = n4202 & n4527 ;
  assign n5912 = ~n5903 & ~n5911 ;
  assign n5913 = n4062 & ~n5912 ;
  assign n5914 = n4202 & ~n4535 ;
  assign n5915 = ~n5903 & ~n5914 ;
  assign n5916 = n4025 & ~n5915 ;
  assign n5910 = \P1_reg1_reg[27]/NET0131  & ~n4216 ;
  assign n5917 = n4202 & n5733 ;
  assign n5918 = ~n5910 & ~n5917 ;
  assign n5919 = ~n5916 & n5918 ;
  assign n5920 = ~n5913 & n5919 ;
  assign n5921 = ~n5909 & n5920 ;
  assign n5922 = ~n5906 & n5921 ;
  assign n5923 = n2701 & ~n5922 ;
  assign n5924 = \P1_reg1_reg[27]/NET0131  & n4081 ;
  assign n5925 = ~n5923 & ~n5924 ;
  assign n5926 = \P1_state_reg[0]/NET0131  & ~n5925 ;
  assign n5927 = ~n5902 & ~n5926 ;
  assign n5928 = \P1_reg1_reg[28]/NET0131  & ~n4085 ;
  assign n5929 = \P1_reg1_reg[28]/NET0131  & n4081 ;
  assign n5930 = \P1_reg1_reg[28]/NET0131  & ~n4202 ;
  assign n5931 = n4202 & ~n4712 ;
  assign n5932 = ~n5930 & ~n5931 ;
  assign n5933 = n3829 & ~n5932 ;
  assign n5934 = n4202 & ~n4790 ;
  assign n5935 = ~n5930 & ~n5934 ;
  assign n5936 = n3969 & ~n5935 ;
  assign n5937 = n4202 & n4796 ;
  assign n5938 = ~n5930 & ~n5937 ;
  assign n5939 = n4062 & ~n5938 ;
  assign n5940 = n4202 & n4804 ;
  assign n5941 = ~n5930 & ~n5940 ;
  assign n5942 = n4025 & ~n5941 ;
  assign n5943 = \P1_reg1_reg[28]/NET0131  & ~n4216 ;
  assign n5944 = n4202 & n4794 ;
  assign n5945 = ~n5943 & ~n5944 ;
  assign n5946 = ~n5942 & n5945 ;
  assign n5947 = ~n5939 & n5946 ;
  assign n5948 = ~n5936 & n5947 ;
  assign n5949 = ~n5933 & n5948 ;
  assign n5950 = n2701 & ~n5949 ;
  assign n5951 = ~n5929 & ~n5950 ;
  assign n5952 = \P1_state_reg[0]/NET0131  & ~n5951 ;
  assign n5953 = ~n5928 & ~n5952 ;
  assign n5956 = n3633 & n4081 ;
  assign n5964 = n3633 & ~n4449 ;
  assign n5965 = ~n3717 & n4000 ;
  assign n5966 = ~n3613 & n5965 ;
  assign n5967 = ~n3640 & n5966 ;
  assign n5968 = n3587 & ~n5967 ;
  assign n5969 = ~n3587 & n5967 ;
  assign n5970 = ~n5968 & ~n5969 ;
  assign n5971 = ~n2731 & ~n5970 ;
  assign n5972 = n2731 & n3613 ;
  assign n5973 = ~n5971 & ~n5972 ;
  assign n5974 = n4449 & n5973 ;
  assign n5975 = ~n5964 & ~n5974 ;
  assign n5976 = n4025 & ~n5975 ;
  assign n5983 = ~n5009 & n5411 ;
  assign n5984 = n5009 & ~n5411 ;
  assign n5985 = ~n5983 & ~n5984 ;
  assign n5986 = n4449 & n5985 ;
  assign n5987 = ~n5964 & ~n5986 ;
  assign n5988 = n3829 & ~n5987 ;
  assign n5977 = ~n4976 & n5411 ;
  assign n5978 = n4976 & ~n5411 ;
  assign n5979 = ~n5977 & ~n5978 ;
  assign n5980 = n4449 & ~n5979 ;
  assign n5981 = ~n5964 & ~n5980 ;
  assign n5982 = n3969 & ~n5981 ;
  assign n5957 = ~n4046 & n4062 ;
  assign n5958 = ~n3631 & ~n5957 ;
  assign n5959 = n4046 & n4062 ;
  assign n5960 = n3631 & ~n4028 ;
  assign n5961 = ~n5959 & n5960 ;
  assign n5962 = ~n5958 & ~n5961 ;
  assign n5963 = n4449 & n5962 ;
  assign n5989 = n3631 & n4073 ;
  assign n5990 = n4069 & ~n4449 ;
  assign n5991 = ~n4067 & ~n5990 ;
  assign n5992 = n3633 & ~n5991 ;
  assign n5993 = ~n5989 & ~n5992 ;
  assign n5994 = ~n5963 & n5993 ;
  assign n5995 = ~n5982 & n5994 ;
  assign n5996 = ~n5988 & n5995 ;
  assign n5997 = ~n5976 & n5996 ;
  assign n5998 = n2701 & ~n5997 ;
  assign n5999 = ~n5956 & ~n5998 ;
  assign n6000 = \P1_state_reg[0]/NET0131  & ~n5999 ;
  assign n5954 = n3633 & n4552 ;
  assign n5955 = \P1_reg3_reg[18]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6001 = ~n5954 & ~n5955 ;
  assign n6002 = ~n6000 & n6001 ;
  assign n6005 = n3609 & n4081 ;
  assign n6007 = n3609 & ~n4449 ;
  assign n6016 = ~n3884 & n3920 ;
  assign n6017 = n3898 & ~n6016 ;
  assign n6018 = n5423 & ~n6017 ;
  assign n6019 = ~n5423 & n6017 ;
  assign n6020 = ~n6018 & ~n6019 ;
  assign n6021 = n4449 & ~n6020 ;
  assign n6022 = ~n6007 & ~n6021 ;
  assign n6023 = n3969 & ~n6022 ;
  assign n6008 = ~n3540 & n3744 ;
  assign n6009 = n3756 & ~n6008 ;
  assign n6010 = n5423 & n6009 ;
  assign n6011 = ~n5423 & ~n6009 ;
  assign n6012 = ~n6010 & ~n6011 ;
  assign n6013 = n4449 & ~n6012 ;
  assign n6014 = ~n6007 & ~n6013 ;
  assign n6015 = n3829 & ~n6014 ;
  assign n6024 = n3640 & ~n5966 ;
  assign n6025 = ~n5967 & ~n6024 ;
  assign n6026 = ~n2731 & ~n6025 ;
  assign n6027 = n2731 & n3717 ;
  assign n6028 = ~n6026 & ~n6027 ;
  assign n6029 = n4449 & n6028 ;
  assign n6030 = ~n6007 & ~n6029 ;
  assign n6031 = n4025 & ~n6030 ;
  assign n6032 = ~n3656 & n4042 ;
  assign n6033 = ~n3732 & n6032 ;
  assign n6034 = ~n3708 & n6033 ;
  assign n6035 = n3603 & ~n6034 ;
  assign n6036 = ~n4046 & ~n6035 ;
  assign n6037 = n4062 & n6036 ;
  assign n6038 = n4449 & n6037 ;
  assign n6006 = n3609 & ~n4542 ;
  assign n6039 = n3603 & ~n4522 ;
  assign n6040 = ~n6006 & ~n6039 ;
  assign n6041 = ~n6038 & n6040 ;
  assign n6042 = ~n6031 & n6041 ;
  assign n6043 = ~n6015 & n6042 ;
  assign n6044 = ~n6023 & n6043 ;
  assign n6045 = n2701 & ~n6044 ;
  assign n6046 = ~n6005 & ~n6045 ;
  assign n6047 = \P1_state_reg[0]/NET0131  & ~n6046 ;
  assign n6003 = n3609 & n4552 ;
  assign n6004 = \P1_reg3_reg[17]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6048 = ~n6003 & ~n6004 ;
  assign n6049 = ~n6047 & n6048 ;
  assign n6050 = n3580 & n4081 ;
  assign n6059 = n3580 & ~n4449 ;
  assign n6060 = n3561 & ~n5969 ;
  assign n6061 = n3975 & n5966 ;
  assign n6062 = ~n6060 & ~n6061 ;
  assign n6063 = ~n2731 & ~n6062 ;
  assign n6064 = n2731 & n3640 ;
  assign n6065 = ~n6063 & ~n6064 ;
  assign n6066 = n4449 & n6065 ;
  assign n6067 = ~n6059 & ~n6066 ;
  assign n6068 = n4025 & ~n6067 ;
  assign n6069 = n4477 & ~n5412 ;
  assign n6070 = ~n4477 & n5412 ;
  assign n6071 = ~n6069 & ~n6070 ;
  assign n6072 = n4449 & ~n6071 ;
  assign n6073 = ~n6059 & ~n6072 ;
  assign n6074 = n3829 & ~n6073 ;
  assign n6075 = n4503 & ~n5412 ;
  assign n6076 = ~n4503 & n5412 ;
  assign n6077 = ~n6075 & ~n6076 ;
  assign n6078 = n4449 & n6077 ;
  assign n6079 = ~n6059 & ~n6078 ;
  assign n6080 = n3969 & ~n6079 ;
  assign n6051 = n3578 & n4028 ;
  assign n6052 = ~n3631 & n4046 ;
  assign n6054 = n3578 & ~n6052 ;
  assign n6053 = ~n3578 & n6052 ;
  assign n6055 = n4062 & ~n6053 ;
  assign n6056 = ~n6054 & n6055 ;
  assign n6057 = ~n6051 & ~n6056 ;
  assign n6058 = n4449 & ~n6057 ;
  assign n6081 = n3578 & n4073 ;
  assign n6082 = n3580 & ~n5991 ;
  assign n6083 = ~n6081 & ~n6082 ;
  assign n6084 = ~n6058 & n6083 ;
  assign n6085 = ~n6080 & n6084 ;
  assign n6086 = ~n6074 & n6085 ;
  assign n6087 = ~n6068 & n6086 ;
  assign n6088 = n2701 & ~n6087 ;
  assign n6089 = ~n6050 & ~n6088 ;
  assign n6090 = \P1_state_reg[0]/NET0131  & ~n6089 ;
  assign n6091 = \P1_reg3_reg[19]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6092 = n3580 & n4552 ;
  assign n6093 = ~n6091 & ~n6092 ;
  assign n6094 = ~n6090 & n6093 ;
  assign n6097 = ~n1226 & n2035 ;
  assign n6108 = ~n1226 & ~n2053 ;
  assign n6100 = ~n2340 & n2343 ;
  assign n6101 = n2354 & ~n6100 ;
  assign n6102 = n1932 & n6101 ;
  assign n6103 = ~n1932 & ~n6101 ;
  assign n6104 = ~n6102 & ~n6103 ;
  assign n6109 = n2053 & n6104 ;
  assign n6110 = ~n6108 & ~n6109 ;
  assign n6111 = ~n2224 & ~n6110 ;
  assign n6099 = ~n1226 & ~n2124 ;
  assign n6105 = n2124 & n6104 ;
  assign n6106 = ~n6099 & ~n6105 ;
  assign n6107 = n2123 & ~n6106 ;
  assign n6112 = ~n1856 & n1932 ;
  assign n6113 = n1856 & ~n1932 ;
  assign n6114 = ~n6112 & ~n6113 ;
  assign n6115 = n2053 & n6114 ;
  assign n6116 = ~n6108 & ~n6115 ;
  assign n6117 = ~n2120 & ~n6116 ;
  assign n6118 = n1193 & ~n2247 ;
  assign n6119 = n2263 & ~n4261 ;
  assign n6120 = ~n6118 & n6119 ;
  assign n6121 = ~n601 & ~n2263 ;
  assign n6122 = ~n6120 & ~n6121 ;
  assign n6123 = n2124 & ~n6122 ;
  assign n6124 = ~n6099 & ~n6123 ;
  assign n6125 = n1790 & ~n6124 ;
  assign n6098 = ~n1255 & n2229 ;
  assign n6126 = ~n1226 & ~n2274 ;
  assign n6127 = ~n6098 & ~n6126 ;
  assign n6128 = ~n6125 & n6127 ;
  assign n6129 = ~n6117 & n6128 ;
  assign n6130 = ~n6107 & n6129 ;
  assign n6131 = ~n6111 & n6130 ;
  assign n6132 = n2037 & ~n6131 ;
  assign n6133 = ~n6097 & ~n6132 ;
  assign n6134 = \P1_state_reg[0]/NET0131  & ~n6133 ;
  assign n6095 = ~n1226 & n2014 ;
  assign n6096 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[16]/NET0131  ;
  assign n6135 = ~n6095 & ~n6096 ;
  assign n6136 = ~n6134 & n6135 ;
  assign n6137 = n3101 & ~n4449 ;
  assign n6138 = n4449 & ~n5054 ;
  assign n6139 = ~n6137 & ~n6138 ;
  assign n6140 = n3969 & ~n6139 ;
  assign n6141 = n4449 & ~n5068 ;
  assign n6142 = ~n6137 & ~n6141 ;
  assign n6143 = n3829 & ~n6142 ;
  assign n6144 = n4449 & n5080 ;
  assign n6145 = ~n6137 & ~n6144 ;
  assign n6146 = n4025 & ~n6145 ;
  assign n6148 = n4449 & n5090 ;
  assign n6147 = n3101 & ~n4542 ;
  assign n6149 = n3096 & ~n4522 ;
  assign n6150 = ~n6147 & ~n6149 ;
  assign n6151 = ~n6148 & n6150 ;
  assign n6152 = ~n6146 & n6151 ;
  assign n6153 = ~n6143 & n6152 ;
  assign n6154 = ~n6140 & n6153 ;
  assign n6155 = n2701 & ~n6154 ;
  assign n6156 = n3101 & n4081 ;
  assign n6157 = ~n6155 & ~n6156 ;
  assign n6158 = \P1_state_reg[0]/NET0131  & ~n6157 ;
  assign n6159 = \P1_reg3_reg[24]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6160 = n3101 & n4552 ;
  assign n6161 = ~n6159 & ~n6160 ;
  assign n6162 = ~n6158 & n6161 ;
  assign n6163 = \P1_reg2_reg[31]/NET0131  & ~n4085 ;
  assign n6164 = \P1_reg2_reg[31]/NET0131  & n4081 ;
  assign n6165 = \P1_reg2_reg[31]/NET0131  & ~n2717 ;
  assign n6166 = n4059 & ~n5371 ;
  assign n6167 = n5352 & ~n6166 ;
  assign n6168 = ~n5352 & n6166 ;
  assign n6169 = ~n6167 & ~n6168 ;
  assign n6170 = n2717 & n6169 ;
  assign n6171 = ~n6165 & ~n6170 ;
  assign n6172 = n4062 & ~n6171 ;
  assign n6173 = ~n3801 & ~n4015 ;
  assign n6174 = ~n2904 & n6173 ;
  assign n6175 = n4950 & n6174 ;
  assign n6176 = ~n3973 & ~n3984 ;
  assign n6177 = ~n6175 & n6176 ;
  assign n6178 = n2717 & n4025 ;
  assign n6179 = n6177 & n6178 ;
  assign n6180 = n2717 & n5352 ;
  assign n6181 = ~n6165 & ~n6180 ;
  assign n6182 = n4028 & ~n6181 ;
  assign n6183 = ~n3816 & ~n4024 ;
  assign n6184 = ~n2717 & ~n6183 ;
  assign n6185 = ~n4067 & ~n6184 ;
  assign n6186 = \P1_reg2_reg[31]/NET0131  & ~n6185 ;
  assign n6187 = ~n4074 & ~n6186 ;
  assign n6188 = ~n6182 & n6187 ;
  assign n6189 = ~n6179 & n6188 ;
  assign n6190 = ~n6172 & n6189 ;
  assign n6191 = n2701 & ~n6190 ;
  assign n6192 = ~n6164 & ~n6191 ;
  assign n6193 = \P1_state_reg[0]/NET0131  & ~n6192 ;
  assign n6194 = ~n6163 & ~n6193 ;
  assign n6195 = \P2_reg2_reg[23]/NET0131  & ~n2286 ;
  assign n6196 = \P2_reg2_reg[23]/NET0131  & n2035 ;
  assign n6197 = \P2_reg2_reg[23]/NET0131  & ~n2310 ;
  assign n6198 = ~n1549 & ~n4410 ;
  assign n6199 = n1549 & n4410 ;
  assign n6200 = ~n6198 & ~n6199 ;
  assign n6201 = n2263 & ~n6200 ;
  assign n6202 = ~n1474 & ~n2263 ;
  assign n6203 = ~n6201 & ~n6202 ;
  assign n6204 = n2310 & ~n6203 ;
  assign n6205 = ~n6197 & ~n6204 ;
  assign n6206 = n1790 & ~n6205 ;
  assign n6207 = \P2_reg2_reg[23]/NET0131  & ~n2291 ;
  assign n6208 = ~n2172 & n2181 ;
  assign n6209 = n2130 & n2198 ;
  assign n6210 = ~n6208 & n6209 ;
  assign n6211 = ~n2190 & n2198 ;
  assign n6212 = n2212 & ~n6211 ;
  assign n6213 = ~n6210 & n6212 ;
  assign n6214 = n1947 & ~n6213 ;
  assign n6215 = ~n1947 & n6213 ;
  assign n6216 = ~n6214 & ~n6215 ;
  assign n6217 = n2291 & n6216 ;
  assign n6218 = ~n6207 & ~n6217 ;
  assign n6219 = ~n2392 & ~n6218 ;
  assign n6235 = n1434 & n2272 ;
  assign n6236 = n2291 & n6235 ;
  assign n6237 = ~n1441 & n1854 ;
  assign n6238 = \P2_reg2_reg[23]/NET0131  & ~n2407 ;
  assign n6239 = ~n6237 & ~n6238 ;
  assign n6240 = ~n6236 & n6239 ;
  assign n6241 = ~n6219 & n6240 ;
  assign n6220 = ~n2078 & n2084 ;
  assign n6221 = n2057 & n2095 ;
  assign n6222 = ~n6220 & n6221 ;
  assign n6223 = ~n2090 & n2095 ;
  assign n6224 = n2108 & ~n6223 ;
  assign n6225 = ~n6222 & n6224 ;
  assign n6226 = n1947 & ~n6225 ;
  assign n6227 = ~n1947 & n6225 ;
  assign n6228 = ~n6226 & ~n6227 ;
  assign n6229 = n2291 & ~n6228 ;
  assign n6230 = ~n6207 & ~n6229 ;
  assign n6231 = ~n2290 & ~n6230 ;
  assign n6232 = n2310 & ~n6228 ;
  assign n6233 = ~n6197 & ~n6232 ;
  assign n6234 = n2314 & ~n6233 ;
  assign n6242 = ~n6231 & ~n6234 ;
  assign n6243 = n6241 & n6242 ;
  assign n6244 = ~n6206 & n6243 ;
  assign n6245 = n2037 & ~n6244 ;
  assign n6246 = ~n6196 & ~n6245 ;
  assign n6247 = \P1_state_reg[0]/NET0131  & ~n6246 ;
  assign n6248 = ~n6195 & ~n6247 ;
  assign n6249 = ~n1441 & n2035 ;
  assign n6250 = ~n1441 & ~n2124 ;
  assign n6251 = n2124 & ~n6203 ;
  assign n6252 = ~n6250 & ~n6251 ;
  assign n6253 = n1790 & ~n6252 ;
  assign n6254 = n2124 & n6216 ;
  assign n6255 = ~n6250 & ~n6254 ;
  assign n6256 = n2123 & ~n6255 ;
  assign n6257 = ~n1441 & ~n2274 ;
  assign n6258 = n1434 & n2229 ;
  assign n6266 = ~n6257 & ~n6258 ;
  assign n6267 = ~n6256 & n6266 ;
  assign n6259 = ~n1441 & ~n2053 ;
  assign n6260 = n2053 & ~n6228 ;
  assign n6261 = ~n6259 & ~n6260 ;
  assign n6262 = ~n2120 & ~n6261 ;
  assign n6263 = n2053 & n6216 ;
  assign n6264 = ~n6259 & ~n6263 ;
  assign n6265 = ~n2224 & ~n6264 ;
  assign n6268 = ~n6262 & ~n6265 ;
  assign n6269 = n6267 & n6268 ;
  assign n6270 = ~n6253 & n6269 ;
  assign n6271 = n2037 & ~n6270 ;
  assign n6272 = ~n6249 & ~n6271 ;
  assign n6273 = \P1_state_reg[0]/NET0131  & ~n6272 ;
  assign n6274 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[23]/NET0131  ;
  assign n6275 = ~n1441 & n2014 ;
  assign n6276 = ~n6274 & ~n6275 ;
  assign n6277 = ~n6273 & n6276 ;
  assign n6280 = n2970 & n4081 ;
  assign n6281 = n2970 & ~n4449 ;
  assign n6282 = n4449 & ~n5113 ;
  assign n6283 = ~n6281 & ~n6282 ;
  assign n6284 = n4025 & ~n6283 ;
  assign n6292 = n4449 & n5151 ;
  assign n6293 = ~n6281 & ~n6292 ;
  assign n6294 = n4062 & ~n6293 ;
  assign n6291 = n2970 & ~n4540 ;
  assign n6295 = n2964 & ~n4522 ;
  assign n6296 = ~n6291 & ~n6295 ;
  assign n6297 = ~n6294 & n6296 ;
  assign n6298 = ~n6284 & n6297 ;
  assign n6285 = n4449 & ~n5128 ;
  assign n6286 = ~n6281 & ~n6285 ;
  assign n6287 = n3829 & ~n6286 ;
  assign n6288 = n4449 & ~n5143 ;
  assign n6289 = ~n6281 & ~n6288 ;
  assign n6290 = n3969 & ~n6289 ;
  assign n6299 = ~n6287 & ~n6290 ;
  assign n6300 = n6298 & n6299 ;
  assign n6301 = n2701 & ~n6300 ;
  assign n6302 = ~n6280 & ~n6301 ;
  assign n6303 = \P1_state_reg[0]/NET0131  & ~n6302 ;
  assign n6278 = n2970 & n4552 ;
  assign n6279 = \P1_reg3_reg[25]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6304 = ~n6278 & ~n6279 ;
  assign n6305 = ~n6303 & n6304 ;
  assign n6306 = \P2_reg0_reg[22]/NET0131  & ~n2286 ;
  assign n6307 = \P2_reg0_reg[22]/NET0131  & n2035 ;
  assign n6311 = \P2_reg0_reg[22]/NET0131  & ~n2053 ;
  assign n6312 = ~n4400 & ~n6311 ;
  assign n6313 = n2123 & ~n6312 ;
  assign n6308 = \P2_reg0_reg[22]/NET0131  & ~n2124 ;
  assign n6309 = ~n4404 & ~n6308 ;
  assign n6310 = ~n2224 & ~n6309 ;
  assign n6315 = n2053 & ~n4415 ;
  assign n6316 = ~n6311 & ~n6315 ;
  assign n6317 = n1790 & ~n6316 ;
  assign n6318 = n2124 & ~n4433 ;
  assign n6319 = ~n6308 & ~n6318 ;
  assign n6320 = ~n2120 & ~n6319 ;
  assign n6314 = n2124 & n4570 ;
  assign n6321 = \P2_reg0_reg[22]/NET0131  & ~n2614 ;
  assign n6322 = ~n6314 & ~n6321 ;
  assign n6323 = ~n6320 & n6322 ;
  assign n6324 = ~n6317 & n6323 ;
  assign n6325 = ~n6310 & n6324 ;
  assign n6326 = ~n6313 & n6325 ;
  assign n6327 = n2037 & ~n6326 ;
  assign n6328 = ~n6307 & ~n6327 ;
  assign n6329 = \P1_state_reg[0]/NET0131  & ~n6328 ;
  assign n6330 = ~n6306 & ~n6329 ;
  assign n6331 = \P1_reg2_reg[26]/NET0131  & ~n4085 ;
  assign n6332 = \P1_reg2_reg[26]/NET0131  & n4081 ;
  assign n6333 = \P1_reg2_reg[26]/NET0131  & ~n2717 ;
  assign n6334 = n2717 & n4954 ;
  assign n6335 = ~n6333 & ~n6334 ;
  assign n6336 = n4025 & ~n6335 ;
  assign n6345 = n2717 & ~n5841 ;
  assign n6343 = \P1_reg2_reg[26]/NET0131  & ~n4071 ;
  assign n6344 = n3022 & n4073 ;
  assign n6346 = ~n6343 & ~n6344 ;
  assign n6347 = ~n6345 & n6346 ;
  assign n6348 = ~n6336 & n6347 ;
  assign n6337 = n2717 & ~n4990 ;
  assign n6338 = ~n6333 & ~n6337 ;
  assign n6339 = n3969 & ~n6338 ;
  assign n6340 = n2717 & ~n5024 ;
  assign n6341 = ~n6333 & ~n6340 ;
  assign n6342 = n3829 & ~n6341 ;
  assign n6349 = ~n6339 & ~n6342 ;
  assign n6350 = n6348 & n6349 ;
  assign n6351 = n2701 & ~n6350 ;
  assign n6352 = ~n6332 & ~n6351 ;
  assign n6353 = \P1_state_reg[0]/NET0131  & ~n6352 ;
  assign n6354 = ~n6331 & ~n6353 ;
  assign n6355 = \P2_reg1_reg[22]/NET0131  & ~n2286 ;
  assign n6356 = \P2_reg1_reg[22]/NET0131  & n2035 ;
  assign n6357 = n2310 & ~n4399 ;
  assign n6358 = \P2_reg1_reg[22]/NET0131  & ~n2310 ;
  assign n6359 = ~n6357 & ~n6358 ;
  assign n6360 = ~n2392 & ~n6359 ;
  assign n6361 = \P2_reg1_reg[22]/NET0131  & ~n2291 ;
  assign n6362 = n2291 & ~n4415 ;
  assign n6363 = ~n6361 & ~n6362 ;
  assign n6364 = n1790 & ~n6363 ;
  assign n6368 = ~n4567 & ~n6361 ;
  assign n6369 = n2314 & ~n6368 ;
  assign n6365 = ~n4572 & ~n6358 ;
  assign n6366 = ~n2290 & ~n6365 ;
  assign n6367 = n2310 & n4570 ;
  assign n6370 = \P2_reg1_reg[22]/NET0131  & ~n4099 ;
  assign n6371 = ~n6367 & ~n6370 ;
  assign n6372 = ~n6366 & n6371 ;
  assign n6373 = ~n6369 & n6372 ;
  assign n6374 = ~n6364 & n6373 ;
  assign n6375 = ~n6360 & n6374 ;
  assign n6376 = n2037 & ~n6375 ;
  assign n6377 = ~n6356 & ~n6376 ;
  assign n6378 = \P1_state_reg[0]/NET0131  & ~n6377 ;
  assign n6379 = ~n6355 & ~n6378 ;
  assign n6380 = \P1_reg0_reg[22]/NET0131  & ~n4085 ;
  assign n6381 = \P1_reg0_reg[22]/NET0131  & n4081 ;
  assign n6382 = \P1_reg0_reg[22]/NET0131  & ~n4869 ;
  assign n6383 = n3128 & ~n4947 ;
  assign n6384 = ~n3128 & n4947 ;
  assign n6385 = ~n6383 & ~n6384 ;
  assign n6386 = ~n2731 & ~n6385 ;
  assign n6387 = n2731 & n3177 ;
  assign n6388 = ~n6386 & ~n6387 ;
  assign n6389 = n4869 & n6388 ;
  assign n6390 = ~n6382 & ~n6389 ;
  assign n6391 = n4025 & ~n6390 ;
  assign n6416 = n3143 & n4028 ;
  assign n6417 = ~n3168 & n4049 ;
  assign n6418 = n3143 & ~n6417 ;
  assign n6419 = ~n4051 & ~n6418 ;
  assign n6420 = n4062 & n6419 ;
  assign n6421 = ~n6416 & ~n6420 ;
  assign n6422 = n4869 & ~n6421 ;
  assign n6423 = \P1_reg0_reg[22]/NET0131  & ~n5844 ;
  assign n6424 = ~n6422 & ~n6423 ;
  assign n6425 = ~n6391 & n6424 ;
  assign n6393 = ~n5001 & n5004 ;
  assign n6394 = n4994 & n5010 ;
  assign n6395 = ~n6393 & n6394 ;
  assign n6392 = ~n5007 & n5010 ;
  assign n6396 = n5015 & ~n6392 ;
  assign n6397 = ~n6395 & n6396 ;
  assign n6398 = n5410 & n6397 ;
  assign n6399 = ~n5410 & ~n6397 ;
  assign n6400 = ~n6398 & ~n6399 ;
  assign n6401 = n4869 & ~n6400 ;
  assign n6402 = ~n6382 & ~n6401 ;
  assign n6403 = n3829 & ~n6402 ;
  assign n6405 = ~n4968 & n4971 ;
  assign n6406 = n4959 & n4978 ;
  assign n6407 = ~n6405 & n6406 ;
  assign n6404 = ~n4974 & n4978 ;
  assign n6408 = n4982 & ~n6404 ;
  assign n6409 = ~n6407 & n6408 ;
  assign n6410 = n5410 & ~n6409 ;
  assign n6411 = ~n5410 & n6409 ;
  assign n6412 = ~n6410 & ~n6411 ;
  assign n6413 = n4869 & ~n6412 ;
  assign n6414 = ~n6382 & ~n6413 ;
  assign n6415 = n3969 & ~n6414 ;
  assign n6426 = ~n6403 & ~n6415 ;
  assign n6427 = n6425 & n6426 ;
  assign n6428 = n2701 & ~n6427 ;
  assign n6429 = ~n6381 & ~n6428 ;
  assign n6430 = \P1_state_reg[0]/NET0131  & ~n6429 ;
  assign n6431 = ~n6380 & ~n6430 ;
  assign n6432 = \P1_reg0_reg[25]/NET0131  & ~n4085 ;
  assign n6433 = \P1_reg0_reg[25]/NET0131  & n4081 ;
  assign n6434 = \P1_reg0_reg[25]/NET0131  & ~n4869 ;
  assign n6435 = n4869 & ~n5113 ;
  assign n6436 = ~n6434 & ~n6435 ;
  assign n6437 = n4025 & ~n6436 ;
  assign n6445 = n4869 & n5151 ;
  assign n6446 = ~n6434 & ~n6445 ;
  assign n6447 = n4062 & ~n6446 ;
  assign n6444 = \P1_reg0_reg[25]/NET0131  & ~n5864 ;
  assign n6448 = n4869 & n5156 ;
  assign n6449 = ~n6444 & ~n6448 ;
  assign n6450 = ~n6447 & n6449 ;
  assign n6451 = ~n6437 & n6450 ;
  assign n6438 = n4869 & ~n5128 ;
  assign n6439 = ~n6434 & ~n6438 ;
  assign n6440 = n3829 & ~n6439 ;
  assign n6441 = n4869 & ~n5143 ;
  assign n6442 = ~n6434 & ~n6441 ;
  assign n6443 = n3969 & ~n6442 ;
  assign n6452 = ~n6440 & ~n6443 ;
  assign n6453 = n6451 & n6452 ;
  assign n6454 = n2701 & ~n6453 ;
  assign n6455 = ~n6433 & ~n6454 ;
  assign n6456 = \P1_state_reg[0]/NET0131  & ~n6455 ;
  assign n6457 = ~n6432 & ~n6456 ;
  assign n6458 = \P1_reg0_reg[24]/NET0131  & ~n4869 ;
  assign n6459 = n4869 & ~n5054 ;
  assign n6460 = ~n6458 & ~n6459 ;
  assign n6461 = n3969 & ~n6460 ;
  assign n6462 = n4869 & ~n5068 ;
  assign n6463 = ~n6458 & ~n6462 ;
  assign n6464 = n3829 & ~n6463 ;
  assign n6465 = n4869 & n5080 ;
  assign n6466 = ~n6458 & ~n6465 ;
  assign n6467 = n4025 & ~n6466 ;
  assign n6468 = n4869 & ~n5091 ;
  assign n6469 = \P1_reg0_reg[24]/NET0131  & ~n5866 ;
  assign n6470 = ~n6468 & ~n6469 ;
  assign n6471 = ~n6467 & n6470 ;
  assign n6472 = ~n6464 & n6471 ;
  assign n6473 = ~n6461 & n6472 ;
  assign n6474 = n2701 & ~n6473 ;
  assign n6475 = \P1_reg0_reg[24]/NET0131  & n4081 ;
  assign n6476 = ~n6474 & ~n6475 ;
  assign n6477 = \P1_state_reg[0]/NET0131  & ~n6476 ;
  assign n6478 = \P1_reg0_reg[24]/NET0131  & ~n4085 ;
  assign n6479 = ~n6477 & ~n6478 ;
  assign n6480 = \P1_reg1_reg[22]/NET0131  & ~n4085 ;
  assign n6481 = \P1_reg1_reg[22]/NET0131  & n4081 ;
  assign n6482 = \P1_reg1_reg[22]/NET0131  & ~n4202 ;
  assign n6483 = n4202 & n6388 ;
  assign n6484 = ~n6482 & ~n6483 ;
  assign n6485 = n4025 & ~n6484 ;
  assign n6492 = n4202 & ~n6421 ;
  assign n6493 = n4069 & ~n4202 ;
  assign n6494 = n4214 & ~n6493 ;
  assign n6495 = \P1_reg1_reg[22]/NET0131  & ~n6494 ;
  assign n6496 = ~n6492 & ~n6495 ;
  assign n6497 = ~n6485 & n6496 ;
  assign n6486 = n4202 & ~n6412 ;
  assign n6487 = ~n6482 & ~n6486 ;
  assign n6488 = n3969 & ~n6487 ;
  assign n6489 = n4202 & ~n6400 ;
  assign n6490 = ~n6482 & ~n6489 ;
  assign n6491 = n3829 & ~n6490 ;
  assign n6498 = ~n6488 & ~n6491 ;
  assign n6499 = n6497 & n6498 ;
  assign n6500 = n2701 & ~n6499 ;
  assign n6501 = ~n6481 & ~n6500 ;
  assign n6502 = \P1_state_reg[0]/NET0131  & ~n6501 ;
  assign n6503 = ~n6480 & ~n6502 ;
  assign n6504 = \P1_reg1_reg[24]/NET0131  & ~n4202 ;
  assign n6505 = n4202 & ~n5054 ;
  assign n6506 = ~n6504 & ~n6505 ;
  assign n6507 = n3969 & ~n6506 ;
  assign n6508 = n4202 & ~n5068 ;
  assign n6509 = ~n6504 & ~n6508 ;
  assign n6510 = n3829 & ~n6509 ;
  assign n6511 = n4202 & n5080 ;
  assign n6512 = ~n6504 & ~n6511 ;
  assign n6513 = n4025 & ~n6512 ;
  assign n6515 = n4202 & n5089 ;
  assign n6516 = ~n6504 & ~n6515 ;
  assign n6517 = n4062 & ~n6516 ;
  assign n6514 = \P1_reg1_reg[24]/NET0131  & ~n4214 ;
  assign n6518 = n3096 & n4202 ;
  assign n6519 = ~n6504 & ~n6518 ;
  assign n6520 = n4028 & ~n6519 ;
  assign n6521 = ~n6514 & ~n6520 ;
  assign n6522 = ~n6517 & n6521 ;
  assign n6523 = ~n6513 & n6522 ;
  assign n6524 = ~n6510 & n6523 ;
  assign n6525 = ~n6507 & n6524 ;
  assign n6526 = n2701 & ~n6525 ;
  assign n6527 = \P1_reg1_reg[24]/NET0131  & n4081 ;
  assign n6528 = ~n6526 & ~n6527 ;
  assign n6529 = \P1_state_reg[0]/NET0131  & ~n6528 ;
  assign n6530 = \P1_reg1_reg[24]/NET0131  & ~n4085 ;
  assign n6531 = ~n6529 & ~n6530 ;
  assign n6532 = \P1_reg1_reg[25]/NET0131  & ~n4085 ;
  assign n6533 = \P1_reg1_reg[25]/NET0131  & n4081 ;
  assign n6534 = \P1_reg1_reg[25]/NET0131  & ~n4202 ;
  assign n6535 = n4202 & ~n5113 ;
  assign n6536 = ~n6534 & ~n6535 ;
  assign n6537 = n4025 & ~n6536 ;
  assign n6545 = n4202 & n5151 ;
  assign n6546 = ~n6534 & ~n6545 ;
  assign n6547 = n4062 & ~n6546 ;
  assign n6544 = \P1_reg1_reg[25]/NET0131  & ~n4216 ;
  assign n6548 = n4202 & n5156 ;
  assign n6549 = ~n6544 & ~n6548 ;
  assign n6550 = ~n6547 & n6549 ;
  assign n6551 = ~n6537 & n6550 ;
  assign n6538 = n4202 & ~n5128 ;
  assign n6539 = ~n6534 & ~n6538 ;
  assign n6540 = n3829 & ~n6539 ;
  assign n6541 = n4202 & ~n5143 ;
  assign n6542 = ~n6534 & ~n6541 ;
  assign n6543 = n3969 & ~n6542 ;
  assign n6552 = ~n6540 & ~n6543 ;
  assign n6553 = n6551 & n6552 ;
  assign n6554 = n2701 & ~n6553 ;
  assign n6555 = ~n6533 & ~n6554 ;
  assign n6556 = \P1_state_reg[0]/NET0131  & ~n6555 ;
  assign n6557 = ~n6532 & ~n6556 ;
  assign n6558 = \P1_reg1_reg[26]/NET0131  & ~n4085 ;
  assign n6559 = \P1_reg1_reg[26]/NET0131  & n4081 ;
  assign n6560 = \P1_reg1_reg[26]/NET0131  & ~n4202 ;
  assign n6561 = n4202 & n4954 ;
  assign n6562 = ~n6560 & ~n6561 ;
  assign n6563 = n4025 & ~n6562 ;
  assign n6570 = n4202 & ~n5841 ;
  assign n6571 = \P1_reg1_reg[26]/NET0131  & ~n6494 ;
  assign n6572 = ~n6570 & ~n6571 ;
  assign n6573 = ~n6563 & n6572 ;
  assign n6564 = n4202 & ~n5024 ;
  assign n6565 = ~n6560 & ~n6564 ;
  assign n6566 = n3829 & ~n6565 ;
  assign n6567 = n4202 & ~n4990 ;
  assign n6568 = ~n6560 & ~n6567 ;
  assign n6569 = n3969 & ~n6568 ;
  assign n6574 = ~n6566 & ~n6569 ;
  assign n6575 = n6573 & n6574 ;
  assign n6576 = n2701 & ~n6575 ;
  assign n6577 = ~n6559 & ~n6576 ;
  assign n6578 = \P1_state_reg[0]/NET0131  & ~n6577 ;
  assign n6579 = ~n6558 & ~n6578 ;
  assign n6581 = n3244 & n4081 ;
  assign n6583 = n3244 & ~n4449 ;
  assign n6584 = ~n4665 & n5419 ;
  assign n6585 = n4665 & ~n5419 ;
  assign n6586 = ~n6584 & ~n6585 ;
  assign n6587 = n4449 & n6586 ;
  assign n6588 = ~n6583 & ~n6587 ;
  assign n6589 = n3829 & ~n6588 ;
  assign n6590 = n3692 & ~n4942 ;
  assign n6591 = ~n4943 & ~n6590 ;
  assign n6592 = ~n2731 & ~n6591 ;
  assign n6593 = n2731 & n3221 ;
  assign n6594 = ~n6592 & ~n6593 ;
  assign n6595 = n4449 & n6594 ;
  assign n6596 = ~n6583 & ~n6595 ;
  assign n6597 = n4025 & ~n6596 ;
  assign n6604 = ~n3435 & n4036 ;
  assign n6605 = ~n3291 & n6604 ;
  assign n6606 = ~n3263 & n6605 ;
  assign n6607 = ~n3211 & n6606 ;
  assign n6608 = n3239 & ~n6607 ;
  assign n6609 = n4037 & n6606 ;
  assign n6610 = ~n6608 & ~n6609 ;
  assign n6611 = n4062 & n6610 ;
  assign n6612 = n4449 & n6611 ;
  assign n6598 = ~n4744 & n5419 ;
  assign n6599 = n4744 & ~n5419 ;
  assign n6600 = ~n6598 & ~n6599 ;
  assign n6601 = n4449 & ~n6600 ;
  assign n6602 = ~n6583 & ~n6601 ;
  assign n6603 = n3969 & ~n6602 ;
  assign n6582 = n3244 & ~n4542 ;
  assign n6613 = n3239 & ~n4522 ;
  assign n6614 = ~n6582 & ~n6613 ;
  assign n6615 = ~n6603 & n6614 ;
  assign n6616 = ~n6612 & n6615 ;
  assign n6617 = ~n6597 & n6616 ;
  assign n6618 = ~n6589 & n6617 ;
  assign n6619 = n2701 & ~n6618 ;
  assign n6620 = ~n6581 & ~n6619 ;
  assign n6621 = \P1_state_reg[0]/NET0131  & ~n6620 ;
  assign n6580 = \P1_reg3_reg[12]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6622 = n3244 & n4552 ;
  assign n6623 = ~n6580 & ~n6622 ;
  assign n6624 = ~n6621 & n6623 ;
  assign n6627 = n3713 & n4081 ;
  assign n6628 = n3713 & ~n4449 ;
  assign n6643 = ~n4665 & n4668 ;
  assign n6644 = n4679 & ~n6643 ;
  assign n6645 = n5425 & n6644 ;
  assign n6646 = ~n5425 & ~n6644 ;
  assign n6647 = ~n6645 & ~n6646 ;
  assign n6648 = n4449 & ~n6647 ;
  assign n6649 = ~n6628 & ~n6648 ;
  assign n6650 = n3829 & ~n6649 ;
  assign n6637 = ~n5047 & n5425 ;
  assign n6638 = n5047 & ~n5425 ;
  assign n6639 = ~n6637 & ~n6638 ;
  assign n6640 = n4449 & ~n6639 ;
  assign n6641 = ~n6628 & ~n6640 ;
  assign n6642 = n3969 & ~n6641 ;
  assign n6629 = n3613 & ~n5965 ;
  assign n6630 = ~n5966 & ~n6629 ;
  assign n6631 = ~n2731 & ~n6630 ;
  assign n6632 = n2731 & n3741 ;
  assign n6633 = ~n6631 & ~n6632 ;
  assign n6634 = n4449 & n6633 ;
  assign n6635 = ~n6628 & ~n6634 ;
  assign n6636 = n4025 & ~n6635 ;
  assign n6652 = n3708 & ~n6033 ;
  assign n6653 = ~n6034 & ~n6652 ;
  assign n6654 = n4062 & n6653 ;
  assign n6655 = n4449 & n6654 ;
  assign n6651 = n3713 & ~n4542 ;
  assign n6656 = n3708 & ~n4522 ;
  assign n6657 = ~n6651 & ~n6656 ;
  assign n6658 = ~n6655 & n6657 ;
  assign n6659 = ~n6636 & n6658 ;
  assign n6660 = ~n6642 & n6659 ;
  assign n6661 = ~n6650 & n6660 ;
  assign n6662 = n2701 & ~n6661 ;
  assign n6663 = ~n6627 & ~n6662 ;
  assign n6664 = \P1_state_reg[0]/NET0131  & ~n6663 ;
  assign n6625 = \P1_reg3_reg[16]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6626 = n3713 & n4552 ;
  assign n6665 = ~n6625 & ~n6626 ;
  assign n6666 = ~n6664 & n6665 ;
  assign n6667 = n3172 & ~n4449 ;
  assign n6668 = n3917 & ~n6017 ;
  assign n6669 = n3912 & ~n6668 ;
  assign n6670 = n5433 & ~n6669 ;
  assign n6671 = ~n5433 & n6669 ;
  assign n6672 = ~n6670 & ~n6671 ;
  assign n6673 = n4449 & ~n6672 ;
  assign n6674 = ~n6667 & ~n6673 ;
  assign n6675 = n3969 & ~n6674 ;
  assign n6677 = n3769 & n5433 ;
  assign n6678 = ~n3769 & ~n5433 ;
  assign n6679 = ~n6677 & ~n6678 ;
  assign n6680 = n4449 & ~n6679 ;
  assign n6681 = ~n6667 & ~n6680 ;
  assign n6682 = n3829 & ~n6681 ;
  assign n6683 = ~n3153 & n4001 ;
  assign n6684 = n3153 & ~n4001 ;
  assign n6685 = ~n6683 & ~n6684 ;
  assign n6686 = ~n2731 & ~n6685 ;
  assign n6687 = n2731 & n3561 ;
  assign n6688 = n4025 & ~n6687 ;
  assign n6689 = ~n6686 & n6688 ;
  assign n6690 = n3168 & ~n4049 ;
  assign n6691 = n4062 & ~n6417 ;
  assign n6692 = ~n6690 & n6691 ;
  assign n6693 = ~n6689 & ~n6692 ;
  assign n6694 = n4449 & ~n6693 ;
  assign n6676 = n3168 & ~n4522 ;
  assign n6695 = ~n3816 & n4066 ;
  assign n6696 = ~n4028 & ~n6695 ;
  assign n6697 = ~n4449 & ~n6696 ;
  assign n6698 = ~n4067 & ~n6697 ;
  assign n6699 = n3172 & ~n6698 ;
  assign n6700 = ~n6676 & ~n6699 ;
  assign n6701 = ~n6694 & n6700 ;
  assign n6702 = ~n6682 & n6701 ;
  assign n6703 = ~n6675 & n6702 ;
  assign n6704 = n2701 & ~n6703 ;
  assign n6705 = n3172 & n4081 ;
  assign n6706 = ~n6704 & ~n6705 ;
  assign n6707 = \P1_state_reg[0]/NET0131  & ~n6706 ;
  assign n6708 = \P1_reg3_reg[21]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6709 = n3172 & n4552 ;
  assign n6710 = ~n6708 & ~n6709 ;
  assign n6711 = ~n6707 & n6710 ;
  assign n6712 = n3557 & n4081 ;
  assign n6714 = n3557 & ~n4449 ;
  assign n6723 = n4688 & n5432 ;
  assign n6724 = ~n4688 & ~n5432 ;
  assign n6725 = ~n6723 & ~n6724 ;
  assign n6726 = n4449 & ~n6725 ;
  assign n6727 = ~n6714 & ~n6726 ;
  assign n6728 = n3829 & ~n6727 ;
  assign n6715 = n3177 & ~n6061 ;
  assign n6716 = ~n4001 & ~n6715 ;
  assign n6717 = ~n2731 & ~n6716 ;
  assign n6718 = n2731 & n3587 ;
  assign n6719 = ~n6717 & ~n6718 ;
  assign n6720 = n4449 & n6719 ;
  assign n6721 = ~n6714 & ~n6720 ;
  assign n6722 = n4025 & ~n6721 ;
  assign n6729 = ~n4764 & n5432 ;
  assign n6730 = n4764 & ~n5432 ;
  assign n6731 = ~n6729 & ~n6730 ;
  assign n6732 = n4449 & ~n6731 ;
  assign n6733 = ~n6714 & ~n6732 ;
  assign n6734 = n3969 & ~n6733 ;
  assign n6735 = n3548 & ~n6053 ;
  assign n6736 = ~n4049 & ~n6735 ;
  assign n6737 = n4062 & n6736 ;
  assign n6738 = n4449 & n6737 ;
  assign n6713 = n3557 & ~n4542 ;
  assign n6739 = n3548 & ~n4522 ;
  assign n6740 = ~n6713 & ~n6739 ;
  assign n6741 = ~n6738 & n6740 ;
  assign n6742 = ~n6734 & n6741 ;
  assign n6743 = ~n6722 & n6742 ;
  assign n6744 = ~n6728 & n6743 ;
  assign n6745 = n2701 & ~n6744 ;
  assign n6746 = ~n6712 & ~n6745 ;
  assign n6747 = \P1_state_reg[0]/NET0131  & ~n6746 ;
  assign n6748 = n3557 & n4552 ;
  assign n6749 = \P1_reg3_reg[20]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6750 = ~n6748 & ~n6749 ;
  assign n6751 = ~n6747 & n6750 ;
  assign n6752 = \P1_reg2_reg[21]/NET0131  & ~n4085 ;
  assign n6753 = \P1_reg2_reg[21]/NET0131  & ~n2717 ;
  assign n6754 = n2717 & ~n6672 ;
  assign n6755 = ~n6753 & ~n6754 ;
  assign n6756 = n3969 & ~n6755 ;
  assign n6760 = n2717 & ~n6679 ;
  assign n6761 = ~n6753 & ~n6760 ;
  assign n6762 = n3829 & ~n6761 ;
  assign n6757 = n3168 & n4028 ;
  assign n6758 = n6693 & ~n6757 ;
  assign n6759 = n2717 & ~n6758 ;
  assign n6763 = ~n2717 & ~n6696 ;
  assign n6764 = ~n4067 & ~n6763 ;
  assign n6765 = \P1_reg2_reg[21]/NET0131  & ~n6764 ;
  assign n6766 = n3172 & n4073 ;
  assign n6767 = ~n6765 & ~n6766 ;
  assign n6768 = ~n6759 & n6767 ;
  assign n6769 = ~n6762 & n6768 ;
  assign n6770 = ~n6756 & n6769 ;
  assign n6771 = n2701 & ~n6770 ;
  assign n6772 = \P1_reg2_reg[21]/NET0131  & n4081 ;
  assign n6773 = ~n6771 & ~n6772 ;
  assign n6774 = \P1_state_reg[0]/NET0131  & ~n6773 ;
  assign n6775 = ~n6752 & ~n6774 ;
  assign n6776 = \P1_reg2_reg[18]/NET0131  & ~n4085 ;
  assign n6777 = \P1_reg2_reg[18]/NET0131  & n4081 ;
  assign n6779 = \P1_reg2_reg[18]/NET0131  & ~n2717 ;
  assign n6780 = n2717 & n5973 ;
  assign n6781 = ~n6779 & ~n6780 ;
  assign n6782 = n4025 & ~n6781 ;
  assign n6786 = n2717 & ~n5979 ;
  assign n6787 = ~n6779 & ~n6786 ;
  assign n6788 = n3969 & ~n6787 ;
  assign n6783 = n2717 & n5985 ;
  assign n6784 = ~n6779 & ~n6783 ;
  assign n6785 = n3829 & ~n6784 ;
  assign n6778 = n2717 & n5962 ;
  assign n6789 = n3633 & n4073 ;
  assign n6790 = \P1_reg2_reg[18]/NET0131  & ~n4071 ;
  assign n6791 = ~n6789 & ~n6790 ;
  assign n6792 = ~n6778 & n6791 ;
  assign n6793 = ~n6785 & n6792 ;
  assign n6794 = ~n6788 & n6793 ;
  assign n6795 = ~n6782 & n6794 ;
  assign n6796 = n2701 & ~n6795 ;
  assign n6797 = ~n6777 & ~n6796 ;
  assign n6798 = \P1_state_reg[0]/NET0131  & ~n6797 ;
  assign n6799 = ~n6776 & ~n6798 ;
  assign n6800 = \P1_reg2_reg[17]/NET0131  & ~n4085 ;
  assign n6801 = \P1_reg2_reg[17]/NET0131  & n4081 ;
  assign n6803 = \P1_reg2_reg[17]/NET0131  & ~n2717 ;
  assign n6807 = n2717 & ~n6020 ;
  assign n6808 = ~n6803 & ~n6807 ;
  assign n6809 = n3969 & ~n6808 ;
  assign n6804 = n2717 & ~n6012 ;
  assign n6805 = ~n6803 & ~n6804 ;
  assign n6806 = n3829 & ~n6805 ;
  assign n6810 = n2717 & n6028 ;
  assign n6811 = ~n6803 & ~n6810 ;
  assign n6812 = n4025 & ~n6811 ;
  assign n6813 = n2717 & n6036 ;
  assign n6814 = ~n6803 & ~n6813 ;
  assign n6815 = n4062 & ~n6814 ;
  assign n6817 = n3603 & n4028 ;
  assign n6818 = n2717 & n6817 ;
  assign n6802 = \P1_reg2_reg[17]/NET0131  & ~n5148 ;
  assign n6816 = n3609 & n4073 ;
  assign n6819 = ~n6802 & ~n6816 ;
  assign n6820 = ~n6818 & n6819 ;
  assign n6821 = ~n6815 & n6820 ;
  assign n6822 = ~n6812 & n6821 ;
  assign n6823 = ~n6806 & n6822 ;
  assign n6824 = ~n6809 & n6823 ;
  assign n6825 = n2701 & ~n6824 ;
  assign n6826 = ~n6801 & ~n6825 ;
  assign n6827 = \P1_state_reg[0]/NET0131  & ~n6826 ;
  assign n6828 = ~n6800 & ~n6827 ;
  assign n6829 = \P1_reg2_reg[19]/NET0131  & ~n4085 ;
  assign n6830 = \P1_reg2_reg[19]/NET0131  & n4081 ;
  assign n6832 = \P1_reg2_reg[19]/NET0131  & ~n2717 ;
  assign n6833 = n2717 & n6065 ;
  assign n6834 = ~n6832 & ~n6833 ;
  assign n6835 = n4025 & ~n6834 ;
  assign n6836 = n2717 & ~n6071 ;
  assign n6837 = ~n6832 & ~n6836 ;
  assign n6838 = n3829 & ~n6837 ;
  assign n6839 = n2717 & n6077 ;
  assign n6840 = ~n6832 & ~n6839 ;
  assign n6841 = n3969 & ~n6840 ;
  assign n6831 = n2717 & ~n6057 ;
  assign n6842 = n3580 & n4073 ;
  assign n6843 = \P1_reg2_reg[19]/NET0131  & ~n4071 ;
  assign n6844 = ~n6842 & ~n6843 ;
  assign n6845 = ~n6831 & n6844 ;
  assign n6846 = ~n6841 & n6845 ;
  assign n6847 = ~n6838 & n6846 ;
  assign n6848 = ~n6835 & n6847 ;
  assign n6849 = n2701 & ~n6848 ;
  assign n6850 = ~n6830 & ~n6849 ;
  assign n6851 = \P1_state_reg[0]/NET0131  & ~n6850 ;
  assign n6852 = ~n6829 & ~n6851 ;
  assign n6855 = ~n1378 & n2035 ;
  assign n6858 = ~n1378 & ~n2124 ;
  assign n6859 = n2124 & ~n5629 ;
  assign n6860 = ~n6858 & ~n6859 ;
  assign n6861 = n1790 & ~n6860 ;
  assign n6856 = n1371 & n2229 ;
  assign n6857 = ~n1378 & ~n2274 ;
  assign n6872 = ~n6856 & ~n6857 ;
  assign n6873 = ~n6861 & n6872 ;
  assign n6865 = ~n1378 & ~n2053 ;
  assign n6869 = n2053 & ~n5617 ;
  assign n6870 = ~n6865 & ~n6869 ;
  assign n6871 = ~n2120 & ~n6870 ;
  assign n6862 = n2124 & ~n5611 ;
  assign n6863 = ~n6858 & ~n6862 ;
  assign n6864 = n2123 & ~n6863 ;
  assign n6866 = n2053 & ~n5611 ;
  assign n6867 = ~n6865 & ~n6866 ;
  assign n6868 = ~n2224 & ~n6867 ;
  assign n6874 = ~n6864 & ~n6868 ;
  assign n6875 = ~n6871 & n6874 ;
  assign n6876 = n6873 & n6875 ;
  assign n6877 = n2037 & ~n6876 ;
  assign n6878 = ~n6855 & ~n6877 ;
  assign n6879 = \P1_state_reg[0]/NET0131  & ~n6878 ;
  assign n6853 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[21]/NET0131  ;
  assign n6854 = ~n1378 & n2014 ;
  assign n6880 = ~n6853 & ~n6854 ;
  assign n6881 = ~n6879 & n6880 ;
  assign n6884 = n3149 & n4081 ;
  assign n6885 = n3149 & ~n4449 ;
  assign n6886 = n4449 & n6388 ;
  assign n6887 = ~n6885 & ~n6886 ;
  assign n6888 = n4025 & ~n6887 ;
  assign n6896 = n4449 & n6420 ;
  assign n6895 = n3149 & ~n4542 ;
  assign n6897 = n3143 & ~n4522 ;
  assign n6898 = ~n6895 & ~n6897 ;
  assign n6899 = ~n6896 & n6898 ;
  assign n6900 = ~n6888 & n6899 ;
  assign n6889 = n4449 & ~n6400 ;
  assign n6890 = ~n6885 & ~n6889 ;
  assign n6891 = n3829 & ~n6890 ;
  assign n6892 = n4449 & ~n6412 ;
  assign n6893 = ~n6885 & ~n6892 ;
  assign n6894 = n3969 & ~n6893 ;
  assign n6901 = ~n6891 & ~n6894 ;
  assign n6902 = n6900 & n6901 ;
  assign n6903 = n2701 & ~n6902 ;
  assign n6904 = ~n6884 & ~n6903 ;
  assign n6905 = \P1_state_reg[0]/NET0131  & ~n6904 ;
  assign n6882 = \P1_reg3_reg[22]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6883 = n3149 & n4552 ;
  assign n6906 = ~n6882 & ~n6883 ;
  assign n6907 = ~n6905 & n6906 ;
  assign n6908 = \P2_reg0_reg[18]/NET0131  & ~n2286 ;
  assign n6909 = \P2_reg0_reg[18]/NET0131  & n2035 ;
  assign n6910 = \P2_reg0_reg[18]/NET0131  & ~n2124 ;
  assign n6911 = ~n4258 & ~n6910 ;
  assign n6912 = ~n2224 & ~n6911 ;
  assign n6922 = \P2_reg0_reg[18]/NET0131  & ~n2614 ;
  assign n6923 = n2124 & n5214 ;
  assign n6924 = ~n6922 & ~n6923 ;
  assign n6925 = ~n6912 & n6924 ;
  assign n6919 = n2124 & ~n4289 ;
  assign n6920 = ~n6910 & ~n6919 ;
  assign n6921 = ~n2120 & ~n6920 ;
  assign n6913 = \P2_reg0_reg[18]/NET0131  & ~n2053 ;
  assign n6914 = ~n4254 & ~n6913 ;
  assign n6915 = n2123 & ~n6914 ;
  assign n6916 = n2053 & ~n4268 ;
  assign n6917 = ~n6913 & ~n6916 ;
  assign n6918 = n1790 & ~n6917 ;
  assign n6926 = ~n6915 & ~n6918 ;
  assign n6927 = ~n6921 & n6926 ;
  assign n6928 = n6925 & n6927 ;
  assign n6929 = n2037 & ~n6928 ;
  assign n6930 = ~n6909 & ~n6929 ;
  assign n6931 = \P1_state_reg[0]/NET0131  & ~n6930 ;
  assign n6932 = ~n6908 & ~n6931 ;
  assign n6933 = \P1_reg1_reg[31]/NET0131  & ~n4085 ;
  assign n6934 = \P1_reg1_reg[31]/NET0131  & n4081 ;
  assign n6935 = \P1_reg1_reg[31]/NET0131  & ~n4202 ;
  assign n6936 = n4202 & n6169 ;
  assign n6937 = ~n6935 & ~n6936 ;
  assign n6938 = n4062 & ~n6937 ;
  assign n6945 = n4025 & n4202 ;
  assign n6946 = n6177 & n6945 ;
  assign n6939 = n4202 & n5352 ;
  assign n6940 = ~n6935 & ~n6939 ;
  assign n6941 = n4028 & ~n6940 ;
  assign n6942 = ~n4202 & ~n6183 ;
  assign n6943 = n4214 & ~n6942 ;
  assign n6944 = \P1_reg1_reg[31]/NET0131  & ~n6943 ;
  assign n6947 = ~n6941 & ~n6944 ;
  assign n6948 = ~n6946 & n6947 ;
  assign n6949 = ~n6938 & n6948 ;
  assign n6950 = n2701 & ~n6949 ;
  assign n6951 = ~n6934 & ~n6950 ;
  assign n6952 = \P1_state_reg[0]/NET0131  & ~n6951 ;
  assign n6953 = ~n6933 & ~n6952 ;
  assign n6954 = \P2_reg0_reg[19]/NET0131  & ~n2286 ;
  assign n6955 = \P2_reg0_reg[19]/NET0131  & n2035 ;
  assign n6956 = \P2_reg0_reg[19]/NET0131  & ~n2124 ;
  assign n6957 = ~n4325 & ~n6956 ;
  assign n6958 = ~n2224 & ~n6957 ;
  assign n6968 = \P2_reg0_reg[19]/NET0131  & ~n2614 ;
  assign n6969 = n2124 & n5244 ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = ~n6958 & n6970 ;
  assign n6965 = n2124 & n4330 ;
  assign n6966 = ~n6956 & ~n6965 ;
  assign n6967 = ~n2120 & ~n6966 ;
  assign n6959 = \P2_reg0_reg[19]/NET0131  & ~n2053 ;
  assign n6960 = n2053 & ~n4321 ;
  assign n6961 = ~n6959 & ~n6960 ;
  assign n6962 = n1790 & ~n6961 ;
  assign n6963 = ~n4312 & ~n6959 ;
  assign n6964 = n2123 & ~n6963 ;
  assign n6972 = ~n6962 & ~n6964 ;
  assign n6973 = ~n6967 & n6972 ;
  assign n6974 = n6971 & n6973 ;
  assign n6975 = n2037 & ~n6974 ;
  assign n6976 = ~n6955 & ~n6975 ;
  assign n6977 = \P1_state_reg[0]/NET0131  & ~n6976 ;
  assign n6978 = ~n6954 & ~n6977 ;
  assign n6979 = \P2_reg0_reg[17]/NET0131  & ~n2286 ;
  assign n6980 = \P2_reg0_reg[17]/NET0131  & n2035 ;
  assign n6982 = \P2_reg0_reg[17]/NET0131  & ~n2124 ;
  assign n6983 = ~n4358 & ~n6982 ;
  assign n6984 = ~n2224 & ~n6983 ;
  assign n6985 = \P2_reg0_reg[17]/NET0131  & ~n2053 ;
  assign n6991 = n2053 & ~n4373 ;
  assign n6992 = ~n6985 & ~n6991 ;
  assign n6993 = n1790 & ~n6992 ;
  assign n6981 = n2124 & n5184 ;
  assign n6994 = \P2_reg0_reg[17]/NET0131  & ~n2614 ;
  assign n6995 = ~n6981 & ~n6994 ;
  assign n6996 = ~n6993 & n6995 ;
  assign n6997 = ~n6984 & n6996 ;
  assign n6986 = ~n4354 & ~n6985 ;
  assign n6987 = n2123 & ~n6986 ;
  assign n6988 = n2124 & ~n4365 ;
  assign n6989 = ~n6982 & ~n6988 ;
  assign n6990 = ~n2120 & ~n6989 ;
  assign n6998 = ~n6987 & ~n6990 ;
  assign n6999 = n6997 & n6998 ;
  assign n7000 = n2037 & ~n6999 ;
  assign n7001 = ~n6980 & ~n7000 ;
  assign n7002 = \P1_state_reg[0]/NET0131  & ~n7001 ;
  assign n7003 = ~n6979 & ~n7002 ;
  assign n7004 = \P2_reg0_reg[21]/NET0131  & ~n2286 ;
  assign n7005 = \P2_reg0_reg[21]/NET0131  & n2035 ;
  assign n7006 = \P2_reg0_reg[21]/NET0131  & ~n2053 ;
  assign n7007 = n2053 & ~n5629 ;
  assign n7008 = ~n7006 & ~n7007 ;
  assign n7009 = n1790 & ~n7008 ;
  assign n7018 = \P2_reg0_reg[21]/NET0131  & ~n2614 ;
  assign n7019 = n2124 & n5633 ;
  assign n7020 = ~n7018 & ~n7019 ;
  assign n7021 = ~n7009 & n7020 ;
  assign n7012 = \P2_reg0_reg[21]/NET0131  & ~n2124 ;
  assign n7015 = n2124 & ~n5617 ;
  assign n7016 = ~n7012 & ~n7015 ;
  assign n7017 = ~n2120 & ~n7016 ;
  assign n7010 = ~n6866 & ~n7006 ;
  assign n7011 = n2123 & ~n7010 ;
  assign n7013 = ~n6862 & ~n7012 ;
  assign n7014 = ~n2224 & ~n7013 ;
  assign n7022 = ~n7011 & ~n7014 ;
  assign n7023 = ~n7017 & n7022 ;
  assign n7024 = n7021 & n7023 ;
  assign n7025 = n2037 & ~n7024 ;
  assign n7026 = ~n7005 & ~n7025 ;
  assign n7027 = \P1_state_reg[0]/NET0131  & ~n7026 ;
  assign n7028 = ~n7004 & ~n7027 ;
  assign n7029 = \P2_reg0_reg[20]/NET0131  & ~n2286 ;
  assign n7030 = \P2_reg0_reg[20]/NET0131  & n2035 ;
  assign n7032 = \P2_reg0_reg[20]/NET0131  & ~n2124 ;
  assign n7033 = ~n5263 & ~n7032 ;
  assign n7034 = ~n2224 & ~n7033 ;
  assign n7031 = \P2_reg0_reg[20]/NET0131  & ~n2614 ;
  assign n7044 = n1401 & n2616 ;
  assign n7045 = ~n7031 & ~n7044 ;
  assign n7046 = ~n7034 & n7045 ;
  assign n7035 = \P2_reg0_reg[20]/NET0131  & ~n2053 ;
  assign n7041 = n2053 & ~n4905 ;
  assign n7042 = ~n7035 & ~n7041 ;
  assign n7043 = n1790 & ~n7042 ;
  assign n7036 = ~n5267 & ~n7035 ;
  assign n7037 = n2123 & ~n7036 ;
  assign n7038 = n2124 & ~n4918 ;
  assign n7039 = ~n7032 & ~n7038 ;
  assign n7040 = ~n2120 & ~n7039 ;
  assign n7047 = ~n7037 & ~n7040 ;
  assign n7048 = ~n7043 & n7047 ;
  assign n7049 = n7046 & n7048 ;
  assign n7050 = n2037 & ~n7049 ;
  assign n7051 = ~n7030 & ~n7050 ;
  assign n7052 = \P1_state_reg[0]/NET0131  & ~n7051 ;
  assign n7053 = ~n7029 & ~n7052 ;
  assign n7054 = \P1_reg2_reg[20]/NET0131  & ~n4085 ;
  assign n7055 = \P1_reg2_reg[20]/NET0131  & n4081 ;
  assign n7059 = \P1_reg2_reg[20]/NET0131  & ~n2717 ;
  assign n7063 = n2717 & ~n6725 ;
  assign n7064 = ~n7059 & ~n7063 ;
  assign n7065 = n3829 & ~n7064 ;
  assign n7060 = n2717 & n6719 ;
  assign n7061 = ~n7059 & ~n7060 ;
  assign n7062 = n4025 & ~n7061 ;
  assign n7066 = n2717 & ~n6731 ;
  assign n7067 = ~n7059 & ~n7066 ;
  assign n7068 = n3969 & ~n7067 ;
  assign n7069 = n3548 & n4028 ;
  assign n7070 = ~n6737 & ~n7069 ;
  assign n7071 = n2717 & ~n7070 ;
  assign n7056 = ~n2717 & n4062 ;
  assign n7057 = n5148 & ~n7056 ;
  assign n7058 = \P1_reg2_reg[20]/NET0131  & ~n7057 ;
  assign n7072 = n3557 & n4073 ;
  assign n7073 = ~n7058 & ~n7072 ;
  assign n7074 = ~n7071 & n7073 ;
  assign n7075 = ~n7068 & n7074 ;
  assign n7076 = ~n7062 & n7075 ;
  assign n7077 = ~n7065 & n7076 ;
  assign n7078 = n2701 & ~n7077 ;
  assign n7079 = ~n7055 & ~n7078 ;
  assign n7080 = \P1_state_reg[0]/NET0131  & ~n7079 ;
  assign n7081 = ~n7054 & ~n7080 ;
  assign n7082 = \P2_reg1_reg[17]/NET0131  & ~n2286 ;
  assign n7083 = \P2_reg1_reg[17]/NET0131  & n2035 ;
  assign n7085 = \P2_reg1_reg[17]/NET0131  & ~n2310 ;
  assign n7086 = n2310 & n4353 ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7088 = ~n2392 & ~n7087 ;
  assign n7089 = \P2_reg1_reg[17]/NET0131  & ~n2291 ;
  assign n7094 = n2291 & ~n4373 ;
  assign n7095 = ~n7089 & ~n7094 ;
  assign n7096 = n1790 & ~n7095 ;
  assign n7084 = n2310 & n5184 ;
  assign n7097 = \P2_reg1_reg[17]/NET0131  & ~n4099 ;
  assign n7098 = ~n7084 & ~n7097 ;
  assign n7099 = ~n7096 & n7098 ;
  assign n7100 = ~n7088 & n7099 ;
  assign n7090 = ~n5181 & ~n7089 ;
  assign n7091 = n2314 & ~n7090 ;
  assign n7092 = ~n5178 & ~n7085 ;
  assign n7093 = ~n2290 & ~n7092 ;
  assign n7101 = ~n7091 & ~n7093 ;
  assign n7102 = n7100 & n7101 ;
  assign n7103 = n2037 & ~n7102 ;
  assign n7104 = ~n7083 & ~n7103 ;
  assign n7105 = \P1_state_reg[0]/NET0131  & ~n7104 ;
  assign n7106 = ~n7082 & ~n7105 ;
  assign n7107 = \P2_reg1_reg[18]/NET0131  & ~n2286 ;
  assign n7108 = \P2_reg1_reg[18]/NET0131  & n2035 ;
  assign n7109 = \P2_reg1_reg[18]/NET0131  & ~n2310 ;
  assign n7110 = n2310 & n4253 ;
  assign n7111 = ~n7109 & ~n7110 ;
  assign n7112 = ~n2392 & ~n7111 ;
  assign n7121 = \P2_reg1_reg[18]/NET0131  & ~n4099 ;
  assign n7122 = n2310 & n5214 ;
  assign n7123 = ~n7121 & ~n7122 ;
  assign n7124 = ~n7112 & n7123 ;
  assign n7119 = ~n5211 & ~n7109 ;
  assign n7120 = ~n2290 & ~n7119 ;
  assign n7113 = \P2_reg1_reg[18]/NET0131  & ~n2291 ;
  assign n7114 = ~n5208 & ~n7113 ;
  assign n7115 = n2314 & ~n7114 ;
  assign n7116 = n2291 & ~n4268 ;
  assign n7117 = ~n7113 & ~n7116 ;
  assign n7118 = n1790 & ~n7117 ;
  assign n7125 = ~n7115 & ~n7118 ;
  assign n7126 = ~n7120 & n7125 ;
  assign n7127 = n7124 & n7126 ;
  assign n7128 = n2037 & ~n7127 ;
  assign n7129 = ~n7108 & ~n7128 ;
  assign n7130 = \P1_state_reg[0]/NET0131  & ~n7129 ;
  assign n7131 = ~n7107 & ~n7130 ;
  assign n7132 = \P2_reg1_reg[19]/NET0131  & ~n2286 ;
  assign n7133 = \P2_reg1_reg[19]/NET0131  & n2035 ;
  assign n7134 = \P2_reg1_reg[19]/NET0131  & ~n2291 ;
  assign n7135 = n2291 & ~n4321 ;
  assign n7136 = ~n7134 & ~n7135 ;
  assign n7137 = n1790 & ~n7136 ;
  assign n7146 = \P2_reg1_reg[19]/NET0131  & ~n4099 ;
  assign n7147 = n2310 & n5244 ;
  assign n7148 = ~n7146 & ~n7147 ;
  assign n7149 = ~n7137 & n7148 ;
  assign n7140 = \P2_reg1_reg[19]/NET0131  & ~n2310 ;
  assign n7143 = n2310 & ~n4311 ;
  assign n7144 = ~n7140 & ~n7143 ;
  assign n7145 = ~n2392 & ~n7144 ;
  assign n7138 = ~n5238 & ~n7134 ;
  assign n7139 = n2314 & ~n7138 ;
  assign n7141 = ~n5234 & ~n7140 ;
  assign n7142 = ~n2290 & ~n7141 ;
  assign n7150 = ~n7139 & ~n7142 ;
  assign n7151 = ~n7145 & n7150 ;
  assign n7152 = n7149 & n7151 ;
  assign n7153 = n2037 & ~n7152 ;
  assign n7154 = ~n7133 & ~n7153 ;
  assign n7155 = \P1_state_reg[0]/NET0131  & ~n7154 ;
  assign n7156 = ~n7132 & ~n7155 ;
  assign n7157 = \P2_reg1_reg[20]/NET0131  & ~n2286 ;
  assign n7158 = \P2_reg1_reg[20]/NET0131  & n2035 ;
  assign n7160 = \P2_reg1_reg[20]/NET0131  & ~n2310 ;
  assign n7161 = n2310 & ~n4912 ;
  assign n7162 = ~n7160 & ~n7161 ;
  assign n7163 = ~n2392 & ~n7162 ;
  assign n7159 = \P2_reg1_reg[20]/NET0131  & ~n4099 ;
  assign n7172 = n1401 & n4101 ;
  assign n7173 = ~n7159 & ~n7172 ;
  assign n7174 = ~n7163 & n7173 ;
  assign n7166 = \P2_reg1_reg[20]/NET0131  & ~n2291 ;
  assign n7169 = n2291 & ~n4905 ;
  assign n7170 = ~n7166 & ~n7169 ;
  assign n7171 = n1790 & ~n7170 ;
  assign n7164 = ~n4919 & ~n7160 ;
  assign n7165 = ~n2290 & ~n7164 ;
  assign n7167 = ~n4922 & ~n7166 ;
  assign n7168 = n2314 & ~n7167 ;
  assign n7175 = ~n7165 & ~n7168 ;
  assign n7176 = ~n7171 & n7175 ;
  assign n7177 = n7174 & n7176 ;
  assign n7178 = n2037 & ~n7177 ;
  assign n7179 = ~n7158 & ~n7178 ;
  assign n7180 = \P1_state_reg[0]/NET0131  & ~n7179 ;
  assign n7181 = ~n7157 & ~n7180 ;
  assign n7182 = \P2_reg1_reg[21]/NET0131  & ~n2286 ;
  assign n7183 = \P2_reg1_reg[21]/NET0131  & n2035 ;
  assign n7184 = \P2_reg1_reg[21]/NET0131  & ~n2310 ;
  assign n7185 = n2310 & ~n5611 ;
  assign n7186 = ~n7184 & ~n7185 ;
  assign n7187 = ~n2392 & ~n7186 ;
  assign n7196 = \P2_reg1_reg[21]/NET0131  & ~n4099 ;
  assign n7197 = n2310 & n5633 ;
  assign n7198 = ~n7196 & ~n7197 ;
  assign n7199 = ~n7187 & n7198 ;
  assign n7190 = \P2_reg1_reg[21]/NET0131  & ~n2291 ;
  assign n7193 = n2291 & ~n5629 ;
  assign n7194 = ~n7190 & ~n7193 ;
  assign n7195 = n1790 & ~n7194 ;
  assign n7188 = ~n5622 & ~n7184 ;
  assign n7189 = ~n2290 & ~n7188 ;
  assign n7191 = ~n5618 & ~n7190 ;
  assign n7192 = n2314 & ~n7191 ;
  assign n7200 = ~n7189 & ~n7192 ;
  assign n7201 = ~n7195 & n7200 ;
  assign n7202 = n7199 & n7201 ;
  assign n7203 = n2037 & ~n7202 ;
  assign n7204 = ~n7183 & ~n7203 ;
  assign n7205 = \P1_state_reg[0]/NET0131  & ~n7204 ;
  assign n7206 = ~n7182 & ~n7205 ;
  assign n7207 = \P1_reg0_reg[17]/NET0131  & ~n4085 ;
  assign n7208 = \P1_reg0_reg[17]/NET0131  & n4081 ;
  assign n7210 = \P1_reg0_reg[17]/NET0131  & ~n4869 ;
  assign n7214 = n4869 & ~n6020 ;
  assign n7215 = ~n7210 & ~n7214 ;
  assign n7216 = n3969 & ~n7215 ;
  assign n7211 = n4869 & ~n6012 ;
  assign n7212 = ~n7210 & ~n7211 ;
  assign n7213 = n3829 & ~n7212 ;
  assign n7217 = n4869 & n6028 ;
  assign n7218 = ~n7210 & ~n7217 ;
  assign n7219 = n4025 & ~n7218 ;
  assign n7209 = \P1_reg0_reg[17]/NET0131  & ~n5866 ;
  assign n7220 = ~n6037 & ~n6817 ;
  assign n7221 = n4869 & ~n7220 ;
  assign n7222 = ~n7209 & ~n7221 ;
  assign n7223 = ~n7219 & n7222 ;
  assign n7224 = ~n7213 & n7223 ;
  assign n7225 = ~n7216 & n7224 ;
  assign n7226 = n2701 & ~n7225 ;
  assign n7227 = ~n7208 & ~n7226 ;
  assign n7228 = \P1_state_reg[0]/NET0131  & ~n7227 ;
  assign n7229 = ~n7207 & ~n7228 ;
  assign n7230 = \P1_reg0_reg[18]/NET0131  & ~n4085 ;
  assign n7231 = \P1_reg0_reg[18]/NET0131  & n4081 ;
  assign n7233 = \P1_reg0_reg[18]/NET0131  & ~n4869 ;
  assign n7234 = n4869 & n5973 ;
  assign n7235 = ~n7233 & ~n7234 ;
  assign n7236 = n4025 & ~n7235 ;
  assign n7240 = n4869 & ~n5979 ;
  assign n7241 = ~n7233 & ~n7240 ;
  assign n7242 = n3969 & ~n7241 ;
  assign n7237 = n4869 & n5985 ;
  assign n7238 = ~n7233 & ~n7237 ;
  assign n7239 = n3829 & ~n7238 ;
  assign n7232 = n4869 & n5962 ;
  assign n7243 = \P1_reg0_reg[18]/NET0131  & ~n5844 ;
  assign n7244 = ~n7232 & ~n7243 ;
  assign n7245 = ~n7239 & n7244 ;
  assign n7246 = ~n7242 & n7245 ;
  assign n7247 = ~n7236 & n7246 ;
  assign n7248 = n2701 & ~n7247 ;
  assign n7249 = ~n7231 & ~n7248 ;
  assign n7250 = \P1_state_reg[0]/NET0131  & ~n7249 ;
  assign n7251 = ~n7230 & ~n7250 ;
  assign n7252 = \P1_reg0_reg[19]/NET0131  & ~n4085 ;
  assign n7253 = \P1_reg0_reg[19]/NET0131  & n4081 ;
  assign n7255 = \P1_reg0_reg[19]/NET0131  & ~n4869 ;
  assign n7256 = n4869 & n6065 ;
  assign n7257 = ~n7255 & ~n7256 ;
  assign n7258 = n4025 & ~n7257 ;
  assign n7259 = n4869 & ~n6071 ;
  assign n7260 = ~n7255 & ~n7259 ;
  assign n7261 = n3829 & ~n7260 ;
  assign n7262 = n4869 & n6077 ;
  assign n7263 = ~n7255 & ~n7262 ;
  assign n7264 = n3969 & ~n7263 ;
  assign n7254 = n4869 & ~n6057 ;
  assign n7265 = \P1_reg0_reg[19]/NET0131  & ~n5844 ;
  assign n7266 = ~n7254 & ~n7265 ;
  assign n7267 = ~n7264 & n7266 ;
  assign n7268 = ~n7261 & n7267 ;
  assign n7269 = ~n7258 & n7268 ;
  assign n7270 = n2701 & ~n7269 ;
  assign n7271 = ~n7253 & ~n7270 ;
  assign n7272 = \P1_state_reg[0]/NET0131  & ~n7271 ;
  assign n7273 = ~n7252 & ~n7272 ;
  assign n7274 = \P1_reg0_reg[21]/NET0131  & ~n4085 ;
  assign n7275 = \P1_reg0_reg[21]/NET0131  & n4081 ;
  assign n7276 = \P1_reg0_reg[21]/NET0131  & ~n4869 ;
  assign n7277 = n4869 & ~n6672 ;
  assign n7278 = ~n7276 & ~n7277 ;
  assign n7279 = n3969 & ~n7278 ;
  assign n7281 = n4869 & ~n6679 ;
  assign n7282 = ~n7276 & ~n7281 ;
  assign n7283 = n3829 & ~n7282 ;
  assign n7280 = n4869 & ~n6758 ;
  assign n7284 = ~n4869 & ~n6696 ;
  assign n7285 = n4214 & ~n7284 ;
  assign n7286 = \P1_reg0_reg[21]/NET0131  & ~n7285 ;
  assign n7287 = ~n7280 & ~n7286 ;
  assign n7288 = ~n7283 & n7287 ;
  assign n7289 = ~n7279 & n7288 ;
  assign n7290 = n2701 & ~n7289 ;
  assign n7291 = ~n7275 & ~n7290 ;
  assign n7292 = \P1_state_reg[0]/NET0131  & ~n7291 ;
  assign n7293 = ~n7274 & ~n7292 ;
  assign n7294 = \P1_reg0_reg[31]/NET0131  & ~n4085 ;
  assign n7295 = \P1_reg0_reg[31]/NET0131  & n4081 ;
  assign n7296 = \P1_reg0_reg[31]/NET0131  & ~n4869 ;
  assign n7297 = n4869 & n6169 ;
  assign n7298 = ~n7296 & ~n7297 ;
  assign n7299 = n4062 & ~n7298 ;
  assign n7306 = n4025 & n4869 ;
  assign n7307 = n6177 & n7306 ;
  assign n7300 = n4869 & n5352 ;
  assign n7301 = ~n7296 & ~n7300 ;
  assign n7302 = n4028 & ~n7301 ;
  assign n7303 = ~n4869 & ~n6183 ;
  assign n7304 = n4214 & ~n7303 ;
  assign n7305 = \P1_reg0_reg[31]/NET0131  & ~n7304 ;
  assign n7308 = ~n7302 & ~n7305 ;
  assign n7309 = ~n7307 & n7308 ;
  assign n7310 = ~n7299 & n7309 ;
  assign n7311 = n2701 & ~n7310 ;
  assign n7312 = ~n7295 & ~n7311 ;
  assign n7313 = \P1_state_reg[0]/NET0131  & ~n7312 ;
  assign n7314 = ~n7294 & ~n7313 ;
  assign n7315 = \P1_reg1_reg[17]/NET0131  & ~n4085 ;
  assign n7316 = \P1_reg1_reg[17]/NET0131  & n4081 ;
  assign n7318 = \P1_reg1_reg[17]/NET0131  & ~n4202 ;
  assign n7322 = n4202 & ~n6020 ;
  assign n7323 = ~n7318 & ~n7322 ;
  assign n7324 = n3969 & ~n7323 ;
  assign n7319 = n4202 & ~n6012 ;
  assign n7320 = ~n7318 & ~n7319 ;
  assign n7321 = n3829 & ~n7320 ;
  assign n7325 = n4202 & n6028 ;
  assign n7326 = ~n7318 & ~n7325 ;
  assign n7327 = n4025 & ~n7326 ;
  assign n7317 = \P1_reg1_reg[17]/NET0131  & ~n4218 ;
  assign n7328 = n4202 & ~n7220 ;
  assign n7329 = ~n7317 & ~n7328 ;
  assign n7330 = ~n7327 & n7329 ;
  assign n7331 = ~n7321 & n7330 ;
  assign n7332 = ~n7324 & n7331 ;
  assign n7333 = n2701 & ~n7332 ;
  assign n7334 = ~n7316 & ~n7333 ;
  assign n7335 = \P1_state_reg[0]/NET0131  & ~n7334 ;
  assign n7336 = ~n7315 & ~n7335 ;
  assign n7337 = \P1_reg1_reg[18]/NET0131  & ~n4085 ;
  assign n7338 = \P1_reg1_reg[18]/NET0131  & n4081 ;
  assign n7340 = \P1_reg1_reg[18]/NET0131  & ~n4202 ;
  assign n7341 = n4202 & n5973 ;
  assign n7342 = ~n7340 & ~n7341 ;
  assign n7343 = n4025 & ~n7342 ;
  assign n7347 = n4202 & ~n5979 ;
  assign n7348 = ~n7340 & ~n7347 ;
  assign n7349 = n3969 & ~n7348 ;
  assign n7344 = n4202 & n5985 ;
  assign n7345 = ~n7340 & ~n7344 ;
  assign n7346 = n3829 & ~n7345 ;
  assign n7339 = \P1_reg1_reg[18]/NET0131  & ~n6494 ;
  assign n7350 = n4202 & n5962 ;
  assign n7351 = ~n7339 & ~n7350 ;
  assign n7352 = ~n7346 & n7351 ;
  assign n7353 = ~n7349 & n7352 ;
  assign n7354 = ~n7343 & n7353 ;
  assign n7355 = n2701 & ~n7354 ;
  assign n7356 = ~n7338 & ~n7355 ;
  assign n7357 = \P1_state_reg[0]/NET0131  & ~n7356 ;
  assign n7358 = ~n7337 & ~n7357 ;
  assign n7359 = \P1_reg1_reg[19]/NET0131  & ~n4085 ;
  assign n7360 = \P1_reg1_reg[19]/NET0131  & n4081 ;
  assign n7362 = \P1_reg1_reg[19]/NET0131  & ~n4202 ;
  assign n7363 = n4202 & n6065 ;
  assign n7364 = ~n7362 & ~n7363 ;
  assign n7365 = n4025 & ~n7364 ;
  assign n7366 = n4202 & ~n6071 ;
  assign n7367 = ~n7362 & ~n7366 ;
  assign n7368 = n3829 & ~n7367 ;
  assign n7369 = n4202 & n6077 ;
  assign n7370 = ~n7362 & ~n7369 ;
  assign n7371 = n3969 & ~n7370 ;
  assign n7361 = n4202 & ~n6057 ;
  assign n7372 = \P1_reg1_reg[19]/NET0131  & ~n6494 ;
  assign n7373 = ~n7361 & ~n7372 ;
  assign n7374 = ~n7371 & n7373 ;
  assign n7375 = ~n7368 & n7374 ;
  assign n7376 = ~n7365 & n7375 ;
  assign n7377 = n2701 & ~n7376 ;
  assign n7378 = ~n7360 & ~n7377 ;
  assign n7379 = \P1_state_reg[0]/NET0131  & ~n7378 ;
  assign n7380 = ~n7359 & ~n7379 ;
  assign n7381 = \P1_reg1_reg[21]/NET0131  & ~n4085 ;
  assign n7382 = \P1_reg1_reg[21]/NET0131  & n4081 ;
  assign n7383 = \P1_reg1_reg[21]/NET0131  & ~n4202 ;
  assign n7384 = n4202 & ~n6672 ;
  assign n7385 = ~n7383 & ~n7384 ;
  assign n7386 = n3969 & ~n7385 ;
  assign n7388 = n4202 & ~n6679 ;
  assign n7389 = ~n7383 & ~n7388 ;
  assign n7390 = n3829 & ~n7389 ;
  assign n7387 = n4202 & ~n6758 ;
  assign n7391 = ~n4202 & ~n6696 ;
  assign n7392 = n4214 & ~n7391 ;
  assign n7393 = \P1_reg1_reg[21]/NET0131  & ~n7392 ;
  assign n7394 = ~n7387 & ~n7393 ;
  assign n7395 = ~n7390 & n7394 ;
  assign n7396 = ~n7386 & n7395 ;
  assign n7397 = n2701 & ~n7396 ;
  assign n7398 = ~n7382 & ~n7397 ;
  assign n7399 = \P1_state_reg[0]/NET0131  & ~n7398 ;
  assign n7400 = ~n7381 & ~n7399 ;
  assign n7403 = n3271 & n4081 ;
  assign n7405 = n3271 & ~n4449 ;
  assign n7406 = ~n3275 & n3994 ;
  assign n7407 = n3221 & ~n7406 ;
  assign n7408 = n3994 & n3995 ;
  assign n7409 = ~n7407 & ~n7408 ;
  assign n7410 = ~n2731 & ~n7409 ;
  assign n7411 = n2731 & n3300 ;
  assign n7412 = ~n7410 & ~n7411 ;
  assign n7413 = n4449 & n7412 ;
  assign n7414 = ~n7405 & ~n7413 ;
  assign n7415 = n4025 & ~n7414 ;
  assign n7422 = ~n4966 & n5414 ;
  assign n7423 = n4966 & ~n5414 ;
  assign n7424 = ~n7422 & ~n7423 ;
  assign n7425 = n4449 & ~n7424 ;
  assign n7426 = ~n7405 & ~n7425 ;
  assign n7427 = n3969 & ~n7426 ;
  assign n7416 = ~n4999 & n5414 ;
  assign n7417 = n4999 & ~n5414 ;
  assign n7418 = ~n7416 & ~n7417 ;
  assign n7419 = n4449 & n7418 ;
  assign n7420 = ~n7405 & ~n7419 ;
  assign n7421 = n3829 & ~n7420 ;
  assign n7428 = n3263 & ~n6605 ;
  assign n7429 = ~n6606 & ~n7428 ;
  assign n7430 = n4449 & n7429 ;
  assign n7431 = ~n7405 & ~n7430 ;
  assign n7432 = n4062 & ~n7431 ;
  assign n7404 = n3263 & ~n4522 ;
  assign n7433 = n3271 & ~n4540 ;
  assign n7434 = ~n7404 & ~n7433 ;
  assign n7435 = ~n7432 & n7434 ;
  assign n7436 = ~n7421 & n7435 ;
  assign n7437 = ~n7427 & n7436 ;
  assign n7438 = ~n7415 & n7437 ;
  assign n7439 = n2701 & ~n7438 ;
  assign n7440 = ~n7403 & ~n7439 ;
  assign n7441 = \P1_state_reg[0]/NET0131  & ~n7440 ;
  assign n7401 = \P1_reg3_reg[10]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7402 = n3271 & n4552 ;
  assign n7442 = ~n7401 & ~n7402 ;
  assign n7443 = ~n7441 & n7442 ;
  assign n7446 = n3686 & n4081 ;
  assign n7448 = n3686 & ~n4449 ;
  assign n7449 = n3665 & ~n4943 ;
  assign n7450 = ~n4944 & ~n7449 ;
  assign n7451 = ~n2731 & ~n7450 ;
  assign n7452 = n2731 & n3248 ;
  assign n7453 = ~n7451 & ~n7452 ;
  assign n7454 = n4449 & n7453 ;
  assign n7455 = ~n7448 & ~n7454 ;
  assign n7456 = n4025 & ~n7455 ;
  assign n7469 = n3683 & ~n6609 ;
  assign n7470 = ~n4042 & n4062 ;
  assign n7471 = ~n7469 & n7470 ;
  assign n7472 = n4449 & n7471 ;
  assign n7447 = n3686 & ~n4542 ;
  assign n7473 = n3683 & ~n4522 ;
  assign n7474 = ~n7447 & ~n7473 ;
  assign n7475 = ~n7472 & n7474 ;
  assign n7476 = ~n7456 & n7475 ;
  assign n7457 = ~n3884 & n5430 ;
  assign n7458 = n3884 & ~n5430 ;
  assign n7459 = ~n7457 & ~n7458 ;
  assign n7460 = n4449 & ~n7459 ;
  assign n7461 = ~n7448 & ~n7460 ;
  assign n7462 = n3969 & ~n7461 ;
  assign n7463 = ~n3540 & n5430 ;
  assign n7464 = n3540 & ~n5430 ;
  assign n7465 = ~n7463 & ~n7464 ;
  assign n7466 = n4449 & n7465 ;
  assign n7467 = ~n7448 & ~n7466 ;
  assign n7468 = n3829 & ~n7467 ;
  assign n7477 = ~n7462 & ~n7468 ;
  assign n7478 = n7476 & n7477 ;
  assign n7479 = n2701 & ~n7478 ;
  assign n7480 = ~n7446 & ~n7479 ;
  assign n7481 = \P1_state_reg[0]/NET0131  & ~n7480 ;
  assign n7444 = n3686 & n4552 ;
  assign n7445 = \P1_reg3_reg[13]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7482 = ~n7444 & ~n7445 ;
  assign n7483 = ~n7481 & n7482 ;
  assign n7486 = ~n888 & n2035 ;
  assign n7501 = ~n888 & ~n2124 ;
  assign n7505 = ~n921 & n2239 ;
  assign n7506 = ~n893 & n7505 ;
  assign n7508 = ~n868 & n7506 ;
  assign n7507 = n868 & ~n7506 ;
  assign n7509 = n2263 & ~n7507 ;
  assign n7510 = ~n7508 & n7509 ;
  assign n7511 = ~n921 & ~n2263 ;
  assign n7512 = ~n7510 & ~n7511 ;
  assign n7513 = n2124 & ~n7512 ;
  assign n7514 = ~n7501 & ~n7513 ;
  assign n7515 = n1790 & ~n7514 ;
  assign n7488 = ~n888 & ~n2053 ;
  assign n7489 = n1907 & ~n4281 ;
  assign n7490 = ~n1907 & n4281 ;
  assign n7491 = ~n7489 & ~n7490 ;
  assign n7492 = n2053 & ~n7491 ;
  assign n7493 = ~n7488 & ~n7492 ;
  assign n7494 = ~n2120 & ~n7493 ;
  assign n7487 = ~n909 & n2229 ;
  assign n7516 = ~n888 & ~n2274 ;
  assign n7517 = ~n7487 & ~n7516 ;
  assign n7518 = ~n7494 & n7517 ;
  assign n7495 = n1907 & ~n4240 ;
  assign n7496 = ~n1907 & n4240 ;
  assign n7497 = ~n7495 & ~n7496 ;
  assign n7498 = n2053 & n7497 ;
  assign n7499 = ~n7488 & ~n7498 ;
  assign n7500 = ~n2224 & ~n7499 ;
  assign n7502 = n2124 & n7497 ;
  assign n7503 = ~n7501 & ~n7502 ;
  assign n7504 = n2123 & ~n7503 ;
  assign n7519 = ~n7500 & ~n7504 ;
  assign n7520 = n7518 & n7519 ;
  assign n7521 = ~n7515 & n7520 ;
  assign n7522 = n2037 & ~n7521 ;
  assign n7523 = ~n7486 & ~n7522 ;
  assign n7524 = \P1_state_reg[0]/NET0131  & ~n7523 ;
  assign n7484 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[10]/NET0131  ;
  assign n7485 = ~n888 & n2014 ;
  assign n7525 = ~n7484 & ~n7485 ;
  assign n7526 = ~n7524 & n7525 ;
  assign n7529 = ~n815 & n2035 ;
  assign n7531 = ~n815 & ~n2053 ;
  assign n7532 = n1912 & ~n2293 ;
  assign n7533 = ~n1912 & n2293 ;
  assign n7534 = ~n7532 & ~n7533 ;
  assign n7535 = n2053 & ~n7534 ;
  assign n7536 = ~n7531 & ~n7535 ;
  assign n7537 = ~n2120 & ~n7536 ;
  assign n7544 = ~n815 & ~n2124 ;
  assign n7548 = n783 & ~n2243 ;
  assign n7549 = ~n2244 & n2263 ;
  assign n7550 = ~n7548 & n7549 ;
  assign n7551 = ~n868 & ~n2263 ;
  assign n7552 = ~n7550 & ~n7551 ;
  assign n7553 = n2124 & ~n7552 ;
  assign n7554 = ~n7544 & ~n7553 ;
  assign n7555 = n1790 & ~n7554 ;
  assign n7530 = ~n850 & n2229 ;
  assign n7556 = ~n815 & ~n2274 ;
  assign n7557 = ~n7530 & ~n7556 ;
  assign n7558 = ~n7555 & n7557 ;
  assign n7559 = ~n7537 & n7558 ;
  assign n7538 = n1912 & ~n2340 ;
  assign n7539 = ~n1912 & n2340 ;
  assign n7540 = ~n7538 & ~n7539 ;
  assign n7541 = n2053 & n7540 ;
  assign n7542 = ~n7531 & ~n7541 ;
  assign n7543 = ~n2224 & ~n7542 ;
  assign n7545 = n2124 & n7540 ;
  assign n7546 = ~n7544 & ~n7545 ;
  assign n7547 = n2123 & ~n7546 ;
  assign n7560 = ~n7543 & ~n7547 ;
  assign n7561 = n7559 & n7560 ;
  assign n7562 = n2037 & ~n7561 ;
  assign n7563 = ~n7529 & ~n7562 ;
  assign n7564 = \P1_state_reg[0]/NET0131  & ~n7563 ;
  assign n7527 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[12]/NET0131  ;
  assign n7528 = ~n815 & n2014 ;
  assign n7565 = ~n7527 & ~n7528 ;
  assign n7566 = ~n7564 & n7565 ;
  assign n7569 = ~n777 & n2035 ;
  assign n7571 = ~n777 & ~n2124 ;
  assign n7572 = n1913 & ~n2629 ;
  assign n7573 = ~n1913 & n2629 ;
  assign n7574 = ~n7572 & ~n7573 ;
  assign n7575 = n2124 & ~n7574 ;
  assign n7576 = ~n7571 & ~n7575 ;
  assign n7577 = n2123 & ~n7576 ;
  assign n7589 = n772 & ~n2244 ;
  assign n7588 = ~n772 & n2244 ;
  assign n7590 = n2263 & ~n7588 ;
  assign n7591 = ~n7589 & n7590 ;
  assign n7592 = ~n822 & ~n2263 ;
  assign n7593 = ~n7591 & ~n7592 ;
  assign n7594 = n2124 & ~n7593 ;
  assign n7595 = ~n7571 & ~n7594 ;
  assign n7596 = n1790 & ~n7595 ;
  assign n7570 = ~n811 & n2229 ;
  assign n7597 = ~n777 & ~n2274 ;
  assign n7598 = ~n7570 & ~n7597 ;
  assign n7599 = ~n7596 & n7598 ;
  assign n7600 = ~n7577 & n7599 ;
  assign n7578 = ~n777 & ~n2053 ;
  assign n7579 = n2053 & ~n7574 ;
  assign n7580 = ~n7578 & ~n7579 ;
  assign n7581 = ~n2224 & ~n7580 ;
  assign n7582 = n1913 & ~n2571 ;
  assign n7583 = ~n1913 & n2571 ;
  assign n7584 = ~n7582 & ~n7583 ;
  assign n7585 = n2053 & n7584 ;
  assign n7586 = ~n7578 & ~n7585 ;
  assign n7587 = ~n2120 & ~n7586 ;
  assign n7601 = ~n7581 & ~n7587 ;
  assign n7602 = n7600 & n7601 ;
  assign n7603 = n2037 & ~n7602 ;
  assign n7604 = ~n7569 & ~n7603 ;
  assign n7605 = \P1_state_reg[0]/NET0131  & ~n7604 ;
  assign n7567 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[13]/NET0131  ;
  assign n7568 = ~n777 & n2014 ;
  assign n7606 = ~n7567 & ~n7568 ;
  assign n7607 = ~n7605 & n7606 ;
  assign n7610 = n3296 & n4081 ;
  assign n7612 = n3296 & ~n4449 ;
  assign n7613 = n3879 & ~n5421 ;
  assign n7614 = ~n3879 & n5421 ;
  assign n7615 = ~n7613 & ~n7614 ;
  assign n7616 = n4449 & n7615 ;
  assign n7617 = ~n7612 & ~n7616 ;
  assign n7618 = n3969 & ~n7617 ;
  assign n7633 = n3291 & ~n6604 ;
  assign n7634 = ~n6605 & ~n7633 ;
  assign n7635 = n4449 & n7634 ;
  assign n7636 = ~n7612 & ~n7635 ;
  assign n7637 = n4062 & ~n7636 ;
  assign n7611 = n3291 & ~n4522 ;
  assign n7638 = n3296 & ~n4540 ;
  assign n7639 = ~n7611 & ~n7638 ;
  assign n7640 = ~n7637 & n7639 ;
  assign n7641 = ~n7618 & n7640 ;
  assign n7619 = n3535 & ~n5421 ;
  assign n7620 = ~n3535 & n5421 ;
  assign n7621 = ~n7619 & ~n7620 ;
  assign n7622 = n4449 & ~n7621 ;
  assign n7623 = ~n7612 & ~n7622 ;
  assign n7624 = n3829 & ~n7623 ;
  assign n7625 = n3275 & ~n3994 ;
  assign n7626 = ~n7406 & ~n7625 ;
  assign n7627 = ~n2731 & ~n7626 ;
  assign n7628 = n2731 & n3444 ;
  assign n7629 = ~n7627 & ~n7628 ;
  assign n7630 = n4449 & n7629 ;
  assign n7631 = ~n7612 & ~n7630 ;
  assign n7632 = n4025 & ~n7631 ;
  assign n7642 = ~n7624 & ~n7632 ;
  assign n7643 = n7641 & n7642 ;
  assign n7644 = n2701 & ~n7643 ;
  assign n7645 = ~n7610 & ~n7644 ;
  assign n7646 = \P1_state_reg[0]/NET0131  & ~n7645 ;
  assign n7608 = \P1_reg3_reg[9]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7609 = n3296 & n4552 ;
  assign n7647 = ~n7608 & ~n7609 ;
  assign n7648 = ~n7646 & n7647 ;
  assign n7651 = ~n915 & n2035 ;
  assign n7654 = ~n915 & ~n2124 ;
  assign n7655 = n1927 & ~n2626 ;
  assign n7656 = ~n1927 & n2626 ;
  assign n7657 = ~n7655 & ~n7656 ;
  assign n7658 = n2124 & ~n7657 ;
  assign n7659 = ~n7654 & ~n7658 ;
  assign n7660 = n2123 & ~n7659 ;
  assign n7652 = ~n934 & n2229 ;
  assign n7653 = ~n915 & ~n2274 ;
  assign n7679 = ~n7652 & ~n7653 ;
  assign n7680 = ~n7660 & n7679 ;
  assign n7669 = ~n915 & ~n2053 ;
  assign n7673 = n1927 & ~n2568 ;
  assign n7674 = ~n1927 & n2568 ;
  assign n7675 = ~n7673 & ~n7674 ;
  assign n7676 = n2053 & n7675 ;
  assign n7677 = ~n7669 & ~n7676 ;
  assign n7678 = ~n2120 & ~n7677 ;
  assign n7661 = n893 & ~n7505 ;
  assign n7662 = n2263 & ~n7506 ;
  assign n7663 = ~n7661 & n7662 ;
  assign n7664 = ~n944 & ~n2263 ;
  assign n7665 = ~n7663 & ~n7664 ;
  assign n7666 = n2124 & ~n7665 ;
  assign n7667 = ~n7654 & ~n7666 ;
  assign n7668 = n1790 & ~n7667 ;
  assign n7670 = n2053 & ~n7657 ;
  assign n7671 = ~n7669 & ~n7670 ;
  assign n7672 = ~n2224 & ~n7671 ;
  assign n7681 = ~n7668 & ~n7672 ;
  assign n7682 = ~n7678 & n7681 ;
  assign n7683 = n7680 & n7682 ;
  assign n7684 = n2037 & ~n7683 ;
  assign n7685 = ~n7651 & ~n7684 ;
  assign n7686 = \P1_state_reg[0]/NET0131  & ~n7685 ;
  assign n7649 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[9]/NET0131  ;
  assign n7650 = ~n915 & n2014 ;
  assign n7687 = ~n7649 & ~n7650 ;
  assign n7688 = ~n7686 & n7687 ;
  assign n7689 = n3121 & ~n4449 ;
  assign n7690 = ~n4466 & n4467 ;
  assign n7691 = n4472 & ~n7690 ;
  assign n7692 = n4468 & n4478 ;
  assign n7693 = ~n7691 & n7692 ;
  assign n7694 = ~n4475 & n4478 ;
  assign n7695 = n4453 & ~n7694 ;
  assign n7696 = ~n7693 & n7695 ;
  assign n7697 = n5417 & n7696 ;
  assign n7698 = ~n5417 & ~n7696 ;
  assign n7699 = ~n7697 & ~n7698 ;
  assign n7700 = n4449 & ~n7699 ;
  assign n7701 = ~n7689 & ~n7700 ;
  assign n7702 = n3829 & ~n7701 ;
  assign n7703 = ~n4492 & n4493 ;
  assign n7704 = n4498 & ~n7703 ;
  assign n7705 = n4494 & n4504 ;
  assign n7706 = ~n7704 & n7705 ;
  assign n7707 = ~n4501 & n4504 ;
  assign n7708 = n4509 & ~n7707 ;
  assign n7709 = ~n7706 & n7708 ;
  assign n7710 = n5417 & ~n7709 ;
  assign n7711 = ~n5417 & n7709 ;
  assign n7712 = ~n7710 & ~n7711 ;
  assign n7713 = n4449 & ~n7712 ;
  assign n7714 = ~n7689 & ~n7713 ;
  assign n7715 = n3969 & ~n7714 ;
  assign n7722 = n3105 & ~n5073 ;
  assign n7723 = ~n5074 & ~n7722 ;
  assign n7724 = ~n2731 & ~n7723 ;
  assign n7725 = n2731 & n3153 ;
  assign n7726 = ~n7724 & ~n7725 ;
  assign n7727 = n4449 & n7726 ;
  assign n7728 = ~n7689 & ~n7727 ;
  assign n7729 = n4025 & ~n7728 ;
  assign n7716 = n3119 & n4028 ;
  assign n7717 = n3119 & ~n4051 ;
  assign n7718 = n4062 & ~n5086 ;
  assign n7719 = ~n7717 & n7718 ;
  assign n7720 = ~n7716 & ~n7719 ;
  assign n7721 = n4449 & ~n7720 ;
  assign n7730 = n3119 & n4073 ;
  assign n7731 = n3121 & ~n5991 ;
  assign n7732 = ~n7730 & ~n7731 ;
  assign n7733 = ~n7721 & n7732 ;
  assign n7734 = ~n7729 & n7733 ;
  assign n7735 = ~n7715 & n7734 ;
  assign n7736 = ~n7702 & n7735 ;
  assign n7737 = n2701 & ~n7736 ;
  assign n7738 = n3121 & n4081 ;
  assign n7739 = ~n7737 & ~n7738 ;
  assign n7740 = \P1_state_reg[0]/NET0131  & ~n7739 ;
  assign n7741 = \P1_reg3_reg[23]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7742 = n3121 & n4552 ;
  assign n7743 = ~n7741 & ~n7742 ;
  assign n7744 = ~n7740 & n7743 ;
  assign n7745 = \P1_reg2_reg[16]/NET0131  & ~n4085 ;
  assign n7746 = \P1_reg2_reg[16]/NET0131  & n4081 ;
  assign n7747 = \P1_reg2_reg[16]/NET0131  & ~n2717 ;
  assign n7754 = n2717 & ~n6647 ;
  assign n7755 = ~n7747 & ~n7754 ;
  assign n7756 = n3829 & ~n7755 ;
  assign n7751 = n2717 & ~n6639 ;
  assign n7752 = ~n7747 & ~n7751 ;
  assign n7753 = n3969 & ~n7752 ;
  assign n7748 = n2717 & n6633 ;
  assign n7749 = ~n7747 & ~n7748 ;
  assign n7750 = n4025 & ~n7749 ;
  assign n7758 = n2717 & n6653 ;
  assign n7759 = ~n7747 & ~n7758 ;
  assign n7760 = n4062 & ~n7759 ;
  assign n7762 = n3708 & n4028 ;
  assign n7763 = n2717 & n7762 ;
  assign n7757 = \P1_reg2_reg[16]/NET0131  & ~n5148 ;
  assign n7761 = n3713 & n4073 ;
  assign n7764 = ~n7757 & ~n7761 ;
  assign n7765 = ~n7763 & n7764 ;
  assign n7766 = ~n7760 & n7765 ;
  assign n7767 = ~n7750 & n7766 ;
  assign n7768 = ~n7753 & n7767 ;
  assign n7769 = ~n7756 & n7768 ;
  assign n7770 = n2701 & ~n7769 ;
  assign n7771 = ~n7746 & ~n7770 ;
  assign n7772 = \P1_state_reg[0]/NET0131  & ~n7771 ;
  assign n7773 = ~n7745 & ~n7772 ;
  assign n7774 = \P1_reg2_reg[12]/NET0131  & ~n4085 ;
  assign n7775 = \P1_reg2_reg[12]/NET0131  & n4081 ;
  assign n7777 = \P1_reg2_reg[12]/NET0131  & ~n2717 ;
  assign n7778 = n2717 & n6586 ;
  assign n7779 = ~n7777 & ~n7778 ;
  assign n7780 = n3829 & ~n7779 ;
  assign n7787 = n2717 & n6610 ;
  assign n7788 = ~n7777 & ~n7787 ;
  assign n7789 = n4062 & ~n7788 ;
  assign n7784 = n2717 & n6594 ;
  assign n7785 = ~n7777 & ~n7784 ;
  assign n7786 = n4025 & ~n7785 ;
  assign n7781 = n2717 & ~n6600 ;
  assign n7782 = ~n7777 & ~n7781 ;
  assign n7783 = n3969 & ~n7782 ;
  assign n7791 = n3239 & n4028 ;
  assign n7792 = n2717 & n7791 ;
  assign n7776 = \P1_reg2_reg[12]/NET0131  & ~n5148 ;
  assign n7790 = n3244 & n4073 ;
  assign n7793 = ~n7776 & ~n7790 ;
  assign n7794 = ~n7792 & n7793 ;
  assign n7795 = ~n7783 & n7794 ;
  assign n7796 = ~n7786 & n7795 ;
  assign n7797 = ~n7789 & n7796 ;
  assign n7798 = ~n7780 & n7797 ;
  assign n7799 = n2701 & ~n7798 ;
  assign n7800 = ~n7775 & ~n7799 ;
  assign n7801 = \P1_state_reg[0]/NET0131  & ~n7800 ;
  assign n7802 = ~n7774 & ~n7801 ;
  assign n7803 = \P2_reg0_reg[23]/NET0131  & ~n2286 ;
  assign n7804 = \P2_reg0_reg[23]/NET0131  & n2035 ;
  assign n7805 = \P2_reg0_reg[23]/NET0131  & ~n2053 ;
  assign n7806 = n2053 & ~n6203 ;
  assign n7807 = ~n7805 & ~n7806 ;
  assign n7808 = n1790 & ~n7807 ;
  assign n7809 = ~n6263 & ~n7805 ;
  assign n7810 = n2123 & ~n7809 ;
  assign n7811 = \P2_reg0_reg[23]/NET0131  & ~n2614 ;
  assign n7812 = n2124 & n6235 ;
  assign n7819 = ~n7811 & ~n7812 ;
  assign n7820 = ~n7810 & n7819 ;
  assign n7813 = \P2_reg0_reg[23]/NET0131  & ~n2124 ;
  assign n7814 = n2124 & ~n6228 ;
  assign n7815 = ~n7813 & ~n7814 ;
  assign n7816 = ~n2120 & ~n7815 ;
  assign n7817 = ~n6254 & ~n7813 ;
  assign n7818 = ~n2224 & ~n7817 ;
  assign n7821 = ~n7816 & ~n7818 ;
  assign n7822 = n7820 & n7821 ;
  assign n7823 = ~n7808 & n7822 ;
  assign n7824 = n2037 & ~n7823 ;
  assign n7825 = ~n7804 & ~n7824 ;
  assign n7826 = \P1_state_reg[0]/NET0131  & ~n7825 ;
  assign n7827 = ~n7803 & ~n7826 ;
  assign n7828 = \P1_reg0_reg[12]/NET0131  & ~n4085 ;
  assign n7829 = \P1_reg0_reg[12]/NET0131  & n4081 ;
  assign n7832 = \P1_reg0_reg[12]/NET0131  & ~n4869 ;
  assign n7833 = n4869 & n6586 ;
  assign n7834 = ~n7832 & ~n7833 ;
  assign n7835 = n3829 & ~n7834 ;
  assign n7839 = n4869 & n6594 ;
  assign n7840 = ~n7832 & ~n7839 ;
  assign n7841 = n4025 & ~n7840 ;
  assign n7830 = ~n6611 & ~n7791 ;
  assign n7831 = n4869 & ~n7830 ;
  assign n7836 = n4869 & ~n6600 ;
  assign n7837 = ~n7832 & ~n7836 ;
  assign n7838 = n3969 & ~n7837 ;
  assign n7842 = \P1_reg0_reg[12]/NET0131  & ~n5866 ;
  assign n7843 = ~n7838 & ~n7842 ;
  assign n7844 = ~n7831 & n7843 ;
  assign n7845 = ~n7841 & n7844 ;
  assign n7846 = ~n7835 & n7845 ;
  assign n7847 = n2701 & ~n7846 ;
  assign n7848 = ~n7829 & ~n7847 ;
  assign n7849 = \P1_state_reg[0]/NET0131  & ~n7848 ;
  assign n7850 = ~n7828 & ~n7849 ;
  assign n7851 = \P2_reg1_reg[23]/NET0131  & ~n2286 ;
  assign n7852 = \P2_reg1_reg[23]/NET0131  & n2035 ;
  assign n7853 = \P2_reg1_reg[23]/NET0131  & ~n2291 ;
  assign n7854 = n2291 & ~n6203 ;
  assign n7855 = ~n7853 & ~n7854 ;
  assign n7856 = n1790 & ~n7855 ;
  assign n7857 = \P2_reg1_reg[23]/NET0131  & ~n2310 ;
  assign n7858 = n2310 & n6216 ;
  assign n7859 = ~n7857 & ~n7858 ;
  assign n7860 = ~n2392 & ~n7859 ;
  assign n7865 = \P2_reg1_reg[23]/NET0131  & ~n4099 ;
  assign n7866 = n2310 & n6235 ;
  assign n7867 = ~n7865 & ~n7866 ;
  assign n7868 = ~n7860 & n7867 ;
  assign n7861 = ~n6232 & ~n7857 ;
  assign n7862 = ~n2290 & ~n7861 ;
  assign n7863 = ~n6229 & ~n7853 ;
  assign n7864 = n2314 & ~n7863 ;
  assign n7869 = ~n7862 & ~n7864 ;
  assign n7870 = n7868 & n7869 ;
  assign n7871 = ~n7856 & n7870 ;
  assign n7872 = n2037 & ~n7871 ;
  assign n7873 = ~n7852 & ~n7872 ;
  assign n7874 = \P1_state_reg[0]/NET0131  & ~n7873 ;
  assign n7875 = ~n7851 & ~n7874 ;
  assign n7876 = \P1_reg0_reg[16]/NET0131  & ~n4085 ;
  assign n7877 = \P1_reg0_reg[16]/NET0131  & n4081 ;
  assign n7878 = \P1_reg0_reg[16]/NET0131  & ~n4869 ;
  assign n7885 = n4869 & ~n6647 ;
  assign n7886 = ~n7878 & ~n7885 ;
  assign n7887 = n3829 & ~n7886 ;
  assign n7882 = n4869 & ~n6639 ;
  assign n7883 = ~n7878 & ~n7882 ;
  assign n7884 = n3969 & ~n7883 ;
  assign n7879 = n4869 & n6633 ;
  assign n7880 = ~n7878 & ~n7879 ;
  assign n7881 = n4025 & ~n7880 ;
  assign n7888 = ~n6654 & ~n7762 ;
  assign n7889 = n4869 & ~n7888 ;
  assign n7890 = \P1_reg0_reg[16]/NET0131  & ~n5866 ;
  assign n7891 = ~n7889 & ~n7890 ;
  assign n7892 = ~n7881 & n7891 ;
  assign n7893 = ~n7884 & n7892 ;
  assign n7894 = ~n7887 & n7893 ;
  assign n7895 = n2701 & ~n7894 ;
  assign n7896 = ~n7877 & ~n7895 ;
  assign n7897 = \P1_state_reg[0]/NET0131  & ~n7896 ;
  assign n7898 = ~n7876 & ~n7897 ;
  assign n7899 = \P1_reg0_reg[20]/NET0131  & ~n4085 ;
  assign n7900 = \P1_reg0_reg[20]/NET0131  & n4081 ;
  assign n7902 = \P1_reg0_reg[20]/NET0131  & ~n4869 ;
  assign n7906 = n4869 & ~n6725 ;
  assign n7907 = ~n7902 & ~n7906 ;
  assign n7908 = n3829 & ~n7907 ;
  assign n7903 = n4869 & n6719 ;
  assign n7904 = ~n7902 & ~n7903 ;
  assign n7905 = n4025 & ~n7904 ;
  assign n7909 = n4869 & ~n6731 ;
  assign n7910 = ~n7902 & ~n7909 ;
  assign n7911 = n3969 & ~n7910 ;
  assign n7901 = n4869 & ~n7070 ;
  assign n7912 = \P1_reg0_reg[20]/NET0131  & ~n5866 ;
  assign n7913 = ~n7901 & ~n7912 ;
  assign n7914 = ~n7911 & n7913 ;
  assign n7915 = ~n7905 & n7914 ;
  assign n7916 = ~n7908 & n7915 ;
  assign n7917 = n2701 & ~n7916 ;
  assign n7918 = ~n7900 & ~n7917 ;
  assign n7919 = \P1_state_reg[0]/NET0131  & ~n7918 ;
  assign n7920 = ~n7899 & ~n7919 ;
  assign n7921 = \P1_reg1_reg[12]/NET0131  & ~n4085 ;
  assign n7922 = \P1_reg1_reg[12]/NET0131  & n4081 ;
  assign n7924 = \P1_reg1_reg[12]/NET0131  & ~n4202 ;
  assign n7925 = n4202 & n6586 ;
  assign n7926 = ~n7924 & ~n7925 ;
  assign n7927 = n3829 & ~n7926 ;
  assign n7931 = n4202 & n6594 ;
  assign n7932 = ~n7924 & ~n7931 ;
  assign n7933 = n4025 & ~n7932 ;
  assign n7923 = n4202 & ~n7830 ;
  assign n7928 = n4202 & ~n6600 ;
  assign n7929 = ~n7924 & ~n7928 ;
  assign n7930 = n3969 & ~n7929 ;
  assign n7934 = \P1_reg1_reg[12]/NET0131  & ~n4218 ;
  assign n7935 = ~n7930 & ~n7934 ;
  assign n7936 = ~n7923 & n7935 ;
  assign n7937 = ~n7933 & n7936 ;
  assign n7938 = ~n7927 & n7937 ;
  assign n7939 = n2701 & ~n7938 ;
  assign n7940 = ~n7922 & ~n7939 ;
  assign n7941 = \P1_state_reg[0]/NET0131  & ~n7940 ;
  assign n7942 = ~n7921 & ~n7941 ;
  assign n7943 = \P1_reg1_reg[16]/NET0131  & ~n4085 ;
  assign n7944 = \P1_reg1_reg[16]/NET0131  & n4081 ;
  assign n7945 = \P1_reg1_reg[16]/NET0131  & ~n4202 ;
  assign n7952 = n4202 & ~n6647 ;
  assign n7953 = ~n7945 & ~n7952 ;
  assign n7954 = n3829 & ~n7953 ;
  assign n7949 = n4202 & ~n6639 ;
  assign n7950 = ~n7945 & ~n7949 ;
  assign n7951 = n3969 & ~n7950 ;
  assign n7946 = n4202 & n6633 ;
  assign n7947 = ~n7945 & ~n7946 ;
  assign n7948 = n4025 & ~n7947 ;
  assign n7955 = n4202 & ~n7888 ;
  assign n7956 = \P1_reg1_reg[16]/NET0131  & ~n4218 ;
  assign n7957 = ~n7955 & ~n7956 ;
  assign n7958 = ~n7948 & n7957 ;
  assign n7959 = ~n7951 & n7958 ;
  assign n7960 = ~n7954 & n7959 ;
  assign n7961 = n2701 & ~n7960 ;
  assign n7962 = ~n7944 & ~n7961 ;
  assign n7963 = \P1_state_reg[0]/NET0131  & ~n7962 ;
  assign n7964 = ~n7943 & ~n7963 ;
  assign n7965 = \P1_reg1_reg[20]/NET0131  & ~n4085 ;
  assign n7966 = \P1_reg1_reg[20]/NET0131  & n4081 ;
  assign n7968 = \P1_reg1_reg[20]/NET0131  & ~n4202 ;
  assign n7972 = n4202 & ~n6725 ;
  assign n7973 = ~n7968 & ~n7972 ;
  assign n7974 = n3829 & ~n7973 ;
  assign n7969 = n4202 & n6719 ;
  assign n7970 = ~n7968 & ~n7969 ;
  assign n7971 = n4025 & ~n7970 ;
  assign n7975 = n4202 & ~n6731 ;
  assign n7976 = ~n7968 & ~n7975 ;
  assign n7977 = n3969 & ~n7976 ;
  assign n7978 = n4202 & n6736 ;
  assign n7979 = ~n7968 & ~n7978 ;
  assign n7980 = n4062 & ~n7979 ;
  assign n7967 = n4202 & n7069 ;
  assign n7981 = \P1_reg1_reg[20]/NET0131  & ~n4216 ;
  assign n7982 = ~n7967 & ~n7981 ;
  assign n7983 = ~n7980 & n7982 ;
  assign n7984 = ~n7977 & n7983 ;
  assign n7985 = ~n7971 & n7984 ;
  assign n7986 = ~n7974 & n7985 ;
  assign n7987 = n2701 & ~n7986 ;
  assign n7988 = ~n7966 & ~n7987 ;
  assign n7989 = \P1_state_reg[0]/NET0131  & ~n7988 ;
  assign n7990 = ~n7965 & ~n7989 ;
  assign n7993 = n3214 & n4081 ;
  assign n7995 = n3214 & ~n4449 ;
  assign n7996 = n4466 & ~n5424 ;
  assign n7997 = ~n4466 & n5424 ;
  assign n7998 = ~n7996 & ~n7997 ;
  assign n7999 = n4449 & ~n7998 ;
  assign n8000 = ~n7995 & ~n7999 ;
  assign n8001 = n3829 & ~n8000 ;
  assign n8010 = n4492 & ~n5424 ;
  assign n8011 = ~n4492 & n5424 ;
  assign n8012 = ~n8010 & ~n8011 ;
  assign n8013 = n4449 & n8012 ;
  assign n8014 = ~n7995 & ~n8013 ;
  assign n8015 = n3969 & ~n8014 ;
  assign n8002 = n3248 & ~n7408 ;
  assign n8003 = ~n4942 & ~n8002 ;
  assign n8004 = ~n2731 & ~n8003 ;
  assign n8005 = n2731 & n3275 ;
  assign n8006 = ~n8004 & ~n8005 ;
  assign n8007 = n4449 & n8006 ;
  assign n8008 = ~n7995 & ~n8007 ;
  assign n8009 = n4025 & ~n8008 ;
  assign n8016 = n3211 & ~n6606 ;
  assign n8017 = n4062 & ~n6607 ;
  assign n8018 = ~n8016 & n8017 ;
  assign n8019 = n4449 & n8018 ;
  assign n7994 = n3214 & ~n4542 ;
  assign n8020 = n3211 & ~n4522 ;
  assign n8021 = ~n7994 & ~n8020 ;
  assign n8022 = ~n8019 & n8021 ;
  assign n8023 = ~n8009 & n8022 ;
  assign n8024 = ~n8015 & n8023 ;
  assign n8025 = ~n8001 & n8024 ;
  assign n8026 = n2701 & ~n8025 ;
  assign n8027 = ~n7993 & ~n8026 ;
  assign n8028 = \P1_state_reg[0]/NET0131  & ~n8027 ;
  assign n7991 = \P1_reg3_reg[11]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7992 = n3214 & n4552 ;
  assign n8029 = ~n7991 & ~n7992 ;
  assign n8030 = ~n8028 & n8029 ;
  assign n8039 = n3735 & ~n4449 ;
  assign n8040 = n5418 & ~n7691 ;
  assign n8041 = ~n5418 & n7691 ;
  assign n8042 = ~n8040 & ~n8041 ;
  assign n8043 = n4449 & n8042 ;
  assign n8044 = ~n8039 & ~n8043 ;
  assign n8045 = n3829 & ~n8044 ;
  assign n8046 = n5418 & ~n7704 ;
  assign n8047 = ~n5418 & n7704 ;
  assign n8048 = ~n8046 & ~n8047 ;
  assign n8049 = n4449 & ~n8048 ;
  assign n8050 = ~n8039 & ~n8049 ;
  assign n8051 = n3969 & ~n8050 ;
  assign n8052 = n3717 & ~n4000 ;
  assign n8053 = ~n5965 & ~n8052 ;
  assign n8054 = ~n2731 & ~n8053 ;
  assign n8055 = n2731 & n3665 ;
  assign n8056 = ~n8054 & ~n8055 ;
  assign n8057 = n4449 & n8056 ;
  assign n8058 = ~n8039 & ~n8057 ;
  assign n8059 = n4025 & ~n8058 ;
  assign n8032 = n4062 & ~n6032 ;
  assign n8033 = ~n3732 & ~n8032 ;
  assign n8034 = n4062 & n6032 ;
  assign n8035 = n3732 & ~n4028 ;
  assign n8036 = ~n8034 & n8035 ;
  assign n8037 = ~n8033 & ~n8036 ;
  assign n8038 = n4449 & n8037 ;
  assign n8060 = n3732 & n4073 ;
  assign n8061 = n3735 & ~n5991 ;
  assign n8062 = ~n8060 & ~n8061 ;
  assign n8063 = ~n8038 & n8062 ;
  assign n8064 = ~n8059 & n8063 ;
  assign n8065 = ~n8051 & n8064 ;
  assign n8066 = ~n8045 & n8065 ;
  assign n8067 = n2701 & ~n8066 ;
  assign n8068 = n3735 & n4081 ;
  assign n8069 = ~n8067 & ~n8068 ;
  assign n8070 = \P1_state_reg[0]/NET0131  & ~n8069 ;
  assign n8031 = \P1_reg3_reg[15]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8071 = n3735 & n4552 ;
  assign n8072 = ~n8031 & ~n8071 ;
  assign n8073 = ~n8070 & n8072 ;
  assign n8076 = n3659 & n4081 ;
  assign n8082 = n3659 & ~n4449 ;
  assign n8083 = n3741 & ~n4944 ;
  assign n8084 = ~n4000 & ~n8083 ;
  assign n8085 = ~n2731 & ~n8084 ;
  assign n8086 = n2731 & n3692 ;
  assign n8087 = ~n8085 & ~n8086 ;
  assign n8088 = n4449 & n8087 ;
  assign n8089 = ~n8082 & ~n8088 ;
  assign n8090 = n4025 & ~n8089 ;
  assign n8097 = n5413 & ~n6405 ;
  assign n8098 = ~n5413 & n6405 ;
  assign n8099 = ~n8097 & ~n8098 ;
  assign n8100 = n4449 & ~n8099 ;
  assign n8101 = ~n8082 & ~n8100 ;
  assign n8102 = n3969 & ~n8101 ;
  assign n8091 = n5413 & ~n6393 ;
  assign n8092 = ~n5413 & n6393 ;
  assign n8093 = ~n8091 & ~n8092 ;
  assign n8094 = n4449 & n8093 ;
  assign n8095 = ~n8082 & ~n8094 ;
  assign n8096 = n3829 & ~n8095 ;
  assign n8077 = n3656 & n4028 ;
  assign n8078 = n3656 & ~n4042 ;
  assign n8079 = n8032 & ~n8078 ;
  assign n8080 = ~n8077 & ~n8079 ;
  assign n8081 = n4449 & ~n8080 ;
  assign n8103 = n3656 & n4073 ;
  assign n8104 = n3659 & ~n5991 ;
  assign n8105 = ~n8103 & ~n8104 ;
  assign n8106 = ~n8081 & n8105 ;
  assign n8107 = ~n8096 & n8106 ;
  assign n8108 = ~n8102 & n8107 ;
  assign n8109 = ~n8090 & n8108 ;
  assign n8110 = n2701 & ~n8109 ;
  assign n8111 = ~n8076 & ~n8110 ;
  assign n8112 = \P1_state_reg[0]/NET0131  & ~n8111 ;
  assign n8074 = \P1_reg3_reg[14]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8075 = n3659 & n4552 ;
  assign n8113 = ~n8074 & ~n8075 ;
  assign n8114 = ~n8112 & n8113 ;
  assign n8117 = ~n861 & n2035 ;
  assign n8119 = ~n861 & ~n2053 ;
  assign n8120 = n1902 & ~n2074 ;
  assign n8121 = ~n1902 & n2074 ;
  assign n8122 = ~n8120 & ~n8121 ;
  assign n8123 = n2053 & ~n8122 ;
  assign n8124 = ~n8119 & ~n8123 ;
  assign n8125 = ~n2120 & ~n8124 ;
  assign n8118 = ~n882 & n2229 ;
  assign n8144 = ~n861 & ~n2274 ;
  assign n8145 = ~n8118 & ~n8144 ;
  assign n8146 = ~n8125 & n8145 ;
  assign n8132 = ~n861 & ~n2124 ;
  assign n8136 = ~n893 & ~n2263 ;
  assign n8137 = n822 & ~n7508 ;
  assign n8138 = ~n2243 & n2263 ;
  assign n8139 = ~n8137 & n8138 ;
  assign n8140 = ~n8136 & ~n8139 ;
  assign n8141 = n2124 & ~n8140 ;
  assign n8142 = ~n8132 & ~n8141 ;
  assign n8143 = n1790 & ~n8142 ;
  assign n8126 = n1902 & ~n2166 ;
  assign n8127 = ~n1902 & n2166 ;
  assign n8128 = ~n8126 & ~n8127 ;
  assign n8129 = n2053 & n8128 ;
  assign n8130 = ~n8119 & ~n8129 ;
  assign n8131 = ~n2224 & ~n8130 ;
  assign n8133 = n2124 & n8128 ;
  assign n8134 = ~n8132 & ~n8133 ;
  assign n8135 = n2123 & ~n8134 ;
  assign n8147 = ~n8131 & ~n8135 ;
  assign n8148 = ~n8143 & n8147 ;
  assign n8149 = n8146 & n8148 ;
  assign n8150 = n2037 & ~n8149 ;
  assign n8151 = ~n8117 & ~n8150 ;
  assign n8152 = \P1_state_reg[0]/NET0131  & ~n8151 ;
  assign n8115 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[11]/NET0131  ;
  assign n8116 = ~n861 & n2014 ;
  assign n8153 = ~n8115 & ~n8116 ;
  assign n8154 = ~n8152 & n8153 ;
  assign n8157 = ~n767 & n2035 ;
  assign n8160 = ~n767 & ~n2124 ;
  assign n8161 = n1931 & ~n4245 ;
  assign n8162 = ~n1931 & n4245 ;
  assign n8163 = ~n8161 & ~n8162 ;
  assign n8164 = n2124 & ~n8163 ;
  assign n8165 = ~n8160 & ~n8164 ;
  assign n8166 = n2123 & ~n8165 ;
  assign n8177 = n601 & ~n7588 ;
  assign n8178 = n2244 & n2245 ;
  assign n8179 = n2263 & ~n8178 ;
  assign n8180 = ~n8177 & n8179 ;
  assign n8181 = ~n783 & ~n2263 ;
  assign n8182 = ~n8180 & ~n8181 ;
  assign n8183 = n2124 & ~n8182 ;
  assign n8184 = ~n8160 & ~n8183 ;
  assign n8185 = n1790 & ~n8184 ;
  assign n8158 = ~n760 & n2229 ;
  assign n8159 = ~n767 & ~n2274 ;
  assign n8186 = ~n8158 & ~n8159 ;
  assign n8187 = ~n8185 & n8186 ;
  assign n8188 = ~n8166 & n8187 ;
  assign n8167 = ~n767 & ~n2053 ;
  assign n8168 = n2053 & ~n8163 ;
  assign n8169 = ~n8167 & ~n8168 ;
  assign n8170 = ~n2224 & ~n8169 ;
  assign n8171 = n1931 & ~n4284 ;
  assign n8172 = ~n1931 & n4284 ;
  assign n8173 = ~n8171 & ~n8172 ;
  assign n8174 = n2053 & n8173 ;
  assign n8175 = ~n8167 & ~n8174 ;
  assign n8176 = ~n2120 & ~n8175 ;
  assign n8189 = ~n8170 & ~n8176 ;
  assign n8190 = n8188 & n8189 ;
  assign n8191 = n2037 & ~n8190 ;
  assign n8192 = ~n8157 & ~n8191 ;
  assign n8193 = \P1_state_reg[0]/NET0131  & ~n8192 ;
  assign n8155 = ~n767 & n2014 ;
  assign n8156 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[14]/NET0131  ;
  assign n8194 = ~n8155 & ~n8156 ;
  assign n8195 = ~n8193 & n8194 ;
  assign n8198 = ~n595 & n2035 ;
  assign n8201 = ~n595 & ~n2124 ;
  assign n8210 = n1930 & ~n6208 ;
  assign n8211 = ~n1930 & n6208 ;
  assign n8212 = ~n8210 & ~n8211 ;
  assign n8213 = n2124 & n8212 ;
  assign n8214 = ~n8201 & ~n8213 ;
  assign n8215 = n2123 & ~n8214 ;
  assign n8202 = ~n772 & ~n2263 ;
  assign n8203 = n1231 & ~n8178 ;
  assign n8204 = ~n2247 & n2263 ;
  assign n8205 = ~n8203 & n8204 ;
  assign n8206 = ~n8202 & ~n8205 ;
  assign n8207 = n2124 & ~n8206 ;
  assign n8208 = ~n8201 & ~n8207 ;
  assign n8209 = n1790 & ~n8208 ;
  assign n8199 = ~n718 & n2229 ;
  assign n8200 = ~n595 & ~n2274 ;
  assign n8226 = ~n8199 & ~n8200 ;
  assign n8227 = ~n8209 & n8226 ;
  assign n8228 = ~n8215 & n8227 ;
  assign n8216 = ~n595 & ~n2053 ;
  assign n8217 = n2053 & n8212 ;
  assign n8218 = ~n8216 & ~n8217 ;
  assign n8219 = ~n2224 & ~n8218 ;
  assign n8220 = n1930 & ~n6220 ;
  assign n8221 = ~n1930 & n6220 ;
  assign n8222 = ~n8220 & ~n8221 ;
  assign n8223 = n2053 & ~n8222 ;
  assign n8224 = ~n8216 & ~n8223 ;
  assign n8225 = ~n2120 & ~n8224 ;
  assign n8229 = ~n8219 & ~n8225 ;
  assign n8230 = n8228 & n8229 ;
  assign n8231 = n2037 & ~n8230 ;
  assign n8232 = ~n8198 & ~n8231 ;
  assign n8233 = \P1_state_reg[0]/NET0131  & ~n8232 ;
  assign n8196 = ~n595 & n2014 ;
  assign n8197 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[15]/NET0131  ;
  assign n8234 = ~n8196 & ~n8197 ;
  assign n8235 = ~n8233 & n8234 ;
  assign n8238 = n3440 & n4081 ;
  assign n8252 = n2731 & ~n3470 ;
  assign n8253 = ~n3494 & n3990 ;
  assign n8254 = ~n3470 & n8253 ;
  assign n8255 = ~n3444 & n8254 ;
  assign n8256 = n3300 & ~n8255 ;
  assign n8257 = ~n2731 & ~n3994 ;
  assign n8258 = ~n8256 & n8257 ;
  assign n8259 = ~n8252 & ~n8258 ;
  assign n8260 = n4025 & ~n8259 ;
  assign n8244 = ~n4654 & n5420 ;
  assign n8243 = n4654 & ~n5420 ;
  assign n8245 = n3829 & ~n8243 ;
  assign n8246 = ~n8244 & n8245 ;
  assign n8248 = ~n4733 & ~n5420 ;
  assign n8247 = n4733 & n5420 ;
  assign n8249 = n3969 & ~n8247 ;
  assign n8250 = ~n8248 & n8249 ;
  assign n8251 = ~n8246 & ~n8250 ;
  assign n8261 = n3435 & ~n4036 ;
  assign n8262 = n4062 & ~n6604 ;
  assign n8263 = ~n8261 & n8262 ;
  assign n8264 = n8251 & ~n8263 ;
  assign n8265 = ~n8260 & n8264 ;
  assign n8266 = n4449 & ~n8265 ;
  assign n8239 = n3435 & ~n4522 ;
  assign n8240 = ~n4449 & ~n6183 ;
  assign n8241 = n4542 & ~n8240 ;
  assign n8242 = n3440 & ~n8241 ;
  assign n8267 = ~n8239 & ~n8242 ;
  assign n8268 = ~n8266 & n8267 ;
  assign n8269 = n2701 & ~n8268 ;
  assign n8270 = ~n8238 & ~n8269 ;
  assign n8271 = \P1_state_reg[0]/NET0131  & ~n8270 ;
  assign n8236 = \P1_reg3_reg[8]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8237 = n3440 & n4552 ;
  assign n8272 = ~n8236 & ~n8237 ;
  assign n8273 = ~n8271 & n8272 ;
  assign n8276 = ~n939 & n2035 ;
  assign n8278 = ~n939 & ~n2124 ;
  assign n8279 = n1916 & ~n2329 ;
  assign n8280 = ~n1916 & n2329 ;
  assign n8281 = ~n8279 & ~n8280 ;
  assign n8282 = n2124 & n8281 ;
  assign n8283 = ~n8278 & ~n8282 ;
  assign n8284 = n2123 & ~n8283 ;
  assign n8295 = n921 & ~n2239 ;
  assign n8296 = n2263 & ~n7505 ;
  assign n8297 = ~n8295 & n8296 ;
  assign n8298 = ~n1013 & ~n2263 ;
  assign n8299 = ~n8297 & ~n8298 ;
  assign n8300 = n2124 & ~n8299 ;
  assign n8301 = ~n8278 & ~n8300 ;
  assign n8302 = n1790 & ~n8301 ;
  assign n8277 = ~n958 & n2229 ;
  assign n8303 = ~n939 & ~n2274 ;
  assign n8304 = ~n8277 & ~n8303 ;
  assign n8305 = ~n8302 & n8304 ;
  assign n8306 = ~n8284 & n8305 ;
  assign n8285 = ~n939 & ~n2053 ;
  assign n8286 = n2053 & n8281 ;
  assign n8287 = ~n8285 & ~n8286 ;
  assign n8288 = ~n2224 & ~n8287 ;
  assign n8289 = n1815 & ~n1916 ;
  assign n8290 = ~n1815 & n1916 ;
  assign n8291 = ~n8289 & ~n8290 ;
  assign n8292 = n2053 & ~n8291 ;
  assign n8293 = ~n8285 & ~n8292 ;
  assign n8294 = ~n2120 & ~n8293 ;
  assign n8307 = ~n8288 & ~n8294 ;
  assign n8308 = n8306 & n8307 ;
  assign n8309 = n2037 & ~n8308 ;
  assign n8310 = ~n8276 & ~n8309 ;
  assign n8311 = \P1_state_reg[0]/NET0131  & ~n8310 ;
  assign n8274 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[8]/NET0131  ;
  assign n8275 = ~n939 & n2014 ;
  assign n8312 = ~n8274 & ~n8275 ;
  assign n8313 = ~n8311 & n8312 ;
  assign n8314 = \P1_reg2_reg[10]/NET0131  & ~n4085 ;
  assign n8315 = \P1_reg2_reg[10]/NET0131  & n4081 ;
  assign n8317 = \P1_reg2_reg[10]/NET0131  & ~n2717 ;
  assign n8318 = n2717 & n7412 ;
  assign n8319 = ~n8317 & ~n8318 ;
  assign n8320 = n4025 & ~n8319 ;
  assign n8324 = n2717 & ~n7424 ;
  assign n8325 = ~n8317 & ~n8324 ;
  assign n8326 = n3969 & ~n8325 ;
  assign n8321 = n2717 & n7418 ;
  assign n8322 = ~n8317 & ~n8321 ;
  assign n8323 = n3829 & ~n8322 ;
  assign n8327 = n2717 & n7429 ;
  assign n8328 = ~n8317 & ~n8327 ;
  assign n8329 = n4062 & ~n8328 ;
  assign n8316 = \P1_reg2_reg[10]/NET0131  & ~n5148 ;
  assign n8330 = n3271 & n4073 ;
  assign n8331 = n3263 & n4028 ;
  assign n8332 = n2717 & n8331 ;
  assign n8333 = ~n8330 & ~n8332 ;
  assign n8334 = ~n8316 & n8333 ;
  assign n8335 = ~n8329 & n8334 ;
  assign n8336 = ~n8323 & n8335 ;
  assign n8337 = ~n8326 & n8336 ;
  assign n8338 = ~n8320 & n8337 ;
  assign n8339 = n2701 & ~n8338 ;
  assign n8340 = ~n8315 & ~n8339 ;
  assign n8341 = \P1_state_reg[0]/NET0131  & ~n8340 ;
  assign n8342 = ~n8314 & ~n8341 ;
  assign n8343 = \P1_reg2_reg[13]/NET0131  & ~n4085 ;
  assign n8344 = \P1_reg2_reg[13]/NET0131  & n4081 ;
  assign n8350 = \P1_reg2_reg[13]/NET0131  & ~n2717 ;
  assign n8351 = n2717 & ~n7459 ;
  assign n8352 = ~n8350 & ~n8351 ;
  assign n8353 = n3969 & ~n8352 ;
  assign n8345 = n3683 & n4028 ;
  assign n8346 = ~n7471 & ~n8345 ;
  assign n8347 = n2717 & ~n8346 ;
  assign n8348 = \P1_reg2_reg[13]/NET0131  & ~n7057 ;
  assign n8349 = n3686 & n4073 ;
  assign n8360 = ~n8348 & ~n8349 ;
  assign n8361 = ~n8347 & n8360 ;
  assign n8362 = ~n8353 & n8361 ;
  assign n8354 = n2717 & n7465 ;
  assign n8355 = ~n8350 & ~n8354 ;
  assign n8356 = n3829 & ~n8355 ;
  assign n8357 = n2717 & n7453 ;
  assign n8358 = ~n8350 & ~n8357 ;
  assign n8359 = n4025 & ~n8358 ;
  assign n8363 = ~n8356 & ~n8359 ;
  assign n8364 = n8362 & n8363 ;
  assign n8365 = n2701 & ~n8364 ;
  assign n8366 = ~n8344 & ~n8365 ;
  assign n8367 = \P1_state_reg[0]/NET0131  & ~n8366 ;
  assign n8368 = ~n8343 & ~n8367 ;
  assign n8369 = \P1_reg2_reg[9]/NET0131  & ~n4085 ;
  assign n8370 = \P1_reg2_reg[9]/NET0131  & n4081 ;
  assign n8372 = \P1_reg2_reg[9]/NET0131  & ~n2717 ;
  assign n8373 = n2717 & ~n7621 ;
  assign n8374 = ~n8372 & ~n8373 ;
  assign n8375 = n3829 & ~n8374 ;
  assign n8382 = n2717 & n7634 ;
  assign n8383 = ~n8372 & ~n8382 ;
  assign n8384 = n4062 & ~n8383 ;
  assign n8371 = \P1_reg2_reg[9]/NET0131  & ~n5148 ;
  assign n8385 = n3296 & n4073 ;
  assign n8386 = n3291 & n4028 ;
  assign n8387 = n2717 & n8386 ;
  assign n8388 = ~n8385 & ~n8387 ;
  assign n8389 = ~n8371 & n8388 ;
  assign n8390 = ~n8384 & n8389 ;
  assign n8391 = ~n8375 & n8390 ;
  assign n8376 = n2717 & n7629 ;
  assign n8377 = ~n8372 & ~n8376 ;
  assign n8378 = n4025 & ~n8377 ;
  assign n8379 = n2717 & n7615 ;
  assign n8380 = ~n8372 & ~n8379 ;
  assign n8381 = n3969 & ~n8380 ;
  assign n8392 = ~n8378 & ~n8381 ;
  assign n8393 = n8391 & n8392 ;
  assign n8394 = n2701 & ~n8393 ;
  assign n8395 = ~n8370 & ~n8394 ;
  assign n8396 = \P1_state_reg[0]/NET0131  & ~n8395 ;
  assign n8397 = ~n8369 & ~n8396 ;
  assign n8398 = \P2_reg0_reg[16]/NET0131  & ~n2286 ;
  assign n8399 = \P2_reg0_reg[16]/NET0131  & n2035 ;
  assign n8404 = \P2_reg0_reg[16]/NET0131  & ~n2124 ;
  assign n8405 = ~n6105 & ~n8404 ;
  assign n8406 = ~n2224 & ~n8405 ;
  assign n8401 = \P2_reg0_reg[16]/NET0131  & ~n2053 ;
  assign n8402 = ~n6109 & ~n8401 ;
  assign n8403 = n2123 & ~n8402 ;
  assign n8407 = n2124 & n6114 ;
  assign n8408 = ~n8404 & ~n8407 ;
  assign n8409 = ~n2120 & ~n8408 ;
  assign n8410 = n2053 & ~n6122 ;
  assign n8411 = ~n8401 & ~n8410 ;
  assign n8412 = n1790 & ~n8411 ;
  assign n8400 = ~n1255 & n2616 ;
  assign n8413 = \P2_reg0_reg[16]/NET0131  & ~n2614 ;
  assign n8414 = ~n8400 & ~n8413 ;
  assign n8415 = ~n8412 & n8414 ;
  assign n8416 = ~n8409 & n8415 ;
  assign n8417 = ~n8403 & n8416 ;
  assign n8418 = ~n8406 & n8417 ;
  assign n8419 = n2037 & ~n8418 ;
  assign n8420 = ~n8399 & ~n8419 ;
  assign n8421 = \P1_state_reg[0]/NET0131  & ~n8420 ;
  assign n8422 = ~n8398 & ~n8421 ;
  assign n8423 = \P1_reg1_reg[9]/NET0131  & ~n4085 ;
  assign n8424 = \P1_reg1_reg[9]/NET0131  & n4081 ;
  assign n8426 = \P1_reg1_reg[9]/NET0131  & ~n4202 ;
  assign n8427 = n4202 & n7615 ;
  assign n8428 = ~n8426 & ~n8427 ;
  assign n8429 = n3969 & ~n8428 ;
  assign n8436 = n4202 & n7634 ;
  assign n8437 = ~n8426 & ~n8436 ;
  assign n8438 = n4062 & ~n8437 ;
  assign n8425 = n4202 & n8386 ;
  assign n8439 = \P1_reg1_reg[9]/NET0131  & ~n4216 ;
  assign n8440 = ~n8425 & ~n8439 ;
  assign n8441 = ~n8438 & n8440 ;
  assign n8442 = ~n8429 & n8441 ;
  assign n8430 = n4202 & n7629 ;
  assign n8431 = ~n8426 & ~n8430 ;
  assign n8432 = n4025 & ~n8431 ;
  assign n8433 = n4202 & ~n7621 ;
  assign n8434 = ~n8426 & ~n8433 ;
  assign n8435 = n3829 & ~n8434 ;
  assign n8443 = ~n8432 & ~n8435 ;
  assign n8444 = n8442 & n8443 ;
  assign n8445 = n2701 & ~n8444 ;
  assign n8446 = ~n8424 & ~n8445 ;
  assign n8447 = \P1_state_reg[0]/NET0131  & ~n8446 ;
  assign n8448 = ~n8423 & ~n8447 ;
  assign n8449 = \P2_reg0_reg[9]/NET0131  & ~n2286 ;
  assign n8450 = \P2_reg0_reg[9]/NET0131  & n2035 ;
  assign n8454 = \P2_reg0_reg[9]/NET0131  & ~n2053 ;
  assign n8455 = ~n7670 & ~n8454 ;
  assign n8456 = n2123 & ~n8455 ;
  assign n8451 = ~n934 & n2272 ;
  assign n8452 = n2124 & n8451 ;
  assign n8453 = \P2_reg0_reg[9]/NET0131  & ~n2614 ;
  assign n8466 = ~n8452 & ~n8453 ;
  assign n8467 = ~n8456 & n8466 ;
  assign n8460 = \P2_reg0_reg[9]/NET0131  & ~n2124 ;
  assign n8463 = n2124 & n7675 ;
  assign n8464 = ~n8460 & ~n8463 ;
  assign n8465 = ~n2120 & ~n8464 ;
  assign n8457 = n2053 & ~n7665 ;
  assign n8458 = ~n8454 & ~n8457 ;
  assign n8459 = n1790 & ~n8458 ;
  assign n8461 = ~n7658 & ~n8460 ;
  assign n8462 = ~n2224 & ~n8461 ;
  assign n8468 = ~n8459 & ~n8462 ;
  assign n8469 = ~n8465 & n8468 ;
  assign n8470 = n8467 & n8469 ;
  assign n8471 = n2037 & ~n8470 ;
  assign n8472 = ~n8450 & ~n8471 ;
  assign n8473 = \P1_state_reg[0]/NET0131  & ~n8472 ;
  assign n8474 = ~n8449 & ~n8473 ;
  assign n8475 = \P1_reg2_reg[23]/NET0131  & ~n2717 ;
  assign n8476 = n2717 & ~n7699 ;
  assign n8477 = ~n8475 & ~n8476 ;
  assign n8478 = n3829 & ~n8477 ;
  assign n8479 = n2717 & ~n7712 ;
  assign n8480 = ~n8475 & ~n8479 ;
  assign n8481 = n3969 & ~n8480 ;
  assign n8483 = n2717 & n7726 ;
  assign n8484 = ~n8475 & ~n8483 ;
  assign n8485 = n4025 & ~n8484 ;
  assign n8482 = n2717 & ~n7720 ;
  assign n8486 = n3121 & n4073 ;
  assign n8487 = \P1_reg2_reg[23]/NET0131  & ~n4071 ;
  assign n8488 = ~n8486 & ~n8487 ;
  assign n8489 = ~n8482 & n8488 ;
  assign n8490 = ~n8485 & n8489 ;
  assign n8491 = ~n8481 & n8490 ;
  assign n8492 = ~n8478 & n8491 ;
  assign n8493 = n2701 & ~n8492 ;
  assign n8494 = \P1_reg2_reg[23]/NET0131  & n4081 ;
  assign n8495 = ~n8493 & ~n8494 ;
  assign n8496 = \P1_state_reg[0]/NET0131  & ~n8495 ;
  assign n8497 = \P1_reg2_reg[23]/NET0131  & ~n4085 ;
  assign n8498 = ~n8496 & ~n8497 ;
  assign n8499 = \P2_reg1_reg[10]/NET0131  & ~n2286 ;
  assign n8500 = \P2_reg1_reg[10]/NET0131  & n2035 ;
  assign n8507 = \P2_reg1_reg[10]/NET0131  & ~n2291 ;
  assign n8514 = n2291 & ~n7512 ;
  assign n8515 = ~n8507 & ~n8514 ;
  assign n8516 = n1790 & ~n8515 ;
  assign n8503 = \P2_reg1_reg[10]/NET0131  & ~n2310 ;
  assign n8504 = n2310 & n7497 ;
  assign n8505 = ~n8503 & ~n8504 ;
  assign n8506 = ~n2392 & ~n8505 ;
  assign n8501 = ~n909 & n2272 ;
  assign n8502 = n2310 & n8501 ;
  assign n8517 = \P2_reg1_reg[10]/NET0131  & ~n4099 ;
  assign n8518 = ~n8502 & ~n8517 ;
  assign n8519 = ~n8506 & n8518 ;
  assign n8508 = n2291 & ~n7491 ;
  assign n8509 = ~n8507 & ~n8508 ;
  assign n8510 = n2314 & ~n8509 ;
  assign n8511 = n2310 & ~n7491 ;
  assign n8512 = ~n8503 & ~n8511 ;
  assign n8513 = ~n2290 & ~n8512 ;
  assign n8520 = ~n8510 & ~n8513 ;
  assign n8521 = n8519 & n8520 ;
  assign n8522 = ~n8516 & n8521 ;
  assign n8523 = n2037 & ~n8522 ;
  assign n8524 = ~n8500 & ~n8523 ;
  assign n8525 = \P1_state_reg[0]/NET0131  & ~n8524 ;
  assign n8526 = ~n8499 & ~n8525 ;
  assign n8527 = \P2_reg1_reg[12]/NET0131  & ~n2286 ;
  assign n8528 = \P2_reg1_reg[12]/NET0131  & n2035 ;
  assign n8531 = \P2_reg1_reg[12]/NET0131  & ~n2310 ;
  assign n8532 = n2310 & ~n7534 ;
  assign n8533 = ~n8531 & ~n8532 ;
  assign n8534 = ~n2290 & ~n8533 ;
  assign n8535 = \P2_reg1_reg[12]/NET0131  & ~n2291 ;
  assign n8542 = n2291 & ~n7552 ;
  assign n8543 = ~n8535 & ~n8542 ;
  assign n8544 = n1790 & ~n8543 ;
  assign n8529 = ~n850 & n2272 ;
  assign n8530 = n2310 & n8529 ;
  assign n8545 = \P2_reg1_reg[12]/NET0131  & ~n4099 ;
  assign n8546 = ~n8530 & ~n8545 ;
  assign n8547 = ~n8544 & n8546 ;
  assign n8548 = ~n8534 & n8547 ;
  assign n8536 = n2291 & ~n7534 ;
  assign n8537 = ~n8535 & ~n8536 ;
  assign n8538 = n2314 & ~n8537 ;
  assign n8539 = n2310 & n7540 ;
  assign n8540 = ~n8531 & ~n8539 ;
  assign n8541 = ~n2392 & ~n8540 ;
  assign n8549 = ~n8538 & ~n8541 ;
  assign n8550 = n8548 & n8549 ;
  assign n8551 = n2037 & ~n8550 ;
  assign n8552 = ~n8528 & ~n8551 ;
  assign n8553 = \P1_state_reg[0]/NET0131  & ~n8552 ;
  assign n8554 = ~n8527 & ~n8553 ;
  assign n8555 = \P2_reg1_reg[13]/NET0131  & ~n2286 ;
  assign n8556 = \P2_reg1_reg[13]/NET0131  & n2035 ;
  assign n8559 = \P2_reg1_reg[13]/NET0131  & ~n2310 ;
  assign n8560 = n2310 & ~n7574 ;
  assign n8561 = ~n8559 & ~n8560 ;
  assign n8562 = ~n2392 & ~n8561 ;
  assign n8563 = \P2_reg1_reg[13]/NET0131  & ~n2291 ;
  assign n8570 = n2291 & ~n7593 ;
  assign n8571 = ~n8563 & ~n8570 ;
  assign n8572 = n1790 & ~n8571 ;
  assign n8557 = ~n811 & n2272 ;
  assign n8558 = n2310 & n8557 ;
  assign n8573 = \P2_reg1_reg[13]/NET0131  & ~n4099 ;
  assign n8574 = ~n8558 & ~n8573 ;
  assign n8575 = ~n8572 & n8574 ;
  assign n8576 = ~n8562 & n8575 ;
  assign n8564 = n2291 & n7584 ;
  assign n8565 = ~n8563 & ~n8564 ;
  assign n8566 = n2314 & ~n8565 ;
  assign n8567 = n2310 & n7584 ;
  assign n8568 = ~n8559 & ~n8567 ;
  assign n8569 = ~n2290 & ~n8568 ;
  assign n8577 = ~n8566 & ~n8569 ;
  assign n8578 = n8576 & n8577 ;
  assign n8579 = n2037 & ~n8578 ;
  assign n8580 = ~n8556 & ~n8579 ;
  assign n8581 = \P1_state_reg[0]/NET0131  & ~n8580 ;
  assign n8582 = ~n8555 & ~n8581 ;
  assign n8583 = \P2_reg1_reg[16]/NET0131  & ~n2286 ;
  assign n8584 = \P2_reg1_reg[16]/NET0131  & n2035 ;
  assign n8591 = \P2_reg1_reg[16]/NET0131  & ~n2310 ;
  assign n8595 = n2310 & n6104 ;
  assign n8596 = ~n8591 & ~n8595 ;
  assign n8597 = ~n2392 & ~n8596 ;
  assign n8592 = n2310 & n6114 ;
  assign n8593 = ~n8591 & ~n8592 ;
  assign n8594 = ~n2290 & ~n8593 ;
  assign n8585 = \P2_reg1_reg[16]/NET0131  & ~n2291 ;
  assign n8586 = n2291 & n6114 ;
  assign n8587 = ~n8585 & ~n8586 ;
  assign n8588 = n2314 & ~n8587 ;
  assign n8598 = n2291 & ~n6122 ;
  assign n8599 = ~n8585 & ~n8598 ;
  assign n8600 = n1790 & ~n8599 ;
  assign n8589 = \P2_reg1_reg[16]/NET0131  & ~n4099 ;
  assign n8590 = ~n1255 & n4101 ;
  assign n8601 = ~n8589 & ~n8590 ;
  assign n8602 = ~n8600 & n8601 ;
  assign n8603 = ~n8588 & n8602 ;
  assign n8604 = ~n8594 & n8603 ;
  assign n8605 = ~n8597 & n8604 ;
  assign n8606 = n2037 & ~n8605 ;
  assign n8607 = ~n8584 & ~n8606 ;
  assign n8608 = \P1_state_reg[0]/NET0131  & ~n8607 ;
  assign n8609 = ~n8583 & ~n8608 ;
  assign n8610 = \P1_reg2_reg[30]/NET0131  & ~n4085 ;
  assign n8611 = \P1_reg2_reg[30]/NET0131  & n4081 ;
  assign n8618 = ~n4059 & n5371 ;
  assign n8619 = ~n6166 & ~n8618 ;
  assign n8620 = n2717 & ~n8619 ;
  assign n8617 = ~\P1_reg2_reg[30]/NET0131  & ~n2717 ;
  assign n8621 = n4062 & ~n8617 ;
  assign n8622 = ~n8620 & n8621 ;
  assign n8612 = n2717 & n4028 ;
  assign n8613 = n5371 & n8612 ;
  assign n8614 = ~n2717 & ~n4061 ;
  assign n8615 = ~n4067 & ~n8614 ;
  assign n8616 = \P1_reg2_reg[30]/NET0131  & ~n8615 ;
  assign n8623 = ~n4074 & ~n8616 ;
  assign n8624 = ~n8613 & n8623 ;
  assign n8625 = ~n6179 & n8624 ;
  assign n8626 = ~n8622 & n8625 ;
  assign n8627 = n2701 & ~n8626 ;
  assign n8628 = ~n8611 & ~n8627 ;
  assign n8629 = \P1_state_reg[0]/NET0131  & ~n8628 ;
  assign n8630 = ~n8610 & ~n8629 ;
  assign n8631 = \P2_reg1_reg[9]/NET0131  & ~n2286 ;
  assign n8632 = \P2_reg1_reg[9]/NET0131  & n2035 ;
  assign n8635 = \P2_reg1_reg[9]/NET0131  & ~n2291 ;
  assign n8636 = n2291 & ~n7665 ;
  assign n8637 = ~n8635 & ~n8636 ;
  assign n8638 = n1790 & ~n8637 ;
  assign n8633 = n2310 & n8451 ;
  assign n8634 = \P2_reg1_reg[9]/NET0131  & ~n4099 ;
  assign n8649 = ~n8633 & ~n8634 ;
  assign n8650 = ~n8638 & n8649 ;
  assign n8642 = \P2_reg1_reg[9]/NET0131  & ~n2310 ;
  assign n8646 = n2310 & ~n7657 ;
  assign n8647 = ~n8642 & ~n8646 ;
  assign n8648 = ~n2392 & ~n8647 ;
  assign n8639 = n2291 & n7675 ;
  assign n8640 = ~n8635 & ~n8639 ;
  assign n8641 = n2314 & ~n8640 ;
  assign n8643 = n2310 & n7675 ;
  assign n8644 = ~n8642 & ~n8643 ;
  assign n8645 = ~n2290 & ~n8644 ;
  assign n8651 = ~n8641 & ~n8645 ;
  assign n8652 = ~n8648 & n8651 ;
  assign n8653 = n8650 & n8652 ;
  assign n8654 = n2037 & ~n8653 ;
  assign n8655 = ~n8632 & ~n8654 ;
  assign n8656 = \P1_state_reg[0]/NET0131  & ~n8655 ;
  assign n8657 = ~n8631 & ~n8656 ;
  assign n8658 = \P2_reg2_reg[10]/NET0131  & ~n2286 ;
  assign n8659 = \P2_reg2_reg[10]/NET0131  & n2035 ;
  assign n8665 = \P2_reg2_reg[10]/NET0131  & ~n2310 ;
  assign n8670 = n2310 & ~n7512 ;
  assign n8671 = ~n8665 & ~n8670 ;
  assign n8672 = n1790 & ~n8671 ;
  assign n8661 = \P2_reg2_reg[10]/NET0131  & ~n2291 ;
  assign n8662 = n2291 & n7497 ;
  assign n8663 = ~n8661 & ~n8662 ;
  assign n8664 = ~n2392 & ~n8663 ;
  assign n8674 = \P2_reg2_reg[10]/NET0131  & ~n2407 ;
  assign n8660 = n2291 & n8501 ;
  assign n8673 = ~n888 & n1854 ;
  assign n8675 = ~n8660 & ~n8673 ;
  assign n8676 = ~n8674 & n8675 ;
  assign n8677 = ~n8664 & n8676 ;
  assign n8666 = ~n8511 & ~n8665 ;
  assign n8667 = n2314 & ~n8666 ;
  assign n8668 = ~n8508 & ~n8661 ;
  assign n8669 = ~n2290 & ~n8668 ;
  assign n8678 = ~n8667 & ~n8669 ;
  assign n8679 = n8677 & n8678 ;
  assign n8680 = ~n8672 & n8679 ;
  assign n8681 = n2037 & ~n8680 ;
  assign n8682 = ~n8659 & ~n8681 ;
  assign n8683 = \P1_state_reg[0]/NET0131  & ~n8682 ;
  assign n8684 = ~n8658 & ~n8683 ;
  assign n8685 = \P2_reg2_reg[12]/NET0131  & ~n2286 ;
  assign n8686 = \P2_reg2_reg[12]/NET0131  & n2035 ;
  assign n8688 = \P2_reg2_reg[12]/NET0131  & ~n2291 ;
  assign n8689 = n2291 & n7540 ;
  assign n8690 = ~n8688 & ~n8689 ;
  assign n8691 = ~n2392 & ~n8690 ;
  assign n8692 = \P2_reg2_reg[12]/NET0131  & ~n2310 ;
  assign n8697 = n2310 & ~n7552 ;
  assign n8698 = ~n8692 & ~n8697 ;
  assign n8699 = n1790 & ~n8698 ;
  assign n8700 = \P2_reg2_reg[12]/NET0131  & ~n2407 ;
  assign n8687 = n2291 & n8529 ;
  assign n8701 = ~n815 & n1854 ;
  assign n8702 = ~n8687 & ~n8701 ;
  assign n8703 = ~n8700 & n8702 ;
  assign n8704 = ~n8699 & n8703 ;
  assign n8705 = ~n8691 & n8704 ;
  assign n8693 = ~n8532 & ~n8692 ;
  assign n8694 = n2314 & ~n8693 ;
  assign n8695 = ~n8536 & ~n8688 ;
  assign n8696 = ~n2290 & ~n8695 ;
  assign n8706 = ~n8694 & ~n8696 ;
  assign n8707 = n8705 & n8706 ;
  assign n8708 = n2037 & ~n8707 ;
  assign n8709 = ~n8686 & ~n8708 ;
  assign n8710 = \P1_state_reg[0]/NET0131  & ~n8709 ;
  assign n8711 = ~n8685 & ~n8710 ;
  assign n8712 = \P2_reg2_reg[13]/NET0131  & ~n2286 ;
  assign n8713 = \P2_reg2_reg[13]/NET0131  & n2035 ;
  assign n8719 = \P2_reg2_reg[13]/NET0131  & ~n2291 ;
  assign n8720 = n2291 & ~n7574 ;
  assign n8721 = ~n8719 & ~n8720 ;
  assign n8722 = ~n2392 & ~n8721 ;
  assign n8715 = \P2_reg2_reg[13]/NET0131  & ~n2310 ;
  assign n8716 = n2310 & ~n7593 ;
  assign n8717 = ~n8715 & ~n8716 ;
  assign n8718 = n1790 & ~n8717 ;
  assign n8727 = \P2_reg2_reg[13]/NET0131  & ~n2407 ;
  assign n8714 = n2291 & n8557 ;
  assign n8728 = ~n777 & n1854 ;
  assign n8729 = ~n8714 & ~n8728 ;
  assign n8730 = ~n8727 & n8729 ;
  assign n8731 = ~n8718 & n8730 ;
  assign n8732 = ~n8722 & n8731 ;
  assign n8723 = ~n8567 & ~n8715 ;
  assign n8724 = n2314 & ~n8723 ;
  assign n8725 = ~n8564 & ~n8719 ;
  assign n8726 = ~n2290 & ~n8725 ;
  assign n8733 = ~n8724 & ~n8726 ;
  assign n8734 = n8732 & n8733 ;
  assign n8735 = n2037 & ~n8734 ;
  assign n8736 = ~n8713 & ~n8735 ;
  assign n8737 = \P1_state_reg[0]/NET0131  & ~n8736 ;
  assign n8738 = ~n8712 & ~n8737 ;
  assign n8739 = \P2_reg2_reg[16]/NET0131  & ~n2286 ;
  assign n8740 = \P2_reg2_reg[16]/NET0131  & n2035 ;
  assign n8744 = \P2_reg2_reg[16]/NET0131  & ~n2291 ;
  assign n8747 = n2291 & n6104 ;
  assign n8748 = ~n8744 & ~n8747 ;
  assign n8749 = ~n2392 & ~n8748 ;
  assign n8745 = ~n8586 & ~n8744 ;
  assign n8746 = ~n2290 & ~n8745 ;
  assign n8741 = \P2_reg2_reg[16]/NET0131  & ~n2310 ;
  assign n8742 = ~n8592 & ~n8741 ;
  assign n8743 = n2314 & ~n8742 ;
  assign n8750 = n2310 & ~n6122 ;
  assign n8751 = ~n8741 & ~n8750 ;
  assign n8752 = n1790 & ~n8751 ;
  assign n8755 = \P2_reg2_reg[16]/NET0131  & ~n2407 ;
  assign n8753 = ~n1255 & n2394 ;
  assign n8754 = ~n1226 & n1854 ;
  assign n8756 = ~n8753 & ~n8754 ;
  assign n8757 = ~n8755 & n8756 ;
  assign n8758 = ~n8752 & n8757 ;
  assign n8759 = ~n8743 & n8758 ;
  assign n8760 = ~n8746 & n8759 ;
  assign n8761 = ~n8749 & n8760 ;
  assign n8762 = n2037 & ~n8761 ;
  assign n8763 = ~n8740 & ~n8762 ;
  assign n8764 = \P1_state_reg[0]/NET0131  & ~n8763 ;
  assign n8765 = ~n8739 & ~n8764 ;
  assign n8766 = \P1_reg0_reg[10]/NET0131  & ~n4085 ;
  assign n8767 = \P1_reg0_reg[10]/NET0131  & n4081 ;
  assign n8769 = \P1_reg0_reg[10]/NET0131  & ~n4869 ;
  assign n8770 = n4869 & n7412 ;
  assign n8771 = ~n8769 & ~n8770 ;
  assign n8772 = n4025 & ~n8771 ;
  assign n8776 = n4869 & n7418 ;
  assign n8777 = ~n8769 & ~n8776 ;
  assign n8778 = n3829 & ~n8777 ;
  assign n8773 = n4869 & ~n7424 ;
  assign n8774 = ~n8769 & ~n8773 ;
  assign n8775 = n3969 & ~n8774 ;
  assign n8779 = n4869 & n7429 ;
  assign n8780 = ~n8769 & ~n8779 ;
  assign n8781 = n4062 & ~n8780 ;
  assign n8768 = n4869 & n8331 ;
  assign n8782 = \P1_reg0_reg[10]/NET0131  & ~n5864 ;
  assign n8783 = ~n8768 & ~n8782 ;
  assign n8784 = ~n8781 & n8783 ;
  assign n8785 = ~n8775 & n8784 ;
  assign n8786 = ~n8778 & n8785 ;
  assign n8787 = ~n8772 & n8786 ;
  assign n8788 = n2701 & ~n8787 ;
  assign n8789 = ~n8767 & ~n8788 ;
  assign n8790 = \P1_state_reg[0]/NET0131  & ~n8789 ;
  assign n8791 = ~n8766 & ~n8790 ;
  assign n8792 = \P2_reg2_reg[9]/NET0131  & ~n2286 ;
  assign n8793 = \P2_reg2_reg[9]/NET0131  & n2035 ;
  assign n8795 = \P2_reg2_reg[9]/NET0131  & ~n2310 ;
  assign n8796 = n2310 & ~n7665 ;
  assign n8797 = ~n8795 & ~n8796 ;
  assign n8798 = n1790 & ~n8797 ;
  assign n8808 = \P2_reg2_reg[9]/NET0131  & ~n2407 ;
  assign n8794 = n2291 & n8451 ;
  assign n8807 = ~n915 & n1854 ;
  assign n8809 = ~n8794 & ~n8807 ;
  assign n8810 = ~n8808 & n8809 ;
  assign n8811 = ~n8798 & n8810 ;
  assign n8801 = \P2_reg2_reg[9]/NET0131  & ~n2291 ;
  assign n8804 = n2291 & ~n7657 ;
  assign n8805 = ~n8801 & ~n8804 ;
  assign n8806 = ~n2392 & ~n8805 ;
  assign n8799 = ~n8643 & ~n8795 ;
  assign n8800 = n2314 & ~n8799 ;
  assign n8802 = ~n8639 & ~n8801 ;
  assign n8803 = ~n2290 & ~n8802 ;
  assign n8812 = ~n8800 & ~n8803 ;
  assign n8813 = ~n8806 & n8812 ;
  assign n8814 = n8811 & n8813 ;
  assign n8815 = n2037 & ~n8814 ;
  assign n8816 = ~n8793 & ~n8815 ;
  assign n8817 = \P1_state_reg[0]/NET0131  & ~n8816 ;
  assign n8818 = ~n8792 & ~n8817 ;
  assign n8819 = \P1_reg0_reg[13]/NET0131  & ~n4085 ;
  assign n8820 = \P1_reg0_reg[13]/NET0131  & n4081 ;
  assign n8821 = \P1_reg0_reg[13]/NET0131  & ~n4869 ;
  assign n8822 = n4869 & n7453 ;
  assign n8823 = ~n8821 & ~n8822 ;
  assign n8824 = n4025 & ~n8823 ;
  assign n8825 = \P1_reg0_reg[13]/NET0131  & ~n5866 ;
  assign n8829 = n4869 & ~n8346 ;
  assign n8833 = ~n8825 & ~n8829 ;
  assign n8834 = ~n8824 & n8833 ;
  assign n8826 = n4869 & n7465 ;
  assign n8827 = ~n8821 & ~n8826 ;
  assign n8828 = n3829 & ~n8827 ;
  assign n8830 = n4869 & ~n7459 ;
  assign n8831 = ~n8821 & ~n8830 ;
  assign n8832 = n3969 & ~n8831 ;
  assign n8835 = ~n8828 & ~n8832 ;
  assign n8836 = n8834 & n8835 ;
  assign n8837 = n2701 & ~n8836 ;
  assign n8838 = ~n8820 & ~n8837 ;
  assign n8839 = \P1_state_reg[0]/NET0131  & ~n8838 ;
  assign n8840 = ~n8819 & ~n8839 ;
  assign n8841 = \P1_reg0_reg[23]/NET0131  & ~n4085 ;
  assign n8842 = \P1_reg0_reg[23]/NET0131  & ~n4869 ;
  assign n8843 = n4869 & ~n7699 ;
  assign n8844 = ~n8842 & ~n8843 ;
  assign n8845 = n3829 & ~n8844 ;
  assign n8846 = n4869 & ~n7712 ;
  assign n8847 = ~n8842 & ~n8846 ;
  assign n8848 = n3969 & ~n8847 ;
  assign n8850 = n4869 & n7726 ;
  assign n8851 = ~n8842 & ~n8850 ;
  assign n8852 = n4025 & ~n8851 ;
  assign n8849 = \P1_reg0_reg[23]/NET0131  & ~n5844 ;
  assign n8853 = n4869 & ~n7720 ;
  assign n8854 = ~n8849 & ~n8853 ;
  assign n8855 = ~n8852 & n8854 ;
  assign n8856 = ~n8848 & n8855 ;
  assign n8857 = ~n8845 & n8856 ;
  assign n8858 = n2701 & ~n8857 ;
  assign n8859 = \P1_reg0_reg[23]/NET0131  & n4081 ;
  assign n8860 = ~n8858 & ~n8859 ;
  assign n8861 = \P1_state_reg[0]/NET0131  & ~n8860 ;
  assign n8862 = ~n8841 & ~n8861 ;
  assign n8863 = \P1_reg0_reg[30]/NET0131  & ~n4085 ;
  assign n8864 = \P1_reg0_reg[30]/NET0131  & n4081 ;
  assign n8865 = \P1_reg0_reg[30]/NET0131  & ~n4869 ;
  assign n8870 = n4869 & n8619 ;
  assign n8871 = ~n8865 & ~n8870 ;
  assign n8872 = n4062 & ~n8871 ;
  assign n8866 = n4869 & n5371 ;
  assign n8867 = ~n8865 & ~n8866 ;
  assign n8868 = n4028 & ~n8867 ;
  assign n8869 = \P1_reg0_reg[30]/NET0131  & ~n7304 ;
  assign n8873 = ~n8868 & ~n8869 ;
  assign n8874 = ~n7307 & n8873 ;
  assign n8875 = ~n8872 & n8874 ;
  assign n8876 = n2701 & ~n8875 ;
  assign n8877 = ~n8864 & ~n8876 ;
  assign n8878 = \P1_state_reg[0]/NET0131  & ~n8877 ;
  assign n8879 = ~n8863 & ~n8878 ;
  assign n8880 = \P1_reg0_reg[9]/NET0131  & ~n4085 ;
  assign n8881 = \P1_reg0_reg[9]/NET0131  & n4081 ;
  assign n8883 = \P1_reg0_reg[9]/NET0131  & ~n4869 ;
  assign n8884 = n4869 & n7615 ;
  assign n8885 = ~n8883 & ~n8884 ;
  assign n8886 = n3969 & ~n8885 ;
  assign n8893 = n4869 & n7634 ;
  assign n8894 = ~n8883 & ~n8893 ;
  assign n8895 = n4062 & ~n8894 ;
  assign n8882 = n4869 & n8386 ;
  assign n8896 = \P1_reg0_reg[9]/NET0131  & ~n5864 ;
  assign n8897 = ~n8882 & ~n8896 ;
  assign n8898 = ~n8895 & n8897 ;
  assign n8899 = ~n8886 & n8898 ;
  assign n8887 = n4869 & n7629 ;
  assign n8888 = ~n8883 & ~n8887 ;
  assign n8889 = n4025 & ~n8888 ;
  assign n8890 = n4869 & ~n7621 ;
  assign n8891 = ~n8883 & ~n8890 ;
  assign n8892 = n3829 & ~n8891 ;
  assign n8900 = ~n8889 & ~n8892 ;
  assign n8901 = n8899 & n8900 ;
  assign n8902 = n2701 & ~n8901 ;
  assign n8903 = ~n8881 & ~n8902 ;
  assign n8904 = \P1_state_reg[0]/NET0131  & ~n8903 ;
  assign n8905 = ~n8880 & ~n8904 ;
  assign n8906 = \P1_reg1_reg[10]/NET0131  & ~n4085 ;
  assign n8907 = \P1_reg1_reg[10]/NET0131  & n4081 ;
  assign n8909 = \P1_reg1_reg[10]/NET0131  & ~n4202 ;
  assign n8910 = n4202 & n7412 ;
  assign n8911 = ~n8909 & ~n8910 ;
  assign n8912 = n4025 & ~n8911 ;
  assign n8916 = n4202 & n7418 ;
  assign n8917 = ~n8909 & ~n8916 ;
  assign n8918 = n3829 & ~n8917 ;
  assign n8913 = n4202 & ~n7424 ;
  assign n8914 = ~n8909 & ~n8913 ;
  assign n8915 = n3969 & ~n8914 ;
  assign n8919 = n4202 & n7429 ;
  assign n8920 = ~n8909 & ~n8919 ;
  assign n8921 = n4062 & ~n8920 ;
  assign n8908 = n4202 & n8331 ;
  assign n8922 = \P1_reg1_reg[10]/NET0131  & ~n4216 ;
  assign n8923 = ~n8908 & ~n8922 ;
  assign n8924 = ~n8921 & n8923 ;
  assign n8925 = ~n8915 & n8924 ;
  assign n8926 = ~n8918 & n8925 ;
  assign n8927 = ~n8912 & n8926 ;
  assign n8928 = n2701 & ~n8927 ;
  assign n8929 = ~n8907 & ~n8928 ;
  assign n8930 = \P1_state_reg[0]/NET0131  & ~n8929 ;
  assign n8931 = ~n8906 & ~n8930 ;
  assign n8932 = \P1_reg1_reg[13]/NET0131  & ~n4085 ;
  assign n8933 = \P1_reg1_reg[13]/NET0131  & n4081 ;
  assign n8934 = \P1_reg1_reg[13]/NET0131  & ~n4202 ;
  assign n8935 = n4202 & n7465 ;
  assign n8936 = ~n8934 & ~n8935 ;
  assign n8937 = n3829 & ~n8936 ;
  assign n8938 = n4202 & ~n8346 ;
  assign n8942 = \P1_reg1_reg[13]/NET0131  & ~n4218 ;
  assign n8946 = ~n8938 & ~n8942 ;
  assign n8947 = ~n8937 & n8946 ;
  assign n8939 = n4202 & n7453 ;
  assign n8940 = ~n8934 & ~n8939 ;
  assign n8941 = n4025 & ~n8940 ;
  assign n8943 = n4202 & ~n7459 ;
  assign n8944 = ~n8934 & ~n8943 ;
  assign n8945 = n3969 & ~n8944 ;
  assign n8948 = ~n8941 & ~n8945 ;
  assign n8949 = n8947 & n8948 ;
  assign n8950 = n2701 & ~n8949 ;
  assign n8951 = ~n8933 & ~n8950 ;
  assign n8952 = \P1_state_reg[0]/NET0131  & ~n8951 ;
  assign n8953 = ~n8932 & ~n8952 ;
  assign n8954 = \P1_reg1_reg[23]/NET0131  & ~n4202 ;
  assign n8955 = n4202 & ~n7699 ;
  assign n8956 = ~n8954 & ~n8955 ;
  assign n8957 = n3829 & ~n8956 ;
  assign n8958 = n4202 & ~n7712 ;
  assign n8959 = ~n8954 & ~n8958 ;
  assign n8960 = n3969 & ~n8959 ;
  assign n8962 = n4202 & n7726 ;
  assign n8963 = ~n8954 & ~n8962 ;
  assign n8964 = n4025 & ~n8963 ;
  assign n8961 = n4202 & ~n7720 ;
  assign n8965 = \P1_reg1_reg[23]/NET0131  & ~n6494 ;
  assign n8966 = ~n8961 & ~n8965 ;
  assign n8967 = ~n8964 & n8966 ;
  assign n8968 = ~n8960 & n8967 ;
  assign n8969 = ~n8957 & n8968 ;
  assign n8970 = n2701 & ~n8969 ;
  assign n8971 = \P1_reg1_reg[23]/NET0131  & n4081 ;
  assign n8972 = ~n8970 & ~n8971 ;
  assign n8973 = \P1_state_reg[0]/NET0131  & ~n8972 ;
  assign n8974 = \P1_reg1_reg[23]/NET0131  & ~n4085 ;
  assign n8975 = ~n8973 & ~n8974 ;
  assign n8976 = \P2_reg0_reg[10]/NET0131  & ~n2286 ;
  assign n8977 = \P2_reg0_reg[10]/NET0131  & n2035 ;
  assign n8985 = \P2_reg0_reg[10]/NET0131  & ~n2053 ;
  assign n8988 = n2053 & ~n7512 ;
  assign n8989 = ~n8985 & ~n8988 ;
  assign n8990 = n1790 & ~n8989 ;
  assign n8979 = \P2_reg0_reg[10]/NET0131  & ~n2124 ;
  assign n8980 = ~n7502 & ~n8979 ;
  assign n8981 = ~n2224 & ~n8980 ;
  assign n8978 = n2124 & n8501 ;
  assign n8991 = \P2_reg0_reg[10]/NET0131  & ~n2614 ;
  assign n8992 = ~n8978 & ~n8991 ;
  assign n8993 = ~n8981 & n8992 ;
  assign n8982 = n2124 & ~n7491 ;
  assign n8983 = ~n8979 & ~n8982 ;
  assign n8984 = ~n2120 & ~n8983 ;
  assign n8986 = ~n7498 & ~n8985 ;
  assign n8987 = n2123 & ~n8986 ;
  assign n8994 = ~n8984 & ~n8987 ;
  assign n8995 = n8993 & n8994 ;
  assign n8996 = ~n8990 & n8995 ;
  assign n8997 = n2037 & ~n8996 ;
  assign n8998 = ~n8977 & ~n8997 ;
  assign n8999 = \P1_state_reg[0]/NET0131  & ~n8998 ;
  assign n9000 = ~n8976 & ~n8999 ;
  assign n9001 = \P2_reg0_reg[12]/NET0131  & ~n2286 ;
  assign n9002 = \P2_reg0_reg[12]/NET0131  & n2035 ;
  assign n9004 = \P2_reg0_reg[12]/NET0131  & ~n2124 ;
  assign n9005 = n2124 & ~n7534 ;
  assign n9006 = ~n9004 & ~n9005 ;
  assign n9007 = ~n2120 & ~n9006 ;
  assign n9010 = \P2_reg0_reg[12]/NET0131  & ~n2053 ;
  assign n9013 = n2053 & ~n7552 ;
  assign n9014 = ~n9010 & ~n9013 ;
  assign n9015 = n1790 & ~n9014 ;
  assign n9003 = n2124 & n8529 ;
  assign n9016 = \P2_reg0_reg[12]/NET0131  & ~n2614 ;
  assign n9017 = ~n9003 & ~n9016 ;
  assign n9018 = ~n9015 & n9017 ;
  assign n9019 = ~n9007 & n9018 ;
  assign n9008 = ~n7545 & ~n9004 ;
  assign n9009 = ~n2224 & ~n9008 ;
  assign n9011 = ~n7541 & ~n9010 ;
  assign n9012 = n2123 & ~n9011 ;
  assign n9020 = ~n9009 & ~n9012 ;
  assign n9021 = n9019 & n9020 ;
  assign n9022 = n2037 & ~n9021 ;
  assign n9023 = ~n9002 & ~n9022 ;
  assign n9024 = \P1_state_reg[0]/NET0131  & ~n9023 ;
  assign n9025 = ~n9001 & ~n9024 ;
  assign n9026 = \P2_reg0_reg[13]/NET0131  & ~n2286 ;
  assign n9027 = \P2_reg0_reg[13]/NET0131  & n2035 ;
  assign n9029 = \P2_reg0_reg[13]/NET0131  & ~n2124 ;
  assign n9030 = ~n7575 & ~n9029 ;
  assign n9031 = ~n2224 & ~n9030 ;
  assign n9032 = \P2_reg0_reg[13]/NET0131  & ~n2053 ;
  assign n9038 = n2053 & ~n7593 ;
  assign n9039 = ~n9032 & ~n9038 ;
  assign n9040 = n1790 & ~n9039 ;
  assign n9028 = n2124 & n8557 ;
  assign n9041 = \P2_reg0_reg[13]/NET0131  & ~n2614 ;
  assign n9042 = ~n9028 & ~n9041 ;
  assign n9043 = ~n9040 & n9042 ;
  assign n9044 = ~n9031 & n9043 ;
  assign n9033 = ~n7579 & ~n9032 ;
  assign n9034 = n2123 & ~n9033 ;
  assign n9035 = n2124 & n7584 ;
  assign n9036 = ~n9029 & ~n9035 ;
  assign n9037 = ~n2120 & ~n9036 ;
  assign n9045 = ~n9034 & ~n9037 ;
  assign n9046 = n9044 & n9045 ;
  assign n9047 = n2037 & ~n9046 ;
  assign n9048 = ~n9027 & ~n9047 ;
  assign n9049 = \P1_state_reg[0]/NET0131  & ~n9048 ;
  assign n9050 = ~n9026 & ~n9049 ;
  assign n9051 = \P1_reg1_reg[30]/NET0131  & ~n4085 ;
  assign n9052 = \P1_reg1_reg[30]/NET0131  & n4081 ;
  assign n9053 = \P1_reg1_reg[30]/NET0131  & ~n4202 ;
  assign n9058 = n4202 & n8619 ;
  assign n9059 = ~n9053 & ~n9058 ;
  assign n9060 = n4062 & ~n9059 ;
  assign n9054 = n4202 & n5371 ;
  assign n9055 = ~n9053 & ~n9054 ;
  assign n9056 = n4028 & ~n9055 ;
  assign n9057 = \P1_reg1_reg[30]/NET0131  & ~n6943 ;
  assign n9061 = ~n9056 & ~n9057 ;
  assign n9062 = ~n6946 & n9061 ;
  assign n9063 = ~n9060 & n9062 ;
  assign n9064 = n2701 & ~n9063 ;
  assign n9065 = ~n9052 & ~n9064 ;
  assign n9066 = \P1_state_reg[0]/NET0131  & ~n9065 ;
  assign n9067 = ~n9051 & ~n9066 ;
  assign n9070 = n3312 & n4081 ;
  assign n9072 = n3312 & ~n4449 ;
  assign n9085 = n3520 & ~n3989 ;
  assign n9086 = ~n3990 & ~n9085 ;
  assign n9087 = ~n2731 & ~n9086 ;
  assign n9088 = n523 & n2731 ;
  assign n9089 = ~n9087 & ~n9088 ;
  assign n9090 = n4449 & n9089 ;
  assign n9091 = ~n9072 & ~n9090 ;
  assign n9092 = n4025 & ~n9091 ;
  assign n9079 = ~n4729 & n5416 ;
  assign n9080 = n4729 & ~n5416 ;
  assign n9081 = ~n9079 & ~n9080 ;
  assign n9082 = n4449 & n9081 ;
  assign n9083 = ~n9072 & ~n9082 ;
  assign n9084 = n3969 & ~n9083 ;
  assign n9073 = ~n4645 & n5416 ;
  assign n9074 = n4645 & ~n5416 ;
  assign n9075 = ~n9073 & ~n9074 ;
  assign n9076 = n4449 & ~n9075 ;
  assign n9077 = ~n9072 & ~n9076 ;
  assign n9078 = n3829 & ~n9077 ;
  assign n9093 = ~n3332 & ~n4032 ;
  assign n9094 = ~n4033 & ~n9093 ;
  assign n9095 = n4449 & n9094 ;
  assign n9096 = ~n9072 & ~n9095 ;
  assign n9097 = n4062 & ~n9096 ;
  assign n9071 = ~n3332 & ~n4522 ;
  assign n9098 = n3312 & ~n4540 ;
  assign n9099 = ~n9071 & ~n9098 ;
  assign n9100 = ~n9097 & n9099 ;
  assign n9101 = ~n9078 & n9100 ;
  assign n9102 = ~n9084 & n9101 ;
  assign n9103 = ~n9092 & n9102 ;
  assign n9104 = n2701 & ~n9103 ;
  assign n9105 = ~n9070 & ~n9104 ;
  assign n9106 = \P1_state_reg[0]/NET0131  & ~n9105 ;
  assign n9068 = \P1_reg3_reg[4]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9069 = n3312 & n4552 ;
  assign n9107 = ~n9068 & ~n9069 ;
  assign n9108 = ~n9106 & n9107 ;
  assign n9111 = n3516 & ~n4449 ;
  assign n9112 = n3494 & ~n3990 ;
  assign n9113 = ~n8253 & ~n9112 ;
  assign n9114 = ~n2731 & ~n9113 ;
  assign n9115 = n2731 & n3318 ;
  assign n9116 = ~n9114 & ~n9115 ;
  assign n9117 = n4449 & n9116 ;
  assign n9118 = ~n9111 & ~n9117 ;
  assign n9119 = n4025 & ~n9118 ;
  assign n9120 = n3421 & ~n5422 ;
  assign n9121 = ~n3421 & n5422 ;
  assign n9122 = ~n9120 & ~n9121 ;
  assign n9123 = n4449 & ~n9122 ;
  assign n9124 = ~n9111 & ~n9123 ;
  assign n9125 = n3829 & ~n9124 ;
  assign n9126 = ~n3859 & ~n3861 ;
  assign n9127 = n5422 & ~n9126 ;
  assign n9128 = ~n5422 & n9126 ;
  assign n9129 = ~n9127 & ~n9128 ;
  assign n9130 = n4449 & n9129 ;
  assign n9131 = ~n9111 & ~n9130 ;
  assign n9132 = n3969 & ~n9131 ;
  assign n9134 = ~n3511 & ~n4033 ;
  assign n9133 = n3511 & n4033 ;
  assign n9135 = n4062 & ~n9133 ;
  assign n9136 = ~n9134 & n9135 ;
  assign n9137 = n4449 & n9136 ;
  assign n9110 = n3516 & ~n4542 ;
  assign n9138 = ~n3511 & ~n4522 ;
  assign n9139 = ~n9110 & ~n9138 ;
  assign n9140 = ~n9137 & n9139 ;
  assign n9141 = ~n9132 & n9140 ;
  assign n9142 = ~n9125 & n9141 ;
  assign n9143 = ~n9119 & n9142 ;
  assign n9144 = n2701 & ~n9143 ;
  assign n9145 = n3516 & n4081 ;
  assign n9146 = ~n9144 & ~n9145 ;
  assign n9147 = \P1_state_reg[0]/NET0131  & ~n9146 ;
  assign n9109 = \P1_reg3_reg[5]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9148 = n3516 & n4552 ;
  assign n9149 = ~n9109 & ~n9148 ;
  assign n9150 = ~n9147 & n9149 ;
  assign n9153 = ~n1030 & n2035 ;
  assign n9164 = ~n1030 & ~n2124 ;
  assign n9171 = ~n1062 & ~n2263 ;
  assign n9172 = ~n1086 & n2233 ;
  assign n9173 = ~n1062 & n9172 ;
  assign n9174 = ~n1037 & n9173 ;
  assign n9175 = n986 & ~n9174 ;
  assign n9176 = ~n2237 & n2263 ;
  assign n9177 = ~n9175 & n9176 ;
  assign n9178 = ~n9171 & ~n9177 ;
  assign n9179 = n2124 & ~n9178 ;
  assign n9180 = ~n9164 & ~n9179 ;
  assign n9181 = n1790 & ~n9180 ;
  assign n9155 = ~n1030 & ~n2053 ;
  assign n9156 = ~n1077 & ~n2061 ;
  assign n9157 = n1909 & n9156 ;
  assign n9158 = ~n1909 & ~n9156 ;
  assign n9159 = ~n9157 & ~n9158 ;
  assign n9160 = n2053 & n9159 ;
  assign n9161 = ~n9155 & ~n9160 ;
  assign n9162 = ~n2120 & ~n9161 ;
  assign n9165 = n1909 & ~n2145 ;
  assign n9166 = ~n1909 & n2145 ;
  assign n9167 = ~n9165 & ~n9166 ;
  assign n9182 = n2053 & ~n9167 ;
  assign n9183 = ~n9155 & ~n9182 ;
  assign n9184 = ~n2224 & ~n9183 ;
  assign n9168 = n2124 & ~n9167 ;
  assign n9169 = ~n9164 & ~n9168 ;
  assign n9170 = n2123 & ~n9169 ;
  assign n9154 = ~n1050 & n2229 ;
  assign n9163 = ~n1030 & ~n2274 ;
  assign n9185 = ~n9154 & ~n9163 ;
  assign n9186 = ~n9170 & n9185 ;
  assign n9187 = ~n9184 & n9186 ;
  assign n9188 = ~n9162 & n9187 ;
  assign n9189 = ~n9181 & n9188 ;
  assign n9190 = n2037 & ~n9189 ;
  assign n9191 = ~n9153 & ~n9190 ;
  assign n9192 = \P1_state_reg[0]/NET0131  & ~n9191 ;
  assign n9151 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[5]/NET0131  ;
  assign n9152 = ~n1030 & n2014 ;
  assign n9193 = ~n9151 & ~n9152 ;
  assign n9194 = ~n9192 & n9193 ;
  assign n9197 = ~n981 & n2035 ;
  assign n9200 = ~n981 & ~n2053 ;
  assign n9201 = n1920 & ~n2325 ;
  assign n9202 = ~n1920 & n2325 ;
  assign n9203 = ~n9201 & ~n9202 ;
  assign n9204 = n2053 & n9203 ;
  assign n9205 = ~n9200 & ~n9204 ;
  assign n9206 = ~n2224 & ~n9205 ;
  assign n9198 = ~n1003 & n2229 ;
  assign n9199 = ~n981 & ~n2274 ;
  assign n9226 = ~n9198 & ~n9199 ;
  assign n9227 = ~n9206 & n9226 ;
  assign n9220 = n1811 & ~n1920 ;
  assign n9221 = ~n1811 & n1920 ;
  assign n9222 = ~n9220 & ~n9221 ;
  assign n9223 = n2053 & ~n9222 ;
  assign n9224 = ~n9200 & ~n9223 ;
  assign n9225 = ~n2120 & ~n9224 ;
  assign n9207 = ~n981 & ~n2124 ;
  assign n9208 = n2124 & n9203 ;
  assign n9209 = ~n9207 & ~n9208 ;
  assign n9210 = n2123 & ~n9209 ;
  assign n9212 = n1013 & ~n2237 ;
  assign n9211 = ~n1013 & n2237 ;
  assign n9213 = n2263 & ~n9211 ;
  assign n9214 = ~n9212 & n9213 ;
  assign n9215 = ~n1037 & ~n2263 ;
  assign n9216 = ~n9214 & ~n9215 ;
  assign n9217 = n2124 & ~n9216 ;
  assign n9218 = ~n9207 & ~n9217 ;
  assign n9219 = n1790 & ~n9218 ;
  assign n9228 = ~n9210 & ~n9219 ;
  assign n9229 = ~n9225 & n9228 ;
  assign n9230 = n9227 & n9229 ;
  assign n9231 = n2037 & ~n9230 ;
  assign n9232 = ~n9197 & ~n9231 ;
  assign n9233 = \P1_state_reg[0]/NET0131  & ~n9232 ;
  assign n9195 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[6]/NET0131  ;
  assign n9196 = ~n981 & n2014 ;
  assign n9234 = ~n9195 & ~n9196 ;
  assign n9235 = ~n9233 & n9234 ;
  assign n9238 = ~n1007 & n2035 ;
  assign n9240 = ~n1007 & ~n2053 ;
  assign n9241 = n1903 & ~n2151 ;
  assign n9242 = ~n1903 & n2151 ;
  assign n9243 = ~n9241 & ~n9242 ;
  assign n9244 = n2053 & ~n9243 ;
  assign n9245 = ~n9240 & ~n9244 ;
  assign n9246 = ~n2224 & ~n9245 ;
  assign n9247 = ~n1007 & ~n2124 ;
  assign n9257 = ~n986 & ~n2263 ;
  assign n9258 = n944 & ~n9211 ;
  assign n9259 = ~n2239 & n2263 ;
  assign n9260 = ~n9258 & n9259 ;
  assign n9261 = ~n9257 & ~n9260 ;
  assign n9262 = n2124 & ~n9261 ;
  assign n9263 = ~n9247 & ~n9262 ;
  assign n9264 = n1790 & ~n9263 ;
  assign n9239 = ~n1026 & n2229 ;
  assign n9265 = ~n1007 & ~n2274 ;
  assign n9266 = ~n9239 & ~n9265 ;
  assign n9267 = ~n9264 & n9266 ;
  assign n9268 = ~n9246 & n9267 ;
  assign n9248 = n2124 & ~n9243 ;
  assign n9249 = ~n9247 & ~n9248 ;
  assign n9250 = n2123 & ~n9249 ;
  assign n9251 = n1903 & ~n2064 ;
  assign n9252 = ~n1903 & n2064 ;
  assign n9253 = ~n9251 & ~n9252 ;
  assign n9254 = n2053 & n9253 ;
  assign n9255 = ~n9240 & ~n9254 ;
  assign n9256 = ~n2120 & ~n9255 ;
  assign n9269 = ~n9250 & ~n9256 ;
  assign n9270 = n9268 & n9269 ;
  assign n9271 = n2037 & ~n9270 ;
  assign n9272 = ~n9238 & ~n9271 ;
  assign n9273 = \P1_state_reg[0]/NET0131  & ~n9272 ;
  assign n9236 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[7]/NET0131  ;
  assign n9237 = ~n1007 & n2014 ;
  assign n9274 = ~n9236 & ~n9237 ;
  assign n9275 = ~n9273 & n9274 ;
  assign n9276 = \P1_reg1_reg[4]/NET0131  & ~n4085 ;
  assign n9277 = \P1_reg1_reg[4]/NET0131  & n4081 ;
  assign n9280 = \P1_reg1_reg[4]/NET0131  & ~n4202 ;
  assign n9287 = n4202 & n9089 ;
  assign n9288 = ~n9280 & ~n9287 ;
  assign n9289 = n4025 & ~n9288 ;
  assign n9284 = n4202 & n9081 ;
  assign n9285 = ~n9280 & ~n9284 ;
  assign n9286 = n3969 & ~n9285 ;
  assign n9281 = n4202 & ~n9075 ;
  assign n9282 = ~n9280 & ~n9281 ;
  assign n9283 = n3829 & ~n9282 ;
  assign n9290 = n4202 & n9094 ;
  assign n9291 = ~n9280 & ~n9290 ;
  assign n9292 = n4062 & ~n9291 ;
  assign n9278 = ~n3332 & n4028 ;
  assign n9279 = n4202 & n9278 ;
  assign n9293 = \P1_reg1_reg[4]/NET0131  & ~n4216 ;
  assign n9294 = ~n9279 & ~n9293 ;
  assign n9295 = ~n9292 & n9294 ;
  assign n9296 = ~n9283 & n9295 ;
  assign n9297 = ~n9286 & n9296 ;
  assign n9298 = ~n9289 & n9297 ;
  assign n9299 = n2701 & ~n9298 ;
  assign n9300 = ~n9277 & ~n9299 ;
  assign n9301 = \P1_state_reg[0]/NET0131  & ~n9300 ;
  assign n9302 = ~n9276 & ~n9301 ;
  assign n9303 = \P1_reg0_reg[4]/NET0131  & ~n4085 ;
  assign n9304 = \P1_reg0_reg[4]/NET0131  & n4081 ;
  assign n9306 = \P1_reg0_reg[4]/NET0131  & ~n4869 ;
  assign n9313 = n4869 & n9089 ;
  assign n9314 = ~n9306 & ~n9313 ;
  assign n9315 = n4025 & ~n9314 ;
  assign n9310 = n4869 & n9081 ;
  assign n9311 = ~n9306 & ~n9310 ;
  assign n9312 = n3969 & ~n9311 ;
  assign n9307 = n4869 & ~n9075 ;
  assign n9308 = ~n9306 & ~n9307 ;
  assign n9309 = n3829 & ~n9308 ;
  assign n9316 = n4869 & n9094 ;
  assign n9317 = ~n9306 & ~n9316 ;
  assign n9318 = n4062 & ~n9317 ;
  assign n9305 = n4869 & n9278 ;
  assign n9319 = \P1_reg0_reg[4]/NET0131  & ~n5864 ;
  assign n9320 = ~n9305 & ~n9319 ;
  assign n9321 = ~n9318 & n9320 ;
  assign n9322 = ~n9309 & n9321 ;
  assign n9323 = ~n9312 & n9322 ;
  assign n9324 = ~n9315 & n9323 ;
  assign n9325 = n2701 & ~n9324 ;
  assign n9326 = ~n9304 & ~n9325 ;
  assign n9327 = \P1_state_reg[0]/NET0131  & ~n9326 ;
  assign n9328 = ~n9303 & ~n9327 ;
  assign n9330 = ~\P1_reg2_reg[8]/NET0131  & ~n2717 ;
  assign n9331 = \P1_state_reg[0]/NET0131  & n2701 ;
  assign n9332 = n8251 & n9331 ;
  assign n9333 = ~n8260 & n9332 ;
  assign n9334 = ~n9330 & ~n9333 ;
  assign n9335 = ~n4036 & n4062 ;
  assign n9336 = ~n3435 & ~n9335 ;
  assign n9337 = n4036 & n4062 ;
  assign n9338 = n3435 & ~n4028 ;
  assign n9339 = ~n9337 & n9338 ;
  assign n9340 = ~n9336 & ~n9339 ;
  assign n9341 = n2717 & n9340 ;
  assign n9329 = n3440 & n4073 ;
  assign n9342 = n4071 & ~n6184 ;
  assign n9343 = \P1_reg2_reg[8]/NET0131  & ~n9342 ;
  assign n9344 = ~n9329 & ~n9343 ;
  assign n9345 = ~n9341 & n9344 ;
  assign n9346 = ~n9334 & n9345 ;
  assign n9347 = ~\P1_reg2_reg[8]/NET0131  & ~n9331 ;
  assign n9348 = ~n9346 & ~n9347 ;
  assign n9349 = \P2_reg0_reg[15]/NET0131  & ~n2286 ;
  assign n9350 = \P2_reg0_reg[15]/NET0131  & n2035 ;
  assign n9354 = \P2_reg0_reg[15]/NET0131  & ~n2053 ;
  assign n9358 = ~n8217 & ~n9354 ;
  assign n9359 = n2123 & ~n9358 ;
  assign n9355 = n2053 & ~n8206 ;
  assign n9356 = ~n9354 & ~n9355 ;
  assign n9357 = n1790 & ~n9356 ;
  assign n9351 = ~n718 & n2272 ;
  assign n9352 = n2124 & n9351 ;
  assign n9353 = \P2_reg0_reg[15]/NET0131  & ~n2614 ;
  assign n9366 = ~n9352 & ~n9353 ;
  assign n9367 = ~n9357 & n9366 ;
  assign n9368 = ~n9359 & n9367 ;
  assign n9360 = \P2_reg0_reg[15]/NET0131  & ~n2124 ;
  assign n9361 = ~n8213 & ~n9360 ;
  assign n9362 = ~n2224 & ~n9361 ;
  assign n9363 = n2124 & ~n8222 ;
  assign n9364 = ~n9360 & ~n9363 ;
  assign n9365 = ~n2120 & ~n9364 ;
  assign n9369 = ~n9362 & ~n9365 ;
  assign n9370 = n9368 & n9369 ;
  assign n9371 = n2037 & ~n9370 ;
  assign n9372 = ~n9350 & ~n9371 ;
  assign n9373 = \P1_state_reg[0]/NET0131  & ~n9372 ;
  assign n9374 = ~n9349 & ~n9373 ;
  assign n9376 = n4202 & n8259 ;
  assign n9377 = n4025 & ~n9376 ;
  assign n9375 = n4202 & n9340 ;
  assign n9378 = n3816 & ~n4202 ;
  assign n9379 = ~n9375 & ~n9378 ;
  assign n9380 = n9332 & n9379 ;
  assign n9381 = ~n9377 & n9380 ;
  assign n9382 = n6494 & n9381 ;
  assign n9383 = n4202 & n9331 ;
  assign n9384 = ~n9381 & n9383 ;
  assign n9385 = ~\P1_reg1_reg[8]/NET0131  & ~n9384 ;
  assign n9386 = ~n9382 & ~n9385 ;
  assign n9387 = \P1_reg2_reg[11]/NET0131  & ~n4085 ;
  assign n9388 = \P1_reg2_reg[11]/NET0131  & n4081 ;
  assign n9392 = \P1_reg2_reg[11]/NET0131  & ~n2717 ;
  assign n9393 = n2717 & ~n7998 ;
  assign n9394 = ~n9392 & ~n9393 ;
  assign n9395 = n3829 & ~n9394 ;
  assign n9399 = n2717 & n8012 ;
  assign n9400 = ~n9392 & ~n9399 ;
  assign n9401 = n3969 & ~n9400 ;
  assign n9396 = n2717 & n8006 ;
  assign n9397 = ~n9392 & ~n9396 ;
  assign n9398 = n4025 & ~n9397 ;
  assign n9389 = n3211 & n4028 ;
  assign n9390 = ~n8018 & ~n9389 ;
  assign n9391 = n2717 & ~n9390 ;
  assign n9402 = n3214 & n4073 ;
  assign n9403 = \P1_reg2_reg[11]/NET0131  & ~n4071 ;
  assign n9404 = ~n9402 & ~n9403 ;
  assign n9405 = ~n9391 & n9404 ;
  assign n9406 = ~n9398 & n9405 ;
  assign n9407 = ~n9401 & n9406 ;
  assign n9408 = ~n9395 & n9407 ;
  assign n9409 = n2701 & ~n9408 ;
  assign n9410 = ~n9388 & ~n9409 ;
  assign n9411 = \P1_state_reg[0]/NET0131  & ~n9410 ;
  assign n9412 = ~n9387 & ~n9411 ;
  assign n9414 = \P1_reg2_reg[15]/NET0131  & ~n2717 ;
  assign n9415 = n2717 & n8042 ;
  assign n9416 = ~n9414 & ~n9415 ;
  assign n9417 = n3829 & ~n9416 ;
  assign n9418 = n2717 & ~n8048 ;
  assign n9419 = ~n9414 & ~n9418 ;
  assign n9420 = n3969 & ~n9419 ;
  assign n9421 = n2717 & n8056 ;
  assign n9422 = ~n9414 & ~n9421 ;
  assign n9423 = n4025 & ~n9422 ;
  assign n9413 = n2717 & n8037 ;
  assign n9424 = n3735 & n4073 ;
  assign n9425 = \P1_reg2_reg[15]/NET0131  & ~n4071 ;
  assign n9426 = ~n9424 & ~n9425 ;
  assign n9427 = ~n9413 & n9426 ;
  assign n9428 = ~n9423 & n9427 ;
  assign n9429 = ~n9420 & n9428 ;
  assign n9430 = ~n9417 & n9429 ;
  assign n9431 = n2701 & ~n9430 ;
  assign n9432 = \P1_reg2_reg[15]/NET0131  & n4081 ;
  assign n9433 = ~n9431 & ~n9432 ;
  assign n9434 = \P1_state_reg[0]/NET0131  & ~n9433 ;
  assign n9435 = \P1_reg2_reg[15]/NET0131  & ~n4085 ;
  assign n9436 = ~n9434 & ~n9435 ;
  assign n9437 = \P1_reg2_reg[14]/NET0131  & ~n4085 ;
  assign n9438 = \P1_reg2_reg[14]/NET0131  & n4081 ;
  assign n9440 = \P1_reg2_reg[14]/NET0131  & ~n2717 ;
  assign n9441 = n2717 & n8087 ;
  assign n9442 = ~n9440 & ~n9441 ;
  assign n9443 = n4025 & ~n9442 ;
  assign n9447 = n2717 & n8093 ;
  assign n9448 = ~n9440 & ~n9447 ;
  assign n9449 = n3829 & ~n9448 ;
  assign n9444 = n2717 & ~n8099 ;
  assign n9445 = ~n9440 & ~n9444 ;
  assign n9446 = n3969 & ~n9445 ;
  assign n9439 = n2717 & ~n8080 ;
  assign n9450 = n3659 & n4073 ;
  assign n9451 = \P1_reg2_reg[14]/NET0131  & ~n4071 ;
  assign n9452 = ~n9450 & ~n9451 ;
  assign n9453 = ~n9439 & n9452 ;
  assign n9454 = ~n9446 & n9453 ;
  assign n9455 = ~n9449 & n9454 ;
  assign n9456 = ~n9443 & n9455 ;
  assign n9457 = n2701 & ~n9456 ;
  assign n9458 = ~n9438 & ~n9457 ;
  assign n9459 = \P1_state_reg[0]/NET0131  & ~n9458 ;
  assign n9460 = ~n9437 & ~n9459 ;
  assign n9461 = \P2_reg1_reg[11]/NET0131  & ~n2286 ;
  assign n9462 = \P2_reg1_reg[11]/NET0131  & n2035 ;
  assign n9464 = \P2_reg1_reg[11]/NET0131  & ~n2310 ;
  assign n9465 = n2310 & n8128 ;
  assign n9466 = ~n9464 & ~n9465 ;
  assign n9467 = ~n2392 & ~n9466 ;
  assign n9463 = ~n882 & n4101 ;
  assign n9478 = \P2_reg1_reg[11]/NET0131  & ~n4099 ;
  assign n9479 = ~n9463 & ~n9478 ;
  assign n9480 = ~n9467 & n9479 ;
  assign n9468 = \P2_reg1_reg[11]/NET0131  & ~n2291 ;
  assign n9475 = n2291 & ~n8140 ;
  assign n9476 = ~n9468 & ~n9475 ;
  assign n9477 = n1790 & ~n9476 ;
  assign n9469 = n2291 & ~n8122 ;
  assign n9470 = ~n9468 & ~n9469 ;
  assign n9471 = n2314 & ~n9470 ;
  assign n9472 = n2310 & ~n8122 ;
  assign n9473 = ~n9464 & ~n9472 ;
  assign n9474 = ~n2290 & ~n9473 ;
  assign n9481 = ~n9471 & ~n9474 ;
  assign n9482 = ~n9477 & n9481 ;
  assign n9483 = n9480 & n9482 ;
  assign n9484 = n2037 & ~n9483 ;
  assign n9485 = ~n9462 & ~n9484 ;
  assign n9486 = \P1_state_reg[0]/NET0131  & ~n9485 ;
  assign n9487 = ~n9461 & ~n9486 ;
  assign n9488 = \P2_reg1_reg[14]/NET0131  & ~n2286 ;
  assign n9489 = \P2_reg1_reg[14]/NET0131  & n2035 ;
  assign n9493 = \P2_reg1_reg[14]/NET0131  & ~n2291 ;
  assign n9494 = n2291 & n8173 ;
  assign n9495 = ~n9493 & ~n9494 ;
  assign n9496 = n2314 & ~n9495 ;
  assign n9504 = n2291 & ~n8182 ;
  assign n9505 = ~n9493 & ~n9504 ;
  assign n9506 = n1790 & ~n9505 ;
  assign n9490 = ~n760 & n2272 ;
  assign n9491 = n2310 & n9490 ;
  assign n9492 = \P2_reg1_reg[14]/NET0131  & ~n4099 ;
  assign n9507 = ~n9491 & ~n9492 ;
  assign n9508 = ~n9506 & n9507 ;
  assign n9509 = ~n9496 & n9508 ;
  assign n9497 = \P2_reg1_reg[14]/NET0131  & ~n2310 ;
  assign n9498 = n2310 & n8173 ;
  assign n9499 = ~n9497 & ~n9498 ;
  assign n9500 = ~n2290 & ~n9499 ;
  assign n9501 = n2310 & ~n8163 ;
  assign n9502 = ~n9497 & ~n9501 ;
  assign n9503 = ~n2392 & ~n9502 ;
  assign n9510 = ~n9500 & ~n9503 ;
  assign n9511 = n9509 & n9510 ;
  assign n9512 = n2037 & ~n9511 ;
  assign n9513 = ~n9489 & ~n9512 ;
  assign n9514 = \P1_state_reg[0]/NET0131  & ~n9513 ;
  assign n9515 = ~n9488 & ~n9514 ;
  assign n9516 = \P2_reg1_reg[15]/NET0131  & ~n2286 ;
  assign n9517 = \P2_reg1_reg[15]/NET0131  & n2035 ;
  assign n9520 = \P2_reg1_reg[15]/NET0131  & ~n2291 ;
  assign n9524 = n2291 & ~n8222 ;
  assign n9525 = ~n9520 & ~n9524 ;
  assign n9526 = n2314 & ~n9525 ;
  assign n9521 = n2291 & ~n8206 ;
  assign n9522 = ~n9520 & ~n9521 ;
  assign n9523 = n1790 & ~n9522 ;
  assign n9518 = n2310 & n9351 ;
  assign n9519 = \P2_reg1_reg[15]/NET0131  & ~n4099 ;
  assign n9534 = ~n9518 & ~n9519 ;
  assign n9535 = ~n9523 & n9534 ;
  assign n9536 = ~n9526 & n9535 ;
  assign n9527 = \P2_reg1_reg[15]/NET0131  & ~n2310 ;
  assign n9528 = n2310 & n8212 ;
  assign n9529 = ~n9527 & ~n9528 ;
  assign n9530 = ~n2392 & ~n9529 ;
  assign n9531 = n2310 & ~n8222 ;
  assign n9532 = ~n9527 & ~n9531 ;
  assign n9533 = ~n2290 & ~n9532 ;
  assign n9537 = ~n9530 & ~n9533 ;
  assign n9538 = n9536 & n9537 ;
  assign n9539 = n2037 & ~n9538 ;
  assign n9540 = ~n9517 & ~n9539 ;
  assign n9541 = \P1_state_reg[0]/NET0131  & ~n9540 ;
  assign n9542 = ~n9516 & ~n9541 ;
  assign n9543 = \P2_reg2_reg[11]/NET0131  & ~n2286 ;
  assign n9544 = \P2_reg2_reg[11]/NET0131  & n2035 ;
  assign n9546 = \P2_reg2_reg[11]/NET0131  & ~n2291 ;
  assign n9547 = n2291 & n8128 ;
  assign n9548 = ~n9546 & ~n9547 ;
  assign n9549 = ~n2392 & ~n9548 ;
  assign n9545 = \P2_reg2_reg[11]/NET0131  & ~n2407 ;
  assign n9558 = ~n861 & n1854 ;
  assign n9559 = ~n882 & n2394 ;
  assign n9560 = ~n9558 & ~n9559 ;
  assign n9561 = ~n9545 & n9560 ;
  assign n9562 = ~n9549 & n9561 ;
  assign n9550 = \P2_reg2_reg[11]/NET0131  & ~n2310 ;
  assign n9555 = n2310 & ~n8140 ;
  assign n9556 = ~n9550 & ~n9555 ;
  assign n9557 = n1790 & ~n9556 ;
  assign n9551 = ~n9472 & ~n9550 ;
  assign n9552 = n2314 & ~n9551 ;
  assign n9553 = ~n9469 & ~n9546 ;
  assign n9554 = ~n2290 & ~n9553 ;
  assign n9563 = ~n9552 & ~n9554 ;
  assign n9564 = ~n9557 & n9563 ;
  assign n9565 = n9562 & n9564 ;
  assign n9566 = n2037 & ~n9565 ;
  assign n9567 = ~n9544 & ~n9566 ;
  assign n9568 = \P1_state_reg[0]/NET0131  & ~n9567 ;
  assign n9569 = ~n9543 & ~n9568 ;
  assign n9570 = \P2_reg2_reg[14]/NET0131  & ~n2286 ;
  assign n9571 = \P2_reg2_reg[14]/NET0131  & n2035 ;
  assign n9573 = \P2_reg2_reg[14]/NET0131  & ~n2310 ;
  assign n9574 = ~n9498 & ~n9573 ;
  assign n9575 = n2314 & ~n9574 ;
  assign n9582 = n2310 & ~n8182 ;
  assign n9583 = ~n9573 & ~n9582 ;
  assign n9584 = n1790 & ~n9583 ;
  assign n9572 = n2291 & n9490 ;
  assign n9585 = ~n767 & n1854 ;
  assign n9586 = \P2_reg2_reg[14]/NET0131  & ~n2407 ;
  assign n9587 = ~n9585 & ~n9586 ;
  assign n9588 = ~n9572 & n9587 ;
  assign n9589 = ~n9584 & n9588 ;
  assign n9590 = ~n9575 & n9589 ;
  assign n9576 = \P2_reg2_reg[14]/NET0131  & ~n2291 ;
  assign n9577 = ~n9494 & ~n9576 ;
  assign n9578 = ~n2290 & ~n9577 ;
  assign n9579 = n2291 & ~n8163 ;
  assign n9580 = ~n9576 & ~n9579 ;
  assign n9581 = ~n2392 & ~n9580 ;
  assign n9591 = ~n9578 & ~n9581 ;
  assign n9592 = n9590 & n9591 ;
  assign n9593 = n2037 & ~n9592 ;
  assign n9594 = ~n9571 & ~n9593 ;
  assign n9595 = \P1_state_reg[0]/NET0131  & ~n9594 ;
  assign n9596 = ~n9570 & ~n9595 ;
  assign n9597 = \P2_reg2_reg[15]/NET0131  & ~n2286 ;
  assign n9598 = \P2_reg2_reg[15]/NET0131  & n2035 ;
  assign n9600 = \P2_reg2_reg[15]/NET0131  & ~n2310 ;
  assign n9604 = ~n9531 & ~n9600 ;
  assign n9605 = n2314 & ~n9604 ;
  assign n9601 = n2310 & ~n8206 ;
  assign n9602 = ~n9600 & ~n9601 ;
  assign n9603 = n1790 & ~n9602 ;
  assign n9599 = n2291 & n9351 ;
  assign n9612 = ~n595 & n1854 ;
  assign n9613 = \P2_reg2_reg[15]/NET0131  & ~n2407 ;
  assign n9614 = ~n9612 & ~n9613 ;
  assign n9615 = ~n9599 & n9614 ;
  assign n9616 = ~n9603 & n9615 ;
  assign n9617 = ~n9605 & n9616 ;
  assign n9606 = \P2_reg2_reg[15]/NET0131  & ~n2291 ;
  assign n9607 = n2291 & n8212 ;
  assign n9608 = ~n9606 & ~n9607 ;
  assign n9609 = ~n2392 & ~n9608 ;
  assign n9610 = ~n9524 & ~n9606 ;
  assign n9611 = ~n2290 & ~n9610 ;
  assign n9618 = ~n9609 & ~n9611 ;
  assign n9619 = n9617 & n9618 ;
  assign n9620 = n2037 & ~n9619 ;
  assign n9621 = ~n9598 & ~n9620 ;
  assign n9622 = \P1_state_reg[0]/NET0131  & ~n9621 ;
  assign n9623 = ~n9597 & ~n9622 ;
  assign n9624 = \P1_reg0_reg[15]/NET0131  & ~n4085 ;
  assign n9626 = \P1_reg0_reg[15]/NET0131  & ~n4869 ;
  assign n9627 = n4869 & n8042 ;
  assign n9628 = ~n9626 & ~n9627 ;
  assign n9629 = n3829 & ~n9628 ;
  assign n9630 = n4869 & ~n8048 ;
  assign n9631 = ~n9626 & ~n9630 ;
  assign n9632 = n3969 & ~n9631 ;
  assign n9633 = n4869 & n8056 ;
  assign n9634 = ~n9626 & ~n9633 ;
  assign n9635 = n4025 & ~n9634 ;
  assign n9625 = n4869 & n8037 ;
  assign n9636 = \P1_reg0_reg[15]/NET0131  & ~n5844 ;
  assign n9637 = ~n9625 & ~n9636 ;
  assign n9638 = ~n9635 & n9637 ;
  assign n9639 = ~n9632 & n9638 ;
  assign n9640 = ~n9629 & n9639 ;
  assign n9641 = n2701 & ~n9640 ;
  assign n9642 = \P1_reg0_reg[15]/NET0131  & n4081 ;
  assign n9643 = ~n9641 & ~n9642 ;
  assign n9644 = \P1_state_reg[0]/NET0131  & ~n9643 ;
  assign n9645 = ~n9624 & ~n9644 ;
  assign n9646 = n9333 & ~n9340 ;
  assign n9647 = n4869 & ~n9646 ;
  assign n9648 = n9331 & n9647 ;
  assign n9649 = ~\P1_reg0_reg[8]/NET0131  & ~n9648 ;
  assign n9650 = ~n7303 & n9333 ;
  assign n9651 = \P1_reg0_reg[8]/NET0131  & ~n9650 ;
  assign n9652 = n5844 & ~n9647 ;
  assign n9653 = ~n9651 & n9652 ;
  assign n9654 = ~n9649 & ~n9653 ;
  assign n9656 = \P1_reg1_reg[15]/NET0131  & ~n4202 ;
  assign n9657 = n4202 & n8042 ;
  assign n9658 = ~n9656 & ~n9657 ;
  assign n9659 = n3829 & ~n9658 ;
  assign n9660 = n4202 & ~n8048 ;
  assign n9661 = ~n9656 & ~n9660 ;
  assign n9662 = n3969 & ~n9661 ;
  assign n9663 = n4202 & n8056 ;
  assign n9664 = ~n9656 & ~n9663 ;
  assign n9665 = n4025 & ~n9664 ;
  assign n9655 = \P1_reg1_reg[15]/NET0131  & ~n6494 ;
  assign n9666 = n4202 & n8037 ;
  assign n9667 = ~n9655 & ~n9666 ;
  assign n9668 = ~n9665 & n9667 ;
  assign n9669 = ~n9662 & n9668 ;
  assign n9670 = ~n9659 & n9669 ;
  assign n9671 = n2701 & ~n9670 ;
  assign n9672 = \P1_reg1_reg[15]/NET0131  & n4081 ;
  assign n9673 = ~n9671 & ~n9672 ;
  assign n9674 = \P1_state_reg[0]/NET0131  & ~n9673 ;
  assign n9675 = \P1_reg1_reg[15]/NET0131  & ~n4085 ;
  assign n9676 = ~n9674 & ~n9675 ;
  assign n9677 = \P2_reg0_reg[11]/NET0131  & ~n2286 ;
  assign n9678 = \P2_reg0_reg[11]/NET0131  & n2035 ;
  assign n9680 = \P2_reg0_reg[11]/NET0131  & ~n2124 ;
  assign n9681 = n2124 & ~n8122 ;
  assign n9682 = ~n9680 & ~n9681 ;
  assign n9683 = ~n2120 & ~n9682 ;
  assign n9679 = ~n882 & n2616 ;
  assign n9692 = \P2_reg0_reg[11]/NET0131  & ~n2614 ;
  assign n9693 = ~n9679 & ~n9692 ;
  assign n9694 = ~n9683 & n9693 ;
  assign n9686 = \P2_reg0_reg[11]/NET0131  & ~n2053 ;
  assign n9689 = n2053 & ~n8140 ;
  assign n9690 = ~n9686 & ~n9689 ;
  assign n9691 = n1790 & ~n9690 ;
  assign n9684 = ~n8133 & ~n9680 ;
  assign n9685 = ~n2224 & ~n9684 ;
  assign n9687 = ~n8129 & ~n9686 ;
  assign n9688 = n2123 & ~n9687 ;
  assign n9695 = ~n9685 & ~n9688 ;
  assign n9696 = ~n9691 & n9695 ;
  assign n9697 = n9694 & n9696 ;
  assign n9698 = n2037 & ~n9697 ;
  assign n9699 = ~n9678 & ~n9698 ;
  assign n9700 = \P1_state_reg[0]/NET0131  & ~n9699 ;
  assign n9701 = ~n9677 & ~n9700 ;
  assign n9702 = \P2_reg0_reg[14]/NET0131  & ~n2286 ;
  assign n9703 = \P2_reg0_reg[14]/NET0131  & n2035 ;
  assign n9706 = \P2_reg0_reg[14]/NET0131  & ~n2053 ;
  assign n9707 = ~n8168 & ~n9706 ;
  assign n9708 = n2123 & ~n9707 ;
  assign n9715 = n2053 & ~n8182 ;
  assign n9716 = ~n9706 & ~n9715 ;
  assign n9717 = n1790 & ~n9716 ;
  assign n9704 = n2124 & n9490 ;
  assign n9705 = \P2_reg0_reg[14]/NET0131  & ~n2614 ;
  assign n9718 = ~n9704 & ~n9705 ;
  assign n9719 = ~n9717 & n9718 ;
  assign n9720 = ~n9708 & n9719 ;
  assign n9709 = \P2_reg0_reg[14]/NET0131  & ~n2124 ;
  assign n9710 = ~n8164 & ~n9709 ;
  assign n9711 = ~n2224 & ~n9710 ;
  assign n9712 = n2124 & n8173 ;
  assign n9713 = ~n9709 & ~n9712 ;
  assign n9714 = ~n2120 & ~n9713 ;
  assign n9721 = ~n9711 & ~n9714 ;
  assign n9722 = n9720 & n9721 ;
  assign n9723 = n2037 & ~n9722 ;
  assign n9724 = ~n9703 & ~n9723 ;
  assign n9725 = \P1_state_reg[0]/NET0131  & ~n9724 ;
  assign n9726 = ~n9702 & ~n9725 ;
  assign n9729 = ~\P1_reg3_reg[3]/NET0131  & ~n4449 ;
  assign n9730 = n3318 & ~n3988 ;
  assign n9731 = ~n3989 & ~n9730 ;
  assign n9732 = ~n2731 & ~n9731 ;
  assign n9733 = n2731 & n3340 ;
  assign n9734 = ~n9732 & ~n9733 ;
  assign n9735 = n4449 & n9734 ;
  assign n9736 = ~n9729 & ~n9735 ;
  assign n9737 = n4025 & ~n9736 ;
  assign n9738 = ~n3355 & ~n3415 ;
  assign n9739 = ~n5426 & n9738 ;
  assign n9740 = n5426 & ~n9738 ;
  assign n9741 = ~n9739 & ~n9740 ;
  assign n9742 = n4449 & ~n9741 ;
  assign n9743 = ~n9729 & ~n9742 ;
  assign n9744 = n3829 & ~n9743 ;
  assign n9745 = ~n3854 & ~n3855 ;
  assign n9746 = n5426 & ~n9745 ;
  assign n9747 = ~n5426 & n9745 ;
  assign n9748 = ~n9746 & ~n9747 ;
  assign n9749 = n4449 & n9748 ;
  assign n9750 = ~n9729 & ~n9749 ;
  assign n9751 = n3969 & ~n9750 ;
  assign n9753 = ~n3371 & ~n4031 ;
  assign n9754 = ~n4032 & n4062 ;
  assign n9755 = ~n9753 & n9754 ;
  assign n9756 = n4449 & n9755 ;
  assign n9728 = ~\P1_reg3_reg[3]/NET0131  & ~n4542 ;
  assign n9752 = ~n3371 & ~n4522 ;
  assign n9757 = ~n9728 & ~n9752 ;
  assign n9758 = ~n9756 & n9757 ;
  assign n9759 = ~n9751 & n9758 ;
  assign n9760 = ~n9744 & n9759 ;
  assign n9761 = ~n9737 & n9760 ;
  assign n9762 = n2701 & ~n9761 ;
  assign n9763 = ~\P1_reg3_reg[3]/NET0131  & n4081 ;
  assign n9764 = ~n9762 & ~n9763 ;
  assign n9765 = \P1_state_reg[0]/NET0131  & ~n9764 ;
  assign n9727 = \P1_reg3_reg[3]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9766 = ~\P1_reg3_reg[3]/NET0131  & n4552 ;
  assign n9767 = ~n9727 & ~n9766 ;
  assign n9768 = ~n9765 & n9767 ;
  assign n9771 = n3490 & n4081 ;
  assign n9773 = n3490 & ~n4449 ;
  assign n9786 = n3470 & ~n8253 ;
  assign n9787 = ~n8254 & ~n9786 ;
  assign n9788 = ~n2731 & ~n9787 ;
  assign n9789 = n2731 & n3520 ;
  assign n9790 = ~n9788 & ~n9789 ;
  assign n9791 = n4449 & n9790 ;
  assign n9792 = ~n9773 & ~n9791 ;
  assign n9793 = n4025 & ~n9792 ;
  assign n9780 = n4650 & ~n5431 ;
  assign n9781 = ~n4650 & n5431 ;
  assign n9782 = ~n9780 & ~n9781 ;
  assign n9783 = n4449 & n9782 ;
  assign n9784 = ~n9773 & ~n9783 ;
  assign n9785 = n3829 & ~n9784 ;
  assign n9774 = n4961 & ~n5431 ;
  assign n9775 = ~n4961 & n5431 ;
  assign n9776 = ~n9774 & ~n9775 ;
  assign n9777 = n4449 & ~n9776 ;
  assign n9778 = ~n9773 & ~n9777 ;
  assign n9779 = n3969 & ~n9778 ;
  assign n9794 = ~n3485 & ~n9133 ;
  assign n9795 = ~n4035 & ~n9794 ;
  assign n9796 = n4449 & n9795 ;
  assign n9797 = ~n9773 & ~n9796 ;
  assign n9798 = n4062 & ~n9797 ;
  assign n9772 = ~n3485 & ~n4522 ;
  assign n9799 = n3490 & ~n4540 ;
  assign n9800 = ~n9772 & ~n9799 ;
  assign n9801 = ~n9798 & n9800 ;
  assign n9802 = ~n9779 & n9801 ;
  assign n9803 = ~n9785 & n9802 ;
  assign n9804 = ~n9793 & n9803 ;
  assign n9805 = n2701 & ~n9804 ;
  assign n9806 = ~n9771 & ~n9805 ;
  assign n9807 = \P1_state_reg[0]/NET0131  & ~n9806 ;
  assign n9769 = \P1_reg3_reg[6]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9770 = n3490 & n4552 ;
  assign n9808 = ~n9769 & ~n9770 ;
  assign n9809 = ~n9807 & n9808 ;
  assign n9814 = n3463 & ~n4449 ;
  assign n9815 = n3444 & ~n8254 ;
  assign n9816 = ~n8255 & ~n9815 ;
  assign n9817 = ~n2731 & ~n9816 ;
  assign n9818 = n2731 & n3494 ;
  assign n9819 = ~n9817 & ~n9818 ;
  assign n9820 = n4449 & n9819 ;
  assign n9821 = ~n9814 & ~n9820 ;
  assign n9822 = n4025 & ~n9821 ;
  assign n9823 = ~n4461 & n5428 ;
  assign n9824 = n4461 & ~n5428 ;
  assign n9825 = ~n9823 & ~n9824 ;
  assign n9826 = n4449 & n9825 ;
  assign n9827 = ~n9814 & ~n9826 ;
  assign n9828 = n3829 & ~n9827 ;
  assign n9829 = ~n3870 & n5428 ;
  assign n9830 = n3870 & ~n5428 ;
  assign n9831 = ~n9829 & ~n9830 ;
  assign n9832 = n4449 & ~n9831 ;
  assign n9833 = ~n9814 & ~n9832 ;
  assign n9834 = n3969 & ~n9833 ;
  assign n9811 = n3461 & ~n4035 ;
  assign n9812 = n9335 & ~n9811 ;
  assign n9813 = n4449 & n9812 ;
  assign n9835 = n3463 & ~n4542 ;
  assign n9836 = n3461 & ~n4522 ;
  assign n9837 = ~n9835 & ~n9836 ;
  assign n9838 = ~n9813 & n9837 ;
  assign n9839 = ~n9834 & n9838 ;
  assign n9840 = ~n9828 & n9839 ;
  assign n9841 = ~n9822 & n9840 ;
  assign n9842 = n2701 & ~n9841 ;
  assign n9843 = n3463 & n4081 ;
  assign n9844 = ~n9842 & ~n9843 ;
  assign n9845 = \P1_state_reg[0]/NET0131  & ~n9844 ;
  assign n9810 = \P1_reg3_reg[7]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9846 = n3463 & n4552 ;
  assign n9847 = ~n9810 & ~n9846 ;
  assign n9848 = ~n9845 & n9847 ;
  assign n9851 = ~n1055 & n2035 ;
  assign n9867 = ~n1055 & ~n2124 ;
  assign n9868 = n1037 & ~n9173 ;
  assign n9869 = n2263 & ~n9174 ;
  assign n9870 = ~n9868 & n9869 ;
  assign n9871 = ~n1086 & ~n2263 ;
  assign n9872 = ~n9870 & ~n9871 ;
  assign n9873 = n2124 & ~n9872 ;
  assign n9874 = ~n9867 & ~n9873 ;
  assign n9875 = n1790 & ~n9874 ;
  assign n9853 = ~n1055 & ~n2053 ;
  assign n9854 = n1807 & ~n1923 ;
  assign n9855 = ~n1807 & n1923 ;
  assign n9856 = ~n9854 & ~n9855 ;
  assign n9857 = n2053 & ~n9856 ;
  assign n9858 = ~n9853 & ~n9857 ;
  assign n9859 = ~n2120 & ~n9858 ;
  assign n9852 = ~n1076 & n2229 ;
  assign n9860 = ~n1055 & ~n2274 ;
  assign n9879 = ~n9852 & ~n9860 ;
  assign n9880 = ~n9859 & n9879 ;
  assign n9861 = n1923 & ~n2320 ;
  assign n9862 = ~n1923 & n2320 ;
  assign n9863 = ~n9861 & ~n9862 ;
  assign n9864 = n2053 & n9863 ;
  assign n9865 = ~n9853 & ~n9864 ;
  assign n9866 = ~n2224 & ~n9865 ;
  assign n9876 = n2124 & n9863 ;
  assign n9877 = ~n9867 & ~n9876 ;
  assign n9878 = n2123 & ~n9877 ;
  assign n9881 = ~n9866 & ~n9878 ;
  assign n9882 = n9880 & n9881 ;
  assign n9883 = ~n9875 & n9882 ;
  assign n9884 = n2037 & ~n9883 ;
  assign n9885 = ~n9851 & ~n9884 ;
  assign n9886 = \P1_state_reg[0]/NET0131  & ~n9885 ;
  assign n9849 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n9850 = ~n1055 & n2014 ;
  assign n9887 = ~n9849 & ~n9850 ;
  assign n9888 = ~n9886 & n9887 ;
  assign n9889 = \P1_reg2_reg[5]/NET0131  & ~n4085 ;
  assign n9893 = \P1_reg2_reg[5]/NET0131  & ~n2717 ;
  assign n9894 = n2717 & n9116 ;
  assign n9895 = ~n9893 & ~n9894 ;
  assign n9896 = n4025 & ~n9895 ;
  assign n9897 = n2717 & ~n9122 ;
  assign n9898 = ~n9893 & ~n9897 ;
  assign n9899 = n3829 & ~n9898 ;
  assign n9900 = n2717 & n9129 ;
  assign n9901 = ~n9893 & ~n9900 ;
  assign n9902 = n3969 & ~n9901 ;
  assign n9890 = ~n3511 & n4028 ;
  assign n9891 = ~n9136 & ~n9890 ;
  assign n9892 = n2717 & ~n9891 ;
  assign n9903 = n3516 & n4073 ;
  assign n9904 = \P1_reg2_reg[5]/NET0131  & ~n4071 ;
  assign n9905 = ~n9903 & ~n9904 ;
  assign n9906 = ~n9892 & n9905 ;
  assign n9907 = ~n9902 & n9906 ;
  assign n9908 = ~n9899 & n9907 ;
  assign n9909 = ~n9896 & n9908 ;
  assign n9910 = n2701 & ~n9909 ;
  assign n9911 = \P1_reg2_reg[5]/NET0131  & n4081 ;
  assign n9912 = ~n9910 & ~n9911 ;
  assign n9913 = \P1_state_reg[0]/NET0131  & ~n9912 ;
  assign n9914 = ~n9889 & ~n9913 ;
  assign n9916 = \P1_reg1_reg[5]/NET0131  & ~n4202 ;
  assign n9917 = n4202 & n9116 ;
  assign n9918 = ~n9916 & ~n9917 ;
  assign n9919 = n4025 & ~n9918 ;
  assign n9920 = n4202 & ~n9122 ;
  assign n9921 = ~n9916 & ~n9920 ;
  assign n9922 = n3829 & ~n9921 ;
  assign n9923 = n4202 & n9129 ;
  assign n9924 = ~n9916 & ~n9923 ;
  assign n9925 = n3969 & ~n9924 ;
  assign n9915 = \P1_reg1_reg[5]/NET0131  & ~n4218 ;
  assign n9926 = n4202 & ~n9891 ;
  assign n9927 = ~n9915 & ~n9926 ;
  assign n9928 = ~n9925 & n9927 ;
  assign n9929 = ~n9922 & n9928 ;
  assign n9930 = ~n9919 & n9929 ;
  assign n9931 = n2701 & ~n9930 ;
  assign n9932 = \P1_reg1_reg[5]/NET0131  & n4081 ;
  assign n9933 = ~n9931 & ~n9932 ;
  assign n9934 = \P1_state_reg[0]/NET0131  & ~n9933 ;
  assign n9935 = \P1_reg1_reg[5]/NET0131  & ~n4085 ;
  assign n9936 = ~n9934 & ~n9935 ;
  assign n9937 = \P2_reg0_reg[5]/NET0131  & ~n2286 ;
  assign n9938 = \P2_reg0_reg[5]/NET0131  & n2035 ;
  assign n9946 = \P2_reg0_reg[5]/NET0131  & ~n2053 ;
  assign n9949 = n2053 & ~n9178 ;
  assign n9950 = ~n9946 & ~n9949 ;
  assign n9951 = n1790 & ~n9950 ;
  assign n9941 = \P2_reg0_reg[5]/NET0131  & ~n2124 ;
  assign n9942 = n2124 & n9159 ;
  assign n9943 = ~n9941 & ~n9942 ;
  assign n9944 = ~n2120 & ~n9943 ;
  assign n9952 = ~n9168 & ~n9941 ;
  assign n9953 = ~n2224 & ~n9952 ;
  assign n9947 = ~n9182 & ~n9946 ;
  assign n9948 = n2123 & ~n9947 ;
  assign n9939 = ~n1050 & n2272 ;
  assign n9940 = n2124 & n9939 ;
  assign n9945 = \P2_reg0_reg[5]/NET0131  & ~n2614 ;
  assign n9954 = ~n9940 & ~n9945 ;
  assign n9955 = ~n9948 & n9954 ;
  assign n9956 = ~n9953 & n9955 ;
  assign n9957 = ~n9944 & n9956 ;
  assign n9958 = ~n9951 & n9957 ;
  assign n9959 = n2037 & ~n9958 ;
  assign n9960 = ~n9938 & ~n9959 ;
  assign n9961 = \P1_state_reg[0]/NET0131  & ~n9960 ;
  assign n9962 = ~n9937 & ~n9961 ;
  assign n9963 = \P2_reg0_reg[6]/NET0131  & ~n2286 ;
  assign n9964 = \P2_reg0_reg[6]/NET0131  & n2035 ;
  assign n9968 = \P2_reg0_reg[6]/NET0131  & ~n2124 ;
  assign n9969 = n2124 & ~n9222 ;
  assign n9970 = ~n9968 & ~n9969 ;
  assign n9971 = ~n2120 & ~n9970 ;
  assign n9965 = ~n1003 & n2272 ;
  assign n9966 = n2124 & n9965 ;
  assign n9967 = \P2_reg0_reg[6]/NET0131  & ~n2614 ;
  assign n9980 = ~n9966 & ~n9967 ;
  assign n9981 = ~n9971 & n9980 ;
  assign n9978 = ~n9208 & ~n9968 ;
  assign n9979 = ~n2224 & ~n9978 ;
  assign n9972 = \P2_reg0_reg[6]/NET0131  & ~n2053 ;
  assign n9973 = ~n9204 & ~n9972 ;
  assign n9974 = n2123 & ~n9973 ;
  assign n9975 = n2053 & ~n9216 ;
  assign n9976 = ~n9972 & ~n9975 ;
  assign n9977 = n1790 & ~n9976 ;
  assign n9982 = ~n9974 & ~n9977 ;
  assign n9983 = ~n9979 & n9982 ;
  assign n9984 = n9981 & n9983 ;
  assign n9985 = n2037 & ~n9984 ;
  assign n9986 = ~n9964 & ~n9985 ;
  assign n9987 = \P1_state_reg[0]/NET0131  & ~n9986 ;
  assign n9988 = ~n9963 & ~n9987 ;
  assign n9989 = \P2_reg0_reg[7]/NET0131  & ~n2286 ;
  assign n9990 = \P2_reg0_reg[7]/NET0131  & n2035 ;
  assign n9993 = \P2_reg0_reg[7]/NET0131  & ~n2124 ;
  assign n9994 = n2124 & n9253 ;
  assign n9995 = ~n9993 & ~n9994 ;
  assign n9996 = ~n2120 & ~n9995 ;
  assign n9997 = \P2_reg0_reg[7]/NET0131  & ~n2053 ;
  assign n10002 = n2053 & ~n9261 ;
  assign n10003 = ~n9997 & ~n10002 ;
  assign n10004 = n1790 & ~n10003 ;
  assign n9991 = ~n1026 & n2272 ;
  assign n9992 = n2124 & n9991 ;
  assign n10005 = \P2_reg0_reg[7]/NET0131  & ~n2614 ;
  assign n10006 = ~n9992 & ~n10005 ;
  assign n10007 = ~n10004 & n10006 ;
  assign n10008 = ~n9996 & n10007 ;
  assign n9998 = ~n9244 & ~n9997 ;
  assign n9999 = n2123 & ~n9998 ;
  assign n10000 = ~n9248 & ~n9993 ;
  assign n10001 = ~n2224 & ~n10000 ;
  assign n10009 = ~n9999 & ~n10001 ;
  assign n10010 = n10008 & n10009 ;
  assign n10011 = n2037 & ~n10010 ;
  assign n10012 = ~n9990 & ~n10011 ;
  assign n10013 = \P1_state_reg[0]/NET0131  & ~n10012 ;
  assign n10014 = ~n9989 & ~n10013 ;
  assign n10015 = \P2_reg0_reg[8]/NET0131  & ~n2286 ;
  assign n10016 = \P2_reg0_reg[8]/NET0131  & n2035 ;
  assign n10019 = \P2_reg0_reg[8]/NET0131  & ~n2053 ;
  assign n10020 = ~n8286 & ~n10019 ;
  assign n10021 = n2123 & ~n10020 ;
  assign n10028 = n2053 & ~n8299 ;
  assign n10029 = ~n10019 & ~n10028 ;
  assign n10030 = n1790 & ~n10029 ;
  assign n10017 = ~n958 & n2272 ;
  assign n10018 = n2124 & n10017 ;
  assign n10031 = \P2_reg0_reg[8]/NET0131  & ~n2614 ;
  assign n10032 = ~n10018 & ~n10031 ;
  assign n10033 = ~n10030 & n10032 ;
  assign n10034 = ~n10021 & n10033 ;
  assign n10022 = \P2_reg0_reg[8]/NET0131  & ~n2124 ;
  assign n10023 = ~n8282 & ~n10022 ;
  assign n10024 = ~n2224 & ~n10023 ;
  assign n10025 = n2124 & ~n8291 ;
  assign n10026 = ~n10022 & ~n10025 ;
  assign n10027 = ~n2120 & ~n10026 ;
  assign n10035 = ~n10024 & ~n10027 ;
  assign n10036 = n10034 & n10035 ;
  assign n10037 = n2037 & ~n10036 ;
  assign n10038 = ~n10016 & ~n10037 ;
  assign n10039 = \P1_state_reg[0]/NET0131  & ~n10038 ;
  assign n10040 = ~n10015 & ~n10039 ;
  assign n10041 = \P1_reg2_reg[4]/NET0131  & ~n4085 ;
  assign n10042 = \P1_reg2_reg[4]/NET0131  & n4081 ;
  assign n10044 = \P1_reg2_reg[4]/NET0131  & ~n2717 ;
  assign n10051 = n2717 & n9089 ;
  assign n10052 = ~n10044 & ~n10051 ;
  assign n10053 = n4025 & ~n10052 ;
  assign n10048 = n2717 & n9081 ;
  assign n10049 = ~n10044 & ~n10048 ;
  assign n10050 = n3969 & ~n10049 ;
  assign n10045 = n2717 & ~n9075 ;
  assign n10046 = ~n10044 & ~n10045 ;
  assign n10047 = n3829 & ~n10046 ;
  assign n10054 = n2717 & n9094 ;
  assign n10055 = ~n10044 & ~n10054 ;
  assign n10056 = n4062 & ~n10055 ;
  assign n10043 = \P1_reg2_reg[4]/NET0131  & ~n5148 ;
  assign n10057 = n3312 & n4073 ;
  assign n10058 = n2717 & n9278 ;
  assign n10059 = ~n10057 & ~n10058 ;
  assign n10060 = ~n10043 & n10059 ;
  assign n10061 = ~n10056 & n10060 ;
  assign n10062 = ~n10047 & n10061 ;
  assign n10063 = ~n10050 & n10062 ;
  assign n10064 = ~n10053 & n10063 ;
  assign n10065 = n2701 & ~n10064 ;
  assign n10066 = ~n10042 & ~n10065 ;
  assign n10067 = \P1_state_reg[0]/NET0131  & ~n10066 ;
  assign n10068 = ~n10041 & ~n10067 ;
  assign n10069 = \P2_reg1_reg[5]/NET0131  & ~n2286 ;
  assign n10070 = \P2_reg1_reg[5]/NET0131  & n2035 ;
  assign n10076 = \P2_reg1_reg[5]/NET0131  & ~n2291 ;
  assign n10080 = n2291 & ~n9178 ;
  assign n10081 = ~n10076 & ~n10080 ;
  assign n10082 = n1790 & ~n10081 ;
  assign n10077 = n2291 & n9159 ;
  assign n10078 = ~n10076 & ~n10077 ;
  assign n10079 = n2314 & ~n10078 ;
  assign n10072 = \P2_reg1_reg[5]/NET0131  & ~n2310 ;
  assign n10073 = n2310 & n9159 ;
  assign n10074 = ~n10072 & ~n10073 ;
  assign n10075 = ~n2290 & ~n10074 ;
  assign n10083 = n2310 & ~n9167 ;
  assign n10084 = ~n10072 & ~n10083 ;
  assign n10085 = ~n2392 & ~n10084 ;
  assign n10071 = n2310 & n9939 ;
  assign n10086 = \P2_reg1_reg[5]/NET0131  & ~n4099 ;
  assign n10087 = ~n10071 & ~n10086 ;
  assign n10088 = ~n10085 & n10087 ;
  assign n10089 = ~n10075 & n10088 ;
  assign n10090 = ~n10079 & n10089 ;
  assign n10091 = ~n10082 & n10090 ;
  assign n10092 = n2037 & ~n10091 ;
  assign n10093 = ~n10070 & ~n10092 ;
  assign n10094 = \P1_state_reg[0]/NET0131  & ~n10093 ;
  assign n10095 = ~n10069 & ~n10094 ;
  assign n10096 = \P2_reg1_reg[6]/NET0131  & ~n2286 ;
  assign n10097 = \P2_reg1_reg[6]/NET0131  & n2035 ;
  assign n10100 = \P2_reg1_reg[6]/NET0131  & ~n2310 ;
  assign n10101 = n2310 & n9203 ;
  assign n10102 = ~n10100 & ~n10101 ;
  assign n10103 = ~n2392 & ~n10102 ;
  assign n10098 = n2310 & n9965 ;
  assign n10099 = \P2_reg1_reg[6]/NET0131  & ~n4099 ;
  assign n10114 = ~n10098 & ~n10099 ;
  assign n10115 = ~n10103 & n10114 ;
  assign n10111 = n2310 & ~n9222 ;
  assign n10112 = ~n10100 & ~n10111 ;
  assign n10113 = ~n2290 & ~n10112 ;
  assign n10104 = \P2_reg1_reg[6]/NET0131  & ~n2291 ;
  assign n10105 = n2291 & ~n9222 ;
  assign n10106 = ~n10104 & ~n10105 ;
  assign n10107 = n2314 & ~n10106 ;
  assign n10108 = n2291 & ~n9216 ;
  assign n10109 = ~n10104 & ~n10108 ;
  assign n10110 = n1790 & ~n10109 ;
  assign n10116 = ~n10107 & ~n10110 ;
  assign n10117 = ~n10113 & n10116 ;
  assign n10118 = n10115 & n10117 ;
  assign n10119 = n2037 & ~n10118 ;
  assign n10120 = ~n10097 & ~n10119 ;
  assign n10121 = \P1_state_reg[0]/NET0131  & ~n10120 ;
  assign n10122 = ~n10096 & ~n10121 ;
  assign n10123 = \P2_reg1_reg[7]/NET0131  & ~n2286 ;
  assign n10124 = \P2_reg1_reg[7]/NET0131  & n2035 ;
  assign n10126 = \P2_reg1_reg[7]/NET0131  & ~n2310 ;
  assign n10127 = n2310 & ~n9243 ;
  assign n10128 = ~n10126 & ~n10127 ;
  assign n10129 = ~n2392 & ~n10128 ;
  assign n10130 = \P2_reg1_reg[7]/NET0131  & ~n2291 ;
  assign n10137 = n2291 & ~n9261 ;
  assign n10138 = ~n10130 & ~n10137 ;
  assign n10139 = n1790 & ~n10138 ;
  assign n10125 = n2310 & n9991 ;
  assign n10140 = \P2_reg1_reg[7]/NET0131  & ~n4099 ;
  assign n10141 = ~n10125 & ~n10140 ;
  assign n10142 = ~n10139 & n10141 ;
  assign n10143 = ~n10129 & n10142 ;
  assign n10131 = n2291 & n9253 ;
  assign n10132 = ~n10130 & ~n10131 ;
  assign n10133 = n2314 & ~n10132 ;
  assign n10134 = n2310 & n9253 ;
  assign n10135 = ~n10126 & ~n10134 ;
  assign n10136 = ~n2290 & ~n10135 ;
  assign n10144 = ~n10133 & ~n10136 ;
  assign n10145 = n10143 & n10144 ;
  assign n10146 = n2037 & ~n10145 ;
  assign n10147 = ~n10124 & ~n10146 ;
  assign n10148 = \P1_state_reg[0]/NET0131  & ~n10147 ;
  assign n10149 = ~n10123 & ~n10148 ;
  assign n10150 = \P2_reg1_reg[8]/NET0131  & ~n2286 ;
  assign n10151 = \P2_reg1_reg[8]/NET0131  & n2035 ;
  assign n10153 = \P2_reg1_reg[8]/NET0131  & ~n2310 ;
  assign n10154 = n2310 & n8281 ;
  assign n10155 = ~n10153 & ~n10154 ;
  assign n10156 = ~n2392 & ~n10155 ;
  assign n10160 = \P2_reg1_reg[8]/NET0131  & ~n2291 ;
  assign n10164 = n2291 & ~n8299 ;
  assign n10165 = ~n10160 & ~n10164 ;
  assign n10166 = n1790 & ~n10165 ;
  assign n10152 = n2310 & n10017 ;
  assign n10167 = \P2_reg1_reg[8]/NET0131  & ~n4099 ;
  assign n10168 = ~n10152 & ~n10167 ;
  assign n10169 = ~n10166 & n10168 ;
  assign n10170 = ~n10156 & n10169 ;
  assign n10157 = n2310 & ~n8291 ;
  assign n10158 = ~n10153 & ~n10157 ;
  assign n10159 = ~n2290 & ~n10158 ;
  assign n10161 = n2291 & ~n8291 ;
  assign n10162 = ~n10160 & ~n10161 ;
  assign n10163 = n2314 & ~n10162 ;
  assign n10171 = ~n10159 & ~n10163 ;
  assign n10172 = n10170 & n10171 ;
  assign n10173 = n2037 & ~n10172 ;
  assign n10174 = ~n10151 & ~n10173 ;
  assign n10175 = \P1_state_reg[0]/NET0131  & ~n10174 ;
  assign n10176 = ~n10150 & ~n10175 ;
  assign n10177 = \P1_reg0_reg[11]/NET0131  & ~n4085 ;
  assign n10178 = \P1_reg0_reg[11]/NET0131  & n4081 ;
  assign n10180 = \P1_reg0_reg[11]/NET0131  & ~n4869 ;
  assign n10181 = n4869 & ~n7998 ;
  assign n10182 = ~n10180 & ~n10181 ;
  assign n10183 = n3829 & ~n10182 ;
  assign n10187 = n4869 & n8012 ;
  assign n10188 = ~n10180 & ~n10187 ;
  assign n10189 = n3969 & ~n10188 ;
  assign n10184 = n4869 & n8006 ;
  assign n10185 = ~n10180 & ~n10184 ;
  assign n10186 = n4025 & ~n10185 ;
  assign n10179 = \P1_reg0_reg[11]/NET0131  & ~n5866 ;
  assign n10190 = n4869 & ~n9390 ;
  assign n10191 = ~n10179 & ~n10190 ;
  assign n10192 = ~n10186 & n10191 ;
  assign n10193 = ~n10189 & n10192 ;
  assign n10194 = ~n10183 & n10193 ;
  assign n10195 = n2701 & ~n10194 ;
  assign n10196 = ~n10178 & ~n10195 ;
  assign n10197 = \P1_state_reg[0]/NET0131  & ~n10196 ;
  assign n10198 = ~n10177 & ~n10197 ;
  assign n10199 = \P2_reg2_reg[5]/NET0131  & ~n2286 ;
  assign n10200 = \P2_reg2_reg[5]/NET0131  & n2035 ;
  assign n10205 = \P2_reg2_reg[5]/NET0131  & ~n2310 ;
  assign n10208 = n2310 & ~n9178 ;
  assign n10209 = ~n10205 & ~n10208 ;
  assign n10210 = n1790 & ~n10209 ;
  assign n10206 = ~n10073 & ~n10205 ;
  assign n10207 = n2314 & ~n10206 ;
  assign n10202 = \P2_reg2_reg[5]/NET0131  & ~n2291 ;
  assign n10203 = ~n10077 & ~n10202 ;
  assign n10204 = ~n2290 & ~n10203 ;
  assign n10211 = n2291 & ~n9167 ;
  assign n10212 = ~n10202 & ~n10211 ;
  assign n10213 = ~n2392 & ~n10212 ;
  assign n10214 = \P2_reg2_reg[5]/NET0131  & ~n2407 ;
  assign n10201 = n2291 & n9939 ;
  assign n10215 = ~n1030 & n1854 ;
  assign n10216 = ~n10201 & ~n10215 ;
  assign n10217 = ~n10214 & n10216 ;
  assign n10218 = ~n10213 & n10217 ;
  assign n10219 = ~n10204 & n10218 ;
  assign n10220 = ~n10207 & n10219 ;
  assign n10221 = ~n10210 & n10220 ;
  assign n10222 = n2037 & ~n10221 ;
  assign n10223 = ~n10200 & ~n10222 ;
  assign n10224 = \P1_state_reg[0]/NET0131  & ~n10223 ;
  assign n10225 = ~n10199 & ~n10224 ;
  assign n10226 = \P2_reg2_reg[6]/NET0131  & ~n2286 ;
  assign n10227 = \P2_reg2_reg[6]/NET0131  & n2035 ;
  assign n10229 = \P2_reg2_reg[6]/NET0131  & ~n2291 ;
  assign n10230 = ~n10105 & ~n10229 ;
  assign n10231 = ~n2290 & ~n10230 ;
  assign n10242 = \P2_reg2_reg[6]/NET0131  & ~n2407 ;
  assign n10228 = n2291 & n9965 ;
  assign n10241 = ~n981 & n1854 ;
  assign n10243 = ~n10228 & ~n10241 ;
  assign n10244 = ~n10242 & n10243 ;
  assign n10245 = ~n10231 & n10244 ;
  assign n10238 = n2291 & n9203 ;
  assign n10239 = ~n10229 & ~n10238 ;
  assign n10240 = ~n2392 & ~n10239 ;
  assign n10232 = \P2_reg2_reg[6]/NET0131  & ~n2310 ;
  assign n10233 = ~n10111 & ~n10232 ;
  assign n10234 = n2314 & ~n10233 ;
  assign n10235 = n2310 & ~n9216 ;
  assign n10236 = ~n10232 & ~n10235 ;
  assign n10237 = n1790 & ~n10236 ;
  assign n10246 = ~n10234 & ~n10237 ;
  assign n10247 = ~n10240 & n10246 ;
  assign n10248 = n10245 & n10247 ;
  assign n10249 = n2037 & ~n10248 ;
  assign n10250 = ~n10227 & ~n10249 ;
  assign n10251 = \P1_state_reg[0]/NET0131  & ~n10250 ;
  assign n10252 = ~n10226 & ~n10251 ;
  assign n10253 = \P2_reg2_reg[7]/NET0131  & ~n2286 ;
  assign n10254 = \P2_reg2_reg[7]/NET0131  & n2035 ;
  assign n10260 = \P2_reg2_reg[7]/NET0131  & ~n2291 ;
  assign n10261 = n2291 & ~n9243 ;
  assign n10262 = ~n10260 & ~n10261 ;
  assign n10263 = ~n2392 & ~n10262 ;
  assign n10256 = \P2_reg2_reg[7]/NET0131  & ~n2310 ;
  assign n10257 = n2310 & ~n9261 ;
  assign n10258 = ~n10256 & ~n10257 ;
  assign n10259 = n1790 & ~n10258 ;
  assign n10268 = \P2_reg2_reg[7]/NET0131  & ~n2407 ;
  assign n10255 = n2291 & n9991 ;
  assign n10269 = ~n1007 & n1854 ;
  assign n10270 = ~n10255 & ~n10269 ;
  assign n10271 = ~n10268 & n10270 ;
  assign n10272 = ~n10259 & n10271 ;
  assign n10273 = ~n10263 & n10272 ;
  assign n10264 = ~n10134 & ~n10256 ;
  assign n10265 = n2314 & ~n10264 ;
  assign n10266 = ~n10131 & ~n10260 ;
  assign n10267 = ~n2290 & ~n10266 ;
  assign n10274 = ~n10265 & ~n10267 ;
  assign n10275 = n10273 & n10274 ;
  assign n10276 = n2037 & ~n10275 ;
  assign n10277 = ~n10254 & ~n10276 ;
  assign n10278 = \P1_state_reg[0]/NET0131  & ~n10277 ;
  assign n10279 = ~n10253 & ~n10278 ;
  assign n10280 = \P2_reg2_reg[8]/NET0131  & ~n2286 ;
  assign n10281 = \P2_reg2_reg[8]/NET0131  & n2035 ;
  assign n10287 = \P2_reg2_reg[8]/NET0131  & ~n2291 ;
  assign n10288 = n2291 & n8281 ;
  assign n10289 = ~n10287 & ~n10288 ;
  assign n10290 = ~n2392 & ~n10289 ;
  assign n10283 = \P2_reg2_reg[8]/NET0131  & ~n2310 ;
  assign n10284 = n2310 & ~n8299 ;
  assign n10285 = ~n10283 & ~n10284 ;
  assign n10286 = n1790 & ~n10285 ;
  assign n10295 = \P2_reg2_reg[8]/NET0131  & ~n2407 ;
  assign n10282 = n2291 & n10017 ;
  assign n10296 = ~n939 & n1854 ;
  assign n10297 = ~n10282 & ~n10296 ;
  assign n10298 = ~n10295 & n10297 ;
  assign n10299 = ~n10286 & n10298 ;
  assign n10300 = ~n10290 & n10299 ;
  assign n10291 = ~n10157 & ~n10283 ;
  assign n10292 = n2314 & ~n10291 ;
  assign n10293 = ~n10161 & ~n10287 ;
  assign n10294 = ~n2290 & ~n10293 ;
  assign n10301 = ~n10292 & ~n10294 ;
  assign n10302 = n10300 & n10301 ;
  assign n10303 = n2037 & ~n10302 ;
  assign n10304 = ~n10281 & ~n10303 ;
  assign n10305 = \P1_state_reg[0]/NET0131  & ~n10304 ;
  assign n10306 = ~n10280 & ~n10305 ;
  assign n10307 = \P1_reg0_reg[14]/NET0131  & ~n4085 ;
  assign n10308 = \P1_reg0_reg[14]/NET0131  & n4081 ;
  assign n10310 = \P1_reg0_reg[14]/NET0131  & ~n4869 ;
  assign n10311 = n4869 & n8087 ;
  assign n10312 = ~n10310 & ~n10311 ;
  assign n10313 = n4025 & ~n10312 ;
  assign n10317 = n4869 & n8093 ;
  assign n10318 = ~n10310 & ~n10317 ;
  assign n10319 = n3829 & ~n10318 ;
  assign n10314 = n4869 & ~n8099 ;
  assign n10315 = ~n10310 & ~n10314 ;
  assign n10316 = n3969 & ~n10315 ;
  assign n10309 = n4869 & ~n8080 ;
  assign n10320 = \P1_reg0_reg[14]/NET0131  & ~n5844 ;
  assign n10321 = ~n10309 & ~n10320 ;
  assign n10322 = ~n10316 & n10321 ;
  assign n10323 = ~n10319 & n10322 ;
  assign n10324 = ~n10313 & n10323 ;
  assign n10325 = n2701 & ~n10324 ;
  assign n10326 = ~n10308 & ~n10325 ;
  assign n10327 = \P1_state_reg[0]/NET0131  & ~n10326 ;
  assign n10328 = ~n10307 & ~n10327 ;
  assign n10329 = \P1_reg0_reg[5]/NET0131  & ~n4085 ;
  assign n10331 = \P1_reg0_reg[5]/NET0131  & ~n4869 ;
  assign n10332 = n4869 & n9116 ;
  assign n10333 = ~n10331 & ~n10332 ;
  assign n10334 = n4025 & ~n10333 ;
  assign n10335 = n4869 & ~n9122 ;
  assign n10336 = ~n10331 & ~n10335 ;
  assign n10337 = n3829 & ~n10336 ;
  assign n10338 = n4869 & n9129 ;
  assign n10339 = ~n10331 & ~n10338 ;
  assign n10340 = n3969 & ~n10339 ;
  assign n10330 = n4869 & ~n9891 ;
  assign n10341 = \P1_reg0_reg[5]/NET0131  & ~n5844 ;
  assign n10342 = ~n10330 & ~n10341 ;
  assign n10343 = ~n10340 & n10342 ;
  assign n10344 = ~n10337 & n10343 ;
  assign n10345 = ~n10334 & n10344 ;
  assign n10346 = n2701 & ~n10345 ;
  assign n10347 = \P1_reg0_reg[5]/NET0131  & n4081 ;
  assign n10348 = ~n10346 & ~n10347 ;
  assign n10349 = \P1_state_reg[0]/NET0131  & ~n10348 ;
  assign n10350 = ~n10329 & ~n10349 ;
  assign n10351 = \P1_reg1_reg[11]/NET0131  & ~n4085 ;
  assign n10352 = \P1_reg1_reg[11]/NET0131  & n4081 ;
  assign n10354 = \P1_reg1_reg[11]/NET0131  & ~n4202 ;
  assign n10355 = n4202 & ~n7998 ;
  assign n10356 = ~n10354 & ~n10355 ;
  assign n10357 = n3829 & ~n10356 ;
  assign n10361 = n4202 & n8012 ;
  assign n10362 = ~n10354 & ~n10361 ;
  assign n10363 = n3969 & ~n10362 ;
  assign n10358 = n4202 & n8006 ;
  assign n10359 = ~n10354 & ~n10358 ;
  assign n10360 = n4025 & ~n10359 ;
  assign n10353 = n4202 & ~n9390 ;
  assign n10364 = \P1_reg1_reg[11]/NET0131  & ~n6494 ;
  assign n10365 = ~n10353 & ~n10364 ;
  assign n10366 = ~n10360 & n10365 ;
  assign n10367 = ~n10363 & n10366 ;
  assign n10368 = ~n10357 & n10367 ;
  assign n10369 = n2701 & ~n10368 ;
  assign n10370 = ~n10352 & ~n10369 ;
  assign n10371 = \P1_state_reg[0]/NET0131  & ~n10370 ;
  assign n10372 = ~n10351 & ~n10371 ;
  assign n10373 = \P1_reg1_reg[14]/NET0131  & ~n4085 ;
  assign n10374 = \P1_reg1_reg[14]/NET0131  & n4081 ;
  assign n10376 = \P1_reg1_reg[14]/NET0131  & ~n4202 ;
  assign n10377 = n4202 & n8087 ;
  assign n10378 = ~n10376 & ~n10377 ;
  assign n10379 = n4025 & ~n10378 ;
  assign n10383 = n4202 & ~n8099 ;
  assign n10384 = ~n10376 & ~n10383 ;
  assign n10385 = n3969 & ~n10384 ;
  assign n10380 = n4202 & n8093 ;
  assign n10381 = ~n10376 & ~n10380 ;
  assign n10382 = n3829 & ~n10381 ;
  assign n10375 = \P1_reg1_reg[14]/NET0131  & ~n6494 ;
  assign n10386 = n4202 & ~n8080 ;
  assign n10387 = ~n10375 & ~n10386 ;
  assign n10388 = ~n10382 & n10387 ;
  assign n10389 = ~n10385 & n10388 ;
  assign n10390 = ~n10379 & n10389 ;
  assign n10391 = n2701 & ~n10390 ;
  assign n10392 = ~n10374 & ~n10391 ;
  assign n10393 = \P1_state_reg[0]/NET0131  & ~n10392 ;
  assign n10394 = ~n10373 & ~n10393 ;
  assign n10397 = ~\P2_reg3_reg[3]/NET0131  & n2035 ;
  assign n10399 = ~\P2_reg3_reg[3]/NET0131  & ~n2124 ;
  assign n10415 = n1062 & ~n9172 ;
  assign n10416 = n2263 & ~n9173 ;
  assign n10417 = ~n10415 & n10416 ;
  assign n10418 = ~n1110 & ~n2263 ;
  assign n10419 = ~n10417 & ~n10418 ;
  assign n10420 = n2124 & ~n10419 ;
  assign n10421 = ~n10399 & ~n10420 ;
  assign n10422 = n1790 & ~n10421 ;
  assign n10407 = ~n1125 & ~n2059 ;
  assign n10408 = n1926 & ~n10407 ;
  assign n10409 = ~n1926 & n10407 ;
  assign n10410 = ~n10408 & ~n10409 ;
  assign n10411 = ~n2120 & n10410 ;
  assign n10400 = ~n2138 & ~n2139 ;
  assign n10401 = n1926 & ~n10400 ;
  assign n10402 = ~n1926 & n10400 ;
  assign n10403 = ~n10401 & ~n10402 ;
  assign n10412 = ~n2224 & ~n10403 ;
  assign n10413 = ~n10411 & ~n10412 ;
  assign n10414 = n2053 & ~n10413 ;
  assign n10404 = n2124 & ~n10403 ;
  assign n10405 = ~n10399 & ~n10404 ;
  assign n10406 = n2123 & ~n10405 ;
  assign n10398 = ~n1100 & n2229 ;
  assign n10423 = n2120 & n2224 ;
  assign n10424 = ~n2053 & ~n10423 ;
  assign n10425 = n2274 & ~n10424 ;
  assign n10426 = ~\P2_reg3_reg[3]/NET0131  & ~n10425 ;
  assign n10427 = ~n10398 & ~n10426 ;
  assign n10428 = ~n10406 & n10427 ;
  assign n10429 = ~n10414 & n10428 ;
  assign n10430 = ~n10422 & n10429 ;
  assign n10431 = n2037 & ~n10430 ;
  assign n10432 = ~n10397 & ~n10431 ;
  assign n10433 = \P1_state_reg[0]/NET0131  & ~n10432 ;
  assign n10395 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[3]/NET0131  ;
  assign n10396 = ~\P2_reg3_reg[3]/NET0131  & n2014 ;
  assign n10434 = ~n10395 & ~n10396 ;
  assign n10435 = ~n10433 & n10434 ;
  assign n10437 = \P1_reg1_reg[3]/NET0131  & ~n4202 ;
  assign n10438 = n4202 & n9734 ;
  assign n10439 = ~n10437 & ~n10438 ;
  assign n10440 = n4025 & ~n10439 ;
  assign n10441 = n4202 & ~n9741 ;
  assign n10442 = ~n10437 & ~n10441 ;
  assign n10443 = n3829 & ~n10442 ;
  assign n10444 = n4202 & n9748 ;
  assign n10445 = ~n10437 & ~n10444 ;
  assign n10446 = n3969 & ~n10445 ;
  assign n10436 = \P1_reg1_reg[3]/NET0131  & ~n4218 ;
  assign n10447 = ~n3371 & n4028 ;
  assign n10448 = ~n9755 & ~n10447 ;
  assign n10449 = n4202 & ~n10448 ;
  assign n10450 = ~n10436 & ~n10449 ;
  assign n10451 = ~n10446 & n10450 ;
  assign n10452 = ~n10443 & n10451 ;
  assign n10453 = ~n10440 & n10452 ;
  assign n10454 = n2701 & ~n10453 ;
  assign n10455 = \P1_reg1_reg[3]/NET0131  & n4081 ;
  assign n10456 = ~n10454 & ~n10455 ;
  assign n10457 = \P1_state_reg[0]/NET0131  & ~n10456 ;
  assign n10458 = \P1_reg1_reg[3]/NET0131  & ~n4085 ;
  assign n10459 = ~n10457 & ~n10458 ;
  assign n10461 = \P1_reg1_reg[7]/NET0131  & ~n4202 ;
  assign n10462 = n4202 & n9819 ;
  assign n10463 = ~n10461 & ~n10462 ;
  assign n10464 = n4025 & ~n10463 ;
  assign n10465 = n4202 & n9825 ;
  assign n10466 = ~n10461 & ~n10465 ;
  assign n10467 = n3829 & ~n10466 ;
  assign n10468 = n4202 & ~n9831 ;
  assign n10469 = ~n10461 & ~n10468 ;
  assign n10470 = n3969 & ~n10469 ;
  assign n10460 = \P1_reg1_reg[7]/NET0131  & ~n4218 ;
  assign n10471 = n3461 & n4028 ;
  assign n10472 = ~n9812 & ~n10471 ;
  assign n10473 = n4202 & ~n10472 ;
  assign n10474 = ~n10460 & ~n10473 ;
  assign n10475 = ~n10470 & n10474 ;
  assign n10476 = ~n10467 & n10475 ;
  assign n10477 = ~n10464 & n10476 ;
  assign n10478 = n2701 & ~n10477 ;
  assign n10479 = \P1_reg1_reg[7]/NET0131  & n4081 ;
  assign n10480 = ~n10478 & ~n10479 ;
  assign n10481 = \P1_state_reg[0]/NET0131  & ~n10480 ;
  assign n10482 = \P1_reg1_reg[7]/NET0131  & ~n4085 ;
  assign n10483 = ~n10481 & ~n10482 ;
  assign n10485 = n2717 & n9734 ;
  assign n10486 = \P1_reg2_reg[3]/NET0131  & ~n2717 ;
  assign n10487 = ~n10485 & ~n10486 ;
  assign n10488 = n4025 & ~n10487 ;
  assign n10489 = n2717 & ~n9741 ;
  assign n10490 = ~n10486 & ~n10489 ;
  assign n10491 = n3829 & ~n10490 ;
  assign n10492 = n2717 & n9748 ;
  assign n10493 = ~n10486 & ~n10492 ;
  assign n10494 = n3969 & ~n10493 ;
  assign n10496 = n2717 & ~n10448 ;
  assign n10484 = \P1_reg2_reg[3]/NET0131  & ~n4071 ;
  assign n10495 = ~\P1_reg3_reg[3]/NET0131  & n4073 ;
  assign n10497 = ~n10484 & ~n10495 ;
  assign n10498 = ~n10496 & n10497 ;
  assign n10499 = ~n10494 & n10498 ;
  assign n10500 = ~n10491 & n10499 ;
  assign n10501 = ~n10488 & n10500 ;
  assign n10502 = n2701 & ~n10501 ;
  assign n10503 = \P1_reg2_reg[3]/NET0131  & n4081 ;
  assign n10504 = ~n10502 & ~n10503 ;
  assign n10505 = \P1_state_reg[0]/NET0131  & ~n10504 ;
  assign n10506 = \P1_reg2_reg[3]/NET0131  & ~n4085 ;
  assign n10507 = ~n10505 & ~n10506 ;
  assign n10508 = \P1_reg2_reg[6]/NET0131  & ~n4085 ;
  assign n10509 = \P1_reg2_reg[6]/NET0131  & n4081 ;
  assign n10511 = \P1_reg2_reg[6]/NET0131  & ~n2717 ;
  assign n10518 = n2717 & n9790 ;
  assign n10519 = ~n10511 & ~n10518 ;
  assign n10520 = n4025 & ~n10519 ;
  assign n10515 = n2717 & n9782 ;
  assign n10516 = ~n10511 & ~n10515 ;
  assign n10517 = n3829 & ~n10516 ;
  assign n10512 = n2717 & ~n9776 ;
  assign n10513 = ~n10511 & ~n10512 ;
  assign n10514 = n3969 & ~n10513 ;
  assign n10521 = n2717 & n9795 ;
  assign n10522 = ~n10511 & ~n10521 ;
  assign n10523 = n4062 & ~n10522 ;
  assign n10510 = \P1_reg2_reg[6]/NET0131  & ~n5148 ;
  assign n10524 = n3490 & n4073 ;
  assign n10525 = ~n3485 & n4028 ;
  assign n10526 = n2717 & n10525 ;
  assign n10527 = ~n10524 & ~n10526 ;
  assign n10528 = ~n10510 & n10527 ;
  assign n10529 = ~n10523 & n10528 ;
  assign n10530 = ~n10514 & n10529 ;
  assign n10531 = ~n10517 & n10530 ;
  assign n10532 = ~n10520 & n10531 ;
  assign n10533 = n2701 & ~n10532 ;
  assign n10534 = ~n10509 & ~n10533 ;
  assign n10535 = \P1_state_reg[0]/NET0131  & ~n10534 ;
  assign n10536 = ~n10508 & ~n10535 ;
  assign n10538 = \P1_reg2_reg[7]/NET0131  & ~n2717 ;
  assign n10539 = n2717 & n9819 ;
  assign n10540 = ~n10538 & ~n10539 ;
  assign n10541 = n4025 & ~n10540 ;
  assign n10542 = n2717 & n9825 ;
  assign n10543 = ~n10538 & ~n10542 ;
  assign n10544 = n3829 & ~n10543 ;
  assign n10545 = n2717 & ~n9831 ;
  assign n10546 = ~n10538 & ~n10545 ;
  assign n10547 = n3969 & ~n10546 ;
  assign n10537 = n2717 & ~n10472 ;
  assign n10548 = n3463 & n4073 ;
  assign n10549 = \P1_reg2_reg[7]/NET0131  & ~n4071 ;
  assign n10550 = ~n10548 & ~n10549 ;
  assign n10551 = ~n10537 & n10550 ;
  assign n10552 = ~n10547 & n10551 ;
  assign n10553 = ~n10544 & n10552 ;
  assign n10554 = ~n10541 & n10553 ;
  assign n10555 = n2701 & ~n10554 ;
  assign n10556 = \P1_reg2_reg[7]/NET0131  & n4081 ;
  assign n10557 = ~n10555 & ~n10556 ;
  assign n10558 = \P1_state_reg[0]/NET0131  & ~n10557 ;
  assign n10559 = \P1_reg2_reg[7]/NET0131  & ~n4085 ;
  assign n10560 = ~n10558 & ~n10559 ;
  assign n10561 = \P1_reg0_reg[3]/NET0131  & ~n4085 ;
  assign n10563 = \P1_reg0_reg[3]/NET0131  & ~n4869 ;
  assign n10564 = n4869 & n9734 ;
  assign n10565 = ~n10563 & ~n10564 ;
  assign n10566 = n4025 & ~n10565 ;
  assign n10567 = n4869 & ~n9741 ;
  assign n10568 = ~n10563 & ~n10567 ;
  assign n10569 = n3829 & ~n10568 ;
  assign n10570 = n4869 & n9748 ;
  assign n10571 = ~n10563 & ~n10570 ;
  assign n10572 = n3969 & ~n10571 ;
  assign n10562 = n4869 & ~n10448 ;
  assign n10573 = \P1_reg0_reg[3]/NET0131  & ~n5844 ;
  assign n10574 = ~n10562 & ~n10573 ;
  assign n10575 = ~n10572 & n10574 ;
  assign n10576 = ~n10569 & n10575 ;
  assign n10577 = ~n10566 & n10576 ;
  assign n10578 = n2701 & ~n10577 ;
  assign n10579 = \P1_reg0_reg[3]/NET0131  & n4081 ;
  assign n10580 = ~n10578 & ~n10579 ;
  assign n10581 = \P1_state_reg[0]/NET0131  & ~n10580 ;
  assign n10582 = ~n10561 & ~n10581 ;
  assign n10583 = \P1_reg0_reg[7]/NET0131  & ~n4085 ;
  assign n10585 = \P1_reg0_reg[7]/NET0131  & ~n4869 ;
  assign n10586 = n4869 & n9819 ;
  assign n10587 = ~n10585 & ~n10586 ;
  assign n10588 = n4025 & ~n10587 ;
  assign n10589 = n4869 & n9825 ;
  assign n10590 = ~n10585 & ~n10589 ;
  assign n10591 = n3829 & ~n10590 ;
  assign n10592 = n4869 & ~n9831 ;
  assign n10593 = ~n10585 & ~n10592 ;
  assign n10594 = n3969 & ~n10593 ;
  assign n10584 = n4869 & ~n10472 ;
  assign n10595 = \P1_reg0_reg[7]/NET0131  & ~n5844 ;
  assign n10596 = ~n10584 & ~n10595 ;
  assign n10597 = ~n10594 & n10596 ;
  assign n10598 = ~n10591 & n10597 ;
  assign n10599 = ~n10588 & n10598 ;
  assign n10600 = n2701 & ~n10599 ;
  assign n10601 = \P1_reg0_reg[7]/NET0131  & n4081 ;
  assign n10602 = ~n10600 & ~n10601 ;
  assign n10603 = \P1_state_reg[0]/NET0131  & ~n10602 ;
  assign n10604 = ~n10583 & ~n10603 ;
  assign n10605 = \P2_reg3_reg[2]/NET0131  & ~n2286 ;
  assign n10606 = \P2_reg3_reg[2]/NET0131  & n2035 ;
  assign n10616 = \P2_reg3_reg[2]/NET0131  & ~n2124 ;
  assign n10623 = n1086 & ~n2233 ;
  assign n10624 = n2263 & ~n9172 ;
  assign n10625 = ~n10623 & n10624 ;
  assign n10626 = ~n1134 & ~n2263 ;
  assign n10627 = ~n10625 & ~n10626 ;
  assign n10628 = n2124 & ~n10627 ;
  assign n10629 = ~n10616 & ~n10628 ;
  assign n10630 = n1790 & ~n10629 ;
  assign n10608 = \P2_reg3_reg[2]/NET0131  & ~n2053 ;
  assign n10609 = n1803 & ~n1917 ;
  assign n10610 = ~n1803 & n1917 ;
  assign n10611 = ~n10609 & ~n10610 ;
  assign n10612 = n2053 & ~n10611 ;
  assign n10613 = ~n10608 & ~n10612 ;
  assign n10614 = ~n2120 & ~n10613 ;
  assign n10607 = \P2_reg3_reg[2]/NET0131  & ~n2274 ;
  assign n10615 = ~n1124 & n2229 ;
  assign n10634 = ~n10607 & ~n10615 ;
  assign n10635 = ~n10614 & n10634 ;
  assign n10617 = n1917 & ~n2137 ;
  assign n10618 = ~n1917 & n2137 ;
  assign n10619 = ~n10617 & ~n10618 ;
  assign n10620 = n2124 & ~n10619 ;
  assign n10621 = ~n10616 & ~n10620 ;
  assign n10622 = n2123 & ~n10621 ;
  assign n10631 = n2053 & ~n10619 ;
  assign n10632 = ~n10608 & ~n10631 ;
  assign n10633 = ~n2224 & ~n10632 ;
  assign n10636 = ~n10622 & ~n10633 ;
  assign n10637 = n10635 & n10636 ;
  assign n10638 = ~n10630 & n10637 ;
  assign n10639 = n2037 & ~n10638 ;
  assign n10640 = ~n10606 & ~n10639 ;
  assign n10641 = \P1_state_reg[0]/NET0131  & ~n10640 ;
  assign n10642 = ~n10605 & ~n10641 ;
  assign n10643 = \P1_reg1_reg[6]/NET0131  & ~n4085 ;
  assign n10644 = \P1_reg1_reg[6]/NET0131  & n4081 ;
  assign n10646 = \P1_reg1_reg[6]/NET0131  & ~n4202 ;
  assign n10653 = n4202 & n9790 ;
  assign n10654 = ~n10646 & ~n10653 ;
  assign n10655 = n4025 & ~n10654 ;
  assign n10650 = n4202 & ~n9776 ;
  assign n10651 = ~n10646 & ~n10650 ;
  assign n10652 = n3969 & ~n10651 ;
  assign n10647 = n4202 & n9782 ;
  assign n10648 = ~n10646 & ~n10647 ;
  assign n10649 = n3829 & ~n10648 ;
  assign n10656 = n4202 & n9795 ;
  assign n10657 = ~n10646 & ~n10656 ;
  assign n10658 = n4062 & ~n10657 ;
  assign n10645 = n4202 & n10525 ;
  assign n10659 = \P1_reg1_reg[6]/NET0131  & ~n4216 ;
  assign n10660 = ~n10645 & ~n10659 ;
  assign n10661 = ~n10658 & n10660 ;
  assign n10662 = ~n10649 & n10661 ;
  assign n10663 = ~n10652 & n10662 ;
  assign n10664 = ~n10655 & n10663 ;
  assign n10665 = n2701 & ~n10664 ;
  assign n10666 = ~n10644 & ~n10665 ;
  assign n10667 = \P1_state_reg[0]/NET0131  & ~n10666 ;
  assign n10668 = ~n10643 & ~n10667 ;
  assign n10669 = \P2_reg0_reg[3]/NET0131  & ~n2286 ;
  assign n10670 = \P2_reg0_reg[3]/NET0131  & n2035 ;
  assign n10676 = n2053 & n10419 ;
  assign n10677 = ~\P2_reg0_reg[3]/NET0131  & ~n2053 ;
  assign n10678 = n1790 & ~n10677 ;
  assign n10679 = ~n10676 & n10678 ;
  assign n10673 = \P2_reg0_reg[3]/NET0131  & ~n2124 ;
  assign n10680 = n2124 & n10410 ;
  assign n10681 = ~n10673 & ~n10680 ;
  assign n10682 = ~n2120 & ~n10681 ;
  assign n10674 = ~n10404 & ~n10673 ;
  assign n10675 = ~n2224 & ~n10674 ;
  assign n10684 = n2053 & n10403 ;
  assign n10685 = n2123 & ~n10677 ;
  assign n10686 = ~n10684 & n10685 ;
  assign n10671 = ~n1100 & n2272 ;
  assign n10672 = n2124 & n10671 ;
  assign n10683 = \P2_reg0_reg[3]/NET0131  & ~n2614 ;
  assign n10687 = ~n10672 & ~n10683 ;
  assign n10688 = ~n10686 & n10687 ;
  assign n10689 = ~n10675 & n10688 ;
  assign n10690 = ~n10682 & n10689 ;
  assign n10691 = ~n10679 & n10690 ;
  assign n10692 = n2037 & ~n10691 ;
  assign n10693 = ~n10670 & ~n10692 ;
  assign n10694 = \P1_state_reg[0]/NET0131  & ~n10693 ;
  assign n10695 = ~n10669 & ~n10694 ;
  assign n10696 = \P2_reg0_reg[4]/NET0131  & ~n2286 ;
  assign n10697 = \P2_reg0_reg[4]/NET0131  & n2035 ;
  assign n10707 = \P2_reg0_reg[4]/NET0131  & ~n2053 ;
  assign n10708 = n2053 & ~n9872 ;
  assign n10709 = ~n10707 & ~n10708 ;
  assign n10710 = n1790 & ~n10709 ;
  assign n10700 = \P2_reg0_reg[4]/NET0131  & ~n2124 ;
  assign n10701 = n2124 & ~n9856 ;
  assign n10702 = ~n10700 & ~n10701 ;
  assign n10703 = ~n2120 & ~n10702 ;
  assign n10698 = ~n1076 & n2272 ;
  assign n10699 = n2124 & n10698 ;
  assign n10704 = \P2_reg0_reg[4]/NET0131  & ~n2614 ;
  assign n10713 = ~n10699 & ~n10704 ;
  assign n10714 = ~n10703 & n10713 ;
  assign n10705 = ~n9876 & ~n10700 ;
  assign n10706 = ~n2224 & ~n10705 ;
  assign n10711 = ~n9864 & ~n10707 ;
  assign n10712 = n2123 & ~n10711 ;
  assign n10715 = ~n10706 & ~n10712 ;
  assign n10716 = n10714 & n10715 ;
  assign n10717 = ~n10710 & n10716 ;
  assign n10718 = n2037 & ~n10717 ;
  assign n10719 = ~n10697 & ~n10718 ;
  assign n10720 = \P1_state_reg[0]/NET0131  & ~n10719 ;
  assign n10721 = ~n10696 & ~n10720 ;
  assign n10722 = \P2_reg1_reg[3]/NET0131  & ~n2286 ;
  assign n10723 = \P2_reg1_reg[3]/NET0131  & n2035 ;
  assign n10733 = \P2_reg1_reg[3]/NET0131  & ~n2291 ;
  assign n10734 = n2291 & ~n10419 ;
  assign n10735 = ~n10733 & ~n10734 ;
  assign n10736 = n1790 & ~n10735 ;
  assign n10725 = \P2_reg1_reg[3]/NET0131  & ~n2310 ;
  assign n10726 = n2310 & ~n10403 ;
  assign n10727 = ~n10725 & ~n10726 ;
  assign n10728 = ~n2392 & ~n10727 ;
  assign n10724 = n2310 & n10671 ;
  assign n10729 = \P2_reg1_reg[3]/NET0131  & ~n4099 ;
  assign n10740 = ~n10724 & ~n10729 ;
  assign n10741 = ~n10728 & n10740 ;
  assign n10730 = n2310 & n10410 ;
  assign n10731 = ~n10725 & ~n10730 ;
  assign n10732 = ~n2290 & ~n10731 ;
  assign n10737 = n2291 & n10410 ;
  assign n10738 = ~n10733 & ~n10737 ;
  assign n10739 = n2314 & ~n10738 ;
  assign n10742 = ~n10732 & ~n10739 ;
  assign n10743 = n10741 & n10742 ;
  assign n10744 = ~n10736 & n10743 ;
  assign n10745 = n2037 & ~n10744 ;
  assign n10746 = ~n10723 & ~n10745 ;
  assign n10747 = \P1_state_reg[0]/NET0131  & ~n10746 ;
  assign n10748 = ~n10722 & ~n10747 ;
  assign n10749 = \P2_reg1_reg[4]/NET0131  & ~n2286 ;
  assign n10750 = \P2_reg1_reg[4]/NET0131  & n2035 ;
  assign n10752 = \P2_reg1_reg[4]/NET0131  & ~n2291 ;
  assign n10761 = n2291 & ~n9872 ;
  assign n10762 = ~n10752 & ~n10761 ;
  assign n10763 = n1790 & ~n10762 ;
  assign n10753 = n2291 & ~n9856 ;
  assign n10754 = ~n10752 & ~n10753 ;
  assign n10755 = n2314 & ~n10754 ;
  assign n10751 = n2310 & n10698 ;
  assign n10756 = \P2_reg1_reg[4]/NET0131  & ~n4099 ;
  assign n10767 = ~n10751 & ~n10756 ;
  assign n10768 = ~n10755 & n10767 ;
  assign n10757 = \P2_reg1_reg[4]/NET0131  & ~n2310 ;
  assign n10758 = n2310 & ~n9856 ;
  assign n10759 = ~n10757 & ~n10758 ;
  assign n10760 = ~n2290 & ~n10759 ;
  assign n10764 = n2310 & n9863 ;
  assign n10765 = ~n10757 & ~n10764 ;
  assign n10766 = ~n2392 & ~n10765 ;
  assign n10769 = ~n10760 & ~n10766 ;
  assign n10770 = n10768 & n10769 ;
  assign n10771 = ~n10763 & n10770 ;
  assign n10772 = n2037 & ~n10771 ;
  assign n10773 = ~n10750 & ~n10772 ;
  assign n10774 = \P1_state_reg[0]/NET0131  & ~n10773 ;
  assign n10775 = ~n10749 & ~n10774 ;
  assign n10776 = \P2_reg2_reg[3]/NET0131  & ~n2286 ;
  assign n10777 = \P2_reg2_reg[3]/NET0131  & n2035 ;
  assign n10779 = \P2_reg2_reg[3]/NET0131  & ~n2310 ;
  assign n10788 = n2310 & ~n10419 ;
  assign n10789 = ~n10779 & ~n10788 ;
  assign n10790 = n1790 & ~n10789 ;
  assign n10780 = ~n10730 & ~n10779 ;
  assign n10781 = n2314 & ~n10780 ;
  assign n10792 = \P2_reg2_reg[3]/NET0131  & ~n2407 ;
  assign n10778 = n2291 & n10671 ;
  assign n10791 = ~\P2_reg3_reg[3]/NET0131  & n1854 ;
  assign n10793 = ~n10778 & ~n10791 ;
  assign n10794 = ~n10792 & n10793 ;
  assign n10795 = ~n10781 & n10794 ;
  assign n10782 = \P2_reg2_reg[3]/NET0131  & ~n2291 ;
  assign n10783 = n2291 & ~n10403 ;
  assign n10784 = ~n10782 & ~n10783 ;
  assign n10785 = ~n2392 & ~n10784 ;
  assign n10786 = ~n10737 & ~n10782 ;
  assign n10787 = ~n2290 & ~n10786 ;
  assign n10796 = ~n10785 & ~n10787 ;
  assign n10797 = n10795 & n10796 ;
  assign n10798 = ~n10790 & n10797 ;
  assign n10799 = n2037 & ~n10798 ;
  assign n10800 = ~n10777 & ~n10799 ;
  assign n10801 = \P1_state_reg[0]/NET0131  & ~n10800 ;
  assign n10802 = ~n10776 & ~n10801 ;
  assign n10803 = \P2_reg2_reg[4]/NET0131  & ~n2286 ;
  assign n10804 = \P2_reg2_reg[4]/NET0131  & n2035 ;
  assign n10809 = \P2_reg2_reg[4]/NET0131  & ~n2310 ;
  assign n10812 = n2310 & ~n9872 ;
  assign n10813 = ~n10809 & ~n10812 ;
  assign n10814 = n1790 & ~n10813 ;
  assign n10806 = \P2_reg2_reg[4]/NET0131  & ~n2291 ;
  assign n10807 = ~n10753 & ~n10806 ;
  assign n10808 = ~n2290 & ~n10807 ;
  assign n10819 = \P2_reg2_reg[4]/NET0131  & ~n2407 ;
  assign n10805 = n2291 & n10698 ;
  assign n10818 = ~n1055 & n1854 ;
  assign n10820 = ~n10805 & ~n10818 ;
  assign n10821 = ~n10819 & n10820 ;
  assign n10822 = ~n10808 & n10821 ;
  assign n10810 = ~n10758 & ~n10809 ;
  assign n10811 = n2314 & ~n10810 ;
  assign n10815 = n2291 & n9863 ;
  assign n10816 = ~n10806 & ~n10815 ;
  assign n10817 = ~n2392 & ~n10816 ;
  assign n10823 = ~n10811 & ~n10817 ;
  assign n10824 = n10822 & n10823 ;
  assign n10825 = ~n10814 & n10824 ;
  assign n10826 = n2037 & ~n10825 ;
  assign n10827 = ~n10804 & ~n10826 ;
  assign n10828 = \P1_state_reg[0]/NET0131  & ~n10827 ;
  assign n10829 = ~n10803 & ~n10828 ;
  assign n10830 = \P1_reg0_reg[6]/NET0131  & ~n4085 ;
  assign n10831 = \P1_reg0_reg[6]/NET0131  & n4081 ;
  assign n10833 = \P1_reg0_reg[6]/NET0131  & ~n4869 ;
  assign n10840 = n4869 & n9790 ;
  assign n10841 = ~n10833 & ~n10840 ;
  assign n10842 = n4025 & ~n10841 ;
  assign n10837 = n4869 & ~n9776 ;
  assign n10838 = ~n10833 & ~n10837 ;
  assign n10839 = n3969 & ~n10838 ;
  assign n10834 = n4869 & n9782 ;
  assign n10835 = ~n10833 & ~n10834 ;
  assign n10836 = n3829 & ~n10835 ;
  assign n10843 = n4869 & n9795 ;
  assign n10844 = ~n10833 & ~n10843 ;
  assign n10845 = n4062 & ~n10844 ;
  assign n10832 = n4869 & n10525 ;
  assign n10846 = \P1_reg0_reg[6]/NET0131  & ~n5864 ;
  assign n10847 = ~n10832 & ~n10846 ;
  assign n10848 = ~n10845 & n10847 ;
  assign n10849 = ~n10836 & n10848 ;
  assign n10850 = ~n10839 & n10849 ;
  assign n10851 = ~n10842 & n10850 ;
  assign n10852 = n2701 & ~n10851 ;
  assign n10853 = ~n10831 & ~n10852 ;
  assign n10854 = \P1_state_reg[0]/NET0131  & ~n10853 ;
  assign n10855 = ~n10830 & ~n10854 ;
  assign n10856 = \P1_reg3_reg[1]/NET0131  & ~n4085 ;
  assign n10857 = \P1_reg3_reg[1]/NET0131  & n4081 ;
  assign n10868 = ~n3412 & n5427 ;
  assign n10869 = n3412 & ~n5427 ;
  assign n10870 = ~n10868 & ~n10869 ;
  assign n10872 = ~n3411 & n10870 ;
  assign n10873 = n3411 & n5427 ;
  assign n10874 = ~n10872 & ~n10873 ;
  assign n10875 = n3969 & n10874 ;
  assign n10871 = n3829 & n10870 ;
  assign n10876 = ~n3395 & ~n3411 ;
  assign n10877 = ~n4030 & n4062 ;
  assign n10878 = ~n10876 & n10877 ;
  assign n10879 = ~n10871 & ~n10878 ;
  assign n10880 = ~n10875 & n10879 ;
  assign n10881 = n4449 & ~n10880 ;
  assign n10859 = \P1_reg3_reg[1]/NET0131  & ~n4449 ;
  assign n10860 = n3340 & ~n3986 ;
  assign n10861 = ~n3987 & ~n10860 ;
  assign n10862 = ~n2731 & ~n10861 ;
  assign n10863 = n2731 & n3404 ;
  assign n10864 = ~n10862 & ~n10863 ;
  assign n10865 = n4449 & n10864 ;
  assign n10866 = ~n10859 & ~n10865 ;
  assign n10867 = n4025 & ~n10866 ;
  assign n10886 = ~n3395 & n4449 ;
  assign n10887 = ~n10859 & ~n10886 ;
  assign n10888 = n4028 & ~n10887 ;
  assign n10858 = ~n3395 & n4073 ;
  assign n10882 = ~n3816 & ~n5408 ;
  assign n10883 = ~n4449 & ~n10882 ;
  assign n10884 = ~n4067 & ~n10883 ;
  assign n10885 = \P1_reg3_reg[1]/NET0131  & ~n10884 ;
  assign n10889 = ~n10858 & ~n10885 ;
  assign n10890 = ~n10888 & n10889 ;
  assign n10891 = ~n10867 & n10890 ;
  assign n10892 = ~n10881 & n10891 ;
  assign n10893 = n2701 & ~n10892 ;
  assign n10894 = ~n10857 & ~n10893 ;
  assign n10895 = \P1_state_reg[0]/NET0131  & ~n10894 ;
  assign n10896 = ~n10856 & ~n10895 ;
  assign n10897 = \P2_reg3_reg[1]/NET0131  & ~n2286 ;
  assign n10898 = \P2_reg3_reg[1]/NET0131  & n2035 ;
  assign n10910 = \P2_reg3_reg[1]/NET0131  & ~n2124 ;
  assign n10911 = n1110 & ~n2232 ;
  assign n10912 = ~n2233 & n2263 ;
  assign n10913 = ~n10911 & n10912 ;
  assign n10914 = ~n1158 & ~n2263 ;
  assign n10915 = ~n10913 & ~n10914 ;
  assign n10916 = n2124 & ~n10915 ;
  assign n10917 = ~n10910 & ~n10916 ;
  assign n10918 = n1790 & ~n10917 ;
  assign n10900 = \P2_reg3_reg[1]/NET0131  & ~n2053 ;
  assign n10904 = ~n1801 & ~n1904 ;
  assign n10905 = n1801 & n1904 ;
  assign n10906 = ~n10904 & ~n10905 ;
  assign n10907 = n2053 & ~n10906 ;
  assign n10908 = ~n10900 & ~n10907 ;
  assign n10909 = ~n2120 & ~n10908 ;
  assign n10901 = ~n1148 & n2053 ;
  assign n10902 = ~n10900 & ~n10901 ;
  assign n10903 = n2272 & ~n10902 ;
  assign n10899 = \P2_reg3_reg[1]/NET0131  & n2271 ;
  assign n10928 = ~n1148 & n1854 ;
  assign n10929 = ~n10899 & ~n10928 ;
  assign n10930 = ~n10903 & n10929 ;
  assign n10931 = ~n10909 & n10930 ;
  assign n10919 = n1904 & ~n2135 ;
  assign n10920 = ~n1904 & n2135 ;
  assign n10921 = ~n10919 & ~n10920 ;
  assign n10922 = n2053 & n10921 ;
  assign n10923 = ~n10900 & ~n10922 ;
  assign n10924 = ~n2224 & ~n10923 ;
  assign n10925 = n2124 & n10921 ;
  assign n10926 = ~n10910 & ~n10925 ;
  assign n10927 = n2123 & ~n10926 ;
  assign n10932 = ~n10924 & ~n10927 ;
  assign n10933 = n10931 & n10932 ;
  assign n10934 = ~n10918 & n10933 ;
  assign n10935 = n2037 & ~n10934 ;
  assign n10936 = ~n10898 & ~n10935 ;
  assign n10937 = \P1_state_reg[0]/NET0131  & ~n10936 ;
  assign n10938 = ~n10897 & ~n10937 ;
  assign n10939 = \P1_reg3_reg[2]/NET0131  & ~n4085 ;
  assign n10940 = \P1_reg3_reg[2]/NET0131  & n4081 ;
  assign n10942 = \P1_reg3_reg[2]/NET0131  & ~n4449 ;
  assign n10955 = n523 & ~n3987 ;
  assign n10956 = ~n3988 & ~n10955 ;
  assign n10957 = ~n2731 & ~n10956 ;
  assign n10958 = n2731 & n3381 ;
  assign n10959 = ~n10957 & ~n10958 ;
  assign n10960 = n4449 & n10959 ;
  assign n10961 = ~n10942 & ~n10960 ;
  assign n10962 = n4025 & ~n10961 ;
  assign n10949 = n4725 & ~n5429 ;
  assign n10950 = ~n4725 & n5429 ;
  assign n10951 = ~n10949 & ~n10950 ;
  assign n10952 = n4449 & n10951 ;
  assign n10953 = ~n10942 & ~n10952 ;
  assign n10954 = n3969 & ~n10953 ;
  assign n10943 = ~n3414 & n5429 ;
  assign n10944 = n3414 & ~n5429 ;
  assign n10945 = ~n10943 & ~n10944 ;
  assign n10946 = n4449 & ~n10945 ;
  assign n10947 = ~n10942 & ~n10946 ;
  assign n10948 = n3829 & ~n10947 ;
  assign n10963 = ~n3354 & ~n4030 ;
  assign n10964 = ~n4031 & ~n10963 ;
  assign n10965 = n4449 & n10964 ;
  assign n10966 = ~n10942 & ~n10965 ;
  assign n10967 = n4062 & ~n10966 ;
  assign n10941 = ~n3354 & ~n4522 ;
  assign n10968 = \P1_reg3_reg[2]/NET0131  & ~n4540 ;
  assign n10969 = ~n10941 & ~n10968 ;
  assign n10970 = ~n10967 & n10969 ;
  assign n10971 = ~n10948 & n10970 ;
  assign n10972 = ~n10954 & n10971 ;
  assign n10973 = ~n10962 & n10972 ;
  assign n10974 = n2701 & ~n10973 ;
  assign n10975 = ~n10940 & ~n10974 ;
  assign n10976 = \P1_state_reg[0]/NET0131  & ~n10975 ;
  assign n10977 = ~n10939 & ~n10976 ;
  assign n10978 = \P2_reg0_reg[2]/NET0131  & ~n2286 ;
  assign n10979 = \P2_reg0_reg[2]/NET0131  & n2035 ;
  assign n10986 = \P2_reg0_reg[2]/NET0131  & ~n2053 ;
  assign n10989 = n2053 & ~n10627 ;
  assign n10990 = ~n10986 & ~n10989 ;
  assign n10991 = n1790 & ~n10990 ;
  assign n10982 = \P2_reg0_reg[2]/NET0131  & ~n2124 ;
  assign n10983 = ~n10620 & ~n10982 ;
  assign n10984 = ~n2224 & ~n10983 ;
  assign n10980 = ~n1124 & n2272 ;
  assign n10981 = n2124 & n10980 ;
  assign n10985 = \P2_reg0_reg[2]/NET0131  & ~n2614 ;
  assign n10995 = ~n10981 & ~n10985 ;
  assign n10996 = ~n10984 & n10995 ;
  assign n10987 = ~n10631 & ~n10986 ;
  assign n10988 = n2123 & ~n10987 ;
  assign n10992 = n2124 & ~n10611 ;
  assign n10993 = ~n10982 & ~n10992 ;
  assign n10994 = ~n2120 & ~n10993 ;
  assign n10997 = ~n10988 & ~n10994 ;
  assign n10998 = n10996 & n10997 ;
  assign n10999 = ~n10991 & n10998 ;
  assign n11000 = n2037 & ~n10999 ;
  assign n11001 = ~n10979 & ~n11000 ;
  assign n11002 = \P1_state_reg[0]/NET0131  & ~n11001 ;
  assign n11003 = ~n10978 & ~n11002 ;
  assign n11004 = \P2_reg1_reg[2]/NET0131  & ~n2286 ;
  assign n11005 = \P2_reg1_reg[2]/NET0131  & n2035 ;
  assign n11006 = \P2_reg1_reg[2]/NET0131  & ~n2291 ;
  assign n11020 = n2291 & ~n10627 ;
  assign n11021 = ~n11006 & ~n11020 ;
  assign n11022 = n1790 & ~n11021 ;
  assign n11011 = ~n2290 & ~n10611 ;
  assign n11010 = ~n2392 & ~n10619 ;
  assign n11012 = ~n10980 & ~n11010 ;
  assign n11013 = ~n11011 & n11012 ;
  assign n11014 = n2310 & ~n11013 ;
  assign n11007 = n2291 & ~n10611 ;
  assign n11008 = ~n11006 & ~n11007 ;
  assign n11009 = n2314 & ~n11008 ;
  assign n11015 = ~n1989 & ~n2122 ;
  assign n11016 = ~n2289 & n11015 ;
  assign n11017 = ~n2310 & ~n11016 ;
  assign n11018 = n4099 & ~n11017 ;
  assign n11019 = \P2_reg1_reg[2]/NET0131  & ~n11018 ;
  assign n11023 = ~n11009 & ~n11019 ;
  assign n11024 = ~n11014 & n11023 ;
  assign n11025 = ~n11022 & n11024 ;
  assign n11026 = n2037 & ~n11025 ;
  assign n11027 = ~n11005 & ~n11026 ;
  assign n11028 = \P1_state_reg[0]/NET0131  & ~n11027 ;
  assign n11029 = ~n11004 & ~n11028 ;
  assign n11030 = \P2_reg2_reg[2]/NET0131  & ~n2286 ;
  assign n11031 = \P2_reg2_reg[2]/NET0131  & n2035 ;
  assign n11040 = \P2_reg2_reg[2]/NET0131  & ~n2310 ;
  assign n11044 = n2310 & ~n10627 ;
  assign n11045 = ~n11040 & ~n11044 ;
  assign n11046 = n1790 & ~n11045 ;
  assign n11033 = \P2_reg2_reg[2]/NET0131  & ~n2291 ;
  assign n11034 = ~n11007 & ~n11033 ;
  assign n11035 = ~n2290 & ~n11034 ;
  assign n11047 = \P2_reg2_reg[2]/NET0131  & ~n2407 ;
  assign n11032 = n2291 & n10980 ;
  assign n11039 = \P2_reg3_reg[2]/NET0131  & n1854 ;
  assign n11048 = ~n11032 & ~n11039 ;
  assign n11049 = ~n11047 & n11048 ;
  assign n11050 = ~n11035 & n11049 ;
  assign n11036 = n2291 & ~n10619 ;
  assign n11037 = ~n11033 & ~n11036 ;
  assign n11038 = ~n2392 & ~n11037 ;
  assign n11041 = n2310 & ~n10611 ;
  assign n11042 = ~n11040 & ~n11041 ;
  assign n11043 = n2314 & ~n11042 ;
  assign n11051 = ~n11038 & ~n11043 ;
  assign n11052 = n11050 & n11051 ;
  assign n11053 = ~n11046 & n11052 ;
  assign n11054 = n2037 & ~n11053 ;
  assign n11055 = ~n11031 & ~n11054 ;
  assign n11056 = \P1_state_reg[0]/NET0131  & ~n11055 ;
  assign n11057 = ~n11030 & ~n11056 ;
  assign n11058 = \P1_reg0_reg[2]/NET0131  & ~n4085 ;
  assign n11059 = \P1_reg0_reg[2]/NET0131  & n4081 ;
  assign n11062 = \P1_reg0_reg[2]/NET0131  & ~n4869 ;
  assign n11069 = n4869 & n10959 ;
  assign n11070 = ~n11062 & ~n11069 ;
  assign n11071 = n4025 & ~n11070 ;
  assign n11066 = n4869 & ~n10945 ;
  assign n11067 = ~n11062 & ~n11066 ;
  assign n11068 = n3829 & ~n11067 ;
  assign n11063 = n4869 & n10951 ;
  assign n11064 = ~n11062 & ~n11063 ;
  assign n11065 = n3969 & ~n11064 ;
  assign n11072 = n4869 & n10964 ;
  assign n11073 = ~n11062 & ~n11072 ;
  assign n11074 = n4062 & ~n11073 ;
  assign n11060 = ~n3354 & n4028 ;
  assign n11061 = n4869 & n11060 ;
  assign n11075 = \P1_reg0_reg[2]/NET0131  & ~n5864 ;
  assign n11076 = ~n11061 & ~n11075 ;
  assign n11077 = ~n11074 & n11076 ;
  assign n11078 = ~n11065 & n11077 ;
  assign n11079 = ~n11068 & n11078 ;
  assign n11080 = ~n11071 & n11079 ;
  assign n11081 = n2701 & ~n11080 ;
  assign n11082 = ~n11059 & ~n11081 ;
  assign n11083 = \P1_state_reg[0]/NET0131  & ~n11082 ;
  assign n11084 = ~n11058 & ~n11083 ;
  assign n11085 = \P1_reg1_reg[2]/NET0131  & ~n4085 ;
  assign n11086 = \P1_reg1_reg[2]/NET0131  & n4081 ;
  assign n11088 = \P1_reg1_reg[2]/NET0131  & ~n4202 ;
  assign n11095 = n4202 & n10959 ;
  assign n11096 = ~n11088 & ~n11095 ;
  assign n11097 = n4025 & ~n11096 ;
  assign n11092 = n4202 & ~n10945 ;
  assign n11093 = ~n11088 & ~n11092 ;
  assign n11094 = n3829 & ~n11093 ;
  assign n11089 = n4202 & n10951 ;
  assign n11090 = ~n11088 & ~n11089 ;
  assign n11091 = n3969 & ~n11090 ;
  assign n11098 = n4202 & n10964 ;
  assign n11099 = ~n11088 & ~n11098 ;
  assign n11100 = n4062 & ~n11099 ;
  assign n11087 = n4202 & n11060 ;
  assign n11101 = \P1_reg1_reg[2]/NET0131  & ~n4216 ;
  assign n11102 = ~n11087 & ~n11101 ;
  assign n11103 = ~n11100 & n11102 ;
  assign n11104 = ~n11091 & n11103 ;
  assign n11105 = ~n11094 & n11104 ;
  assign n11106 = ~n11097 & n11105 ;
  assign n11107 = n2701 & ~n11106 ;
  assign n11108 = ~n11086 & ~n11107 ;
  assign n11109 = \P1_state_reg[0]/NET0131  & ~n11108 ;
  assign n11110 = ~n11085 & ~n11109 ;
  assign n11111 = \P2_reg0_reg[1]/NET0131  & ~n2286 ;
  assign n11112 = \P2_reg0_reg[1]/NET0131  & n2035 ;
  assign n11114 = \P2_reg0_reg[1]/NET0131  & ~n2053 ;
  assign n11123 = n2053 & ~n10915 ;
  assign n11124 = ~n11114 & ~n11123 ;
  assign n11125 = n1790 & ~n11124 ;
  assign n11115 = ~n10922 & ~n11114 ;
  assign n11116 = n2123 & ~n11115 ;
  assign n11113 = \P2_reg0_reg[1]/NET0131  & ~n2612 ;
  assign n11117 = \P2_reg0_reg[1]/NET0131  & ~n2124 ;
  assign n11126 = ~n1148 & n2124 ;
  assign n11127 = ~n11117 & ~n11126 ;
  assign n11128 = n2272 & ~n11127 ;
  assign n11129 = ~n11113 & ~n11128 ;
  assign n11130 = ~n11116 & n11129 ;
  assign n11118 = ~n10925 & ~n11117 ;
  assign n11119 = ~n2224 & ~n11118 ;
  assign n11120 = n2124 & ~n10906 ;
  assign n11121 = ~n11117 & ~n11120 ;
  assign n11122 = ~n2120 & ~n11121 ;
  assign n11131 = ~n11119 & ~n11122 ;
  assign n11132 = n11130 & n11131 ;
  assign n11133 = ~n11125 & n11132 ;
  assign n11134 = n2037 & ~n11133 ;
  assign n11135 = ~n11112 & ~n11134 ;
  assign n11136 = \P1_state_reg[0]/NET0131  & ~n11135 ;
  assign n11137 = ~n11111 & ~n11136 ;
  assign n11138 = \P2_reg1_reg[1]/NET0131  & ~n2286 ;
  assign n11139 = \P2_reg1_reg[1]/NET0131  & n2035 ;
  assign n11141 = \P2_reg1_reg[1]/NET0131  & ~n2291 ;
  assign n11152 = n2291 & ~n10915 ;
  assign n11153 = ~n11141 & ~n11152 ;
  assign n11154 = n1790 & ~n11153 ;
  assign n11142 = n2291 & ~n10906 ;
  assign n11143 = ~n11141 & ~n11142 ;
  assign n11144 = n2314 & ~n11143 ;
  assign n11140 = \P2_reg1_reg[1]/NET0131  & ~n2612 ;
  assign n11145 = \P2_reg1_reg[1]/NET0131  & ~n2310 ;
  assign n11155 = ~n1148 & n2310 ;
  assign n11156 = ~n11145 & ~n11155 ;
  assign n11157 = n2272 & ~n11156 ;
  assign n11158 = ~n11140 & ~n11157 ;
  assign n11159 = ~n11144 & n11158 ;
  assign n11146 = n2310 & ~n10906 ;
  assign n11147 = ~n11145 & ~n11146 ;
  assign n11148 = ~n2290 & ~n11147 ;
  assign n11149 = n2310 & n10921 ;
  assign n11150 = ~n11145 & ~n11149 ;
  assign n11151 = ~n2392 & ~n11150 ;
  assign n11160 = ~n11148 & ~n11151 ;
  assign n11161 = n11159 & n11160 ;
  assign n11162 = ~n11154 & n11161 ;
  assign n11163 = n2037 & ~n11162 ;
  assign n11164 = ~n11139 & ~n11163 ;
  assign n11165 = \P1_state_reg[0]/NET0131  & ~n11164 ;
  assign n11166 = ~n11138 & ~n11165 ;
  assign n11167 = \P1_reg2_reg[2]/NET0131  & ~n4085 ;
  assign n11168 = \P1_reg2_reg[2]/NET0131  & n4081 ;
  assign n11170 = \P1_reg2_reg[2]/NET0131  & ~n2717 ;
  assign n11171 = n2717 & n10959 ;
  assign n11172 = ~n11170 & ~n11171 ;
  assign n11173 = n4025 & ~n11172 ;
  assign n11175 = n3829 & ~n10945 ;
  assign n11174 = n3969 & n10951 ;
  assign n11176 = n4062 & n10964 ;
  assign n11177 = ~n11174 & ~n11176 ;
  assign n11178 = ~n11175 & n11177 ;
  assign n11179 = n2717 & ~n11178 ;
  assign n11183 = ~n2717 & n3816 ;
  assign n11184 = ~n4067 & ~n7056 ;
  assign n11185 = ~n11183 & n11184 ;
  assign n11186 = \P1_reg2_reg[2]/NET0131  & ~n11185 ;
  assign n11169 = \P1_reg3_reg[2]/NET0131  & n4073 ;
  assign n11180 = n2717 & ~n3354 ;
  assign n11181 = ~n11170 & ~n11180 ;
  assign n11182 = n4028 & ~n11181 ;
  assign n11187 = ~n11169 & ~n11182 ;
  assign n11188 = ~n11186 & n11187 ;
  assign n11189 = ~n11179 & n11188 ;
  assign n11190 = ~n11173 & n11189 ;
  assign n11191 = n2701 & ~n11190 ;
  assign n11192 = ~n11168 & ~n11191 ;
  assign n11193 = \P1_state_reg[0]/NET0131  & ~n11192 ;
  assign n11194 = ~n11167 & ~n11193 ;
  assign n11195 = \P2_reg2_reg[1]/NET0131  & ~n2286 ;
  assign n11196 = \P2_reg2_reg[1]/NET0131  & n2035 ;
  assign n11198 = \P2_reg2_reg[1]/NET0131  & ~n2310 ;
  assign n11204 = n2310 & ~n10915 ;
  assign n11205 = ~n11198 & ~n11204 ;
  assign n11206 = n1790 & ~n11205 ;
  assign n11199 = ~n11146 & ~n11198 ;
  assign n11200 = n2314 & ~n11199 ;
  assign n11201 = \P2_reg2_reg[1]/NET0131  & ~n2291 ;
  assign n11207 = ~n1148 & n2291 ;
  assign n11208 = ~n11201 & ~n11207 ;
  assign n11209 = n2272 & ~n11208 ;
  assign n11197 = \P2_reg3_reg[1]/NET0131  & n1854 ;
  assign n11213 = \P2_reg2_reg[1]/NET0131  & n2271 ;
  assign n11214 = ~n11197 & ~n11213 ;
  assign n11215 = ~n11209 & n11214 ;
  assign n11216 = ~n11200 & n11215 ;
  assign n11202 = ~n11142 & ~n11201 ;
  assign n11203 = ~n2290 & ~n11202 ;
  assign n11210 = n2291 & n10921 ;
  assign n11211 = ~n11201 & ~n11210 ;
  assign n11212 = ~n2392 & ~n11211 ;
  assign n11217 = ~n11203 & ~n11212 ;
  assign n11218 = n11216 & n11217 ;
  assign n11219 = ~n11206 & n11218 ;
  assign n11220 = n2037 & ~n11219 ;
  assign n11221 = ~n11196 & ~n11220 ;
  assign n11222 = \P1_state_reg[0]/NET0131  & ~n11221 ;
  assign n11223 = ~n11195 & ~n11222 ;
  assign n11224 = \P1_reg0_reg[1]/NET0131  & ~n4085 ;
  assign n11225 = \P1_reg0_reg[1]/NET0131  & n4081 ;
  assign n11233 = n4869 & ~n10880 ;
  assign n11226 = \P1_reg0_reg[1]/NET0131  & ~n4869 ;
  assign n11227 = n4869 & n10864 ;
  assign n11228 = ~n11226 & ~n11227 ;
  assign n11229 = n4025 & ~n11228 ;
  assign n11230 = ~n3395 & n4869 ;
  assign n11231 = ~n11226 & ~n11230 ;
  assign n11232 = n4028 & ~n11231 ;
  assign n11234 = ~n4869 & ~n10882 ;
  assign n11235 = n4214 & ~n11234 ;
  assign n11236 = \P1_reg0_reg[1]/NET0131  & ~n11235 ;
  assign n11237 = ~n11232 & ~n11236 ;
  assign n11238 = ~n11229 & n11237 ;
  assign n11239 = ~n11233 & n11238 ;
  assign n11240 = n2701 & ~n11239 ;
  assign n11241 = ~n11225 & ~n11240 ;
  assign n11242 = \P1_state_reg[0]/NET0131  & ~n11241 ;
  assign n11243 = ~n11224 & ~n11242 ;
  assign n11244 = \P1_reg1_reg[1]/NET0131  & ~n4085 ;
  assign n11245 = \P1_reg1_reg[1]/NET0131  & n4081 ;
  assign n11249 = \P1_reg1_reg[1]/NET0131  & ~n4202 ;
  assign n11253 = n4202 & n10864 ;
  assign n11254 = ~n11249 & ~n11253 ;
  assign n11255 = n4025 & ~n11254 ;
  assign n11250 = n4202 & n10874 ;
  assign n11251 = ~n11249 & ~n11250 ;
  assign n11252 = n3969 & ~n11251 ;
  assign n11256 = n4202 & n10870 ;
  assign n11257 = ~n11249 & ~n11256 ;
  assign n11258 = n3829 & ~n11257 ;
  assign n11246 = ~n3395 & n4028 ;
  assign n11247 = ~n10878 & ~n11246 ;
  assign n11248 = n4202 & ~n11247 ;
  assign n11259 = \P1_reg1_reg[1]/NET0131  & ~n4218 ;
  assign n11260 = ~n11248 & ~n11259 ;
  assign n11261 = ~n11258 & n11260 ;
  assign n11262 = ~n11252 & n11261 ;
  assign n11263 = ~n11255 & n11262 ;
  assign n11264 = n2701 & ~n11263 ;
  assign n11265 = ~n11245 & ~n11264 ;
  assign n11266 = \P1_state_reg[0]/NET0131  & ~n11265 ;
  assign n11267 = ~n11244 & ~n11266 ;
  assign n11268 = \P2_reg3_reg[0]/NET0131  & ~n2286 ;
  assign n11269 = \P2_reg3_reg[0]/NET0131  & n2035 ;
  assign n11271 = \P2_reg3_reg[0]/NET0131  & ~n2124 ;
  assign n11280 = n1134 & ~n2231 ;
  assign n11281 = ~n2232 & n2263 ;
  assign n11282 = ~n11280 & n11281 ;
  assign n11283 = n2124 & n11282 ;
  assign n11284 = ~n11271 & ~n11283 ;
  assign n11285 = n1790 & ~n11284 ;
  assign n11272 = ~n1908 & n2124 ;
  assign n11273 = ~n11271 & ~n11272 ;
  assign n11274 = n2123 & ~n11273 ;
  assign n11270 = \P2_reg3_reg[0]/NET0131  & n2271 ;
  assign n11275 = ~n1165 & n1854 ;
  assign n11289 = ~n11270 & ~n11275 ;
  assign n11290 = ~n11274 & n11289 ;
  assign n11276 = \P2_reg3_reg[0]/NET0131  & ~n2053 ;
  assign n11277 = ~n1165 & n2053 ;
  assign n11278 = ~n11276 & ~n11277 ;
  assign n11279 = n2272 & ~n11278 ;
  assign n11286 = ~n1908 & n2053 ;
  assign n11287 = ~n11276 & ~n11286 ;
  assign n11288 = ~n10423 & ~n11287 ;
  assign n11291 = ~n11279 & ~n11288 ;
  assign n11292 = n11290 & n11291 ;
  assign n11293 = ~n11285 & n11292 ;
  assign n11294 = n2037 & ~n11293 ;
  assign n11295 = ~n11269 & ~n11294 ;
  assign n11296 = \P1_state_reg[0]/NET0131  & ~n11295 ;
  assign n11297 = ~n11268 & ~n11296 ;
  assign n11298 = \P1_reg2_reg[1]/NET0131  & ~n4085 ;
  assign n11299 = \P1_reg2_reg[1]/NET0131  & n4081 ;
  assign n11301 = \P1_reg2_reg[1]/NET0131  & ~n2717 ;
  assign n11305 = n2717 & n10864 ;
  assign n11306 = ~n11301 & ~n11305 ;
  assign n11307 = n4025 & ~n11306 ;
  assign n11302 = n2717 & n10874 ;
  assign n11303 = ~n11301 & ~n11302 ;
  assign n11304 = n3969 & ~n11303 ;
  assign n11308 = n2717 & n10870 ;
  assign n11309 = ~n11301 & ~n11308 ;
  assign n11310 = n3829 & ~n11309 ;
  assign n11311 = n2717 & ~n11247 ;
  assign n11300 = \P1_reg2_reg[1]/NET0131  & ~n4071 ;
  assign n11312 = \P1_reg3_reg[1]/NET0131  & n4073 ;
  assign n11313 = ~n11300 & ~n11312 ;
  assign n11314 = ~n11311 & n11313 ;
  assign n11315 = ~n11310 & n11314 ;
  assign n11316 = ~n11304 & n11315 ;
  assign n11317 = ~n11307 & n11316 ;
  assign n11318 = n2701 & ~n11317 ;
  assign n11319 = ~n11299 & ~n11318 ;
  assign n11320 = \P1_state_reg[0]/NET0131  & ~n11319 ;
  assign n11321 = ~n11298 & ~n11320 ;
  assign n11322 = \P2_reg1_reg[0]/NET0131  & ~n2286 ;
  assign n11323 = \P2_reg1_reg[0]/NET0131  & n2035 ;
  assign n11329 = n2291 & ~n11282 ;
  assign n11328 = ~\P2_reg1_reg[0]/NET0131  & ~n2291 ;
  assign n11330 = n1790 & ~n11328 ;
  assign n11331 = ~n11329 & n11330 ;
  assign n11324 = \P2_reg1_reg[0]/NET0131  & ~n2310 ;
  assign n11325 = ~n1908 & n2310 ;
  assign n11326 = ~n11324 & ~n11325 ;
  assign n11327 = ~n11016 & ~n11326 ;
  assign n11332 = \P2_reg1_reg[0]/NET0131  & ~n2612 ;
  assign n11339 = ~n11327 & ~n11332 ;
  assign n11333 = ~n1165 & n2310 ;
  assign n11334 = ~n11324 & ~n11333 ;
  assign n11335 = n2272 & ~n11334 ;
  assign n11336 = n1908 & n2291 ;
  assign n11337 = n2314 & ~n11328 ;
  assign n11338 = ~n11336 & n11337 ;
  assign n11340 = ~n11335 & ~n11338 ;
  assign n11341 = n11339 & n11340 ;
  assign n11342 = ~n11331 & n11341 ;
  assign n11343 = n2037 & ~n11342 ;
  assign n11344 = ~n11323 & ~n11343 ;
  assign n11345 = \P1_state_reg[0]/NET0131  & ~n11344 ;
  assign n11346 = ~n11322 & ~n11345 ;
  assign n11347 = \P2_reg2_reg[0]/NET0131  & ~n2286 ;
  assign n11348 = \P2_reg2_reg[0]/NET0131  & n2035 ;
  assign n11357 = \P2_reg2_reg[0]/NET0131  & ~n2310 ;
  assign n11358 = n2310 & n11282 ;
  assign n11359 = ~n11357 & ~n11358 ;
  assign n11360 = n1790 & ~n11359 ;
  assign n11351 = ~\P2_reg2_reg[0]/NET0131  & ~n2291 ;
  assign n11352 = n1165 & n2291 ;
  assign n11353 = n2272 & ~n11352 ;
  assign n11354 = ~n11016 & ~n11336 ;
  assign n11355 = ~n11353 & ~n11354 ;
  assign n11356 = ~n11351 & ~n11355 ;
  assign n11361 = ~n11325 & ~n11357 ;
  assign n11362 = n2314 & ~n11361 ;
  assign n11349 = \P2_reg3_reg[0]/NET0131  & n1854 ;
  assign n11350 = \P2_reg2_reg[0]/NET0131  & n2271 ;
  assign n11363 = ~n11349 & ~n11350 ;
  assign n11364 = ~n11362 & n11363 ;
  assign n11365 = ~n11356 & n11364 ;
  assign n11366 = ~n11360 & n11365 ;
  assign n11367 = n2037 & ~n11366 ;
  assign n11368 = ~n11348 & ~n11367 ;
  assign n11369 = \P1_state_reg[0]/NET0131  & ~n11368 ;
  assign n11370 = ~n11347 & ~n11369 ;
  assign n11371 = \P2_reg0_reg[0]/NET0131  & ~n2286 ;
  assign n11372 = \P2_reg0_reg[0]/NET0131  & n2035 ;
  assign n11378 = \P2_reg0_reg[0]/NET0131  & ~n2053 ;
  assign n11381 = n2053 & n11282 ;
  assign n11382 = ~n11378 & ~n11381 ;
  assign n11383 = n1790 & ~n11382 ;
  assign n11373 = \P2_reg0_reg[0]/NET0131  & ~n2124 ;
  assign n11374 = ~n1165 & n2124 ;
  assign n11375 = ~n11373 & ~n11374 ;
  assign n11376 = n2272 & ~n11375 ;
  assign n11377 = \P2_reg0_reg[0]/NET0131  & ~n2612 ;
  assign n11386 = ~n11376 & ~n11377 ;
  assign n11379 = ~n11286 & ~n11378 ;
  assign n11380 = n2123 & ~n11379 ;
  assign n11384 = ~n11272 & ~n11373 ;
  assign n11385 = ~n10423 & ~n11384 ;
  assign n11387 = ~n11380 & ~n11385 ;
  assign n11388 = n11386 & n11387 ;
  assign n11389 = ~n11383 & n11388 ;
  assign n11390 = n2037 & ~n11389 ;
  assign n11391 = ~n11372 & ~n11390 ;
  assign n11392 = \P1_state_reg[0]/NET0131  & ~n11391 ;
  assign n11393 = ~n11371 & ~n11392 ;
  assign n11394 = n3816 & ~n5415 ;
  assign n11395 = n3381 & ~n3985 ;
  assign n11396 = ~n2731 & n4025 ;
  assign n11397 = ~n3986 & n11396 ;
  assign n11398 = ~n11395 & n11397 ;
  assign n11399 = ~n11394 & ~n11398 ;
  assign n11400 = n4449 & ~n11399 ;
  assign n11401 = ~n4068 & ~n4449 ;
  assign n11402 = ~n3411 & n3815 ;
  assign n11403 = ~n11401 & n11402 ;
  assign n11404 = ~n11400 & ~n11403 ;
  assign n11405 = n9331 & ~n11404 ;
  assign n11406 = ~n8240 & n9331 ;
  assign n11407 = n5991 & n11406 ;
  assign n11408 = \P1_reg3_reg[0]/NET0131  & ~n11407 ;
  assign n11409 = ~n11405 & ~n11408 ;
  assign n11410 = \P1_reg3_reg[0]/NET0131  & n4073 ;
  assign n11411 = ~n3411 & n4069 ;
  assign n11412 = n11399 & ~n11411 ;
  assign n11413 = n2717 & ~n11412 ;
  assign n11414 = ~n11410 & ~n11413 ;
  assign n11415 = n9331 & ~n11414 ;
  assign n11416 = n9331 & n9342 ;
  assign n11417 = \P1_reg2_reg[0]/NET0131  & ~n11416 ;
  assign n11418 = ~n11415 & ~n11417 ;
  assign n11419 = n9331 & ~n11412 ;
  assign n11420 = n4869 & n11419 ;
  assign n11421 = ~n7303 & n9331 ;
  assign n11422 = n5844 & n11421 ;
  assign n11423 = \P1_reg0_reg[0]/NET0131  & ~n11422 ;
  assign n11424 = ~n11420 & ~n11423 ;
  assign n11425 = n4202 & n11419 ;
  assign n11426 = ~n6942 & n9331 ;
  assign n11427 = n6494 & n11426 ;
  assign n11428 = \P1_reg1_reg[0]/NET0131  & ~n11427 ;
  assign n11429 = ~n11425 & ~n11428 ;
  assign n11430 = ~n1744 & n2124 ;
  assign n11431 = n2272 & ~n11430 ;
  assign n11434 = ~n1790 & ~n2123 ;
  assign n11435 = ~n2053 & ~n11434 ;
  assign n11432 = ~n2124 & ~n10423 ;
  assign n11433 = ~n2034 & n2286 ;
  assign n11436 = ~n1854 & n11433 ;
  assign n11437 = ~n11432 & n11436 ;
  assign n11438 = ~n11435 & n11437 ;
  assign n11439 = ~n11431 & n11438 ;
  assign n11440 = \P2_reg0_reg[30]/NET0131  & ~n11439 ;
  assign n11441 = ~n1701 & n1790 ;
  assign n11442 = n2606 & n11441 ;
  assign n11443 = n2053 & n11442 ;
  assign n11444 = n2124 & n11431 ;
  assign n11445 = ~n11443 & ~n11444 ;
  assign n11446 = n11433 & ~n11445 ;
  assign n11447 = ~n11440 & ~n11446 ;
  assign n11448 = ~n1723 & n2124 ;
  assign n11449 = n2272 & ~n11448 ;
  assign n11450 = n11438 & ~n11449 ;
  assign n11451 = \P2_reg0_reg[31]/NET0131  & ~n11450 ;
  assign n11452 = n2124 & n11449 ;
  assign n11453 = ~n11443 & ~n11452 ;
  assign n11454 = n11433 & ~n11453 ;
  assign n11455 = ~n11451 & ~n11454 ;
  assign n11456 = n1744 & n4101 ;
  assign n11457 = n2291 & n11442 ;
  assign n11458 = ~n11456 & ~n11457 ;
  assign n11459 = n11433 & ~n11458 ;
  assign n11460 = ~n1790 & ~n2314 ;
  assign n11461 = ~n2291 & ~n11460 ;
  assign n11462 = n11433 & ~n11461 ;
  assign n11463 = n11018 & n11462 ;
  assign n11464 = \P2_reg1_reg[30]/NET0131  & ~n11463 ;
  assign n11465 = ~n11459 & ~n11464 ;
  assign n11471 = n2310 & n11442 ;
  assign n11472 = ~n4191 & ~n11471 ;
  assign n11473 = n11433 & ~n11472 ;
  assign n11467 = ~n2291 & ~n11016 ;
  assign n11466 = ~n2310 & ~n11460 ;
  assign n11468 = n11433 & ~n11466 ;
  assign n11469 = ~n11467 & n11468 ;
  assign n11470 = \P2_reg2_reg[30]/NET0131  & ~n11469 ;
  assign n11474 = \P2_reg2_reg[30]/NET0131  & ~n2291 ;
  assign n11475 = n2291 & n11433 ;
  assign n11476 = n1744 & n11475 ;
  assign n11477 = ~n11474 & ~n11476 ;
  assign n11478 = n2272 & ~n11477 ;
  assign n11479 = ~n11470 & ~n11478 ;
  assign n11480 = ~n11473 & n11479 ;
  assign n11481 = n1723 & n4101 ;
  assign n11482 = ~n11457 & ~n11481 ;
  assign n11483 = n11433 & ~n11482 ;
  assign n11484 = \P2_reg1_reg[31]/NET0131  & ~n11463 ;
  assign n11485 = ~n11483 & ~n11484 ;
  assign n11486 = \P2_reg2_reg[31]/NET0131  & ~n11469 ;
  assign n11487 = \P2_reg2_reg[31]/NET0131  & ~n2291 ;
  assign n11488 = n1723 & n11475 ;
  assign n11489 = ~n11487 & ~n11488 ;
  assign n11490 = n2272 & ~n11489 ;
  assign n11491 = ~n11486 & ~n11490 ;
  assign n11492 = ~n11473 & n11491 ;
  assign n11493 = ~\P1_state_reg[0]/NET0131  & ~n3068 ;
  assign n11494 = \P1_state_reg[0]/NET0131  & n2725 ;
  assign n11495 = ~n11493 & ~n11494 ;
  assign n11496 = \P1_state_reg[0]/NET0131  & ~n2024 ;
  assign n11497 = ~\P1_state_reg[0]/NET0131  & n1512 ;
  assign n11498 = ~n11496 & ~n11497 ;
  assign n11499 = \P1_state_reg[0]/NET0131  & ~n2032 ;
  assign n11500 = ~\P1_state_reg[0]/NET0131  & n1572 ;
  assign n11501 = ~n11499 & ~n11500 ;
  assign n11502 = ~\P1_state_reg[0]/NET0131  & ~n1607 ;
  assign n11503 = \P1_state_reg[0]/NET0131  & n633 ;
  assign n11504 = ~n11502 & ~n11503 ;
  assign n11505 = ~\P1_state_reg[0]/NET0131  & ~n2963 ;
  assign n11506 = \P1_state_reg[0]/NET0131  & ~n2686 ;
  assign n11507 = ~n11505 & ~n11506 ;
  assign n11508 = ~\P1_state_reg[0]/NET0131  & ~n3016 ;
  assign n11509 = \P1_state_reg[0]/NET0131  & n2689 ;
  assign n11510 = ~n11508 & ~n11509 ;
  assign n11511 = ~\P1_state_reg[0]/NET0131  & n1722 ;
  assign n11512 = \P1_state_reg[0]/NET0131  & ~\P2_IR_reg[27]/NET0131  ;
  assign n11513 = ~\P2_IR_reg[30]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n11514 = n11512 & n11513 ;
  assign n11515 = n568 & n11514 ;
  assign n11516 = n628 & n11515 ;
  assign n11517 = n624 & n11516 ;
  assign n11518 = ~n11511 & ~n11517 ;
  assign n11519 = ~\P1_state_reg[0]/NET0131  & ~n1248 ;
  assign n11520 = \P1_state_reg[0]/NET0131  & n1253 ;
  assign n11521 = ~n11519 & ~n11520 ;
  assign n11522 = ~\P1_state_reg[0]/NET0131  & n1433 ;
  assign n11523 = ~n2286 & ~n11522 ;
  assign n11524 = ~\P1_state_reg[0]/NET0131  & ~n900 ;
  assign n11525 = \P1_state_reg[0]/NET0131  & n907 ;
  assign n11526 = ~n11524 & ~n11525 ;
  assign n11527 = ~\P1_state_reg[0]/NET0131  & ~n875 ;
  assign n11528 = \P1_state_reg[0]/NET0131  & n880 ;
  assign n11529 = ~n11527 & ~n11528 ;
  assign n11530 = ~\P1_state_reg[0]/NET0131  & ~n841 ;
  assign n11531 = \P1_state_reg[0]/NET0131  & n848 ;
  assign n11532 = ~n11530 & ~n11531 ;
  assign n11533 = ~\P1_state_reg[0]/NET0131  & ~n805 ;
  assign n11534 = \P1_state_reg[0]/NET0131  & n809 ;
  assign n11535 = ~n11533 & ~n11534 ;
  assign n11536 = ~\P1_state_reg[0]/NET0131  & ~n754 ;
  assign n11537 = \P1_state_reg[0]/NET0131  & n758 ;
  assign n11538 = ~n11536 & ~n11537 ;
  assign n11539 = ~\P1_state_reg[0]/NET0131  & ~n711 ;
  assign n11540 = \P1_state_reg[0]/NET0131  & n716 ;
  assign n11541 = ~n11539 & ~n11540 ;
  assign n11542 = ~\P1_state_reg[0]/NET0131  & ~n1213 ;
  assign n11543 = \P1_state_reg[0]/NET0131  & n1219 ;
  assign n11544 = ~n11542 & ~n11543 ;
  assign n11545 = ~\P1_state_reg[0]/NET0131  & ~n1326 ;
  assign n11546 = \P1_state_reg[0]/NET0131  & n1332 ;
  assign n11547 = ~n11545 & ~n11546 ;
  assign n11548 = ~\P1_state_reg[0]/NET0131  & ~n1293 ;
  assign n11549 = \P1_state_reg[0]/NET0131  & ~n1297 ;
  assign n11550 = ~n11548 & ~n11549 ;
  assign n11551 = \P1_state_reg[0]/NET0131  & ~n1138 ;
  assign n11552 = ~\P1_state_reg[0]/NET0131  & n1146 ;
  assign n11553 = ~n11551 & ~n11552 ;
  assign n11554 = \P1_state_reg[0]/NET0131  & ~n1777 ;
  assign n11555 = ~\P1_state_reg[0]/NET0131  & n1400 ;
  assign n11556 = ~n11554 & ~n11555 ;
  assign n11557 = \P1_state_reg[0]/NET0131  & ~n1771 ;
  assign n11558 = ~\P1_state_reg[0]/NET0131  & n1370 ;
  assign n11559 = ~n11557 & ~n11558 ;
  assign n11560 = ~\P1_state_reg[0]/NET0131  & ~n1464 ;
  assign n11561 = \P1_state_reg[0]/NET0131  & n1783 ;
  assign n11562 = ~n11560 & ~n11561 ;
  assign n11563 = ~\P1_state_reg[0]/NET0131  & ~n1539 ;
  assign n11564 = \P1_state_reg[0]/NET0131  & n2027 ;
  assign n11565 = ~n11563 & ~n11564 ;
  assign n11566 = ~\P1_state_reg[0]/NET0131  & ~n1683 ;
  assign n11567 = \P1_state_reg[0]/NET0131  & n615 ;
  assign n11568 = ~n11566 & ~n11567 ;
  assign n11569 = ~\P1_state_reg[0]/NET0131  & ~n1655 ;
  assign n11570 = \P1_state_reg[0]/NET0131  & n556 ;
  assign n11571 = ~n11569 & ~n11570 ;
  assign n11572 = ~\P1_state_reg[0]/NET0131  & ~n1117 ;
  assign n11573 = \P1_state_reg[0]/NET0131  & ~n1122 ;
  assign n11574 = ~n11572 & ~n11573 ;
  assign n11575 = ~\P1_state_reg[0]/NET0131  & ~n1743 ;
  assign n11576 = \P1_state_reg[0]/NET0131  & n576 ;
  assign n11577 = ~n11575 & ~n11576 ;
  assign n11578 = \P1_state_reg[0]/NET0131  & n1090 ;
  assign n11579 = ~\P1_state_reg[0]/NET0131  & n1098 ;
  assign n11580 = ~n11578 & ~n11579 ;
  assign n11581 = ~\P1_state_reg[0]/NET0131  & ~n1069 ;
  assign n11582 = \P1_state_reg[0]/NET0131  & n1074 ;
  assign n11583 = ~n11581 & ~n11582 ;
  assign n11584 = ~\P1_state_reg[0]/NET0131  & ~n1044 ;
  assign n11585 = \P1_state_reg[0]/NET0131  & ~n1048 ;
  assign n11586 = ~n11584 & ~n11585 ;
  assign n11587 = ~\P1_state_reg[0]/NET0131  & ~n993 ;
  assign n11588 = \P1_state_reg[0]/NET0131  & n1001 ;
  assign n11589 = ~n11587 & ~n11588 ;
  assign n11590 = ~\P1_state_reg[0]/NET0131  & ~n1020 ;
  assign n11591 = \P1_state_reg[0]/NET0131  & n1024 ;
  assign n11592 = ~n11590 & ~n11591 ;
  assign n11593 = ~\P1_state_reg[0]/NET0131  & ~n951 ;
  assign n11594 = \P1_state_reg[0]/NET0131  & n956 ;
  assign n11595 = ~n11593 & ~n11594 ;
  assign n11596 = ~\P1_state_reg[0]/NET0131  & ~n928 ;
  assign n11597 = \P1_state_reg[0]/NET0131  & ~n932 ;
  assign n11598 = ~n11596 & ~n11597 ;
  assign n11599 = ~\P1_state_reg[0]/NET0131  & ~n3261 ;
  assign n11600 = \P1_state_reg[0]/NET0131  & ~n3253 ;
  assign n11601 = ~n11599 & ~n11600 ;
  assign n11602 = ~\P1_state_reg[0]/NET0131  & ~n3209 ;
  assign n11603 = \P1_state_reg[0]/NET0131  & ~n3201 ;
  assign n11604 = ~n11602 & ~n11603 ;
  assign n11605 = \P1_state_reg[0]/NET0131  & ~n3228 ;
  assign n11606 = ~\P1_state_reg[0]/NET0131  & n3237 ;
  assign n11607 = ~n11605 & ~n11606 ;
  assign n11608 = \P1_state_reg[0]/NET0131  & ~n3673 ;
  assign n11609 = ~\P1_state_reg[0]/NET0131  & n3681 ;
  assign n11610 = ~n11608 & ~n11609 ;
  assign n11611 = ~\P1_state_reg[0]/NET0131  & ~n3654 ;
  assign n11612 = \P1_state_reg[0]/NET0131  & n3646 ;
  assign n11613 = ~n11611 & ~n11612 ;
  assign n11614 = ~\P1_state_reg[0]/NET0131  & ~n3730 ;
  assign n11615 = \P1_state_reg[0]/NET0131  & n3722 ;
  assign n11616 = ~n11614 & ~n11615 ;
  assign n11617 = ~\P1_state_reg[0]/NET0131  & ~n3706 ;
  assign n11618 = \P1_state_reg[0]/NET0131  & n3698 ;
  assign n11619 = ~n11617 & ~n11618 ;
  assign n11620 = \P1_state_reg[0]/NET0131  & n3593 ;
  assign n11621 = ~\P1_state_reg[0]/NET0131  & n3601 ;
  assign n11622 = ~n11620 & ~n11621 ;
  assign n11623 = \P1_state_reg[0]/NET0131  & ~n3621 ;
  assign n11624 = ~\P1_state_reg[0]/NET0131  & n3629 ;
  assign n11625 = ~n11623 & ~n11624 ;
  assign n11626 = ~\P1_state_reg[0]/NET0131  & ~n3576 ;
  assign n11627 = \P1_state_reg[0]/NET0131  & ~n3566 ;
  assign n11628 = ~n11626 & ~n11627 ;
  assign n11629 = \P1_state_reg[0]/NET0131  & n3385 ;
  assign n11630 = ~\P1_state_reg[0]/NET0131  & n3393 ;
  assign n11631 = ~n11629 & ~n11630 ;
  assign n11632 = ~\P1_state_reg[0]/NET0131  & ~n3547 ;
  assign n11633 = \P1_state_reg[0]/NET0131  & ~n3826 ;
  assign n11634 = ~n11632 & ~n11633 ;
  assign n11635 = \P1_state_reg[0]/NET0131  & ~n3821 ;
  assign n11636 = ~\P1_state_reg[0]/NET0131  & n3167 ;
  assign n11637 = ~n11635 & ~n11636 ;
  assign n11638 = ~\P1_state_reg[0]/NET0131  & ~n3142 ;
  assign n11639 = \P1_state_reg[0]/NET0131  & n3813 ;
  assign n11640 = ~n11638 & ~n11639 ;
  assign n11641 = ~\P1_state_reg[0]/NET0131  & ~n3118 ;
  assign n11642 = ~n4552 & ~n11641 ;
  assign n11643 = ~\P1_state_reg[0]/NET0131  & ~n3095 ;
  assign n11644 = \P1_state_reg[0]/NET0131  & n2698 ;
  assign n11645 = ~n11643 & ~n11644 ;
  assign n11646 = ~\P1_state_reg[0]/NET0131  & ~n2867 ;
  assign n11647 = \P1_state_reg[0]/NET0131  & n2731 ;
  assign n11648 = ~n11646 & ~n11647 ;
  assign n11649 = ~\P1_state_reg[0]/NET0131  & ~n3793 ;
  assign n11650 = \P1_state_reg[0]/NET0131  & n494 ;
  assign n11651 = ~n11649 & ~n11650 ;
  assign n11652 = ~\P1_state_reg[0]/NET0131  & ~n3347 ;
  assign n11653 = \P1_state_reg[0]/NET0131  & n3352 ;
  assign n11654 = ~n11652 & ~n11653 ;
  assign n11655 = ~\P1_state_reg[0]/NET0131  & ~n5370 ;
  assign n11656 = \P1_state_reg[0]/NET0131  & n512 ;
  assign n11657 = ~n11655 & ~n11656 ;
  assign n11658 = ~\P1_state_reg[0]/NET0131  & n5351 ;
  assign n11659 = ~\P1_IR_reg[30]/NET0131  & \P1_IR_reg[31]/NET0131  ;
  assign n11660 = \P1_state_reg[0]/NET0131  & n11659 ;
  assign n11661 = n506 & n11660 ;
  assign n11662 = n2720 & n11661 ;
  assign n11663 = n2679 & n11662 ;
  assign n11664 = ~n11658 & ~n11663 ;
  assign n11665 = ~\P1_state_reg[0]/NET0131  & ~n3363 ;
  assign n11666 = \P1_state_reg[0]/NET0131  & n3369 ;
  assign n11667 = ~n11665 & ~n11666 ;
  assign n11668 = ~\P1_state_reg[0]/NET0131  & ~n3325 ;
  assign n11669 = \P1_state_reg[0]/NET0131  & ~n3330 ;
  assign n11670 = ~n11668 & ~n11669 ;
  assign n11671 = ~\P1_state_reg[0]/NET0131  & ~n3503 ;
  assign n11672 = \P1_state_reg[0]/NET0131  & n3509 ;
  assign n11673 = ~n11671 & ~n11672 ;
  assign n11674 = \P1_state_reg[0]/NET0131  & ~n3451 ;
  assign n11675 = ~\P1_state_reg[0]/NET0131  & n3459 ;
  assign n11676 = ~n11674 & ~n11675 ;
  assign n11677 = ~\P1_state_reg[0]/NET0131  & ~n3479 ;
  assign n11678 = \P1_state_reg[0]/NET0131  & n3483 ;
  assign n11679 = ~n11677 & ~n11678 ;
  assign n11680 = \P1_state_reg[0]/NET0131  & ~n3425 ;
  assign n11681 = ~\P1_state_reg[0]/NET0131  & n3433 ;
  assign n11682 = ~n11680 & ~n11681 ;
  assign n11683 = ~\P1_state_reg[0]/NET0131  & ~n3289 ;
  assign n11684 = \P1_state_reg[0]/NET0131  & ~n3281 ;
  assign n11685 = ~n11683 & ~n11684 ;
  assign n11729 = \P1_reg1_reg[8]/NET0131  & n3425 ;
  assign n11730 = ~\P1_reg1_reg[8]/NET0131  & ~n3425 ;
  assign n11731 = ~n11729 & ~n11730 ;
  assign n11732 = \P1_reg1_reg[7]/NET0131  & n3451 ;
  assign n11733 = ~\P1_reg1_reg[7]/NET0131  & ~n3451 ;
  assign n11734 = \P1_reg1_reg[6]/NET0131  & n3483 ;
  assign n11735 = ~\P1_reg1_reg[6]/NET0131  & ~n3483 ;
  assign n11736 = \P1_reg1_reg[5]/NET0131  & n3509 ;
  assign n11737 = ~\P1_reg1_reg[5]/NET0131  & ~n3509 ;
  assign n11738 = \P1_reg1_reg[4]/NET0131  & ~n3330 ;
  assign n11739 = ~\P1_reg1_reg[4]/NET0131  & n3330 ;
  assign n11740 = ~\P1_reg1_reg[3]/NET0131  & ~n3369 ;
  assign n11741 = \P1_reg1_reg[3]/NET0131  & n3369 ;
  assign n11742 = ~\P1_reg1_reg[2]/NET0131  & ~n3352 ;
  assign n11743 = \P1_reg1_reg[2]/NET0131  & n3352 ;
  assign n11744 = ~\P1_reg1_reg[1]/NET0131  & ~n3385 ;
  assign n11745 = \P1_reg1_reg[1]/NET0131  & n3385 ;
  assign n11746 = \P1_IR_reg[0]/NET0131  & \P1_reg1_reg[0]/NET0131  ;
  assign n11747 = ~n11745 & ~n11746 ;
  assign n11748 = ~n11744 & ~n11747 ;
  assign n11749 = ~n11743 & ~n11748 ;
  assign n11750 = ~n11742 & ~n11749 ;
  assign n11751 = ~n11741 & ~n11750 ;
  assign n11752 = ~n11740 & ~n11751 ;
  assign n11753 = ~n11739 & n11752 ;
  assign n11754 = ~n11738 & ~n11753 ;
  assign n11755 = ~n11737 & ~n11754 ;
  assign n11756 = ~n11736 & ~n11755 ;
  assign n11757 = ~n11735 & ~n11756 ;
  assign n11758 = ~n11734 & ~n11757 ;
  assign n11759 = ~n11733 & ~n11758 ;
  assign n11760 = ~n11732 & ~n11759 ;
  assign n11762 = n11731 & ~n11760 ;
  assign n11728 = ~n2725 & n2731 ;
  assign n11761 = ~n11731 & n11760 ;
  assign n11763 = n11728 & ~n11761 ;
  assign n11764 = ~n11762 & n11763 ;
  assign n11687 = \P1_reg2_reg[8]/NET0131  & n3425 ;
  assign n11688 = ~\P1_reg2_reg[8]/NET0131  & ~n3425 ;
  assign n11689 = ~n11687 & ~n11688 ;
  assign n11690 = \P1_reg2_reg[7]/NET0131  & n3451 ;
  assign n11691 = ~\P1_reg2_reg[7]/NET0131  & ~n3451 ;
  assign n11692 = \P1_reg2_reg[6]/NET0131  & n3483 ;
  assign n11693 = ~\P1_reg2_reg[6]/NET0131  & ~n3483 ;
  assign n11694 = \P1_reg2_reg[5]/NET0131  & n3509 ;
  assign n11695 = ~\P1_reg2_reg[5]/NET0131  & ~n3509 ;
  assign n11696 = \P1_reg2_reg[4]/NET0131  & ~n3330 ;
  assign n11697 = ~\P1_reg2_reg[4]/NET0131  & n3330 ;
  assign n11698 = ~\P1_reg2_reg[3]/NET0131  & ~n3369 ;
  assign n11699 = \P1_reg2_reg[3]/NET0131  & n3369 ;
  assign n11700 = ~\P1_reg2_reg[2]/NET0131  & ~n3352 ;
  assign n11701 = \P1_reg2_reg[2]/NET0131  & n3352 ;
  assign n11702 = ~\P1_reg2_reg[1]/NET0131  & ~n3385 ;
  assign n11703 = \P1_reg2_reg[1]/NET0131  & n3385 ;
  assign n11704 = \P1_IR_reg[0]/NET0131  & \P1_reg2_reg[0]/NET0131  ;
  assign n11705 = ~n11703 & ~n11704 ;
  assign n11706 = ~n11702 & ~n11705 ;
  assign n11707 = ~n11701 & ~n11706 ;
  assign n11708 = ~n11700 & ~n11707 ;
  assign n11709 = ~n11699 & ~n11708 ;
  assign n11710 = ~n11698 & ~n11709 ;
  assign n11711 = ~n11697 & n11710 ;
  assign n11712 = ~n11696 & ~n11711 ;
  assign n11713 = ~n11695 & ~n11712 ;
  assign n11714 = ~n11694 & ~n11713 ;
  assign n11715 = ~n11693 & ~n11714 ;
  assign n11716 = ~n11692 & ~n11715 ;
  assign n11717 = ~n11691 & ~n11716 ;
  assign n11718 = ~n11690 & ~n11717 ;
  assign n11720 = n11689 & ~n11718 ;
  assign n11686 = n2725 & n2731 ;
  assign n11719 = ~n11689 & n11718 ;
  assign n11721 = n11686 & ~n11719 ;
  assign n11722 = ~n11720 & n11721 ;
  assign n11723 = ~n2725 & ~n4081 ;
  assign n11725 = ~n3425 & ~n11723 ;
  assign n11724 = ~\P1_addr_reg[8]/NET0131  & n11723 ;
  assign n11726 = ~n2731 & ~n11724 ;
  assign n11727 = ~n11725 & n11726 ;
  assign n11765 = ~n11722 & ~n11727 ;
  assign n11766 = ~n11764 & n11765 ;
  assign n11767 = \P1_state_reg[0]/NET0131  & ~n11766 ;
  assign n11768 = ~n8236 & ~n11767 ;
  assign n11769 = \P1_reg1_reg[12]/NET0131  & n3228 ;
  assign n11770 = ~\P1_reg1_reg[12]/NET0131  & ~n3228 ;
  assign n11771 = ~n11769 & ~n11770 ;
  assign n11772 = \P1_reg1_reg[11]/NET0131  & ~n3201 ;
  assign n11773 = \P1_reg1_reg[10]/NET0131  & ~n3253 ;
  assign n11774 = \P1_reg1_reg[9]/NET0131  & ~n3281 ;
  assign n11775 = ~n11730 & ~n11760 ;
  assign n11776 = ~n11729 & ~n11775 ;
  assign n11777 = ~n11774 & n11776 ;
  assign n11778 = ~\P1_reg1_reg[10]/NET0131  & n3253 ;
  assign n11779 = ~\P1_reg1_reg[9]/NET0131  & n3281 ;
  assign n11780 = ~n11778 & ~n11779 ;
  assign n11781 = ~n11777 & n11780 ;
  assign n11782 = ~n11773 & ~n11781 ;
  assign n11783 = ~n11772 & n11782 ;
  assign n11784 = ~\P1_reg1_reg[11]/NET0131  & n3201 ;
  assign n11785 = ~n11783 & ~n11784 ;
  assign n11787 = n11771 & n11785 ;
  assign n11786 = ~n11771 & ~n11785 ;
  assign n11788 = n11728 & ~n11786 ;
  assign n11789 = ~n11787 & n11788 ;
  assign n11791 = ~n3228 & ~n11723 ;
  assign n11790 = ~\P1_addr_reg[12]/NET0131  & n11723 ;
  assign n11792 = ~n2731 & ~n11790 ;
  assign n11793 = ~n11791 & n11792 ;
  assign n11794 = \P1_reg2_reg[12]/NET0131  & n3228 ;
  assign n11795 = ~\P1_reg2_reg[12]/NET0131  & ~n3228 ;
  assign n11796 = ~n11794 & ~n11795 ;
  assign n11797 = ~\P1_reg2_reg[11]/NET0131  & n3201 ;
  assign n11798 = ~\P1_reg2_reg[10]/NET0131  & n3253 ;
  assign n11799 = ~\P1_reg2_reg[9]/NET0131  & n3281 ;
  assign n11801 = ~n11688 & ~n11799 ;
  assign n11802 = ~n11718 & n11801 ;
  assign n11800 = n11687 & ~n11799 ;
  assign n11803 = \P1_reg2_reg[9]/NET0131  & ~n3281 ;
  assign n11804 = ~n11800 & ~n11803 ;
  assign n11805 = ~n11802 & n11804 ;
  assign n11806 = ~n11798 & ~n11805 ;
  assign n11807 = \P1_reg2_reg[11]/NET0131  & ~n3201 ;
  assign n11808 = \P1_reg2_reg[10]/NET0131  & ~n3253 ;
  assign n11809 = ~n11807 & ~n11808 ;
  assign n11810 = ~n11806 & n11809 ;
  assign n11811 = ~n11797 & ~n11810 ;
  assign n11813 = n11796 & n11811 ;
  assign n11812 = ~n11796 & ~n11811 ;
  assign n11814 = n11686 & ~n11812 ;
  assign n11815 = ~n11813 & n11814 ;
  assign n11816 = ~n11793 & ~n11815 ;
  assign n11817 = ~n11789 & n11816 ;
  assign n11818 = \P1_state_reg[0]/NET0131  & ~n11817 ;
  assign n11819 = ~n6580 & ~n11818 ;
  assign n11829 = ~n11799 & ~n11803 ;
  assign n11830 = ~n11687 & n11718 ;
  assign n11831 = ~n11688 & ~n11830 ;
  assign n11833 = n11829 & n11831 ;
  assign n11832 = ~n11829 & ~n11831 ;
  assign n11834 = n11686 & ~n11832 ;
  assign n11835 = ~n11833 & n11834 ;
  assign n11820 = ~n11774 & ~n11779 ;
  assign n11822 = ~n11776 & n11820 ;
  assign n11821 = n11776 & ~n11820 ;
  assign n11823 = n11728 & ~n11821 ;
  assign n11824 = ~n11822 & n11823 ;
  assign n11826 = n3281 & ~n11723 ;
  assign n11825 = ~\P1_addr_reg[9]/NET0131  & n11723 ;
  assign n11827 = ~n2731 & ~n11825 ;
  assign n11828 = ~n11826 & n11827 ;
  assign n11836 = ~n11824 & ~n11828 ;
  assign n11837 = ~n11835 & n11836 ;
  assign n11838 = \P1_state_reg[0]/NET0131  & ~n11837 ;
  assign n11839 = ~n7608 & ~n11838 ;
  assign n11849 = ~n11732 & ~n11733 ;
  assign n11851 = ~n11758 & n11849 ;
  assign n11850 = n11758 & ~n11849 ;
  assign n11852 = n11728 & ~n11850 ;
  assign n11853 = ~n11851 & n11852 ;
  assign n11841 = ~n3451 & ~n11723 ;
  assign n11840 = ~\P1_addr_reg[7]/NET0131  & n11723 ;
  assign n11842 = ~n2731 & ~n11840 ;
  assign n11843 = ~n11841 & n11842 ;
  assign n11844 = ~n11690 & ~n11691 ;
  assign n11846 = ~n11716 & n11844 ;
  assign n11845 = n11716 & ~n11844 ;
  assign n11847 = n11686 & ~n11845 ;
  assign n11848 = ~n11846 & n11847 ;
  assign n11854 = ~n11843 & ~n11848 ;
  assign n11855 = ~n11853 & n11854 ;
  assign n11856 = \P1_state_reg[0]/NET0131  & ~n11855 ;
  assign n11857 = ~n9810 & ~n11856 ;
  assign n11875 = \P1_reg1_reg[14]/NET0131  & n3646 ;
  assign n11876 = ~\P1_reg1_reg[14]/NET0131  & ~n3646 ;
  assign n11877 = ~n11875 & ~n11876 ;
  assign n11878 = \P1_reg1_reg[13]/NET0131  & n3673 ;
  assign n11879 = ~\P1_reg1_reg[13]/NET0131  & ~n3673 ;
  assign n11880 = ~n11770 & ~n11784 ;
  assign n11881 = ~n11783 & n11880 ;
  assign n11882 = ~n11769 & ~n11881 ;
  assign n11883 = ~n11879 & ~n11882 ;
  assign n11884 = ~n11878 & ~n11883 ;
  assign n11886 = n11877 & ~n11884 ;
  assign n11885 = ~n11877 & n11884 ;
  assign n11887 = n11728 & ~n11885 ;
  assign n11888 = ~n11886 & n11887 ;
  assign n11859 = ~n3646 & ~n11723 ;
  assign n11858 = ~\P1_addr_reg[14]/NET0131  & n11723 ;
  assign n11860 = ~n2731 & ~n11858 ;
  assign n11861 = ~n11859 & n11860 ;
  assign n11862 = \P1_reg2_reg[14]/NET0131  & n3646 ;
  assign n11863 = ~\P1_reg2_reg[14]/NET0131  & ~n3646 ;
  assign n11864 = ~n11862 & ~n11863 ;
  assign n11865 = ~\P1_reg2_reg[13]/NET0131  & ~n3673 ;
  assign n11867 = ~n11795 & n11811 ;
  assign n11866 = \P1_reg2_reg[13]/NET0131  & n3673 ;
  assign n11868 = ~n11794 & ~n11866 ;
  assign n11869 = ~n11867 & n11868 ;
  assign n11870 = ~n11865 & ~n11869 ;
  assign n11872 = n11864 & n11870 ;
  assign n11871 = ~n11864 & ~n11870 ;
  assign n11873 = n11686 & ~n11871 ;
  assign n11874 = ~n11872 & n11873 ;
  assign n11889 = ~n11861 & ~n11874 ;
  assign n11890 = ~n11888 & n11889 ;
  assign n11891 = \P1_state_reg[0]/NET0131  & ~n11890 ;
  assign n11892 = ~n8074 & ~n11891 ;
  assign n11894 = ~\P2_reg1_reg[9]/NET0131  & ~n932 ;
  assign n11895 = \P2_reg1_reg[9]/NET0131  & n932 ;
  assign n11896 = ~n11894 & ~n11895 ;
  assign n11928 = \P2_reg1_reg[8]/NET0131  & ~n956 ;
  assign n11897 = ~\P2_reg1_reg[8]/NET0131  & n956 ;
  assign n11899 = \P2_reg1_reg[7]/NET0131  & ~n1024 ;
  assign n11898 = ~\P2_reg1_reg[7]/NET0131  & n1024 ;
  assign n11901 = \P2_reg1_reg[6]/NET0131  & ~n1001 ;
  assign n11900 = ~\P2_reg1_reg[6]/NET0131  & n1001 ;
  assign n11902 = ~\P2_reg1_reg[5]/NET0131  & ~n1048 ;
  assign n11918 = \P2_reg1_reg[5]/NET0131  & n1048 ;
  assign n11919 = \P2_reg1_reg[4]/NET0131  & ~n1074 ;
  assign n11903 = ~\P2_reg1_reg[4]/NET0131  & n1074 ;
  assign n11905 = \P2_reg1_reg[3]/NET0131  & ~n1090 ;
  assign n11904 = ~\P2_reg1_reg[3]/NET0131  & n1090 ;
  assign n11907 = \P2_reg1_reg[2]/NET0131  & n1122 ;
  assign n11906 = ~\P2_reg1_reg[2]/NET0131  & ~n1122 ;
  assign n11909 = \P2_reg1_reg[1]/NET0131  & n1138 ;
  assign n11908 = ~\P2_reg1_reg[1]/NET0131  & ~n1138 ;
  assign n12002 = \P2_IR_reg[0]/NET0131  & ~\P2_reg1_reg[0]/NET0131  ;
  assign n12003 = ~n11908 & ~n12002 ;
  assign n12004 = ~n11909 & ~n12003 ;
  assign n12005 = ~n11906 & ~n12004 ;
  assign n12006 = ~n11907 & ~n12005 ;
  assign n12007 = ~n11904 & ~n12006 ;
  assign n12008 = ~n11905 & ~n12007 ;
  assign n12009 = ~n11903 & ~n12008 ;
  assign n12010 = ~n11919 & ~n12009 ;
  assign n12011 = ~n11918 & n12010 ;
  assign n12012 = ~n11902 & ~n12011 ;
  assign n12013 = ~n11900 & n12012 ;
  assign n12014 = ~n11901 & ~n12013 ;
  assign n12015 = ~n11898 & ~n12014 ;
  assign n12016 = ~n11899 & ~n12015 ;
  assign n12017 = ~n11897 & ~n12016 ;
  assign n12018 = ~n11928 & ~n12017 ;
  assign n12020 = ~n11896 & n12018 ;
  assign n12019 = n11896 & ~n12018 ;
  assign n12021 = n634 & ~n12019 ;
  assign n12022 = ~n12020 & n12021 ;
  assign n11934 = \P2_reg2_reg[9]/NET0131  & n932 ;
  assign n11935 = ~\P2_reg2_reg[9]/NET0131  & ~n932 ;
  assign n11936 = ~n11934 & ~n11935 ;
  assign n11937 = \P2_reg2_reg[8]/NET0131  & ~n956 ;
  assign n11965 = ~\P2_reg2_reg[8]/NET0131  & n956 ;
  assign n11938 = \P2_reg2_reg[7]/NET0131  & ~n1024 ;
  assign n11966 = ~\P2_reg2_reg[7]/NET0131  & n1024 ;
  assign n11939 = \P2_reg2_reg[6]/NET0131  & ~n1001 ;
  assign n11959 = ~\P2_reg2_reg[6]/NET0131  & n1001 ;
  assign n11940 = \P2_reg2_reg[5]/NET0131  & n1048 ;
  assign n11960 = ~\P2_reg2_reg[5]/NET0131  & ~n1048 ;
  assign n11941 = \P2_reg2_reg[4]/NET0131  & ~n1074 ;
  assign n11942 = ~\P2_reg2_reg[4]/NET0131  & n1074 ;
  assign n11943 = \P2_reg2_reg[3]/NET0131  & ~n1090 ;
  assign n11944 = ~\P2_reg2_reg[3]/NET0131  & n1090 ;
  assign n11946 = \P2_reg2_reg[2]/NET0131  & n1122 ;
  assign n11945 = ~\P2_reg2_reg[2]/NET0131  & ~n1122 ;
  assign n11948 = \P2_reg2_reg[1]/NET0131  & n1138 ;
  assign n11947 = ~\P2_reg2_reg[1]/NET0131  & ~n1138 ;
  assign n11981 = \P2_IR_reg[0]/NET0131  & ~\P2_reg2_reg[0]/NET0131  ;
  assign n11982 = ~n11947 & ~n11981 ;
  assign n11983 = ~n11948 & ~n11982 ;
  assign n11984 = ~n11945 & ~n11983 ;
  assign n11985 = ~n11946 & ~n11984 ;
  assign n11986 = ~n11944 & ~n11985 ;
  assign n11987 = ~n11943 & ~n11986 ;
  assign n11988 = ~n11942 & ~n11987 ;
  assign n11989 = ~n11941 & ~n11988 ;
  assign n11990 = ~n11960 & ~n11989 ;
  assign n11991 = ~n11940 & ~n11990 ;
  assign n11992 = ~n11959 & ~n11991 ;
  assign n11993 = ~n11939 & ~n11992 ;
  assign n11994 = ~n11966 & ~n11993 ;
  assign n11995 = ~n11938 & ~n11994 ;
  assign n11996 = ~n11965 & ~n11995 ;
  assign n11997 = ~n11937 & ~n11996 ;
  assign n11999 = n11936 & ~n11997 ;
  assign n11998 = ~n11936 & n11997 ;
  assign n12000 = n2262 & ~n11998 ;
  assign n12001 = ~n11999 & n12000 ;
  assign n11980 = n615 & ~n932 ;
  assign n12023 = n2035 & ~n11980 ;
  assign n12024 = ~n12001 & n12023 ;
  assign n12025 = ~n12022 & n12024 ;
  assign n11910 = ~\P2_IR_reg[0]/NET0131  & \P2_reg1_reg[0]/NET0131  ;
  assign n11911 = ~n11909 & ~n11910 ;
  assign n11912 = ~n11908 & ~n11911 ;
  assign n11913 = ~n11907 & ~n11912 ;
  assign n11914 = ~n11906 & ~n11913 ;
  assign n11915 = ~n11905 & ~n11914 ;
  assign n11916 = ~n11904 & ~n11915 ;
  assign n11917 = ~n11903 & n11916 ;
  assign n11920 = ~n11918 & ~n11919 ;
  assign n11921 = ~n11917 & n11920 ;
  assign n11922 = ~n11902 & ~n11921 ;
  assign n11923 = ~n11901 & ~n11922 ;
  assign n11924 = ~n11900 & ~n11923 ;
  assign n11925 = ~n11899 & ~n11924 ;
  assign n11926 = ~n11898 & ~n11925 ;
  assign n11927 = ~n11897 & n11926 ;
  assign n11929 = ~n11927 & ~n11928 ;
  assign n11931 = n11896 & n11929 ;
  assign n11930 = ~n11896 & ~n11929 ;
  assign n11932 = n2261 & ~n11930 ;
  assign n11933 = ~n11931 & n11932 ;
  assign n11949 = ~\P2_IR_reg[0]/NET0131  & \P2_reg2_reg[0]/NET0131  ;
  assign n11950 = ~n11948 & ~n11949 ;
  assign n11951 = ~n11947 & ~n11950 ;
  assign n11952 = ~n11946 & ~n11951 ;
  assign n11953 = ~n11945 & ~n11952 ;
  assign n11954 = ~n11944 & n11953 ;
  assign n11955 = ~n11943 & ~n11954 ;
  assign n11956 = ~n11942 & ~n11955 ;
  assign n11957 = ~n11941 & ~n11956 ;
  assign n11958 = ~n11940 & n11957 ;
  assign n11961 = ~n11959 & ~n11960 ;
  assign n11962 = ~n11958 & n11961 ;
  assign n11963 = ~n11939 & ~n11962 ;
  assign n11964 = ~n11938 & n11963 ;
  assign n11967 = ~n11965 & ~n11966 ;
  assign n11968 = ~n11964 & n11967 ;
  assign n11969 = ~n11937 & ~n11968 ;
  assign n11972 = n11936 & n11969 ;
  assign n11970 = ~n11936 & ~n11969 ;
  assign n11971 = n615 & n633 ;
  assign n11973 = ~n11970 & n11971 ;
  assign n11974 = ~n11972 & n11973 ;
  assign n11975 = \P2_addr_reg[9]/NET0131  & n634 ;
  assign n11893 = ~n932 & n2262 ;
  assign n11976 = ~n2035 & ~n11893 ;
  assign n11977 = ~n11975 & n11976 ;
  assign n11978 = ~n11974 & n11977 ;
  assign n11979 = ~n11933 & n11978 ;
  assign n12026 = \P1_state_reg[0]/NET0131  & ~n11979 ;
  assign n12027 = ~n12025 & n12026 ;
  assign n12028 = ~n7649 & ~n12027 ;
  assign n12029 = \P1_reg3_reg[0]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12038 = ~\P1_reg2_reg[0]/NET0131  & n2725 ;
  assign n12039 = n2731 & ~n12038 ;
  assign n12040 = ~\P1_IR_reg[0]/NET0131  & ~n11723 ;
  assign n12041 = ~n12039 & n12040 ;
  assign n12035 = n2725 & ~n11704 ;
  assign n12032 = ~\P1_IR_reg[0]/NET0131  & ~\P1_reg1_reg[0]/NET0131  ;
  assign n12033 = ~n11746 & ~n12032 ;
  assign n12034 = ~n2725 & n12033 ;
  assign n12036 = n2731 & ~n12034 ;
  assign n12037 = ~n12035 & n12036 ;
  assign n12030 = ~\P1_addr_reg[0]/NET0131  & ~n2731 ;
  assign n12031 = n11723 & n12030 ;
  assign n12042 = \P1_state_reg[0]/NET0131  & ~n12031 ;
  assign n12043 = ~n12037 & n12042 ;
  assign n12044 = ~n12041 & n12043 ;
  assign n12045 = ~n12029 & ~n12044 ;
  assign n12046 = ~n11773 & ~n11778 ;
  assign n12047 = ~n11777 & ~n11779 ;
  assign n12049 = n12046 & n12047 ;
  assign n12048 = ~n12046 & ~n12047 ;
  assign n12050 = n11728 & ~n12048 ;
  assign n12051 = ~n12049 & n12050 ;
  assign n12053 = n3253 & ~n11723 ;
  assign n12052 = ~\P1_addr_reg[10]/NET0131  & n11723 ;
  assign n12054 = ~n2731 & ~n12052 ;
  assign n12055 = ~n12053 & n12054 ;
  assign n12056 = ~n11798 & ~n11808 ;
  assign n12058 = ~n11805 & n12056 ;
  assign n12057 = n11805 & ~n12056 ;
  assign n12059 = n11686 & ~n12057 ;
  assign n12060 = ~n12058 & n12059 ;
  assign n12061 = ~n12055 & ~n12060 ;
  assign n12062 = ~n12051 & n12061 ;
  assign n12063 = \P1_state_reg[0]/NET0131  & ~n12062 ;
  assign n12064 = ~n7401 & ~n12063 ;
  assign n12079 = ~n11772 & ~n11784 ;
  assign n12081 = n11782 & ~n12079 ;
  assign n12080 = ~n11782 & n12079 ;
  assign n12082 = n11728 & ~n12080 ;
  assign n12083 = ~n12081 & n12082 ;
  assign n12065 = ~n11797 & ~n11807 ;
  assign n12066 = ~n11798 & n11801 ;
  assign n12067 = ~n11830 & n12066 ;
  assign n12068 = ~n11798 & n11803 ;
  assign n12069 = ~n11808 & ~n12068 ;
  assign n12070 = ~n12067 & n12069 ;
  assign n12072 = ~n12065 & n12070 ;
  assign n12071 = n12065 & ~n12070 ;
  assign n12073 = n11686 & ~n12071 ;
  assign n12074 = ~n12072 & n12073 ;
  assign n12076 = n3201 & ~n11723 ;
  assign n12075 = ~\P1_addr_reg[11]/NET0131  & n11723 ;
  assign n12077 = ~n2731 & ~n12075 ;
  assign n12078 = ~n12076 & n12077 ;
  assign n12084 = ~n12074 & ~n12078 ;
  assign n12085 = ~n12083 & n12084 ;
  assign n12086 = \P1_state_reg[0]/NET0131  & ~n12085 ;
  assign n12087 = ~n7991 & ~n12086 ;
  assign n12101 = ~n11878 & ~n11879 ;
  assign n12103 = ~n11882 & n12101 ;
  assign n12102 = n11882 & ~n12101 ;
  assign n12104 = n11728 & ~n12102 ;
  assign n12105 = ~n12103 & n12104 ;
  assign n12089 = ~n3673 & ~n11723 ;
  assign n12088 = ~\P1_addr_reg[13]/NET0131  & n11723 ;
  assign n12090 = ~n2731 & ~n12088 ;
  assign n12091 = ~n12089 & n12090 ;
  assign n12092 = ~n11865 & ~n11866 ;
  assign n12093 = ~n11807 & n12070 ;
  assign n12094 = ~n11795 & ~n11797 ;
  assign n12095 = ~n12093 & n12094 ;
  assign n12096 = ~n11794 & ~n12095 ;
  assign n12098 = n12092 & ~n12096 ;
  assign n12097 = ~n12092 & n12096 ;
  assign n12099 = n11686 & ~n12097 ;
  assign n12100 = ~n12098 & n12099 ;
  assign n12106 = ~n12091 & ~n12100 ;
  assign n12107 = ~n12105 & n12106 ;
  assign n12108 = \P1_state_reg[0]/NET0131  & ~n12107 ;
  assign n12109 = ~n7445 & ~n12108 ;
  assign n12110 = ~\P1_state_reg[0]/NET0131  & ~\P2_reg3_reg[0]/NET0131  ;
  assign n12113 = \P2_IR_reg[0]/NET0131  & n615 ;
  assign n12116 = n2035 & ~n12113 ;
  assign n12111 = ~n11949 & ~n11981 ;
  assign n12112 = n2262 & ~n12111 ;
  assign n12114 = ~n11910 & ~n12002 ;
  assign n12115 = n634 & ~n12114 ;
  assign n12117 = ~n12112 & ~n12115 ;
  assign n12118 = n12116 & n12117 ;
  assign n12119 = \P2_addr_reg[0]/NET0131  & n634 ;
  assign n12123 = ~n2035 & ~n12119 ;
  assign n12122 = n2261 & ~n12114 ;
  assign n12120 = \P2_IR_reg[0]/NET0131  & n2262 ;
  assign n12121 = n11971 & ~n12111 ;
  assign n12124 = ~n12120 & ~n12121 ;
  assign n12125 = ~n12122 & n12124 ;
  assign n12126 = n12123 & n12125 ;
  assign n12127 = ~n12118 & ~n12126 ;
  assign n12128 = \P1_state_reg[0]/NET0131  & ~n12127 ;
  assign n12129 = ~n12110 & ~n12128 ;
  assign n12146 = \P1_reg1_reg[15]/NET0131  & n3722 ;
  assign n12147 = ~\P1_reg1_reg[15]/NET0131  & ~n3722 ;
  assign n12148 = ~n12146 & ~n12147 ;
  assign n12149 = ~n11876 & ~n11884 ;
  assign n12150 = ~n11875 & ~n12149 ;
  assign n12152 = n12148 & ~n12150 ;
  assign n12151 = ~n12148 & n12150 ;
  assign n12153 = n11728 & ~n12151 ;
  assign n12154 = ~n12152 & n12153 ;
  assign n12134 = \P1_reg2_reg[15]/NET0131  & n3722 ;
  assign n12130 = ~n11865 & ~n12096 ;
  assign n12131 = ~n11862 & ~n11866 ;
  assign n12132 = ~n12130 & n12131 ;
  assign n12133 = ~n11863 & ~n12132 ;
  assign n12135 = ~\P1_reg2_reg[15]/NET0131  & ~n3722 ;
  assign n12138 = n12133 & ~n12135 ;
  assign n12139 = ~n12134 & n12138 ;
  assign n12136 = ~n12134 & ~n12135 ;
  assign n12137 = ~n12133 & ~n12136 ;
  assign n12140 = n11686 & ~n12137 ;
  assign n12141 = ~n12139 & n12140 ;
  assign n12143 = ~n3722 & ~n11723 ;
  assign n12142 = ~\P1_addr_reg[15]/NET0131  & n11723 ;
  assign n12144 = ~n2731 & ~n12142 ;
  assign n12145 = ~n12143 & n12144 ;
  assign n12155 = ~n12141 & ~n12145 ;
  assign n12156 = ~n12154 & n12155 ;
  assign n12157 = \P1_state_reg[0]/NET0131  & ~n12156 ;
  assign n12158 = ~n8031 & ~n12157 ;
  assign n12178 = ~\P2_reg2_reg[12]/NET0131  & n848 ;
  assign n12179 = \P2_reg2_reg[12]/NET0131  & ~n848 ;
  assign n12180 = ~n12178 & ~n12179 ;
  assign n12181 = \P2_reg2_reg[11]/NET0131  & ~n880 ;
  assign n12193 = ~\P2_reg2_reg[11]/NET0131  & n880 ;
  assign n12182 = \P2_reg2_reg[10]/NET0131  & ~n907 ;
  assign n12194 = ~\P2_reg2_reg[10]/NET0131  & n907 ;
  assign n12218 = ~n11934 & n11997 ;
  assign n12219 = ~n11935 & ~n12218 ;
  assign n12220 = ~n12194 & n12219 ;
  assign n12221 = ~n12182 & ~n12220 ;
  assign n12222 = ~n12193 & ~n12221 ;
  assign n12223 = ~n12181 & ~n12222 ;
  assign n12225 = ~n12180 & n12223 ;
  assign n12224 = n12180 & ~n12223 ;
  assign n12226 = n2262 & ~n12224 ;
  assign n12227 = ~n12225 & n12226 ;
  assign n12160 = ~\P2_reg1_reg[12]/NET0131  & n848 ;
  assign n12161 = \P2_reg1_reg[12]/NET0131  & ~n848 ;
  assign n12162 = ~n12160 & ~n12161 ;
  assign n12164 = \P2_reg1_reg[11]/NET0131  & ~n880 ;
  assign n12163 = ~\P2_reg1_reg[11]/NET0131  & n880 ;
  assign n12166 = \P2_reg1_reg[10]/NET0131  & ~n907 ;
  assign n12165 = ~\P2_reg1_reg[10]/NET0131  & n907 ;
  assign n12208 = ~n11895 & n12018 ;
  assign n12209 = ~n11894 & ~n12208 ;
  assign n12210 = ~n12165 & n12209 ;
  assign n12211 = ~n12166 & ~n12210 ;
  assign n12212 = ~n12163 & ~n12211 ;
  assign n12213 = ~n12164 & ~n12212 ;
  assign n12215 = n12162 & ~n12213 ;
  assign n12214 = ~n12162 & n12213 ;
  assign n12216 = n634 & ~n12214 ;
  assign n12217 = ~n12215 & n12216 ;
  assign n12207 = n615 & n848 ;
  assign n12228 = n2035 & ~n12207 ;
  assign n12229 = ~n12217 & n12228 ;
  assign n12230 = ~n12227 & n12229 ;
  assign n12167 = ~n11895 & ~n11928 ;
  assign n12168 = ~n11927 & n12167 ;
  assign n12169 = ~n11894 & ~n12168 ;
  assign n12170 = ~n12166 & ~n12169 ;
  assign n12171 = ~n12165 & ~n12170 ;
  assign n12172 = ~n12164 & ~n12171 ;
  assign n12173 = ~n12163 & ~n12172 ;
  assign n12175 = n12162 & ~n12173 ;
  assign n12174 = ~n12162 & n12173 ;
  assign n12176 = n2261 & ~n12174 ;
  assign n12177 = ~n12175 & n12176 ;
  assign n12183 = ~n11958 & ~n11960 ;
  assign n12184 = ~n11939 & ~n12183 ;
  assign n12185 = ~n11959 & ~n11966 ;
  assign n12186 = ~n12184 & n12185 ;
  assign n12187 = ~n11938 & ~n12186 ;
  assign n12188 = ~n11937 & n12187 ;
  assign n12189 = ~n11935 & ~n11965 ;
  assign n12190 = ~n12188 & n12189 ;
  assign n12191 = ~n11934 & ~n12190 ;
  assign n12192 = ~n12182 & n12191 ;
  assign n12195 = ~n12193 & ~n12194 ;
  assign n12196 = ~n12192 & n12195 ;
  assign n12197 = ~n12181 & ~n12196 ;
  assign n12199 = n12180 & n12197 ;
  assign n12198 = ~n12180 & ~n12197 ;
  assign n12200 = n11971 & ~n12198 ;
  assign n12201 = ~n12199 & n12200 ;
  assign n12202 = \P2_addr_reg[12]/NET0131  & n634 ;
  assign n12159 = n848 & n2262 ;
  assign n12203 = ~n2035 & ~n12159 ;
  assign n12204 = ~n12202 & n12203 ;
  assign n12205 = ~n12201 & n12204 ;
  assign n12206 = ~n12177 & n12205 ;
  assign n12231 = \P1_state_reg[0]/NET0131  & ~n12206 ;
  assign n12232 = ~n12230 & n12231 ;
  assign n12233 = ~n7527 & ~n12232 ;
  assign n12249 = \P1_reg1_reg[16]/NET0131  & n3698 ;
  assign n12250 = ~\P1_reg1_reg[16]/NET0131  & ~n3698 ;
  assign n12251 = ~n12249 & ~n12250 ;
  assign n12252 = ~n11875 & ~n12146 ;
  assign n12253 = ~n12149 & n12252 ;
  assign n12254 = ~n12147 & ~n12253 ;
  assign n12256 = n12251 & n12254 ;
  assign n12255 = ~n12251 & ~n12254 ;
  assign n12257 = n11728 & ~n12255 ;
  assign n12258 = ~n12256 & n12257 ;
  assign n12235 = ~n3698 & ~n11723 ;
  assign n12234 = ~\P1_addr_reg[16]/NET0131  & n11723 ;
  assign n12236 = ~n2731 & ~n12234 ;
  assign n12237 = ~n12235 & n12236 ;
  assign n12238 = \P1_reg2_reg[16]/NET0131  & n3698 ;
  assign n12239 = ~\P1_reg2_reg[16]/NET0131  & ~n3698 ;
  assign n12240 = ~n12238 & ~n12239 ;
  assign n12241 = ~n11863 & n11870 ;
  assign n12242 = ~n11862 & ~n12134 ;
  assign n12243 = ~n12241 & n12242 ;
  assign n12244 = ~n12135 & ~n12243 ;
  assign n12246 = n12240 & n12244 ;
  assign n12245 = ~n12240 & ~n12244 ;
  assign n12247 = n11686 & ~n12245 ;
  assign n12248 = ~n12246 & n12247 ;
  assign n12259 = ~n12237 & ~n12248 ;
  assign n12260 = ~n12258 & n12259 ;
  assign n12261 = \P1_state_reg[0]/NET0131  & ~n12260 ;
  assign n12262 = ~n6625 & ~n12261 ;
  assign n12264 = ~\P2_reg1_reg[13]/NET0131  & n809 ;
  assign n12265 = \P2_reg1_reg[13]/NET0131  & ~n809 ;
  assign n12266 = ~n12264 & ~n12265 ;
  assign n12295 = ~n12161 & ~n12164 ;
  assign n12296 = ~n12212 & n12295 ;
  assign n12297 = ~n12160 & ~n12296 ;
  assign n12299 = n12266 & n12297 ;
  assign n12298 = ~n12266 & ~n12297 ;
  assign n12300 = n634 & ~n12298 ;
  assign n12301 = ~n12299 & n12300 ;
  assign n12274 = ~\P2_reg2_reg[13]/NET0131  & n809 ;
  assign n12275 = \P2_reg2_reg[13]/NET0131  & ~n809 ;
  assign n12276 = ~n12274 & ~n12275 ;
  assign n12277 = ~n12178 & ~n12193 ;
  assign n12302 = ~n12221 & n12277 ;
  assign n12303 = ~n12178 & n12181 ;
  assign n12304 = ~n12179 & ~n12303 ;
  assign n12305 = ~n12302 & n12304 ;
  assign n12307 = ~n12276 & n12305 ;
  assign n12306 = n12276 & ~n12305 ;
  assign n12308 = n2262 & ~n12306 ;
  assign n12309 = ~n12307 & n12308 ;
  assign n12294 = n615 & n809 ;
  assign n12310 = n2035 & ~n12294 ;
  assign n12311 = ~n12309 & n12310 ;
  assign n12312 = ~n12301 & n12311 ;
  assign n12267 = ~n12160 & ~n12163 ;
  assign n12268 = ~n12172 & n12267 ;
  assign n12269 = ~n12161 & ~n12268 ;
  assign n12271 = n12266 & n12269 ;
  assign n12270 = ~n12266 & ~n12269 ;
  assign n12272 = n2261 & ~n12270 ;
  assign n12273 = ~n12271 & n12272 ;
  assign n12278 = ~n11934 & n11969 ;
  assign n12279 = ~n11935 & ~n12194 ;
  assign n12280 = ~n12278 & n12279 ;
  assign n12281 = ~n12182 & ~n12280 ;
  assign n12282 = ~n12181 & n12281 ;
  assign n12283 = n12277 & ~n12282 ;
  assign n12284 = ~n12179 & ~n12283 ;
  assign n12286 = n12276 & n12284 ;
  assign n12285 = ~n12276 & ~n12284 ;
  assign n12287 = n11971 & ~n12285 ;
  assign n12288 = ~n12286 & n12287 ;
  assign n12289 = n809 & n2262 ;
  assign n12263 = \P2_addr_reg[13]/NET0131  & n634 ;
  assign n12290 = ~n2035 & ~n12263 ;
  assign n12291 = ~n12289 & n12290 ;
  assign n12292 = ~n12288 & n12291 ;
  assign n12293 = ~n12273 & n12292 ;
  assign n12313 = \P1_state_reg[0]/NET0131  & ~n12293 ;
  assign n12314 = ~n12312 & n12313 ;
  assign n12315 = ~n7567 & ~n12314 ;
  assign n12330 = ~\P1_reg1_reg[17]/NET0131  & n3593 ;
  assign n12331 = \P1_reg1_reg[17]/NET0131  & ~n3593 ;
  assign n12332 = ~n12330 & ~n12331 ;
  assign n12333 = ~n11875 & ~n11878 ;
  assign n12334 = ~n11883 & n12333 ;
  assign n12335 = ~n11876 & ~n12147 ;
  assign n12336 = ~n12334 & n12335 ;
  assign n12337 = ~n12146 & ~n12249 ;
  assign n12338 = ~n12336 & n12337 ;
  assign n12339 = ~n12250 & ~n12338 ;
  assign n12341 = ~n12332 & ~n12339 ;
  assign n12340 = n12332 & n12339 ;
  assign n12342 = n11728 & ~n12340 ;
  assign n12343 = ~n12341 & n12342 ;
  assign n12316 = ~\P1_reg2_reg[17]/NET0131  & n3593 ;
  assign n12317 = \P1_reg2_reg[17]/NET0131  & ~n3593 ;
  assign n12318 = ~n12316 & ~n12317 ;
  assign n12319 = ~n12134 & ~n12238 ;
  assign n12320 = ~n12138 & n12319 ;
  assign n12321 = ~n12239 & ~n12320 ;
  assign n12323 = ~n12318 & ~n12321 ;
  assign n12322 = n12318 & n12321 ;
  assign n12324 = n11686 & ~n12322 ;
  assign n12325 = ~n12323 & n12324 ;
  assign n12327 = n3593 & ~n11723 ;
  assign n12326 = ~\P1_addr_reg[17]/NET0131  & n11723 ;
  assign n12328 = ~n2731 & ~n12326 ;
  assign n12329 = ~n12327 & n12328 ;
  assign n12344 = ~n12325 & ~n12329 ;
  assign n12345 = ~n12343 & n12344 ;
  assign n12346 = \P1_state_reg[0]/NET0131  & ~n12345 ;
  assign n12347 = ~n6004 & ~n12346 ;
  assign n12349 = ~\P2_reg1_reg[15]/NET0131  & n716 ;
  assign n12350 = \P2_reg1_reg[15]/NET0131  & ~n716 ;
  assign n12351 = ~n12349 & ~n12350 ;
  assign n12353 = ~\P2_reg1_reg[14]/NET0131  & n758 ;
  assign n12354 = ~n12264 & ~n12353 ;
  assign n12381 = n12297 & n12354 ;
  assign n12352 = \P2_reg1_reg[14]/NET0131  & ~n758 ;
  assign n12382 = n12265 & ~n12353 ;
  assign n12383 = ~n12352 & ~n12382 ;
  assign n12384 = ~n12381 & n12383 ;
  assign n12386 = n12351 & ~n12384 ;
  assign n12385 = ~n12351 & n12384 ;
  assign n12387 = n634 & ~n12385 ;
  assign n12388 = ~n12386 & n12387 ;
  assign n12362 = ~\P2_reg2_reg[15]/NET0131  & n716 ;
  assign n12363 = \P2_reg2_reg[15]/NET0131  & ~n716 ;
  assign n12364 = ~n12362 & ~n12363 ;
  assign n12366 = ~\P2_reg2_reg[14]/NET0131  & n758 ;
  assign n12367 = ~n12274 & ~n12366 ;
  assign n12389 = ~n12305 & n12367 ;
  assign n12365 = \P2_reg2_reg[14]/NET0131  & ~n758 ;
  assign n12390 = n12275 & ~n12366 ;
  assign n12391 = ~n12365 & ~n12390 ;
  assign n12392 = ~n12389 & n12391 ;
  assign n12394 = ~n12364 & n12392 ;
  assign n12393 = n12364 & ~n12392 ;
  assign n12395 = n2262 & ~n12393 ;
  assign n12396 = ~n12394 & n12395 ;
  assign n12380 = n615 & n716 ;
  assign n12397 = n2035 & ~n12380 ;
  assign n12398 = ~n12396 & n12397 ;
  assign n12399 = ~n12388 & n12398 ;
  assign n12355 = ~n12265 & n12269 ;
  assign n12356 = n12354 & ~n12355 ;
  assign n12357 = ~n12352 & ~n12356 ;
  assign n12359 = n12351 & n12357 ;
  assign n12358 = ~n12351 & ~n12357 ;
  assign n12360 = n2261 & ~n12358 ;
  assign n12361 = ~n12359 & n12360 ;
  assign n12368 = ~n12275 & n12284 ;
  assign n12369 = n12367 & ~n12368 ;
  assign n12370 = ~n12365 & ~n12369 ;
  assign n12372 = n12364 & n12370 ;
  assign n12371 = ~n12364 & ~n12370 ;
  assign n12373 = n11971 & ~n12371 ;
  assign n12374 = ~n12372 & n12373 ;
  assign n12375 = n716 & n2262 ;
  assign n12348 = \P2_addr_reg[15]/NET0131  & n634 ;
  assign n12376 = ~n2035 & ~n12348 ;
  assign n12377 = ~n12375 & n12376 ;
  assign n12378 = ~n12374 & n12377 ;
  assign n12379 = ~n12361 & n12378 ;
  assign n12400 = \P1_state_reg[0]/NET0131  & ~n12379 ;
  assign n12401 = ~n12399 & n12400 ;
  assign n12402 = ~n8197 & ~n12401 ;
  assign n12419 = ~\P2_reg2_reg[16]/NET0131  & n1253 ;
  assign n12420 = \P2_reg2_reg[16]/NET0131  & ~n1253 ;
  assign n12421 = ~n12419 & ~n12420 ;
  assign n12452 = ~n12363 & ~n12365 ;
  assign n12453 = ~n12178 & ~n12223 ;
  assign n12454 = ~n12179 & ~n12275 ;
  assign n12455 = ~n12453 & n12454 ;
  assign n12456 = ~n12274 & ~n12455 ;
  assign n12457 = ~n12366 & n12456 ;
  assign n12458 = n12452 & ~n12457 ;
  assign n12459 = ~n12362 & ~n12458 ;
  assign n12461 = n12421 & n12459 ;
  assign n12460 = ~n12421 & ~n12459 ;
  assign n12462 = n2262 & ~n12460 ;
  assign n12463 = ~n12461 & n12462 ;
  assign n12404 = ~\P2_reg1_reg[16]/NET0131  & n1253 ;
  assign n12405 = \P2_reg1_reg[16]/NET0131  & ~n1253 ;
  assign n12406 = ~n12404 & ~n12405 ;
  assign n12440 = ~n12350 & ~n12352 ;
  assign n12441 = ~n12160 & ~n12213 ;
  assign n12442 = ~n12161 & ~n12265 ;
  assign n12443 = ~n12441 & n12442 ;
  assign n12444 = ~n12264 & ~n12443 ;
  assign n12445 = ~n12353 & n12444 ;
  assign n12446 = n12440 & ~n12445 ;
  assign n12447 = ~n12349 & ~n12446 ;
  assign n12449 = ~n12406 & ~n12447 ;
  assign n12448 = n12406 & n12447 ;
  assign n12450 = n634 & ~n12448 ;
  assign n12451 = ~n12449 & n12450 ;
  assign n12439 = n615 & n1253 ;
  assign n12464 = n2035 & ~n12439 ;
  assign n12465 = ~n12451 & n12464 ;
  assign n12466 = ~n12463 & n12465 ;
  assign n12407 = ~n12349 & ~n12353 ;
  assign n12408 = ~n12161 & ~n12173 ;
  assign n12409 = ~n12160 & ~n12264 ;
  assign n12410 = ~n12408 & n12409 ;
  assign n12411 = ~n12265 & ~n12410 ;
  assign n12412 = ~n12352 & n12411 ;
  assign n12413 = n12407 & ~n12412 ;
  assign n12414 = ~n12350 & ~n12413 ;
  assign n12416 = n12406 & n12414 ;
  assign n12415 = ~n12406 & ~n12414 ;
  assign n12417 = n2261 & ~n12415 ;
  assign n12418 = ~n12416 & n12417 ;
  assign n12422 = ~n12362 & ~n12366 ;
  assign n12423 = ~n12179 & n12197 ;
  assign n12424 = ~n12178 & ~n12274 ;
  assign n12425 = ~n12423 & n12424 ;
  assign n12426 = ~n12275 & ~n12425 ;
  assign n12427 = ~n12365 & n12426 ;
  assign n12428 = n12422 & ~n12427 ;
  assign n12429 = ~n12363 & ~n12428 ;
  assign n12431 = n12421 & n12429 ;
  assign n12430 = ~n12421 & ~n12429 ;
  assign n12432 = n11971 & ~n12430 ;
  assign n12433 = ~n12431 & n12432 ;
  assign n12434 = n1253 & n2262 ;
  assign n12403 = \P2_addr_reg[16]/NET0131  & n634 ;
  assign n12435 = ~n2035 & ~n12403 ;
  assign n12436 = ~n12434 & n12435 ;
  assign n12437 = ~n12433 & n12436 ;
  assign n12438 = ~n12418 & n12437 ;
  assign n12467 = \P1_state_reg[0]/NET0131  & ~n12438 ;
  assign n12468 = ~n12466 & n12467 ;
  assign n12469 = ~n6096 & ~n12468 ;
  assign n12471 = ~\P2_reg1_reg[17]/NET0131  & n1219 ;
  assign n12472 = \P2_reg1_reg[17]/NET0131  & ~n1219 ;
  assign n12473 = ~n12471 & ~n12472 ;
  assign n12474 = ~n12349 & ~n12404 ;
  assign n12499 = ~n12265 & ~n12297 ;
  assign n12500 = n12354 & ~n12499 ;
  assign n12501 = ~n12352 & ~n12500 ;
  assign n12502 = n12474 & ~n12501 ;
  assign n12503 = n12350 & ~n12404 ;
  assign n12504 = ~n12405 & ~n12503 ;
  assign n12505 = ~n12502 & n12504 ;
  assign n12507 = n12473 & ~n12505 ;
  assign n12506 = ~n12473 & n12505 ;
  assign n12508 = n634 & ~n12506 ;
  assign n12509 = ~n12507 & n12508 ;
  assign n12482 = ~\P2_reg2_reg[17]/NET0131  & n1219 ;
  assign n12483 = \P2_reg2_reg[17]/NET0131  & ~n1219 ;
  assign n12484 = ~n12482 & ~n12483 ;
  assign n12485 = ~n12362 & ~n12419 ;
  assign n12510 = ~n12275 & n12305 ;
  assign n12511 = n12367 & ~n12510 ;
  assign n12512 = ~n12365 & ~n12511 ;
  assign n12513 = n12485 & ~n12512 ;
  assign n12514 = n12363 & ~n12419 ;
  assign n12515 = ~n12420 & ~n12514 ;
  assign n12516 = ~n12513 & n12515 ;
  assign n12518 = n12484 & ~n12516 ;
  assign n12517 = ~n12484 & n12516 ;
  assign n12519 = n2262 & ~n12517 ;
  assign n12520 = ~n12518 & n12519 ;
  assign n12498 = n615 & n1219 ;
  assign n12521 = n2035 & ~n12498 ;
  assign n12522 = ~n12520 & n12521 ;
  assign n12523 = ~n12509 & n12522 ;
  assign n12475 = ~n12350 & n12357 ;
  assign n12476 = n12474 & ~n12475 ;
  assign n12477 = ~n12405 & ~n12476 ;
  assign n12479 = n12473 & n12477 ;
  assign n12478 = ~n12473 & ~n12477 ;
  assign n12480 = n2261 & ~n12478 ;
  assign n12481 = ~n12479 & n12480 ;
  assign n12486 = ~n12363 & n12370 ;
  assign n12487 = n12485 & ~n12486 ;
  assign n12488 = ~n12420 & ~n12487 ;
  assign n12490 = n12484 & n12488 ;
  assign n12489 = ~n12484 & ~n12488 ;
  assign n12491 = n11971 & ~n12489 ;
  assign n12492 = ~n12490 & n12491 ;
  assign n12493 = n1219 & n2262 ;
  assign n12470 = \P2_addr_reg[17]/NET0131  & n634 ;
  assign n12494 = ~n2035 & ~n12470 ;
  assign n12495 = ~n12493 & n12494 ;
  assign n12496 = ~n12492 & n12495 ;
  assign n12497 = ~n12481 & n12496 ;
  assign n12524 = \P1_state_reg[0]/NET0131  & ~n12497 ;
  assign n12525 = ~n12523 & n12524 ;
  assign n12526 = ~n4344 & ~n12525 ;
  assign n12528 = ~\P2_reg1_reg[18]/NET0131  & n1332 ;
  assign n12529 = \P2_reg1_reg[18]/NET0131  & ~n1332 ;
  assign n12530 = ~n12528 & ~n12529 ;
  assign n12535 = ~n12404 & ~n12471 ;
  assign n12568 = ~n12405 & n12414 ;
  assign n12569 = n12535 & ~n12568 ;
  assign n12570 = ~n12472 & ~n12569 ;
  assign n12572 = ~n12530 & ~n12570 ;
  assign n12571 = n12530 & n12570 ;
  assign n12573 = n2261 & ~n12571 ;
  assign n12574 = ~n12572 & n12573 ;
  assign n12543 = ~\P2_reg2_reg[18]/NET0131  & n1332 ;
  assign n12544 = \P2_reg2_reg[18]/NET0131  & ~n1332 ;
  assign n12545 = ~n12543 & ~n12544 ;
  assign n12550 = ~n12419 & ~n12482 ;
  assign n12561 = ~n12420 & n12429 ;
  assign n12562 = n12550 & ~n12561 ;
  assign n12563 = ~n12483 & ~n12562 ;
  assign n12565 = ~n12545 & ~n12563 ;
  assign n12564 = n12545 & n12563 ;
  assign n12566 = n11971 & ~n12564 ;
  assign n12567 = ~n12565 & n12566 ;
  assign n12576 = \P2_addr_reg[18]/NET0131  & n634 ;
  assign n12575 = n1332 & n2262 ;
  assign n12577 = ~n2035 & ~n12575 ;
  assign n12578 = ~n12576 & n12577 ;
  assign n12579 = ~n12567 & n12578 ;
  assign n12580 = ~n12574 & n12579 ;
  assign n12546 = ~n12452 & n12485 ;
  assign n12547 = ~n12420 & ~n12483 ;
  assign n12548 = ~n12546 & n12547 ;
  assign n12549 = ~n12482 & ~n12548 ;
  assign n12551 = n12422 & n12550 ;
  assign n12552 = n12456 & n12551 ;
  assign n12553 = ~n12549 & ~n12552 ;
  assign n12555 = n12545 & ~n12553 ;
  assign n12554 = ~n12545 & n12553 ;
  assign n12556 = n2262 & ~n12554 ;
  assign n12557 = ~n12555 & n12556 ;
  assign n12531 = ~n12440 & n12474 ;
  assign n12532 = ~n12405 & ~n12472 ;
  assign n12533 = ~n12531 & n12532 ;
  assign n12534 = ~n12471 & ~n12533 ;
  assign n12536 = n12407 & n12535 ;
  assign n12537 = n12444 & n12536 ;
  assign n12538 = ~n12534 & ~n12537 ;
  assign n12540 = ~n12530 & n12538 ;
  assign n12539 = n12530 & ~n12538 ;
  assign n12541 = n634 & ~n12539 ;
  assign n12542 = ~n12540 & n12541 ;
  assign n12527 = n615 & n1332 ;
  assign n12558 = n2035 & ~n12527 ;
  assign n12559 = ~n12542 & n12558 ;
  assign n12560 = ~n12557 & n12559 ;
  assign n12581 = \P1_state_reg[0]/NET0131  & ~n12560 ;
  assign n12582 = ~n12580 & n12581 ;
  assign n12583 = ~n4231 & ~n12582 ;
  assign n12590 = ~n11900 & ~n11901 ;
  assign n12592 = ~n12012 & ~n12590 ;
  assign n12591 = n12012 & n12590 ;
  assign n12593 = n634 & ~n12591 ;
  assign n12594 = ~n12592 & n12593 ;
  assign n12585 = ~n11939 & ~n11959 ;
  assign n12587 = ~n11991 & n12585 ;
  assign n12586 = n11991 & ~n12585 ;
  assign n12588 = n2262 & ~n12586 ;
  assign n12589 = ~n12587 & n12588 ;
  assign n12584 = n615 & n1001 ;
  assign n12595 = n2035 & ~n12584 ;
  assign n12596 = ~n12589 & n12595 ;
  assign n12597 = ~n12594 & n12596 ;
  assign n12604 = ~n12183 & n12585 ;
  assign n12603 = n12183 & ~n12585 ;
  assign n12605 = n11971 & ~n12603 ;
  assign n12606 = ~n12604 & n12605 ;
  assign n12600 = ~n11922 & n12590 ;
  assign n12599 = n11922 & ~n12590 ;
  assign n12601 = n2261 & ~n12599 ;
  assign n12602 = ~n12600 & n12601 ;
  assign n12607 = \P2_addr_reg[6]/NET0131  & n634 ;
  assign n12598 = n1001 & n2262 ;
  assign n12608 = ~n2035 & ~n12598 ;
  assign n12609 = ~n12607 & n12608 ;
  assign n12610 = ~n12602 & n12609 ;
  assign n12611 = ~n12606 & n12610 ;
  assign n12612 = \P1_state_reg[0]/NET0131  & ~n12611 ;
  assign n12613 = ~n12597 & n12612 ;
  assign n12614 = ~n9195 & ~n12613 ;
  assign n12620 = ~n11702 & ~n11703 ;
  assign n12621 = ~n11704 & ~n12620 ;
  assign n12622 = n11704 & n12620 ;
  assign n12623 = ~n12621 & ~n12622 ;
  assign n12624 = n2725 & n12623 ;
  assign n12615 = ~n11744 & ~n11745 ;
  assign n12616 = n11746 & ~n12615 ;
  assign n12617 = ~n11746 & n12615 ;
  assign n12618 = ~n12616 & ~n12617 ;
  assign n12619 = ~n2725 & ~n12618 ;
  assign n12625 = n2731 & ~n12619 ;
  assign n12626 = ~n12624 & n12625 ;
  assign n12628 = n3385 & ~n11723 ;
  assign n12627 = \P1_addr_reg[1]/NET0131  & n11723 ;
  assign n12629 = ~n2731 & ~n12627 ;
  assign n12630 = ~n12628 & n12629 ;
  assign n12631 = ~n12626 & ~n12630 ;
  assign n12632 = \P1_state_reg[0]/NET0131  & ~n12631 ;
  assign n12633 = ~\P1_reg3_reg[1]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12634 = ~n12632 & ~n12633 ;
  assign n12640 = ~n11700 & ~n11701 ;
  assign n12641 = ~n11706 & ~n12640 ;
  assign n12642 = n11706 & n12640 ;
  assign n12643 = ~n12641 & ~n12642 ;
  assign n12644 = n2725 & n12643 ;
  assign n12635 = ~n11742 & ~n11743 ;
  assign n12636 = ~n11748 & n12635 ;
  assign n12637 = n11748 & ~n12635 ;
  assign n12638 = ~n12636 & ~n12637 ;
  assign n12639 = ~n2725 & ~n12638 ;
  assign n12645 = n2731 & ~n12639 ;
  assign n12646 = ~n12644 & n12645 ;
  assign n12648 = n3352 & ~n11723 ;
  assign n12647 = \P1_addr_reg[2]/NET0131  & n11723 ;
  assign n12649 = ~n2731 & ~n12647 ;
  assign n12650 = ~n12648 & n12649 ;
  assign n12651 = ~n12646 & ~n12650 ;
  assign n12652 = \P1_state_reg[0]/NET0131  & ~n12651 ;
  assign n12653 = ~\P1_reg3_reg[2]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12654 = ~n12652 & ~n12653 ;
  assign n12666 = ~n3369 & ~n11723 ;
  assign n12665 = ~\P1_addr_reg[3]/NET0131  & n11723 ;
  assign n12667 = ~n2731 & ~n12665 ;
  assign n12668 = ~n12666 & n12667 ;
  assign n12655 = ~n11740 & ~n11741 ;
  assign n12656 = ~n11750 & ~n12655 ;
  assign n12657 = n11750 & n12655 ;
  assign n12658 = ~n12656 & ~n12657 ;
  assign n12659 = n11728 & n12658 ;
  assign n12660 = ~n11698 & ~n11699 ;
  assign n12661 = ~n11708 & ~n12660 ;
  assign n12662 = n11708 & n12660 ;
  assign n12663 = ~n12661 & ~n12662 ;
  assign n12664 = n11686 & n12663 ;
  assign n12669 = ~n12659 & ~n12664 ;
  assign n12670 = ~n12668 & n12669 ;
  assign n12671 = \P1_state_reg[0]/NET0131  & ~n12670 ;
  assign n12672 = ~n9727 & ~n12671 ;
  assign n12684 = n3330 & ~n11723 ;
  assign n12683 = ~\P1_addr_reg[4]/NET0131  & n11723 ;
  assign n12685 = ~n2731 & ~n12683 ;
  assign n12686 = ~n12684 & n12685 ;
  assign n12673 = ~n11738 & ~n11739 ;
  assign n12674 = n11752 & n12673 ;
  assign n12675 = ~n11752 & ~n12673 ;
  assign n12676 = ~n12674 & ~n12675 ;
  assign n12677 = n11728 & n12676 ;
  assign n12678 = ~n11696 & ~n11697 ;
  assign n12679 = ~n11710 & ~n12678 ;
  assign n12680 = n11710 & n12678 ;
  assign n12681 = ~n12679 & ~n12680 ;
  assign n12682 = n11686 & n12681 ;
  assign n12687 = ~n12677 & ~n12682 ;
  assign n12688 = ~n12686 & n12687 ;
  assign n12689 = \P1_state_reg[0]/NET0131  & ~n12688 ;
  assign n12690 = ~n9068 & ~n12689 ;
  assign n12702 = ~n3509 & ~n11723 ;
  assign n12701 = ~\P1_addr_reg[5]/NET0131  & n11723 ;
  assign n12703 = ~n2731 & ~n12701 ;
  assign n12704 = ~n12702 & n12703 ;
  assign n12691 = ~n11694 & ~n11695 ;
  assign n12693 = ~n11712 & n12691 ;
  assign n12692 = n11712 & ~n12691 ;
  assign n12694 = n11686 & ~n12692 ;
  assign n12695 = ~n12693 & n12694 ;
  assign n12696 = ~n11736 & ~n11737 ;
  assign n12698 = ~n11754 & n12696 ;
  assign n12697 = n11754 & ~n12696 ;
  assign n12699 = n11728 & ~n12697 ;
  assign n12700 = ~n12698 & n12699 ;
  assign n12705 = ~n12695 & ~n12700 ;
  assign n12706 = ~n12704 & n12705 ;
  assign n12707 = \P1_state_reg[0]/NET0131  & ~n12706 ;
  assign n12708 = ~n9109 & ~n12707 ;
  assign n12718 = ~n11692 & ~n11693 ;
  assign n12720 = ~n11714 & n12718 ;
  assign n12719 = n11714 & ~n12718 ;
  assign n12721 = n11686 & ~n12719 ;
  assign n12722 = ~n12720 & n12721 ;
  assign n12710 = ~n3483 & ~n11723 ;
  assign n12709 = ~\P1_addr_reg[6]/NET0131  & n11723 ;
  assign n12711 = ~n2731 & ~n12709 ;
  assign n12712 = ~n12710 & n12711 ;
  assign n12713 = ~n11734 & ~n11735 ;
  assign n12715 = ~n11756 & n12713 ;
  assign n12714 = n11756 & ~n12713 ;
  assign n12716 = n11728 & ~n12714 ;
  assign n12717 = ~n12715 & n12716 ;
  assign n12723 = ~n12712 & ~n12717 ;
  assign n12724 = ~n12722 & n12723 ;
  assign n12725 = \P1_state_reg[0]/NET0131  & ~n12724 ;
  assign n12726 = ~n9769 & ~n12725 ;
  assign n12728 = ~n12165 & ~n12166 ;
  assign n12749 = ~n12209 & ~n12728 ;
  assign n12748 = n12209 & n12728 ;
  assign n12750 = n634 & ~n12748 ;
  assign n12751 = ~n12749 & n12750 ;
  assign n12733 = ~n12182 & ~n12194 ;
  assign n12745 = n12219 & n12733 ;
  assign n12744 = ~n12219 & ~n12733 ;
  assign n12746 = n2262 & ~n12744 ;
  assign n12747 = ~n12745 & n12746 ;
  assign n12743 = n615 & n907 ;
  assign n12752 = n2035 & ~n12743 ;
  assign n12753 = ~n12747 & n12752 ;
  assign n12754 = ~n12751 & n12753 ;
  assign n12735 = n12191 & n12733 ;
  assign n12734 = ~n12191 & ~n12733 ;
  assign n12736 = n11971 & ~n12734 ;
  assign n12737 = ~n12735 & n12736 ;
  assign n12730 = n12169 & ~n12728 ;
  assign n12729 = ~n12169 & n12728 ;
  assign n12731 = n2261 & ~n12729 ;
  assign n12732 = ~n12730 & n12731 ;
  assign n12738 = \P2_addr_reg[10]/NET0131  & n634 ;
  assign n12727 = n907 & n2262 ;
  assign n12739 = ~n2035 & ~n12727 ;
  assign n12740 = ~n12738 & n12739 ;
  assign n12741 = ~n12732 & n12740 ;
  assign n12742 = ~n12737 & n12741 ;
  assign n12755 = \P1_state_reg[0]/NET0131  & ~n12742 ;
  assign n12756 = ~n12754 & n12755 ;
  assign n12757 = ~n7484 & ~n12756 ;
  assign n12764 = ~n12181 & ~n12193 ;
  assign n12780 = n12221 & ~n12764 ;
  assign n12779 = ~n12221 & n12764 ;
  assign n12781 = n2262 & ~n12779 ;
  assign n12782 = ~n12780 & n12781 ;
  assign n12759 = ~n12163 & ~n12164 ;
  assign n12776 = ~n12211 & n12759 ;
  assign n12775 = n12211 & ~n12759 ;
  assign n12777 = n634 & ~n12775 ;
  assign n12778 = ~n12776 & n12777 ;
  assign n12774 = n615 & n880 ;
  assign n12783 = n2035 & ~n12774 ;
  assign n12784 = ~n12778 & n12783 ;
  assign n12785 = ~n12782 & n12784 ;
  assign n12761 = ~n12171 & n12759 ;
  assign n12760 = n12171 & ~n12759 ;
  assign n12762 = n2261 & ~n12760 ;
  assign n12763 = ~n12761 & n12762 ;
  assign n12766 = n12281 & n12764 ;
  assign n12765 = ~n12281 & ~n12764 ;
  assign n12767 = n11971 & ~n12765 ;
  assign n12768 = ~n12766 & n12767 ;
  assign n12769 = \P2_addr_reg[11]/NET0131  & n634 ;
  assign n12758 = n880 & n2262 ;
  assign n12770 = ~n2035 & ~n12758 ;
  assign n12771 = ~n12769 & n12770 ;
  assign n12772 = ~n12768 & n12771 ;
  assign n12773 = ~n12763 & n12772 ;
  assign n12786 = \P1_state_reg[0]/NET0131  & ~n12773 ;
  assign n12787 = ~n12785 & n12786 ;
  assign n12788 = ~n8115 & ~n12787 ;
  assign n12795 = ~n12365 & ~n12366 ;
  assign n12811 = ~n12456 & ~n12795 ;
  assign n12810 = n12456 & n12795 ;
  assign n12812 = n2262 & ~n12810 ;
  assign n12813 = ~n12811 & n12812 ;
  assign n12790 = ~n12352 & ~n12353 ;
  assign n12807 = n12444 & n12790 ;
  assign n12806 = ~n12444 & ~n12790 ;
  assign n12808 = n634 & ~n12806 ;
  assign n12809 = ~n12807 & n12808 ;
  assign n12805 = n615 & n758 ;
  assign n12814 = n2035 & ~n12805 ;
  assign n12815 = ~n12809 & n12814 ;
  assign n12816 = ~n12813 & n12815 ;
  assign n12792 = n12411 & n12790 ;
  assign n12791 = ~n12411 & ~n12790 ;
  assign n12793 = n2261 & ~n12791 ;
  assign n12794 = ~n12792 & n12793 ;
  assign n12797 = n12426 & n12795 ;
  assign n12796 = ~n12426 & ~n12795 ;
  assign n12798 = n11971 & ~n12796 ;
  assign n12799 = ~n12797 & n12798 ;
  assign n12800 = n758 & n2262 ;
  assign n12789 = \P2_addr_reg[14]/NET0131  & n634 ;
  assign n12801 = ~n2035 & ~n12789 ;
  assign n12802 = ~n12800 & n12801 ;
  assign n12803 = ~n12799 & n12802 ;
  assign n12804 = ~n12794 & n12803 ;
  assign n12817 = \P1_state_reg[0]/NET0131  & ~n12804 ;
  assign n12818 = ~n12816 & n12817 ;
  assign n12819 = ~n8156 & ~n12818 ;
  assign n12821 = ~n11940 & ~n11960 ;
  assign n12842 = ~n11957 & ~n12821 ;
  assign n12841 = n11957 & n12821 ;
  assign n12843 = n11971 & ~n12841 ;
  assign n12844 = ~n12842 & n12843 ;
  assign n12826 = ~n11902 & ~n11918 ;
  assign n12836 = ~n11917 & ~n11919 ;
  assign n12838 = n12826 & n12836 ;
  assign n12837 = ~n12826 & ~n12836 ;
  assign n12839 = n2261 & ~n12837 ;
  assign n12840 = ~n12838 & n12839 ;
  assign n12835 = ~n1048 & n2262 ;
  assign n12834 = \P2_addr_reg[5]/NET0131  & n634 ;
  assign n12845 = ~n2035 & ~n12834 ;
  assign n12846 = ~n12835 & n12845 ;
  assign n12847 = ~n12840 & n12846 ;
  assign n12848 = ~n12844 & n12847 ;
  assign n12828 = n12010 & ~n12826 ;
  assign n12827 = ~n12010 & n12826 ;
  assign n12829 = n634 & ~n12827 ;
  assign n12830 = ~n12828 & n12829 ;
  assign n12823 = ~n11989 & n12821 ;
  assign n12822 = n11989 & ~n12821 ;
  assign n12824 = n2262 & ~n12822 ;
  assign n12825 = ~n12823 & n12824 ;
  assign n12820 = n615 & ~n1048 ;
  assign n12831 = n2035 & ~n12820 ;
  assign n12832 = ~n12825 & n12831 ;
  assign n12833 = ~n12830 & n12832 ;
  assign n12849 = \P1_state_reg[0]/NET0131  & ~n12833 ;
  assign n12850 = ~n12848 & n12849 ;
  assign n12851 = ~n9151 & ~n12850 ;
  assign n12858 = ~n11898 & ~n11899 ;
  assign n12860 = n12014 & ~n12858 ;
  assign n12859 = ~n12014 & n12858 ;
  assign n12861 = n634 & ~n12859 ;
  assign n12862 = ~n12860 & n12861 ;
  assign n12853 = ~n11938 & ~n11966 ;
  assign n12855 = ~n11993 & n12853 ;
  assign n12854 = n11993 & ~n12853 ;
  assign n12856 = n2262 & ~n12854 ;
  assign n12857 = ~n12855 & n12856 ;
  assign n12852 = n615 & n1024 ;
  assign n12863 = n2035 & ~n12852 ;
  assign n12864 = ~n12857 & n12863 ;
  assign n12865 = ~n12862 & n12864 ;
  assign n12872 = n11963 & n12853 ;
  assign n12871 = ~n11963 & ~n12853 ;
  assign n12873 = n11971 & ~n12871 ;
  assign n12874 = ~n12872 & n12873 ;
  assign n12868 = ~n11924 & n12858 ;
  assign n12867 = n11924 & ~n12858 ;
  assign n12869 = n2261 & ~n12867 ;
  assign n12870 = ~n12868 & n12869 ;
  assign n12875 = n1024 & n2262 ;
  assign n12866 = \P2_addr_reg[7]/NET0131  & n634 ;
  assign n12876 = ~n2035 & ~n12866 ;
  assign n12877 = ~n12875 & n12876 ;
  assign n12878 = ~n12870 & n12877 ;
  assign n12879 = ~n12874 & n12878 ;
  assign n12880 = \P1_state_reg[0]/NET0131  & ~n12879 ;
  assign n12881 = ~n12865 & n12880 ;
  assign n12882 = ~n9236 & ~n12881 ;
  assign n12889 = ~n11937 & ~n11965 ;
  assign n12891 = n11995 & ~n12889 ;
  assign n12890 = ~n11995 & n12889 ;
  assign n12892 = n2262 & ~n12890 ;
  assign n12893 = ~n12891 & n12892 ;
  assign n12886 = ~n11928 & n12017 ;
  assign n12884 = ~n11897 & ~n11928 ;
  assign n12885 = n12016 & ~n12884 ;
  assign n12887 = n634 & ~n12885 ;
  assign n12888 = ~n12886 & n12887 ;
  assign n12883 = n615 & n956 ;
  assign n12894 = n2035 & ~n12883 ;
  assign n12895 = ~n12888 & n12894 ;
  assign n12896 = ~n12893 & n12895 ;
  assign n12903 = ~n11926 & n12884 ;
  assign n12902 = n11926 & ~n12884 ;
  assign n12904 = n2261 & ~n12902 ;
  assign n12905 = ~n12903 & n12904 ;
  assign n12899 = n12187 & n12889 ;
  assign n12898 = ~n12187 & ~n12889 ;
  assign n12900 = n11971 & ~n12898 ;
  assign n12901 = ~n12899 & n12900 ;
  assign n12906 = \P2_addr_reg[8]/NET0131  & n634 ;
  assign n12897 = n956 & n2262 ;
  assign n12907 = ~n2035 & ~n12897 ;
  assign n12908 = ~n12906 & n12907 ;
  assign n12909 = ~n12901 & n12908 ;
  assign n12910 = ~n12905 & n12909 ;
  assign n12911 = \P1_state_reg[0]/NET0131  & ~n12910 ;
  assign n12912 = ~n12896 & n12911 ;
  assign n12913 = ~n8274 & ~n12912 ;
  assign n12927 = ~n12471 & ~n12528 ;
  assign n12928 = ~n12472 & n12477 ;
  assign n12929 = n12927 & ~n12928 ;
  assign n12930 = ~n12529 & ~n12929 ;
  assign n12931 = ~\P2_reg1_reg[19]/NET0131  & ~n1297 ;
  assign n12932 = \P2_reg1_reg[19]/NET0131  & n1297 ;
  assign n12933 = ~n12931 & ~n12932 ;
  assign n12935 = ~n12930 & ~n12933 ;
  assign n12934 = n12930 & n12933 ;
  assign n12936 = n2261 & ~n12934 ;
  assign n12937 = ~n12935 & n12936 ;
  assign n12914 = ~n12482 & ~n12543 ;
  assign n12915 = ~n12483 & n12488 ;
  assign n12916 = n12914 & ~n12915 ;
  assign n12917 = ~n12544 & ~n12916 ;
  assign n12918 = ~\P2_reg2_reg[19]/NET0131  & ~n1297 ;
  assign n12919 = \P2_reg2_reg[19]/NET0131  & n1297 ;
  assign n12920 = ~n12918 & ~n12919 ;
  assign n12922 = ~n12917 & ~n12920 ;
  assign n12921 = n12917 & n12920 ;
  assign n12923 = n11971 & ~n12921 ;
  assign n12924 = ~n12922 & n12923 ;
  assign n12926 = \P2_addr_reg[19]/NET0131  & n634 ;
  assign n12925 = ~n1297 & n2262 ;
  assign n12938 = ~n2035 & ~n12925 ;
  assign n12939 = ~n12926 & n12938 ;
  assign n12940 = ~n12924 & n12939 ;
  assign n12941 = ~n12937 & n12940 ;
  assign n12952 = ~n12384 & n12474 ;
  assign n12953 = ~n12472 & n12504 ;
  assign n12954 = ~n12952 & n12953 ;
  assign n12955 = n12927 & ~n12954 ;
  assign n12956 = ~n12529 & ~n12955 ;
  assign n12958 = n12933 & ~n12956 ;
  assign n12957 = ~n12933 & n12956 ;
  assign n12959 = n634 & ~n12957 ;
  assign n12960 = ~n12958 & n12959 ;
  assign n12943 = ~n12392 & n12485 ;
  assign n12944 = ~n12483 & n12515 ;
  assign n12945 = ~n12943 & n12944 ;
  assign n12946 = n12914 & ~n12945 ;
  assign n12947 = ~n12544 & ~n12946 ;
  assign n12949 = n12920 & ~n12947 ;
  assign n12948 = ~n12920 & n12947 ;
  assign n12950 = n2262 & ~n12948 ;
  assign n12951 = ~n12949 & n12950 ;
  assign n12942 = n615 & ~n1297 ;
  assign n12961 = n2035 & ~n12942 ;
  assign n12962 = ~n12951 & n12961 ;
  assign n12963 = ~n12960 & n12962 ;
  assign n12964 = \P1_state_reg[0]/NET0131  & ~n12963 ;
  assign n12965 = ~n12941 & n12964 ;
  assign n12966 = ~n4304 & ~n12965 ;
  assign n12967 = ~\P1_state_reg[0]/NET0131  & ~\P2_reg3_reg[1]/NET0131  ;
  assign n12968 = n615 & ~n1138 ;
  assign n12979 = n2035 & ~n12968 ;
  assign n12969 = ~n11947 & ~n11948 ;
  assign n12970 = n11981 & ~n12969 ;
  assign n12971 = ~n11981 & n12969 ;
  assign n12972 = ~n12970 & ~n12971 ;
  assign n12973 = n2262 & n12972 ;
  assign n12974 = ~n11908 & ~n11909 ;
  assign n12975 = ~n12002 & n12974 ;
  assign n12976 = n12002 & ~n12974 ;
  assign n12977 = ~n12975 & ~n12976 ;
  assign n12978 = n634 & n12977 ;
  assign n12980 = ~n12973 & ~n12978 ;
  assign n12981 = n12979 & n12980 ;
  assign n12982 = \P2_addr_reg[1]/NET0131  & n634 ;
  assign n12992 = ~n2035 & ~n12982 ;
  assign n12988 = ~n11949 & n12969 ;
  assign n12989 = n11949 & ~n12969 ;
  assign n12990 = ~n12988 & ~n12989 ;
  assign n12991 = n11971 & n12990 ;
  assign n12983 = ~n1138 & n2262 ;
  assign n12984 = n11910 & ~n12974 ;
  assign n12985 = ~n11910 & n12974 ;
  assign n12986 = ~n12984 & ~n12985 ;
  assign n12987 = n2261 & n12986 ;
  assign n12993 = ~n12983 & ~n12987 ;
  assign n12994 = ~n12991 & n12993 ;
  assign n12995 = n12992 & n12994 ;
  assign n12996 = ~n12981 & ~n12995 ;
  assign n12997 = \P1_state_reg[0]/NET0131  & ~n12996 ;
  assign n12998 = ~n12967 & ~n12997 ;
  assign n13000 = ~n11904 & ~n11905 ;
  assign n13013 = ~n11914 & n13000 ;
  assign n13014 = n11914 & ~n13000 ;
  assign n13015 = ~n13013 & ~n13014 ;
  assign n13016 = n2261 & n13015 ;
  assign n13023 = ~n2035 & ~n13016 ;
  assign n13005 = ~n11943 & ~n11944 ;
  assign n13019 = n11953 & ~n13005 ;
  assign n13020 = ~n11953 & n13005 ;
  assign n13021 = ~n13019 & ~n13020 ;
  assign n13022 = n11971 & n13021 ;
  assign n13017 = \P2_addr_reg[3]/NET0131  & n634 ;
  assign n13018 = n1090 & n2262 ;
  assign n13024 = ~n13017 & ~n13018 ;
  assign n13025 = ~n13022 & n13024 ;
  assign n13026 = n13023 & n13025 ;
  assign n12999 = n615 & n1090 ;
  assign n13010 = n2035 & ~n12999 ;
  assign n13001 = n12006 & ~n13000 ;
  assign n13002 = ~n12006 & n13000 ;
  assign n13003 = ~n13001 & ~n13002 ;
  assign n13004 = n634 & n13003 ;
  assign n13006 = ~n11985 & n13005 ;
  assign n13007 = n11985 & ~n13005 ;
  assign n13008 = ~n13006 & ~n13007 ;
  assign n13009 = n2262 & n13008 ;
  assign n13011 = ~n13004 & ~n13009 ;
  assign n13012 = n13010 & n13011 ;
  assign n13027 = \P1_state_reg[0]/NET0131  & ~n13012 ;
  assign n13028 = ~n13026 & n13027 ;
  assign n13029 = ~n10395 & ~n13028 ;
  assign n13047 = \P1_reg1_reg[18]/NET0131  & n3621 ;
  assign n13048 = ~n12331 & ~n12339 ;
  assign n13049 = ~\P1_reg1_reg[18]/NET0131  & ~n3621 ;
  assign n13050 = ~n12330 & ~n13049 ;
  assign n13051 = ~n13048 & n13050 ;
  assign n13052 = ~n13047 & ~n13051 ;
  assign n13053 = \P1_reg1_reg[19]/NET0131  & n3566 ;
  assign n13054 = ~\P1_reg1_reg[19]/NET0131  & ~n3566 ;
  assign n13055 = ~n13053 & ~n13054 ;
  assign n13057 = ~n13052 & ~n13055 ;
  assign n13056 = n13052 & n13055 ;
  assign n13058 = n11728 & ~n13056 ;
  assign n13059 = ~n13057 & n13058 ;
  assign n13030 = \P1_reg2_reg[18]/NET0131  & n3621 ;
  assign n13031 = ~n12317 & ~n12321 ;
  assign n13032 = ~\P1_reg2_reg[18]/NET0131  & ~n3621 ;
  assign n13033 = ~n12316 & ~n13032 ;
  assign n13034 = ~n13031 & n13033 ;
  assign n13035 = ~n13030 & ~n13034 ;
  assign n13036 = \P1_reg2_reg[19]/NET0131  & n3566 ;
  assign n13037 = ~\P1_reg2_reg[19]/NET0131  & ~n3566 ;
  assign n13038 = ~n13036 & ~n13037 ;
  assign n13040 = ~n13035 & ~n13038 ;
  assign n13039 = n13035 & n13038 ;
  assign n13041 = n11686 & ~n13039 ;
  assign n13042 = ~n13040 & n13041 ;
  assign n13044 = n3566 & ~n11723 ;
  assign n13043 = ~\P1_addr_reg[19]/NET0131  & n11723 ;
  assign n13045 = ~n2731 & ~n13043 ;
  assign n13046 = ~n13044 & n13045 ;
  assign n13060 = ~n13042 & ~n13046 ;
  assign n13061 = ~n13059 & n13060 ;
  assign n13062 = \P1_state_reg[0]/NET0131  & ~n13061 ;
  assign n13063 = ~n6091 & ~n13062 ;
  assign n13077 = ~n13047 & ~n13049 ;
  assign n13078 = ~n12250 & n12254 ;
  assign n13079 = ~n12249 & ~n12331 ;
  assign n13080 = ~n13078 & n13079 ;
  assign n13081 = ~n12330 & ~n13080 ;
  assign n13083 = n13077 & n13081 ;
  assign n13082 = ~n13077 & ~n13081 ;
  assign n13084 = n11728 & ~n13082 ;
  assign n13085 = ~n13083 & n13084 ;
  assign n13064 = ~n13030 & ~n13032 ;
  assign n13065 = ~n12239 & n12244 ;
  assign n13066 = ~n12238 & ~n12317 ;
  assign n13067 = ~n13065 & n13066 ;
  assign n13068 = ~n12316 & ~n13067 ;
  assign n13070 = n13064 & n13068 ;
  assign n13069 = ~n13064 & ~n13068 ;
  assign n13071 = n11686 & ~n13069 ;
  assign n13072 = ~n13070 & n13071 ;
  assign n13074 = ~n3621 & ~n11723 ;
  assign n13073 = ~\P1_addr_reg[18]/NET0131  & n11723 ;
  assign n13075 = ~n2731 & ~n13073 ;
  assign n13076 = ~n13074 & n13075 ;
  assign n13086 = ~n13072 & ~n13076 ;
  assign n13087 = ~n13085 & n13086 ;
  assign n13088 = \P1_state_reg[0]/NET0131  & ~n13087 ;
  assign n13089 = ~n5955 & ~n13088 ;
  assign n13090 = ~\P1_state_reg[0]/NET0131  & ~\P2_reg3_reg[2]/NET0131  ;
  assign n13091 = n615 & ~n1122 ;
  assign n13102 = n2035 & ~n13091 ;
  assign n13092 = ~n11945 & ~n11946 ;
  assign n13093 = n11983 & ~n13092 ;
  assign n13094 = ~n11983 & n13092 ;
  assign n13095 = ~n13093 & ~n13094 ;
  assign n13096 = n2262 & n13095 ;
  assign n13097 = ~n11906 & ~n11907 ;
  assign n13098 = ~n12004 & n13097 ;
  assign n13099 = n12004 & ~n13097 ;
  assign n13100 = ~n13098 & ~n13099 ;
  assign n13101 = n634 & n13100 ;
  assign n13103 = ~n13096 & ~n13101 ;
  assign n13104 = n13102 & n13103 ;
  assign n13105 = \P2_addr_reg[2]/NET0131  & n634 ;
  assign n13115 = ~n2035 & ~n13105 ;
  assign n13111 = ~n11912 & n13097 ;
  assign n13112 = n11912 & ~n13097 ;
  assign n13113 = ~n13111 & ~n13112 ;
  assign n13114 = n2261 & n13113 ;
  assign n13106 = ~n1122 & n2262 ;
  assign n13107 = n11951 & ~n13092 ;
  assign n13108 = ~n11951 & n13092 ;
  assign n13109 = ~n13107 & ~n13108 ;
  assign n13110 = n11971 & n13109 ;
  assign n13116 = ~n13106 & ~n13110 ;
  assign n13117 = ~n13114 & n13116 ;
  assign n13118 = n13115 & n13117 ;
  assign n13119 = ~n13104 & ~n13118 ;
  assign n13120 = \P1_state_reg[0]/NET0131  & ~n13119 ;
  assign n13121 = ~n13090 & ~n13120 ;
  assign n13136 = \P2_addr_reg[4]/NET0131  & n634 ;
  assign n13146 = ~n2035 & ~n13136 ;
  assign n13128 = ~n11903 & ~n11919 ;
  assign n13142 = ~n11916 & n13128 ;
  assign n13143 = n11916 & ~n13128 ;
  assign n13144 = ~n13142 & ~n13143 ;
  assign n13145 = n2261 & n13144 ;
  assign n13123 = ~n11941 & ~n11942 ;
  assign n13137 = ~n11955 & ~n13123 ;
  assign n13138 = n11955 & n13123 ;
  assign n13139 = ~n13137 & ~n13138 ;
  assign n13140 = n11971 & n13139 ;
  assign n13141 = n1074 & n2262 ;
  assign n13147 = ~n13140 & ~n13141 ;
  assign n13148 = ~n13145 & n13147 ;
  assign n13149 = n13146 & n13148 ;
  assign n13122 = n615 & n1074 ;
  assign n13133 = n2035 & ~n13122 ;
  assign n13124 = n11987 & ~n13123 ;
  assign n13125 = ~n11987 & n13123 ;
  assign n13126 = ~n13124 & ~n13125 ;
  assign n13127 = n2262 & n13126 ;
  assign n13129 = ~n12008 & n13128 ;
  assign n13130 = n12008 & ~n13128 ;
  assign n13131 = ~n13129 & ~n13130 ;
  assign n13132 = n634 & n13131 ;
  assign n13134 = ~n13127 & ~n13132 ;
  assign n13135 = n13133 & n13134 ;
  assign n13150 = \P1_state_reg[0]/NET0131  & ~n13135 ;
  assign n13151 = ~n13149 & n13150 ;
  assign n13152 = ~n9849 & ~n13151 ;
  assign n13153 = ~n2732 & ~n4081 ;
  assign n13154 = \P1_state_reg[0]/NET0131  & ~n13153 ;
  assign n13155 = ~n634 & ~n2035 ;
  assign n13156 = \P1_state_reg[0]/NET0131  & ~n13155 ;
  assign n13157 = \P1_state_reg[0]/NET0131  & n4081 ;
  assign n13158 = \P1_state_reg[0]/NET0131  & n2035 ;
  assign n13159 = \P1_reg2_reg[22]/NET0131  & ~n9331 ;
  assign n13161 = \P1_reg2_reg[22]/NET0131  & ~n2717 ;
  assign n13162 = n2717 & ~n6412 ;
  assign n13163 = ~n13161 & ~n13162 ;
  assign n13164 = n3969 & ~n13163 ;
  assign n13171 = n2717 & n6419 ;
  assign n13172 = ~n13161 & ~n13171 ;
  assign n13173 = n4062 & ~n13172 ;
  assign n13160 = n3149 & n4073 ;
  assign n13174 = n2717 & n3143 ;
  assign n13175 = ~n13161 & ~n13174 ;
  assign n13176 = n4028 & ~n13175 ;
  assign n13177 = ~n13160 & ~n13176 ;
  assign n13178 = ~n13173 & n13177 ;
  assign n13179 = ~n13164 & n13178 ;
  assign n13165 = n2717 & ~n6400 ;
  assign n13166 = ~n13161 & ~n13165 ;
  assign n13167 = n3829 & ~n13166 ;
  assign n13168 = n2717 & n6388 ;
  assign n13169 = ~n13161 & ~n13168 ;
  assign n13170 = n4025 & ~n13169 ;
  assign n13180 = ~n13167 & ~n13170 ;
  assign n13181 = n13179 & n13180 ;
  assign n13182 = n9331 & ~n13181 ;
  assign n13183 = ~n13159 & ~n13182 ;
  assign n13184 = \P2_reg2_reg[26]/NET0131  & ~n2286 ;
  assign n13185 = \P2_reg2_reg[26]/NET0131  & n2035 ;
  assign n13186 = \P2_reg2_reg[26]/NET0131  & ~n2310 ;
  assign n13187 = ~n5778 & ~n13186 ;
  assign n13188 = n2314 & ~n13187 ;
  assign n13189 = n2310 & ~n5570 ;
  assign n13190 = ~n13186 & ~n13189 ;
  assign n13191 = n1790 & ~n13190 ;
  assign n13192 = n1573 & n2394 ;
  assign n13193 = ~n1583 & n1854 ;
  assign n13194 = \P2_reg2_reg[26]/NET0131  & ~n2407 ;
  assign n13201 = ~n13193 & ~n13194 ;
  assign n13202 = ~n13192 & n13201 ;
  assign n13203 = ~n13191 & n13202 ;
  assign n13204 = ~n13188 & n13203 ;
  assign n13195 = \P2_reg2_reg[26]/NET0131  & ~n2291 ;
  assign n13196 = ~n5787 & ~n13195 ;
  assign n13197 = ~n2290 & ~n13196 ;
  assign n13198 = n2291 & ~n5562 ;
  assign n13199 = ~n13195 & ~n13198 ;
  assign n13200 = ~n2392 & ~n13199 ;
  assign n13205 = ~n13197 & ~n13200 ;
  assign n13206 = n13204 & n13205 ;
  assign n13207 = n2037 & ~n13206 ;
  assign n13208 = ~n13185 & ~n13207 ;
  assign n13209 = \P1_state_reg[0]/NET0131  & ~n13208 ;
  assign n13210 = ~n13184 & ~n13209 ;
  assign n13211 = ~\P1_rd_reg/NET0131  & ~\P2_rd_reg/NET0131  ;
  assign n13212 = \P1_rd_reg/NET0131  & \P2_rd_reg/NET0131  ;
  assign n13213 = ~n13211 & ~n13212 ;
  assign n13214 = \P1_addr_reg[0]/NET0131  & \P2_addr_reg[0]/NET0131  ;
  assign n13215 = ~\P1_addr_reg[0]/NET0131  & ~\P2_addr_reg[0]/NET0131  ;
  assign n13216 = ~n13214 & ~n13215 ;
  assign n13217 = \P1_addr_reg[10]/NET0131  & \P2_addr_reg[10]/NET0131  ;
  assign n13218 = ~\P1_addr_reg[10]/NET0131  & ~\P2_addr_reg[10]/NET0131  ;
  assign n13219 = ~n13217 & ~n13218 ;
  assign n13220 = ~\P1_addr_reg[9]/NET0131  & ~\P2_addr_reg[9]/NET0131  ;
  assign n13221 = \P1_addr_reg[9]/NET0131  & \P2_addr_reg[9]/NET0131  ;
  assign n13222 = ~\P1_addr_reg[8]/NET0131  & ~\P2_addr_reg[8]/NET0131  ;
  assign n13223 = \P1_addr_reg[8]/NET0131  & \P2_addr_reg[8]/NET0131  ;
  assign n13224 = ~\P1_addr_reg[7]/NET0131  & ~\P2_addr_reg[7]/NET0131  ;
  assign n13225 = \P1_addr_reg[7]/NET0131  & \P2_addr_reg[7]/NET0131  ;
  assign n13226 = ~\P1_addr_reg[6]/NET0131  & ~\P2_addr_reg[6]/NET0131  ;
  assign n13227 = \P1_addr_reg[6]/NET0131  & \P2_addr_reg[6]/NET0131  ;
  assign n13228 = ~\P1_addr_reg[5]/NET0131  & ~\P2_addr_reg[5]/NET0131  ;
  assign n13229 = \P1_addr_reg[5]/NET0131  & \P2_addr_reg[5]/NET0131  ;
  assign n13230 = ~\P1_addr_reg[4]/NET0131  & ~\P2_addr_reg[4]/NET0131  ;
  assign n13231 = \P1_addr_reg[4]/NET0131  & \P2_addr_reg[4]/NET0131  ;
  assign n13232 = ~\P1_addr_reg[3]/NET0131  & ~\P2_addr_reg[3]/NET0131  ;
  assign n13233 = \P1_addr_reg[3]/NET0131  & \P2_addr_reg[3]/NET0131  ;
  assign n13234 = ~\P1_addr_reg[2]/NET0131  & ~\P2_addr_reg[2]/NET0131  ;
  assign n13235 = \P1_addr_reg[2]/NET0131  & \P2_addr_reg[2]/NET0131  ;
  assign n13236 = ~\P1_addr_reg[1]/NET0131  & ~\P2_addr_reg[1]/NET0131  ;
  assign n13237 = \P1_addr_reg[1]/NET0131  & \P2_addr_reg[1]/NET0131  ;
  assign n13238 = ~n13214 & ~n13237 ;
  assign n13239 = ~n13236 & ~n13238 ;
  assign n13240 = ~n13235 & ~n13239 ;
  assign n13241 = ~n13234 & ~n13240 ;
  assign n13242 = ~n13233 & ~n13241 ;
  assign n13243 = ~n13232 & ~n13242 ;
  assign n13244 = ~n13231 & ~n13243 ;
  assign n13245 = ~n13230 & ~n13244 ;
  assign n13246 = ~n13229 & ~n13245 ;
  assign n13247 = ~n13228 & ~n13246 ;
  assign n13248 = ~n13227 & ~n13247 ;
  assign n13249 = ~n13226 & ~n13248 ;
  assign n13250 = ~n13225 & ~n13249 ;
  assign n13251 = ~n13224 & ~n13250 ;
  assign n13252 = ~n13223 & ~n13251 ;
  assign n13253 = ~n13222 & ~n13252 ;
  assign n13254 = ~n13221 & ~n13253 ;
  assign n13255 = ~n13220 & ~n13254 ;
  assign n13256 = ~n13219 & n13255 ;
  assign n13257 = n13219 & ~n13255 ;
  assign n13258 = ~n13256 & ~n13257 ;
  assign n13259 = \P1_addr_reg[11]/NET0131  & \P2_addr_reg[11]/NET0131  ;
  assign n13260 = ~\P1_addr_reg[11]/NET0131  & ~\P2_addr_reg[11]/NET0131  ;
  assign n13261 = ~n13259 & ~n13260 ;
  assign n13262 = ~n13217 & ~n13255 ;
  assign n13263 = ~n13218 & ~n13262 ;
  assign n13264 = ~n13261 & n13263 ;
  assign n13265 = n13261 & ~n13263 ;
  assign n13266 = ~n13264 & ~n13265 ;
  assign n13267 = \P1_addr_reg[12]/NET0131  & \P2_addr_reg[12]/NET0131  ;
  assign n13268 = ~\P1_addr_reg[12]/NET0131  & ~\P2_addr_reg[12]/NET0131  ;
  assign n13269 = ~n13267 & ~n13268 ;
  assign n13270 = ~n13259 & ~n13263 ;
  assign n13271 = ~n13260 & ~n13270 ;
  assign n13272 = ~n13269 & n13271 ;
  assign n13273 = n13269 & ~n13271 ;
  assign n13274 = ~n13272 & ~n13273 ;
  assign n13275 = \P1_addr_reg[13]/NET0131  & \P2_addr_reg[13]/NET0131  ;
  assign n13276 = ~\P1_addr_reg[13]/NET0131  & ~\P2_addr_reg[13]/NET0131  ;
  assign n13277 = ~n13275 & ~n13276 ;
  assign n13278 = ~n13267 & ~n13271 ;
  assign n13279 = ~n13268 & ~n13278 ;
  assign n13280 = ~n13277 & n13279 ;
  assign n13281 = n13277 & ~n13279 ;
  assign n13282 = ~n13280 & ~n13281 ;
  assign n13283 = \P1_addr_reg[14]/NET0131  & \P2_addr_reg[14]/NET0131  ;
  assign n13284 = ~\P1_addr_reg[14]/NET0131  & ~\P2_addr_reg[14]/NET0131  ;
  assign n13285 = ~n13283 & ~n13284 ;
  assign n13286 = ~n13275 & ~n13279 ;
  assign n13287 = ~n13276 & ~n13286 ;
  assign n13288 = ~n13285 & n13287 ;
  assign n13289 = n13285 & ~n13287 ;
  assign n13290 = ~n13288 & ~n13289 ;
  assign n13291 = \P1_addr_reg[15]/NET0131  & \P2_addr_reg[15]/NET0131  ;
  assign n13292 = ~\P1_addr_reg[15]/NET0131  & ~\P2_addr_reg[15]/NET0131  ;
  assign n13293 = ~n13291 & ~n13292 ;
  assign n13294 = ~n13283 & ~n13287 ;
  assign n13295 = ~n13284 & ~n13294 ;
  assign n13296 = ~n13293 & n13295 ;
  assign n13297 = n13293 & ~n13295 ;
  assign n13298 = ~n13296 & ~n13297 ;
  assign n13299 = \P1_addr_reg[16]/NET0131  & \P2_addr_reg[16]/NET0131  ;
  assign n13300 = ~\P1_addr_reg[16]/NET0131  & ~\P2_addr_reg[16]/NET0131  ;
  assign n13301 = ~n13299 & ~n13300 ;
  assign n13302 = ~n13291 & ~n13295 ;
  assign n13303 = ~n13292 & ~n13302 ;
  assign n13304 = ~n13301 & n13303 ;
  assign n13305 = n13301 & ~n13303 ;
  assign n13306 = ~n13304 & ~n13305 ;
  assign n13307 = \P1_addr_reg[17]/NET0131  & \P2_addr_reg[17]/NET0131  ;
  assign n13308 = ~\P1_addr_reg[17]/NET0131  & ~\P2_addr_reg[17]/NET0131  ;
  assign n13309 = ~n13307 & ~n13308 ;
  assign n13310 = ~n13299 & ~n13303 ;
  assign n13311 = ~n13300 & ~n13310 ;
  assign n13312 = ~n13309 & n13311 ;
  assign n13313 = n13309 & ~n13311 ;
  assign n13314 = ~n13312 & ~n13313 ;
  assign n13315 = \P1_addr_reg[18]/NET0131  & \P2_addr_reg[18]/NET0131  ;
  assign n13316 = ~\P1_addr_reg[18]/NET0131  & ~\P2_addr_reg[18]/NET0131  ;
  assign n13317 = ~n13315 & ~n13316 ;
  assign n13318 = ~n13307 & ~n13311 ;
  assign n13319 = ~n13308 & ~n13318 ;
  assign n13320 = ~n13317 & n13319 ;
  assign n13321 = n13317 & ~n13319 ;
  assign n13322 = ~n13320 & ~n13321 ;
  assign n13323 = ~n635 & ~n637 ;
  assign n13324 = ~n13315 & ~n13319 ;
  assign n13325 = ~n13316 & ~n13324 ;
  assign n13326 = n13323 & ~n13325 ;
  assign n13327 = ~n13323 & n13325 ;
  assign n13328 = ~n13326 & ~n13327 ;
  assign n13329 = ~n13236 & ~n13237 ;
  assign n13330 = n13214 & ~n13329 ;
  assign n13331 = ~n13214 & n13329 ;
  assign n13332 = ~n13330 & ~n13331 ;
  assign n13333 = ~n13234 & ~n13235 ;
  assign n13334 = n13239 & ~n13333 ;
  assign n13335 = ~n13239 & n13333 ;
  assign n13336 = ~n13334 & ~n13335 ;
  assign n13337 = ~n13232 & ~n13233 ;
  assign n13338 = n13241 & ~n13337 ;
  assign n13339 = ~n13241 & n13337 ;
  assign n13340 = ~n13338 & ~n13339 ;
  assign n13341 = ~n13230 & ~n13231 ;
  assign n13342 = n13243 & ~n13341 ;
  assign n13343 = ~n13243 & n13341 ;
  assign n13344 = ~n13342 & ~n13343 ;
  assign n13345 = ~n13228 & ~n13229 ;
  assign n13346 = n13245 & ~n13345 ;
  assign n13347 = ~n13245 & n13345 ;
  assign n13348 = ~n13346 & ~n13347 ;
  assign n13349 = ~n13226 & ~n13227 ;
  assign n13350 = n13247 & ~n13349 ;
  assign n13351 = ~n13247 & n13349 ;
  assign n13352 = ~n13350 & ~n13351 ;
  assign n13353 = ~n13224 & ~n13225 ;
  assign n13354 = n13249 & ~n13353 ;
  assign n13355 = ~n13249 & n13353 ;
  assign n13356 = ~n13354 & ~n13355 ;
  assign n13357 = ~n13222 & ~n13223 ;
  assign n13358 = n13251 & ~n13357 ;
  assign n13359 = ~n13251 & n13357 ;
  assign n13360 = ~n13358 & ~n13359 ;
  assign n13361 = ~n13220 & ~n13221 ;
  assign n13362 = n13253 & ~n13361 ;
  assign n13363 = ~n13253 & n13361 ;
  assign n13364 = ~n13362 & ~n13363 ;
  assign n13365 = ~\P1_wr_reg/NET0131  & ~\P2_wr_reg/NET0131  ;
  assign n13366 = \P1_wr_reg/NET0131  & \P2_wr_reg/NET0131  ;
  assign n13367 = ~n13365 & ~n13366 ;
  assign \P1_state_reg[0]/NET0131_syn_2  = ~\P1_state_reg[0]/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g35/_0_  = ~n523 ;
  assign \g73637/_0_  = ~n2017 ;
  assign \g73647/_0_  = ~n2285 ;
  assign \g73648/_0_  = ~n2419 ;
  assign \g73649/_0_  = ~n2448 ;
  assign \g73650/_0_  = ~n2477 ;
  assign \g73667/_0_  = ~n2527 ;
  assign \g73668/_0_  = ~n2556 ;
  assign \g73669/_0_  = ~n2669 ;
  assign \g73670/_0_  = ~n4087 ;
  assign \g73671/_0_  = ~n4117 ;
  assign \g73672/_0_  = ~n4174 ;
  assign \g73674/_0_  = ~n4201 ;
  assign \g73675/_0_  = ~n4229 ;
  assign \g73709/_0_  = ~n4302 ;
  assign \g73710/_0_  = ~n4343 ;
  assign \g73711/_0_  = ~n4387 ;
  assign \g73716/_0_  = ~n4447 ;
  assign \g73717/_0_  = ~n4556 ;
  assign \g73718/_0_  = ~n4586 ;
  assign \g73719/_0_  = ~n4611 ;
  assign \g73720/_0_  = ~n4637 ;
  assign \g73721/_0_  = ~n4818 ;
  assign \g73722/_0_  = ~n4843 ;
  assign \g73723/_0_  = ~n4868 ;
  assign \g73724/_0_  = ~n4897 ;
  assign \g73765/_0_  = ~n4937 ;
  assign \g73769/_0_  = ~n5044 ;
  assign \g73770/_0_  = ~n5104 ;
  assign \g73771/_0_  = ~n5167 ;
  assign \g73772/_0_  = ~n5197 ;
  assign \g73773/_0_  = ~n5227 ;
  assign \g73774/_0_  = ~n5257 ;
  assign \g73775/_0_  = ~n5286 ;
  assign \g73776/_0_  = ~n5494 ;
  assign \g73777/_0_  = ~n5520 ;
  assign \g73778/_0_  = ~n5549 ;
  assign \g73779/_0_  = ~n5605 ;
  assign \g73780/_0_  = ~n5646 ;
  assign \g73781/_0_  = ~n5672 ;
  assign \g73782/_0_  = ~n5698 ;
  assign \g73783/_0_  = ~n5723 ;
  assign \g73784/_0_  = ~n5749 ;
  assign \g73785/_0_  = ~n5774 ;
  assign \g73786/_0_  = ~n5801 ;
  assign \g73787/_0_  = ~n5826 ;
  assign \g73788/_0_  = ~n5853 ;
  assign \g73789/_0_  = ~n5879 ;
  assign \g73790/_0_  = ~n5901 ;
  assign \g73791/_0_  = ~n5927 ;
  assign \g73792/_0_  = ~n5953 ;
  assign \g73845/_0_  = ~n6002 ;
  assign \g73846/_0_  = ~n6049 ;
  assign \g73847/_0_  = ~n6094 ;
  assign \g73848/_0_  = ~n6136 ;
  assign \g73860/_0_  = ~n6162 ;
  assign \g73863/_0_  = ~n6194 ;
  assign \g73864/_0_  = ~n6248 ;
  assign \g73867/_0_  = ~n6277 ;
  assign \g73870/_0_  = ~n6305 ;
  assign \g73871/_0_  = ~n6330 ;
  assign \g73872/_0_  = ~n6354 ;
  assign \g73873/_0_  = ~n6379 ;
  assign \g73874/_0_  = ~n6431 ;
  assign \g73875/_0_  = ~n6457 ;
  assign \g73876/_0_  = ~n6479 ;
  assign \g73877/_0_  = ~n6503 ;
  assign \g73878/_0_  = ~n6531 ;
  assign \g73879/_0_  = ~n6557 ;
  assign \g73880/_0_  = ~n6579 ;
  assign \g73924/_0_  = ~n6624 ;
  assign \g73925/_0_  = ~n6666 ;
  assign \g73949/_0_  = ~n6711 ;
  assign \g73950/_0_  = ~n6751 ;
  assign \g73953/_0_  = ~n6775 ;
  assign \g73954/_0_  = ~n6799 ;
  assign \g73955/_0_  = ~n6828 ;
  assign \g73956/_0_  = ~n6852 ;
  assign \g73957/_0_  = ~n6881 ;
  assign \g73958/_0_  = ~n6907 ;
  assign \g73960/_0_  = ~n6932 ;
  assign \g73961/_0_  = ~n6953 ;
  assign \g73962/_0_  = ~n6978 ;
  assign \g73963/_0_  = ~n7003 ;
  assign \g73964/_0_  = ~n7028 ;
  assign \g73965/_0_  = ~n7053 ;
  assign \g73966/_0_  = ~n7081 ;
  assign \g73967/_0_  = ~n7106 ;
  assign \g73968/_0_  = ~n7131 ;
  assign \g73969/_0_  = ~n7156 ;
  assign \g73970/_0_  = ~n7181 ;
  assign \g73971/_0_  = ~n7206 ;
  assign \g73972/_0_  = ~n7229 ;
  assign \g73973/_0_  = ~n7251 ;
  assign \g73974/_0_  = ~n7273 ;
  assign \g73975/_0_  = ~n7293 ;
  assign \g73976/_0_  = ~n7314 ;
  assign \g73977/_0_  = ~n7336 ;
  assign \g73978/_0_  = ~n7358 ;
  assign \g73979/_0_  = ~n7380 ;
  assign \g73980/_0_  = ~n7400 ;
  assign \g74062/_0_  = ~n7443 ;
  assign \g74063/_0_  = ~n7483 ;
  assign \g74064/_0_  = ~n7526 ;
  assign \g74065/_0_  = ~n7566 ;
  assign \g74066/_0_  = ~n7607 ;
  assign \g74071/_0_  = ~n7648 ;
  assign \g74072/_0_  = ~n7688 ;
  assign \g74105/_0_  = ~n7744 ;
  assign \g74106/_0_  = ~n7773 ;
  assign \g74107/_0_  = ~n7802 ;
  assign \g74108/_0_  = ~n7827 ;
  assign \g74109/_0_  = ~n7850 ;
  assign \g74110/_0_  = ~n7875 ;
  assign \g74111/_0_  = ~n7898 ;
  assign \g74112/_0_  = ~n7920 ;
  assign \g74113/_0_  = ~n7942 ;
  assign \g74114/_0_  = ~n7964 ;
  assign \g74115/_0_  = ~n7990 ;
  assign \g74167/_0_  = ~n8030 ;
  assign \g74168/_0_  = ~n8073 ;
  assign \g74169/_0_  = ~n8114 ;
  assign \g74170/_0_  = ~n8154 ;
  assign \g74172/_0_  = ~n8195 ;
  assign \g74173/_0_  = ~n8235 ;
  assign \g74174/_0_  = ~n8273 ;
  assign \g74175/_0_  = ~n8313 ;
  assign \g74225/_0_  = ~n8342 ;
  assign \g74226/_0_  = ~n8368 ;
  assign \g74227/_0_  = ~n8397 ;
  assign \g74229/_0_  = ~n8422 ;
  assign \g74230/_0_  = ~n8448 ;
  assign \g74231/_0_  = ~n8474 ;
  assign \g74232/_0_  = ~n8498 ;
  assign \g74233/_0_  = ~n8526 ;
  assign \g74234/_0_  = ~n8554 ;
  assign \g74235/_0_  = ~n8582 ;
  assign \g74236/_0_  = ~n8609 ;
  assign \g74237/_0_  = ~n8630 ;
  assign \g74238/_0_  = ~n8657 ;
  assign \g74239/_0_  = ~n8684 ;
  assign \g74240/_0_  = ~n8711 ;
  assign \g74241/_0_  = ~n8738 ;
  assign \g74242/_0_  = ~n8765 ;
  assign \g74243/_0_  = ~n8791 ;
  assign \g74244/_0_  = ~n8818 ;
  assign \g74245/_0_  = ~n8840 ;
  assign \g74246/_0_  = ~n8862 ;
  assign \g74247/_0_  = ~n8879 ;
  assign \g74248/_0_  = ~n8905 ;
  assign \g74249/_0_  = ~n8931 ;
  assign \g74250/_0_  = ~n8953 ;
  assign \g74251/_0_  = ~n8975 ;
  assign \g74252/_0_  = ~n9000 ;
  assign \g74253/_0_  = ~n9025 ;
  assign \g74254/_0_  = ~n9050 ;
  assign \g74255/_0_  = ~n9067 ;
  assign \g74330/_0_  = ~n9108 ;
  assign \g74331/_0_  = ~n9150 ;
  assign \g74333/_0_  = ~n9194 ;
  assign \g74334/_0_  = ~n9235 ;
  assign \g74335/_0_  = ~n9275 ;
  assign \g74390/_0_  = ~n9302 ;
  assign \g74391/_0_  = ~n9328 ;
  assign \g74405/_0_  = n9348 ;
  assign \g74407/_0_  = ~n9374 ;
  assign \g74408/_0_  = n9386 ;
  assign \g74409/_0_  = ~n9412 ;
  assign \g74410/_0_  = ~n9436 ;
  assign \g74411/_0_  = ~n9460 ;
  assign \g74412/_0_  = ~n9487 ;
  assign \g74413/_0_  = ~n9515 ;
  assign \g74414/_0_  = ~n9542 ;
  assign \g74415/_0_  = ~n9569 ;
  assign \g74416/_0_  = ~n9596 ;
  assign \g74417/_0_  = ~n9623 ;
  assign \g74418/_0_  = ~n9645 ;
  assign \g74419/_0_  = n9654 ;
  assign \g74420/_0_  = ~n9676 ;
  assign \g74421/_0_  = ~n9701 ;
  assign \g74422/_0_  = ~n9726 ;
  assign \g74483/_0_  = ~n9768 ;
  assign \g74485/_0_  = ~n9809 ;
  assign \g74486/_0_  = ~n9848 ;
  assign \g74487/_0_  = ~n9888 ;
  assign \g74576/_0_  = ~n9914 ;
  assign \g74578/_0_  = ~n9936 ;
  assign \g74581/_0_  = ~n9962 ;
  assign \g74582/_0_  = ~n9988 ;
  assign \g74583/_0_  = ~n10014 ;
  assign \g74584/_0_  = ~n10040 ;
  assign \g74585/_0_  = ~n10068 ;
  assign \g74588/_0_  = ~n10095 ;
  assign \g74589/_0_  = ~n10122 ;
  assign \g74590/_0_  = ~n10149 ;
  assign \g74591/_0_  = ~n10176 ;
  assign \g74592/_0_  = ~n10198 ;
  assign \g74595/_0_  = ~n10225 ;
  assign \g74596/_0_  = ~n10252 ;
  assign \g74597/_0_  = ~n10279 ;
  assign \g74598/_0_  = ~n10306 ;
  assign \g74599/_0_  = ~n10328 ;
  assign \g74600/_0_  = ~n10350 ;
  assign \g74601/_0_  = ~n10372 ;
  assign \g74602/_0_  = ~n10394 ;
  assign \g74711/_0_  = ~n10435 ;
  assign \g74835/_0_  = ~n10459 ;
  assign \g74836/_0_  = ~n10483 ;
  assign \g74838/_0_  = ~n10507 ;
  assign \g74840/_0_  = ~n10536 ;
  assign \g74841/_0_  = ~n10560 ;
  assign \g74843/_0_  = ~n10582 ;
  assign \g74844/_0_  = ~n10604 ;
  assign \g74963/_0_  = ~n10642 ;
  assign \g75075/_0_  = ~n10668 ;
  assign \g75078/_0_  = ~n10695 ;
  assign \g75079/_0_  = ~n10721 ;
  assign \g75083/_0_  = ~n10748 ;
  assign \g75084/_0_  = ~n10775 ;
  assign \g75089/_0_  = ~n10802 ;
  assign \g75090/_0_  = ~n10829 ;
  assign \g75091/_0_  = ~n10855 ;
  assign \g75224/_0_  = ~n10896 ;
  assign \g75233/_0_  = ~n10938 ;
  assign \g75234/_0_  = ~n10977 ;
  assign \g75427/_0_  = ~n11003 ;
  assign \g75430/_0_  = ~n11029 ;
  assign \g75434/_0_  = ~n11057 ;
  assign \g75436/_0_  = ~n11084 ;
  assign \g75438/_0_  = ~n11110 ;
  assign \g75844/_0_  = ~n11137 ;
  assign \g75850/_0_  = ~n11166 ;
  assign \g75851/_0_  = ~n11194 ;
  assign \g75860/_0_  = ~n11223 ;
  assign \g75865/_0_  = ~n11243 ;
  assign \g75867/_0_  = ~n11267 ;
  assign \g76076/_0_  = ~n11297 ;
  assign \g76375/_0_  = ~n11321 ;
  assign \g76896/_0_  = ~n11346 ;
  assign \g76901/_0_  = ~n11370 ;
  assign \g76905/_0_  = ~n11393 ;
  assign \g77085/_0_  = ~n11409 ;
  assign \g77892/_0_  = ~n11418 ;
  assign \g77897/_0_  = ~n11424 ;
  assign \g77902/_0_  = ~n11429 ;
  assign \g78635/_0_  = ~n11447 ;
  assign \g78636/_0_  = ~n11455 ;
  assign \g78640/_0_  = ~n11465 ;
  assign \g78642/_0_  = ~n11480 ;
  assign \g78645/_0_  = ~n11485 ;
  assign \g78964/_0_  = ~n11492 ;
  assign \g83163/_3_  = ~n11495 ;
  assign \g83164/_3_  = n11498 ;
  assign \g83165/_3_  = n11501 ;
  assign \g83166/_3_  = ~n11504 ;
  assign \g83167/_3_  = ~n11507 ;
  assign \g83168/_3_  = ~n11510 ;
  assign \g83644/_0_  = ~n11518 ;
  assign \g83645/_0_  = ~n11521 ;
  assign \g83646/_0_  = n11523 ;
  assign \g83647/_0_  = ~n11526 ;
  assign \g83648/_0_  = ~n11529 ;
  assign \g83649/_0_  = ~n11532 ;
  assign \g83650/_0_  = ~n11535 ;
  assign \g83651/_0_  = ~n11538 ;
  assign \g83652/_0_  = ~n11541 ;
  assign \g83653/_0_  = ~n11544 ;
  assign \g83654/_0_  = ~n11547 ;
  assign \g83655/_0_  = ~n11550 ;
  assign \g83656/_0_  = ~n11553 ;
  assign \g83657/_0_  = n11556 ;
  assign \g83658/_0_  = n11559 ;
  assign \g83659/_0_  = ~n11562 ;
  assign \g83660/_0_  = ~n11565 ;
  assign \g83661/_0_  = ~n11568 ;
  assign \g83662/_0_  = ~n11571 ;
  assign \g83663/_0_  = ~n11574 ;
  assign \g83664/_0_  = ~n11577 ;
  assign \g83665/_0_  = ~n11580 ;
  assign \g83666/_0_  = ~n11583 ;
  assign \g83667/_3_  = ~n11586 ;
  assign \g83668/_0_  = ~n11589 ;
  assign \g83669/_0_  = ~n11592 ;
  assign \g83670/_0_  = ~n11595 ;
  assign \g83671/_0_  = ~n11598 ;
  assign \g83715/_3_  = ~n11601 ;
  assign \g83716/_3_  = ~n11604 ;
  assign \g83717/_3_  = n11607 ;
  assign \g83718/_3_  = n11610 ;
  assign \g83719/_3_  = ~n11613 ;
  assign \g83720/_3_  = ~n11616 ;
  assign \g83721/_3_  = ~n11619 ;
  assign \g83722/_3_  = n11622 ;
  assign \g83723/_3_  = n11625 ;
  assign \g83724/_3_  = ~n11628 ;
  assign \g83725/_0_  = ~n11631 ;
  assign \g83726/_3_  = ~n11634 ;
  assign \g83727/_3_  = n11637 ;
  assign \g83728/_3_  = ~n11640 ;
  assign \g83729/_3_  = ~n11642 ;
  assign \g83730/_3_  = ~n11645 ;
  assign \g83731/_3_  = ~n11648 ;
  assign \g83732/_3_  = ~n11651 ;
  assign \g83733/_3_  = ~n11654 ;
  assign \g83734/_3_  = ~n11657 ;
  assign \g83735/_0_  = ~n11664 ;
  assign \g83736/_0_  = ~n11667 ;
  assign \g83737/_0_  = ~n11670 ;
  assign \g83738/_3_  = ~n11673 ;
  assign \g83739/_3_  = n11676 ;
  assign \g83740/_0_  = ~n11679 ;
  assign \g83741/_3_  = n11682 ;
  assign \g83742/_3_  = ~n11685 ;
  assign \g84164/_0_  = n3408 ;
  assign \g84181/_0_  = n1162 ;
  assign \g85146/_0_  = ~n11768 ;
  assign \g85147/_0_  = ~n11819 ;
  assign \g85148/_0_  = ~n11839 ;
  assign \g85149/_0_  = ~n11857 ;
  assign \g85151/_0_  = ~n11892 ;
  assign \g85152/_0_  = ~n12028 ;
  assign \g85154/_0_  = ~n12045 ;
  assign \g85155/_0_  = ~n12064 ;
  assign \g85156/_0_  = ~n12087 ;
  assign \g85157/_0_  = ~n12109 ;
  assign \g85158/_0_  = n12129 ;
  assign \g85159/_0_  = ~n12158 ;
  assign \g85160/_0_  = ~n12233 ;
  assign \g85161/_0_  = ~n12262 ;
  assign \g85162/_0_  = ~n12315 ;
  assign \g85163/_0_  = ~n12347 ;
  assign \g85164/_0_  = ~n12402 ;
  assign \g85165/_0_  = ~n12469 ;
  assign \g85166/_0_  = ~n12526 ;
  assign \g85167/_0_  = ~n12583 ;
  assign \g85168/_0_  = ~n12614 ;
  assign \g85169/_0_  = n12634 ;
  assign \g85171/_0_  = n12654 ;
  assign \g85173/_0_  = ~n12672 ;
  assign \g85174/_0_  = ~n12690 ;
  assign \g85175/_0_  = ~n12708 ;
  assign \g85176/_0_  = ~n12726 ;
  assign \g85178/_0_  = ~n12757 ;
  assign \g85179/_0_  = ~n12788 ;
  assign \g85180/_0_  = ~n12819 ;
  assign \g85181/_0_  = ~n12851 ;
  assign \g85182/_0_  = ~n12882 ;
  assign \g85183/_0_  = ~n12913 ;
  assign \g85184/_0_  = ~n12966 ;
  assign \g85185/_0_  = n12998 ;
  assign \g85186/_0_  = ~n13029 ;
  assign \g85187/_0_  = ~n13063 ;
  assign \g85188/_0_  = ~n13089 ;
  assign \g85189/_0_  = n13121 ;
  assign \g85190/_0_  = ~n13152 ;
  assign \g85510/_0_  = ~n13154 ;
  assign \g85711/u3_syn_4  = n11433 ;
  assign \g85972/_0_  = ~n13156 ;
  assign \g86107/_0_  = ~n2711 ;
  assign \g86200/u3_syn_4  = n9331 ;
  assign \g86477/_0_  = ~n2716 ;
  assign \g86548/_0_  = n2052 ;
  assign \g86652/u3_syn_4  = n13157 ;
  assign \g86807/u3_syn_4  = n13158 ;
  assign \g87581/_0_  = ~n3801 ;
  assign \g88104/_0_  = ~n1665 ;
  assign \g88112/_0_  = ~n3248 ;
  assign \g88136/_0_  = ~n3404 ;
  assign \g88148/_0_  = ~n3520 ;
  assign \g88157/_0_  = ~n3177 ;
  assign \g88171/_0_  = ~n3340 ;
  assign \g88179/_0_  = ~n3444 ;
  assign \g88208/_0_  = ~n3561 ;
  assign \g88217/_0_  = ~n3640 ;
  assign \g88222/_0_  = ~n3587 ;
  assign \g88228/_0_  = ~n3153 ;
  assign \g88236/_0_  = ~n3717 ;
  assign \g88242/_0_  = ~n3613 ;
  assign \g88252_dup/_0_  = ~n1701 ;
  assign \g88253/_2_  = ~n1618 ;
  assign \g88259/_0_  = ~n1750 ;
  assign \g88274/_0_  = ~n3078 ;
  assign \g88286/_0_  = ~n3128 ;
  assign \g88296/_0_  = ~n3105 ;
  assign \g88306/_0_  = ~n2974 ;
  assign \g88319/_0_  = ~n2904 ;
  assign \g88330/_0_  = ~n3318 ;
  assign \g88370/_0_  = ~n3275 ;
  assign \g88375/_0_  = ~n3221 ;
  assign \g88388/_0_  = ~n3494 ;
  assign \g88397/_0_  = ~n3300 ;
  assign \g88404/_0_  = ~n3665 ;
  assign \g88793/_0_  = ~n1269 ;
  assign \g88834/_0_  = ~n944 ;
  assign \g88905/_0_  = ~n921 ;
  assign \g88910/_0_  = ~n1158 ;
  assign \g88936_dup/_0_  = ~n772 ;
  assign \g88953/_0_  = ~n1062 ;
  assign \g88962/_0_  = ~n1693 ;
  assign \g89007/_0_  = ~n1410 ;
  assign \g89018/_0_  = ~n1382 ;
  assign \g89024/_0_  = ~n1474 ;
  assign \g89031/_0_  = ~n1445 ;
  assign \g89066/_0_  = ~n986 ;
  assign \g89082/_0_  = ~n1037 ;
  assign \g89097/_0_  = ~n1134 ;
  assign \g90677/_1__syn_2  = n4085 ;
  assign \g96226/_0_  = ~n3741 ;
  assign \g96236/_0_  = ~n3470 ;
  assign \g96261/_0_  = ~n13183 ;
  assign \g96339/_0_  = ~n3381 ;
  assign \g96380/_1_  = ~n3026 ;
  assign \g96418/_0_  = ~n3692 ;
  assign \g96566/_1_  = ~n4015 ;
  assign \g96574/_0_  = ~n3984 ;
  assign \g96620/_0_  = ~n822 ;
  assign \g96629/_0_  = ~n1309 ;
  assign \g96735/_0_  = ~n2045 ;
  assign \g96866/_0_  = ~n893 ;
  assign \g96875/_0_  = ~n1013 ;
  assign \g96910/_0_  = ~n1193 ;
  assign \g96946/_0_  = ~n1231 ;
  assign \g96965/_0_  = ~n868 ;
  assign \g97098/_0_  = ~n783 ;
  assign \g97228/_0_  = ~n1587 ;
  assign \g97231/_0_  = ~n1525 ;
  assign \g97242/_0_  = ~n1110 ;
  assign \g97384/_0_  = ~n1086 ;
  assign \g97409/_0_  = ~n601 ;
  assign \g97506/_0_  = ~n1549 ;
  assign \g97626/_0_  = ~n13210 ;
  assign rd_pad = ~n13213 ;
  assign \so[0]_pad  = n13216 ;
  assign \so[10]_pad  = ~n13258 ;
  assign \so[11]_pad  = ~n13266 ;
  assign \so[12]_pad  = ~n13274 ;
  assign \so[13]_pad  = ~n13282 ;
  assign \so[14]_pad  = ~n13290 ;
  assign \so[15]_pad  = ~n13298 ;
  assign \so[16]_pad  = ~n13306 ;
  assign \so[17]_pad  = ~n13314 ;
  assign \so[18]_pad  = ~n13322 ;
  assign \so[19]_pad  = ~n13328 ;
  assign \so[1]_pad  = ~n13332 ;
  assign \so[2]_pad  = ~n13336 ;
  assign \so[3]_pad  = ~n13340 ;
  assign \so[4]_pad  = ~n13344 ;
  assign \so[5]_pad  = ~n13348 ;
  assign \so[6]_pad  = ~n13352 ;
  assign \so[7]_pad  = ~n13356 ;
  assign \so[8]_pad  = ~n13360 ;
  assign \so[9]_pad  = ~n13364 ;
  assign wr_pad = ~n13367 ;
endmodule
