module top (\g1002_reg/NET0131 , \g1008_reg/NET0131 , \g10122_pad , \g1018_reg/NET0131 , \g1024_reg/NET0131 , \g10306_pad , \g1030_reg/NET0131 , \g1036_reg/NET0131 , \g1041_reg/NET0131 , \g1046_reg/NET0131 , \g10500_pad , \g10527_pad , \g1052_reg/NET0131 , \g1061_reg/NET0131 , \g1070_reg/NET0131 , \g1087_reg/NET0131 , \g1094_reg/NET0131 , \g1099_reg/NET0131 , \g1105_reg/NET0131 , \g1111_reg/NET0131 , \g1124_reg/NET0131 , \g1129_reg/NET0131 , \g1135_reg/NET0131 , \g1141_reg/NET0131 , \g11447_pad , \g1146_reg/NET0131 , \g1152_reg/NET0131 , \g1171_reg/NET0131 , \g11770_pad , \g1178_reg/NET0131 , \g1183_reg/NET0131 , \g1189_reg/NET0131 , \g1193_reg/NET0131 , \g1199_reg/NET0131 , \g1205_reg/NET0131 , \g1211_reg/NET0131 , \g1216_reg/NET0131 , \g12184_pad , \g1221_reg/NET0131 , \g1236_reg/NET0131 , \g1242_reg/NET0131 , \g1246_reg/NET0131 , \g12919_pad , \g12923_pad , \g1300_reg/NET0131 , \g13039_pad , \g1306_reg/NET0131 , \g1312_reg/NET0131 , \g1319_reg/NET0131 , \g1322_reg/NET0131 , \g13259_pad , \g13272_pad , \g1333_reg/NET0131 , \g1339_reg/NET0131 , \g1345_reg/NET0131 , \g1351_reg/NET0131 , \g1361_reg/NET0131 , \g1367_reg/NET0131 , \g1373_reg/NET0131 , \g1379_reg/NET0131 , \g1384_reg/NET0131 , \g13865_pad , \g13895_pad , \g1389_reg/NET0131 , \g1395_reg/NET0131 , \g1404_reg/NET0131 , \g14096_pad , \g14125_pad , \g1413_reg/NET0131 , \g14147_pad , \g14167_pad , \g14189_pad , \g14201_pad , \g14217_pad , \g142_reg/NET0131 , \g1430_reg/NET0131 , \g1437_reg/NET0131 , \g1442_reg/NET0131 , \g1448_reg/NET0131 , \g1454_reg/NET0131 , \g1467_reg/NET0131 , \g146_reg/NET0131 , \g1472_reg/NET0131 , \g1478_reg/NET0131 , \g1484_reg/NET0131 , \g1489_reg/NET0131 , \g1495_reg/NET0131 , \g150_reg/NET0131 , \g1514_reg/NET0131 , \g1521_reg/NET0131 , \g1526_reg/NET0131 , \g1532_reg/NET0131 , \g1536_reg/NET0131 , \g153_reg/NET0131 , \g1542_reg/NET0131 , \g1548_reg/NET0131 , \g1554_reg/NET0131 , \g1559_reg/NET0131 , \g1564_reg/NET0131 , \g1579_reg/NET0131 , \g157_reg/NET0131 , \g1585_reg/NET0131 , \g1589_reg/NET0131 , \g1592_reg/NET0131 , \g1600_reg/NET0131 , \g1604_reg/NET0131 , \g1608_reg/NET0131 , \g160_reg/NET0131 , \g1612_reg/NET0131 , \g1616_reg/NET0131 , \g1620_reg/NET0131 , \g1624_reg/NET0131 , \g1632_reg/NET0131 , \g1636_reg/NET0131 , \g1644_reg/NET0131 , \g1648_reg/NET0131 , \g164_reg/NET0131 , \g1657_reg/NET0131 , \g16603_pad , \g16624_pad , \g1664_reg/NET0131 , \g16686_pad , \g1668_reg/NET0131 , \g16718_pad , \g1677_reg/NET0131 , \g1682_reg/NET0131 , \g16874_pad , \g1687_reg/NET0131 , \g168_reg/NET0131 , \g1691_reg/NET0131 , \g1696_reg/NET0131 , \g1700_reg/NET0131 , \g1706_reg/NET0131 , \g1710_reg/NET0131 , \g1714_reg/NET0131 , \g1720_reg/NET0131 , \g1724_reg/NET0131 , \g1728_reg/NET0131 , \g17291_pad , \g17316_pad , \g17320_pad , \g1736_reg/NET0131 , \g17400_pad , \g17404_pad , \g1740_reg/NET0131 , \g17423_pad , \g1744_reg/NET0131 , \g1748_reg/NET0131 , \g174_reg/NET0131 , \g1752_reg/NET0131 , \g1756_reg/NET0131 , \g1760_reg/NET0131 , \g1768_reg/NET0131 , \g1772_reg/NET0131 , \g1779_reg/NET0131 , \g1783_reg/NET0131 , \g1792_reg/NET0131 , \g1798_reg/NET0131 , \g1802_reg/NET0131 , \g18094_pad , \g18095_pad , \g18096_pad , \g18098_pad , \g18099_pad , \g1811_reg/NET0131 , \g1816_reg/NET0131 , \g1821_reg/NET0131 , \g1825_reg/NET0131 , \g182_reg/NET0131 , \g1830_reg/NET0131 , \g1834_reg/NET0131 , \g1840_reg/NET0131 , \g1844_reg/NET0131 , \g1848_reg/NET0131 , \g1854_reg/NET0131 , \g1858_reg/NET0131 , \g1862_reg/NET0131 , \g1870_reg/NET0131 , \g1874_reg/NET0131 , \g1878_reg/NET0131 , \g1882_reg/NET0131 , \g1886_reg/NET0131 , \g1890_reg/NET0131 , \g1894_reg/NET0131 , \g1902_reg/NET0131 , \g1906_reg/NET0131 , \g1913_reg/NET0131 , \g1917_reg/NET0131 , \g191_reg/NET0131 , \g1926_reg/NET0131 , \g1932_reg/NET0131 , \g19334_pad , \g19357_pad , \g1936_reg/NET0131 , \g1945_reg/NET0131 , \g1950_reg/NET0131 , \g1955_reg/NET0131 , \g1959_reg/NET0131 , \g1964_reg/NET0131 , \g1968_reg/NET0131 , \g1974_reg/NET0131 , \g1978_reg/NET0131 , \g1982_reg/NET0131 , \g1988_reg/NET0131 , \g1992_reg/NET0131 , \g1996_reg/NET0131 , \g2004_reg/NET0131 , \g2008_reg/NET0131 , \g2012_reg/NET0131 , \g2016_reg/NET0131 , \g2020_reg/NET0131 , \g2024_reg/NET0131 , \g2028_reg/NET0131 , \g2036_reg/NET0131 , \g203_reg/NET0131 , \g2040_reg/NET0131 , \g2047_reg/NET0131 , \g2051_reg/NET0131 , \g2060_reg/NET0131 , \g2066_reg/NET0131 , \g2070_reg/NET0131 , \g2079_reg/NET0131 , \g2084_reg/NET0131 , \g2089_reg/NET0131 , \g2093_reg/NET0131 , \g2098_reg/NET0131 , \g209_reg/NET0131 , \g2102_reg/NET0131 , \g2108_reg/NET0131 , \g2112_reg/NET0131 , \g2116_reg/NET0131 , \g2122_reg/NET0131 , \g2126_reg/NET0131 , \g2153_reg/NET0131 , \g2161_reg/NET0131 , \g2165_reg/NET0131 , \g2169_reg/NET0131 , \g2173_reg/NET0131 , \g2177_reg/NET0131 , \g2181_reg/NET0131 , \g2185_reg/NET0131 , \g218_reg/NET0131 , \g2193_reg/NET0131 , \g2197_reg/NET0131 , \g2204_reg/NET0131 , \g2208_reg/NET0131 , \g2217_reg/NET0131 , \g2223_reg/NET0131 , \g2227_reg/NET0131 , \g222_reg/NET0131 , \g2236_reg/NET0131 , \g2241_reg/NET0131 , \g2246_reg/NET0131 , \g2250_reg/NET0131 , \g2255_reg/NET0131 , \g2259_reg/NET0131 , \g225_reg/NET0131 , \g2265_reg/NET0131 , \g2269_reg/NET0131 , \g2273_reg/NET0131 , \g2279_reg/NET0131 , \g2283_reg/NET0131 , \g2287_reg/NET0131 , \g2295_reg/NET0131 , \g2299_reg/NET0131 , \g2303_reg/NET0131 , \g2307_reg/NET0131 , \g2311_reg/NET0131 , \g2315_reg/NET0131 , \g2319_reg/NET0131 , \g2327_reg/NET0131 , \g232_reg/NET0131 , \g2331_reg/NET0131 , \g2338_reg/NET0131 , \g2342_reg/NET0131 , \g2351_reg/NET0131 , \g2357_reg/NET0131 , \g2361_reg/NET0131 , \g2370_reg/NET0131 , \g2375_reg/NET0131 , \g2380_reg/NET0131 , \g2384_reg/NET0131 , \g2389_reg/NET0131 , \g2393_reg/NET0131 , \g2399_reg/NET0131 , \g239_reg/NET0131 , \g2403_reg/NET0131 , \g2407_reg/NET0131 , \g2413_reg/NET0131 , \g2417_reg/NET0131 , \g2421_reg/NET0131 , \g2429_reg/NET0131 , \g2433_reg/NET0131 , \g2437_reg/NET0131 , \g2441_reg/NET0131 , \g2445_reg/NET0131 , \g2449_reg/NET0131 , \g2453_reg/NET0131 , \g2461_reg/NET0131 , \g2465_reg/NET0131 , \g246_reg/NET0131 , \g2472_reg/NET0131 , \g2476_reg/NET0131 , \g2485_reg/NET0131 , \g2491_reg/NET0131 , \g2495_reg/NET0131 , \g2504_reg/NET0131 , \g2509_reg/NET0131 , \g2514_reg/NET0131 , \g2518_reg/NET0131 , \g2523_reg/NET0131 , \g2527_reg/NET0131 , \g2533_reg/NET0131 , \g2537_reg/NET0131 , \g2541_reg/NET0131 , \g2547_reg/NET0131 , \g2551_reg/NET0131 , \g2555_reg/NET0131 , \g255_reg/NET0131 , \g2563_reg/NET0131 , \g2567_reg/NET0131 , \g2571_reg/NET0131 , \g2575_reg/NET0131 , \g2579_reg/NET0131 , \g2583_reg/NET0131 , \g2587_reg/NET0131 , \g2595_reg/NET0131 , \g2599_reg/NET0131 , \g2606_reg/NET0131 , \g2610_reg/NET0131 , \g2619_reg/NET0131 , \g2625_reg/NET0131 , \g2629_reg/NET0131 , \g262_reg/NET0131 , \g2638_reg/NET0131 , \g2643_reg/NET0131 , \g2648_reg/NET0131 , \g2652_reg/NET0131 , \g2657_reg/NET0131 , \g2661_reg/NET0131 , \g2667_reg/NET0131 , \g2671_reg/NET0131 , \g2675_reg/NET0131 , \g2681_reg/NET0131 , \g2685_reg/NET0131 , \g269_reg/NET0131 , \g2715_reg/NET0131 , \g2719_reg/NET0131 , \g2724_reg/NET0131 , \g2729_reg/NET0131 , \g2735_reg/NET0131 , \g2741_reg/NET0131 , \g2748_reg/NET0131 , \g2756_reg/NET0131 , \g2759_reg/NET0131 , \g2763_reg/NET0131 , \g2767_reg/NET0131 , \g2771_reg/NET0131 , \g2775_reg/NET0131 , \g2779_reg/NET0131 , \g2783_reg/NET0131 , \g2787_reg/NET0131 , \g278_reg/NET0131 , \g2791_reg/NET0131 , \g2795_reg/NET0131 , \g2799_reg/NET0131 , \g2803_reg/NET0131 , \g2807_reg/NET0131 , \g2811_reg/NET0131 , \g2815_reg/NET0131 , \g2819_reg/NET0131 , \g2823_reg/NET0131 , \g2827_reg/NET0131 , \g2831_reg/NET0131 , \g2834_reg/NET0131 , \g283_reg/NET0131 , \g2848_reg/NET0131 , \g2856_reg/NET0131 , \g2864_reg/NET0131 , \g2873_reg/NET0131 , \g2878_reg/NET0131 , \g287_reg/NET0131 , \g2882_reg/NET0131 , \g2886_reg/NET0131 , \g2898_reg/NET0131 , \g2902_reg/NET0131 , \g2907_reg/NET0131 , \g2912_reg/NET0131 , \g2917_reg/NET0131 , \g291_reg/NET0131 , \g29211_pad , \g29212_pad , \g29213_pad , \g29214_pad , \g29215_pad , \g29216_pad , \g29218_pad , \g29219_pad , \g29220_pad , \g29221_pad , \g2922_reg/NET0131 , \g2927_reg/NET0131 , \g2932_reg/NET0131 , \g2936_reg/NET0131 , \g2941_reg/NET0131 , \g2946_reg/NET0131 , \g294_reg/NET0131 , \g2950_reg/NET0131 , \g2955_reg/NET0131 , \g2960_reg/NET0131 , \g2965_reg/NET0131 , \g2970_reg/NET0131 , \g2975_reg/NET0131 , \g2980_reg/NET0131 , \g2984_reg/NET0131 , \g2988_reg/NET0131 , \g298_reg/NET0131 , \g2999_reg/NET0131 , \g3003_reg/NET0131 , \g301_reg/NET0131 , \g3050_reg/NET0131 , \g305_reg/NET0131 , \g3096_reg/NET0131 , \g3100_reg/NET0131 , \g3106_reg/NET0131 , \g3111_reg/NET0131 , \g3115_reg/NET0131 , \g3119_reg/NET0131 , \g311_reg/NET0131 , \g3125_reg/NET0131 , \g3129_reg/NET0131 , \g3133_reg/NET0131 , \g3139_reg/NET0131 , \g3143_reg/NET0131 , \g3147_reg/NET0131 , \g3155_reg/NET0131 , \g3161_reg/NET0131 , \g3167_reg/NET0131 , \g316_reg/NET0131 , \g3171_reg/NET0131 , \g3179_reg/NET0131 , \g3187_reg/NET0131 , \g3191_reg/NET0131 , \g3195_reg/NET0131 , \g3199_reg/NET0131 , \g319_reg/NET0131 , \g3203_reg/NET0131 , \g3207_reg/NET0131 , \g3211_reg/NET0131 , \g3215_reg/NET0131 , \g3219_reg/NET0131 , \g3223_reg/NET0131 , \g3227_reg/NET0131 , \g3231_reg/NET0131 , \g3235_reg/NET0131 , \g3239_reg/NET0131 , \g3243_reg/NET0131 , \g3247_reg/NET0131 , \g324_reg/NET0131 , \g3251_reg/NET0131 , \g3255_reg/NET0131 , \g3259_reg/NET0131 , \g3263_reg/NET0131 , \g3288_reg/NET0131 , \g329_reg/NET0131 , \g3303_reg/NET0131 , \g3329_reg/NET0131 , \g3333_reg/NET0131 , \g3338_reg/NET0131 , \g333_reg/NET0131 , \g3343_reg/NET0131 , \g3347_reg/NET0131 , \g3352_reg/NET0131 , \g336_reg/NET0131 , \g341_reg/NET0131 , \g3457_reg/NET0131 , \g3466_reg/NET0131 , \g3470_reg/NET0131 , \g3476_reg/NET0131 , \g347_reg/NET0131 , \g3480_reg/NET0131 , \g3484_reg/NET0131 , \g3490_reg/NET0131 , \g3494_reg/NET0131 , \g34_reg/NET0131 , \g351_reg/NET0131 , \g355_reg/NET0131 , \g358_reg/NET0131 , \g35_pad , \g3639_reg/NET0131 , \g3684_reg/NET0131 , \g3703_reg/NET0131 , \g370_reg/NET0131 , \g376_reg/NET0131 , \g37_reg/NET0131 , \g3808_reg/NET0131 , \g3817_reg/NET0131 , \g3821_reg/NET0131 , \g3827_reg/NET0131 , \g3831_reg/NET0131 , \g3835_reg/NET0131 , \g3841_reg/NET0131 , \g3845_reg/NET0131 , \g385_reg/NET0131 , \g392_reg/NET0131 , \g3990_reg/NET0131 , \g401_reg/NET0131 , \g4035_reg/NET0131 , \g4054_reg/NET0131 , \g4057_reg/NET0131 , \g405_reg/NET0131 , \g4064_reg/NET0131 , \g4072_reg/NET0131 , \g4076_reg/NET0131 , \g4082_reg/NET0131 , \g4087_reg/NET0131 , \g4093_reg/NET0131 , \g4098_reg/NET0131 , \g4104_reg/NET0131 , \g4108_reg/NET0131 , \g4112_reg/NET0131 , \g4116_reg/NET0131 , \g4119_reg/NET0131 , \g411_reg/NET0131 , \g4122_reg/NET0131 , \g4141_reg/NET0131 , \g4145_reg/NET0131 , \g4146_reg/NET0131 , \g4153_reg/NET0131 , \g4157_reg/NET0131 , \g4164_reg/NET0131 , \g4172_reg/NET0131 , \g4176_reg/NET0131 , \g417_reg/NET0131 , \g4180_reg/NET0131 , \g4235_reg/NET0131 , \g4239_reg/NET0131 , \g4242_reg/NET0131 , \g4245_reg/NET0131 , \g424_reg/NET0131 , \g4253_reg/NET0131 , \g4258_reg/NET0131 , \g4264_reg/NET0131 , \g4269_reg/NET0131 , \g4273_reg/NET0131 , \g4281_reg/NET0131 , \g4284_reg/NET0131 , \g4291_reg/NET0131 , \g4297_reg/NET0131 , \g4300_reg/NET0131 , \g4308_reg/NET0131 , \g4311_reg/NET0131 , \g4322_reg/NET0131 , \g4332_reg/NET0131 , \g433_reg/NET0131 , \g4340_reg/NET0131 , \g4349_reg/NET0131 , \g4358_reg/NET0131 , \g4366_reg/NET0131 , \g4369_reg/NET0131 , \g4372_reg/NET0131 , \g4375_reg/NET0131 , \g437_reg/NET0131 , \g4382_reg/NET0131 , \g4388_reg/NET0131 , \g4392_reg/NET0131 , \g4401_reg/NET0131 , \g4405_reg/NET0131 , \g4411_reg/NET0131 , \g4417_reg/NET0131 , \g441_reg/NET0131 , \g4420_reg/NET0131 , \g4423_reg/NET0131 , \g4427_reg/NET0131 , \g4430_reg/NET0131 , \g4434_reg/NET0131 , \g4438_reg/NET0131 , \g4443_reg/NET0131 , \g4452_reg/NET0131 , \g4455_reg/NET0131 , \g4459_reg/NET0131 , \g4462_reg/NET0131 , \g4467_reg/NET0131 , \g446_reg/NET0131 , \g4473_reg/NET0131 , \g4477_reg/NET0131 , \g4480_reg/NET0131 , \g4483_reg/NET0131 , \g4486_reg/NET0131 , \g4489_reg/NET0131 , \g4492_reg/NET0131 , \g4495_reg/NET0131 , \g4498_reg/NET0131 , \g4501_reg/NET0131 , \g4504_reg/NET0131 , \g4512_reg/NET0131 , \g4515_reg/NET0131 , \g4521_reg/NET0131 , \g4527_reg/NET0131 , \g452_reg/NET0131 , \g4531_reg/NET0131 , \g4534_reg/NET0131 , \g4540_reg/NET0131 , \g4543_reg/NET0131 , \g4546_reg/NET0131 , \g4549_reg/NET0131 , \g4552_reg/NET0131 , \g4555_reg/NET0131 , \g4558_reg/NET0131 , \g4561_reg/NET0131 , \g4564_reg/NET0131 , \g4567_reg/NET0131 , \g4572_reg/NET0131 , \g4575_reg/NET0131 , \g4581_reg/NET0131 , \g4584_reg/NET0131 , \g4593_reg/NET0131 , \g4601_reg/NET0131 , \g4608_reg/NET0131 , \g460_reg/NET0131 , \g4616_reg/NET0131 , \g4621_reg/NET0131 , \g4628_reg/NET0131 , \g4633_reg/NET0131 , \g4639_reg/NET0131 , \g4643_reg/NET0131 , \g4646_reg/NET0131 , \g4653_reg/NET0131 , \g4659_reg/NET0131 , \g4664_reg/NET0131 , \g4669_reg/NET0131 , \g4674_reg/NET0131 , \g4681_reg/NET0131 , \g4688_reg/NET0131 , \g4698_reg/NET0131 , \g4704_reg/NET0131 , \g4709_reg/NET0131 , \g4743_reg/NET0131 , \g4749_reg/NET0131 , \g4754_reg/NET0131 , \g475_reg/NET0131 , \g4760_reg/NET0131 , \g4765_reg/NET0131 , \g4771_reg/NET0131 , \g4776_reg/NET0131 , \g4785_reg/NET0131 , \g4793_reg/NET0131 , \g479_reg/NET0131 , \g4801_reg/NET0131 , \g482_reg/NET0131 , \g490_reg/NET0131 , \g496_reg/NET0131 , \g499_reg/NET0131 , \g5016_reg/NET0131 , \g5022_reg/NET0131 , \g5029_reg/NET0131 , \g5033_reg/NET0131 , \g5037_reg/NET0131 , \g5041_reg/NET0131 , \g5046_reg/NET0131 , \g504_reg/NET0131 , \g5052_reg/NET0131 , \g5057_reg/NET0131 , \g5069_reg/NET0131 , \g5073_reg/NET0131 , \g5077_reg/NET0131 , \g5080_reg/NET0131 , \g5084_reg/NET0131 , \g5092_reg/NET0131 , \g5097_reg/NET0131 , \g5101_reg/NET0131 , \g5112_reg/NET0131 , \g5115_reg/NET0131 , \g5124_reg/NET0131 , \g5128_reg/NET0131 , \g5134_reg/NET0131 , \g5138_reg/NET0131 , \g513_reg/NET0131 , \g5142_reg/NET0131 , \g5148_reg/NET0131 , \g5152_reg/NET0131 , \g518_reg/NET0131 , \g528_reg/NET0131 , \g5297_reg/NET0131 , \g534_reg/NET0131 , \g5357_reg/NET0131 , \g538_reg/NET0131 , \g542_reg/NET0131 , \g546_reg/NET0131 , \g550_reg/NET0131 , \g554_reg/NET0131 , \g645_reg/NET0131 , \g650_reg/NET0131 , \g655_reg/NET0131 , \g661_reg/NET0131 , \g667_reg/NET0131 , \g671_reg/NET0131 , \g676_reg/NET0131 , \g681_reg/NET0131 , \g686_reg/NET0131 , \g691_reg/NET0131 , \g699_reg/NET0131 , \g703_reg/NET0131 , \g714_reg/NET0131 , \g718_reg/NET0131 , \g723_reg/NET0131 , \g7243_pad , \g7245_pad , \g7257_pad , \g7260_pad , \g728_reg/NET0131 , \g732_reg/NET0131 , \g736_reg/NET0131 , \g739_reg/NET0131 , \g744_reg/NET0131 , \g749_reg/NET0131 , \g753_reg/NET0131 , \g7540_pad , \g758_reg/NET0131 , \g763_reg/NET0131 , \g767_reg/NET0131 , \g772_reg/NET0131 , \g776_reg/NET0131 , \g781_reg/NET0131 , \g785_reg/NET0131 , \g790_reg/NET0131 , \g7916_pad , \g7946_pad , \g794_reg/NET0131 , \g802_reg/NET0131 , \g807_reg/NET0131 , \g812_reg/NET0131 , \g817_reg/NET0131 , \g822_reg/NET0131 , \g827_reg/NET0131 , \g8291_pad , \g832_reg/NET0131 , \g8358_pad , \g837_reg/NET0131 , \g8416_pad , \g843_reg/NET0131 , \g8475_pad , \g847_reg/NET0131 , \g854_reg/NET0131 , \g862_reg/NET0131 , \g8719_pad , \g872_reg/NET0131 , \g8783_pad , \g8784_pad , \g8785_pad , \g8786_pad , \g8787_pad , \g8788_pad , \g8789_pad , \g8839_pad , \g8870_pad , \g890_reg/NET0131 , \g8915_pad , \g8916_pad , \g8917_pad , \g8918_pad , \g8919_pad , \g8920_pad , \g896_reg/NET0131 , \g9019_pad , \g9251_pad , \g956_reg/NET0131 , \g962_reg/NET0131 , \g969_reg/NET0131 , \g976_reg/NET0131 , \g979_reg/NET0131 , \g990_reg/NET0131 , \g996_reg/NET0131 , \g136_reg/P0001 , \g21727_pad , \g23190_pad , \g26875_pad , \g26876_pad , \g26877_pad , \g28041_pad , \g28042_pad , \g30327_pad , \g30330_pad , \g30331_pad , \g31793_pad , \g31860_pad , \g31862_pad , \g31863_pad , \g32185_pad , \g33079_pad , \g33435_pad , \g33959_pad , \g34435_pad , \g34788_pad , \g34956_pad , \g34_reg/P0001 , \g35_syn_2 , \g37/_0_ , \g41/_0_ , \g60853/_3_ , \g60856/_3_ , \g60879/_3_ , \g60882/_0_ , \g60888/_0_ , \g60891/_0_ , \g60896/_0_ , \g60899/_0_ , \g60900/_3_ , \g60909/_3_ , \g60911/_0_ , \g60915/_0_ , \g60918/_0_ , \g60919/_0_ , \g60928/_0_ , \g60929/_0_ , \g60936/_0_ , \g60937/_0_ , \g60939/_0_ , \g60940/_0_ , \g60941/_0_ , \g60942/_0_ , \g60943/_0_ , \g60944/_0_ , \g60952/_0_ , \g60954/_0_ , \g60958/_0_ , \g60962/_3_ , \g60972/_0_ , \g60980/_0_ , \g60984/_0_ , \g60986/_0_ , \g60989/_0_ , \g60991/_3_ , \g61006/_0_ , \g61008/_0_ , \g61013/_0_ , \g61014/_0_ , \g61015/_0_ , \g61016/_0_ , \g61017/_0_ , \g61026/_3_ , \g61027/_3_ , \g61030/_0_ , \g61031/_0_ , \g61037/_0_ , \g61038/_0_ , \g61042/_0_ , \g61044/_0_ , \g61045/_0_ , \g61046/_0_ , \g61050/_0_ , \g61051/_0_ , \g61052/_0_ , \g61078/_0_ , \g61131/_0_ , \g61137/_3_ , \g61142/_3_ , \g61143/_3_ , \g61151/_0_ , \g61152/_0_ , \g61161/_0_ , \g61168/_3_ , \g61169/_3_ , \g61170/_0_ , \g61171/_3_ , \g61172/_0_ , \g61173/_0_ , \g61174/_0_ , \g61175/_0_ , \g61176/_0_ , \g61177/_3_ , \g61178/_0_ , \g61179/_0_ , \g61180/_0_ , \g61181/_0_ , \g61182/_3_ , \g61183/_0_ , \g61184/_3_ , \g61185/_0_ , \g61186/_0_ , \g61187/_0_ , \g61188/_0_ , \g61189/_0_ , \g61190/_3_ , \g61191/_0_ , \g61192/_0_ , \g61193/_0_ , \g61194/_0_ , \g61221/_0_ , \g61222/_0_ , \g61223/_3_ , \g61224/_3_ , \g61261/_0_ , \g61295/_3_ , \g61308/_0_ , \g61316/_0_ , \g61327/_0_ , \g61329/_0_ , \g61330/_0_ , \g61331/_0_ , \g61332/_3_ , \g61333/_0_ , \g61334/_0_ , \g61335/_0_ , \g61336/_0_ , \g61337/_0_ , \g61338/_3_ , \g61339/_0_ , \g61340/_0_ , \g61341/_0_ , \g61342/_0_ , \g61343/_0_ , \g61344/_3_ , \g61345/_0_ , \g61346/_0_ , \g61347/_0_ , \g61348/_0_ , \g61349/_0_ , \g61350/_3_ , \g61351/_0_ , \g61352/_0_ , \g61353/_0_ , \g61354/_0_ , \g61367/_0_ , \g61372/_0_ , \g61373/_0_ , \g61375/_0_ , \g61382/_0_ , \g61385/_3_ , \g61386/_0_ , \g61399/_0_ , \g61400/_0_ , \g61402/_0_ , \g61405/_0_ , \g61435/_3_ , \g61449/_0_ , \g61468/_0_ , \g61475/_0_ , \g61480/_0_ , \g61482/_0_ , \g61483/_0_ , \g61484/_0_ , \g61486/_3_ , \g61494/_0_ , \g61496/_0_ , \g61497/_0_ , \g61514/_0_ , \g61517/_0_ , \g61519/_3_ , \g61520/_3_ , \g61527/_0_ , \g61541/_0_ , \g61544/_0_ , \g61550/_0_ , \g61551/_0_ , \g61554/_0_ , \g61556/_3_ , \g61567/_0_ , \g61571/_0_ , \g61574/_0_ , \g61587/_0_ , \g61592/_0_ , \g61632/_0_ , \g61634/_0_ , \g61635/_0_ , \g61639/_0_ , \g61644/_0_ , \g61652/_3_ , \g61709/_0_ , \g61714/_0_ , \g61720/_0_ , \g61721/_0_ , \g61723/_0_ , \g61725/_0_ , \g61726/_0_ , \g61734/_0_ , \g61739/_0_ , \g61744/_0_ , \g61746/_3_ , \g61747/_3_ , \g61748/_3_ , \g61750/u3_syn_7 , \g61802/_0_ , \g61804/_0_ , \g61808/_0_ , \g61811/_0_ , \g61816/_0_ , \g61818/_0_ , \g61820/_0_ , \g61823/_0_ , \g61824/_0_ , \g61841/_0_ , \g61842/_3_ , \g61844/_3_ , \g61845/_3_ , \g61846/_3_ , \g61847/u3_syn_7 , \g61848/_0_ , \g61849/_3_ , \g61850/_0_ , \g61851/u3_syn_7 , \g61852/_0_ , \g61853/_3_ , \g61854/_3_ , \g61855/_0_ , \g61856/u3_syn_7 , \g61857/_0_ , \g61858/_3_ , \g61859/_3_ , \g61860/u3_syn_7 , \g61861/_0_ , \g61862/_3_ , \g61863/_3_ , \g61864/u3_syn_7 , \g61865/_0_ , \g61866/_3_ , \g61867/_3_ , \g61868/u3_syn_7 , \g61869/_0_ , \g61870/_0_ , \g61871/_3_ , \g61872/_3_ , \g61873/u3_syn_7 , \g61874/_0_ , \g61875/_0_ , \g61877/_3_ , \g61878/_3_ , \g61879/u3_syn_7 , \g61880/_0_ , \g61881/_0_ , \g61882/_0_ , \g61883/_0_ , \g61884/_0_ , \g61914/_0_ , \g61915/_0_ , \g61917/_0_ , \g61918/_0_ , \g61922/_0_ , \g61923/_0_ , \g61924/_0_ , \g61932/_0_ , \g61936/_0_ , \g61945/_0_ , \g61947/_0_ , \g61959/_0_ , \g61960/_0_ , \g61962/_0_ , \g61973/_3_ , \g61974/u3_syn_7 , \g61975/_3_ , \g61976/u3_syn_7 , \g61977/_3_ , \g61978/_3_ , \g61979/u3_syn_7 , \g61980/_3_ , \g61981/_3_ , \g61982/_3_ , \g61983/u3_syn_7 , \g61984/_3_ , \g61985/_3_ , \g61986/u3_syn_7 , \g61987/_3_ , \g61988/_3_ , \g61989/u3_syn_7 , \g61990/_3_ , \g61991/_3_ , \g61992/u3_syn_7 , \g61993/_3_ , \g61994/u3_syn_7 , \g61995/_3_ , \g61996/_3_ , \g61997/_3_ , \g62022/_0_ , \g62028/_0_ , \g62029/_0_ , \g62031/_0_ , \g62033/_0_ , \g62038/_0_ , \g62042/_0_ , \g62046/_0_ , \g62048/_0_ , \g62049/_0_ , \g62051/_0_ , \g62053/_0_ , \g62085/_0_ , \g62101/_0_ , \g62102/_0_ , \g62103/_0_ , \g62105/_0_ , \g62108/_3_ , \g62112/_0_ , \g62137/_3_ , \g62207/_0_ , \g62239/_0_ , \g62240/_0_ , \g62267/_0_ , \g62273/_0_ , \g62284/_0_ , \g62291/_0_ , \g62293/_0_ , \g62298/_0_ , \g62303/_3_ , \g62322/_3_ , \g62323/_3_ , \g62324/_3_ , \g62325/_3_ , \g62583/_0_ , \g62598/_0_ , \g62609/_0_ , \g62636/_0_ , \g62646/_0_ , \g62649/_0_ , \g62658/_0_ , \g62663/_0_ , \g62664/_0_ , \g62667/_0_ , \g62676/_0_ , \g62677/_0_ , \g62678/_3_ , \g62679/_0_ , \g62687/u3_syn_7 , \g62688/u3_syn_7 , \g62689/_0_ , \g62690/_3_ , \g62691/_3_ , \g62693/_0_ , \g62694/_3_ , \g62695/_3_ , \g62696/_3_ , \g62697/_3_ , \g62698/_3_ , \g62699/_3_ , \g62700/_3_ , \g62701/_3_ , \g62702/_3_ , \g62703/_3_ , \g62704/u3_syn_7 , \g62705/_0_ , \g62706/_3_ , \g62707/_3_ , \g62708/u3_syn_7 , \g62709/_0_ , \g62710/_3_ , \g62711/_3_ , \g62712/u3_syn_7 , \g62713/_0_ , \g62714/_3_ , \g62715/_0_ , \g62716/u3_syn_7 , \g62717/_0_ , \g62718/_3_ , \g62719/_0_ , \g62720/u3_syn_7 , \g62721/_0_ , \g62722/_3_ , \g62723/_0_ , \g62724/u3_syn_7 , \g62725/_0_ , \g62726/_3_ , \g62728/_0_ , \g62790/_0_ , \g62791/_0_ , \g62793/_0_ , \g62794/_0_ , \g62795/_0_ , \g62796/_0_ , \g62797/_0_ , \g62807/_0_ , \g62823/_0_ , \g62824/_0_ , \g62833/_0_ , \g62846/_0_ , \g62859/_0_ , \g62860/_0_ , \g62897/_0_ , \g62898/_0_ , \g62922/_3_ , \g62923/_0_ , \g62927/_0_ , \g62938/_3_ , \g62939/_3_ , \g62940/_3_ , \g62941/u3_syn_7 , \g62942/_0_ , \g62943/_3_ , \g62987/_3_ , \g62991/_3_ , \g63015/u3_syn_7 , \g63016/_0_ , \g63017/_3_ , \g63018/_3_ , \g63019/_3_ , \g63020/_3_ , \g63021/_3_ , \g63022/_3_ , \g63025/_3_ , \g63026/_3_ , \g63027/_3_ , \g63029/_3_ , \g63030/_3_ , \g63031/_3_ , \g63033/_3_ , \g63034/_3_ , \g63043/_3_ , \g63044/_3_ , \g63051/_3_ , \g63057/_3_ , \g63068/_3_ , \g63070/_3_ , \g63073/_3_ , \g63081/_3_ , \g63082/_3_ , \g63083/u3_syn_7 , \g63084/_3_ , \g63085/_0_ , \g63086/_3_ , \g63107/_3_ , \g63108/u3_syn_7 , \g63109/u3_syn_7 , \g63110/_0_ , \g63111/_3_ , \g63132/_3_ , \g63133/_3_ , \g63134/_3_ , \g63135/_3_ , \g63136/_3_ , \g63137/_3_ , \g63138/_3_ , \g63139/u3_syn_7 , \g63140/_3_ , \g63141/_3_ , \g63142/_3_ , \g63143/_3_ , \g63144/_3_ , \g63145/_3_ , \g63146/u3_syn_7 , \g63198/_0_ , \g63205/_0_ , \g63208/_0_ , \g63212/_0_ , \g63215/_0_ , \g63219/_0_ , \g63244/_0_ , \g63246/_0_ , \g63254/_0_ , \g63255/_0_ , \g63272/_0_ , \g63276/_0_ , \g63278/_0_ , \g63279/_0_ , \g63280/_0_ , \g63327/_0_ , \g63345/_0_ , \g63346/_3_ , \g63347/_3_ , \g63354/_3_ , \g63358/_3_ , \g63359/u3_syn_7 , \g63361/_3_ , \g63365/_3_ , \g63366/_3_ , \g63367/_3_ , \g63368/_3_ , \g63370/_3_ , \g63479/_0_ , \g63484/_0_ , \g63499/_1_ , \g63520/_0_ , \g63523/_0_ , \g63526/_0_ , \g63538/_0_ , \g63539/_0_ , \g63541/_0_ , \g63555/_0_ , \g63642/_0_ , \g63645/_0_ , \g63648/_3_ , \g63777/_3_ , \g63778/_3_ , \g63781/_0_ , \g63786/u3_syn_7 , \g63787/_3_ , \g63788/_3_ , \g63790/_3_ , \g63791/_3_ , \g63792/u3_syn_7 , \g63794/_0_ , \g63795/_0_ , \g63796/_0_ , \g63798/_3_ , \g63800/_3_ , \g63804/_3_ , \g63805/_3_ , \g63806/_3_ , \g63807/_3_ , \g63808/_3_ , \g63809/_3_ , \g63870/_0_ , \g63883/_0_ , \g63934/_0_ , \g63936/_0_ , \g63938/_0_ , \g63939/_0_ , \g63966/_0_ , \g63970/_0_ , \g63999/_0_ , \g64039/_0_ , \g64040/_0_ , \g64043/_0_ , \g64062/_3_ , \g64078/_0_ , \g64091/_0_ , \g64095/_3_ , \g64096/_3_ , \g64097/u3_syn_7 , \g64098/u3_syn_7 , \g64099/u3_syn_7 , \g64100/u3_syn_7 , \g64134/_0_ , \g64135/_0_ , \g64153/_0_ , \g64155/_0_ , \g64179/_0_ , \g64229/_0_ , \g64235/_0_ , \g64236/_0_ , \g64280/_0_ , \g64315/_0_ , \g64365/_0_ , \g64426/_3_ , \g64438/_3_ , \g64442/u3_syn_7 , \g64445/_3_ , \g64447/_3_ , \g64449/_3_ , \g64451/_3_ , \g64453/_3_ , \g64454/_3_ , \g64460/_3_ , \g64461/_3_ , \g64510/_0_ , \g64527/_0_ , \g64528/_0_ , \g64544/_0_ , \g64549/_0_ , \g64566/_0_ , \g64576/_0_ , \g64602/_0_ , \g64691/_0_ , \g64697/_0_ , \g64707/_3_ , \g64778/_3_ , \g64790/_3_ , \g64791/_3_ , \g64792/_3_ , \g64793/_3_ , \g64794/_3_ , \g64795/_3_ , \g64796/_3_ , \g64797/_3_ , \g64877/_0_ , \g64912/_0_ , \g64973/_0_ , \g65047/_3_ , \g65081/_3_ , \g65088/_3_ , \g65097/_3_ , \g65100/_3_ , \g65101/_3_ , \g65104/_3_ , \g65105/_3_ , \g65107/_3_ , \g65110/_3_ , \g65111/_3_ , \g65113/_3_ , \g65114/_3_ , \g65266/_0_ , \g65267/_0_ , \g65294/_1_ , \g65328/_1_ , \g65495/_0_ , \g65499/_0_ , \g65503/_0_ , \g65529/_0_ , \g65530/_3_ , \g65531/_3_ , \g65532/_3_ , \g65533/_3_ , \g65624/_0_ , \g65625/_1_ , \g65641/_0_ , \g65701/_0_ , \g65704/_0_ , \g65853/_0_ , \g65891/_0_ , \g65901/_0_ , \g65986/_0_ , \g66029/_0_ , \g66066/_0_ , \g66067/_0_ , \g66068/_0_ , \g66154/_3_ , \g66362/_0_ , \g66369/_0_ , \g66398/_0_ , \g66409/_0_ , \g66419/_0_ , \g66439/_0_ , \g66443/_0_ , \g66464/_0_ , \g66471/_0_ , \g66512/_0_ , \g66528/_0_ , \g66541/_0_ , \g66558/_0_ , \g66644/_0_ , \g66684/_0_ , \g66697/_0_ , \g66698/_0_ , \g66701/_0_ , \g66714/_0_ , \g66715/_0_ , \g66745/_0_ , \g66750/_0_ , \g66751/_0_ , \g66810/_0_ , \g66844/_0_ , \g66853/_0_ , \g66897/_0_ , \g66905/_0_ , \g69743/_0_ , \g69750/_0_ , \g69773/_1_ , \g69792/_1_ , \g69858/_0_ , \g69938/_0_ , \g69949/_0_ , \g70167/_0_ , \g71190/_0_ , \g71198/_0_ , \g71284/_0_ , \g72369/_1_ , \g72467/_0_ , \g72476/_0_ , \g72477/_1_ , \g72648/_0_ , \g72741/_0_ , \g72772/_0_ , \g8132_pad );
	input \g1002_reg/NET0131  ;
	input \g1008_reg/NET0131  ;
	input \g10122_pad  ;
	input \g1018_reg/NET0131  ;
	input \g1024_reg/NET0131  ;
	input \g10306_pad  ;
	input \g1030_reg/NET0131  ;
	input \g1036_reg/NET0131  ;
	input \g1041_reg/NET0131  ;
	input \g1046_reg/NET0131  ;
	input \g10500_pad  ;
	input \g10527_pad  ;
	input \g1052_reg/NET0131  ;
	input \g1061_reg/NET0131  ;
	input \g1070_reg/NET0131  ;
	input \g1087_reg/NET0131  ;
	input \g1094_reg/NET0131  ;
	input \g1099_reg/NET0131  ;
	input \g1105_reg/NET0131  ;
	input \g1111_reg/NET0131  ;
	input \g1124_reg/NET0131  ;
	input \g1129_reg/NET0131  ;
	input \g1135_reg/NET0131  ;
	input \g1141_reg/NET0131  ;
	input \g11447_pad  ;
	input \g1146_reg/NET0131  ;
	input \g1152_reg/NET0131  ;
	input \g1171_reg/NET0131  ;
	input \g11770_pad  ;
	input \g1178_reg/NET0131  ;
	input \g1183_reg/NET0131  ;
	input \g1189_reg/NET0131  ;
	input \g1193_reg/NET0131  ;
	input \g1199_reg/NET0131  ;
	input \g1205_reg/NET0131  ;
	input \g1211_reg/NET0131  ;
	input \g1216_reg/NET0131  ;
	input \g12184_pad  ;
	input \g1221_reg/NET0131  ;
	input \g1236_reg/NET0131  ;
	input \g1242_reg/NET0131  ;
	input \g1246_reg/NET0131  ;
	input \g12919_pad  ;
	input \g12923_pad  ;
	input \g1300_reg/NET0131  ;
	input \g13039_pad  ;
	input \g1306_reg/NET0131  ;
	input \g1312_reg/NET0131  ;
	input \g1319_reg/NET0131  ;
	input \g1322_reg/NET0131  ;
	input \g13259_pad  ;
	input \g13272_pad  ;
	input \g1333_reg/NET0131  ;
	input \g1339_reg/NET0131  ;
	input \g1345_reg/NET0131  ;
	input \g1351_reg/NET0131  ;
	input \g1361_reg/NET0131  ;
	input \g1367_reg/NET0131  ;
	input \g1373_reg/NET0131  ;
	input \g1379_reg/NET0131  ;
	input \g1384_reg/NET0131  ;
	input \g13865_pad  ;
	input \g13895_pad  ;
	input \g1389_reg/NET0131  ;
	input \g1395_reg/NET0131  ;
	input \g1404_reg/NET0131  ;
	input \g14096_pad  ;
	input \g14125_pad  ;
	input \g1413_reg/NET0131  ;
	input \g14147_pad  ;
	input \g14167_pad  ;
	input \g14189_pad  ;
	input \g14201_pad  ;
	input \g14217_pad  ;
	input \g142_reg/NET0131  ;
	input \g1430_reg/NET0131  ;
	input \g1437_reg/NET0131  ;
	input \g1442_reg/NET0131  ;
	input \g1448_reg/NET0131  ;
	input \g1454_reg/NET0131  ;
	input \g1467_reg/NET0131  ;
	input \g146_reg/NET0131  ;
	input \g1472_reg/NET0131  ;
	input \g1478_reg/NET0131  ;
	input \g1484_reg/NET0131  ;
	input \g1489_reg/NET0131  ;
	input \g1495_reg/NET0131  ;
	input \g150_reg/NET0131  ;
	input \g1514_reg/NET0131  ;
	input \g1521_reg/NET0131  ;
	input \g1526_reg/NET0131  ;
	input \g1532_reg/NET0131  ;
	input \g1536_reg/NET0131  ;
	input \g153_reg/NET0131  ;
	input \g1542_reg/NET0131  ;
	input \g1548_reg/NET0131  ;
	input \g1554_reg/NET0131  ;
	input \g1559_reg/NET0131  ;
	input \g1564_reg/NET0131  ;
	input \g1579_reg/NET0131  ;
	input \g157_reg/NET0131  ;
	input \g1585_reg/NET0131  ;
	input \g1589_reg/NET0131  ;
	input \g1592_reg/NET0131  ;
	input \g1600_reg/NET0131  ;
	input \g1604_reg/NET0131  ;
	input \g1608_reg/NET0131  ;
	input \g160_reg/NET0131  ;
	input \g1612_reg/NET0131  ;
	input \g1616_reg/NET0131  ;
	input \g1620_reg/NET0131  ;
	input \g1624_reg/NET0131  ;
	input \g1632_reg/NET0131  ;
	input \g1636_reg/NET0131  ;
	input \g1644_reg/NET0131  ;
	input \g1648_reg/NET0131  ;
	input \g164_reg/NET0131  ;
	input \g1657_reg/NET0131  ;
	input \g16603_pad  ;
	input \g16624_pad  ;
	input \g1664_reg/NET0131  ;
	input \g16686_pad  ;
	input \g1668_reg/NET0131  ;
	input \g16718_pad  ;
	input \g1677_reg/NET0131  ;
	input \g1682_reg/NET0131  ;
	input \g16874_pad  ;
	input \g1687_reg/NET0131  ;
	input \g168_reg/NET0131  ;
	input \g1691_reg/NET0131  ;
	input \g1696_reg/NET0131  ;
	input \g1700_reg/NET0131  ;
	input \g1706_reg/NET0131  ;
	input \g1710_reg/NET0131  ;
	input \g1714_reg/NET0131  ;
	input \g1720_reg/NET0131  ;
	input \g1724_reg/NET0131  ;
	input \g1728_reg/NET0131  ;
	input \g17291_pad  ;
	input \g17316_pad  ;
	input \g17320_pad  ;
	input \g1736_reg/NET0131  ;
	input \g17400_pad  ;
	input \g17404_pad  ;
	input \g1740_reg/NET0131  ;
	input \g17423_pad  ;
	input \g1744_reg/NET0131  ;
	input \g1748_reg/NET0131  ;
	input \g174_reg/NET0131  ;
	input \g1752_reg/NET0131  ;
	input \g1756_reg/NET0131  ;
	input \g1760_reg/NET0131  ;
	input \g1768_reg/NET0131  ;
	input \g1772_reg/NET0131  ;
	input \g1779_reg/NET0131  ;
	input \g1783_reg/NET0131  ;
	input \g1792_reg/NET0131  ;
	input \g1798_reg/NET0131  ;
	input \g1802_reg/NET0131  ;
	input \g18094_pad  ;
	input \g18095_pad  ;
	input \g18096_pad  ;
	input \g18098_pad  ;
	input \g18099_pad  ;
	input \g1811_reg/NET0131  ;
	input \g1816_reg/NET0131  ;
	input \g1821_reg/NET0131  ;
	input \g1825_reg/NET0131  ;
	input \g182_reg/NET0131  ;
	input \g1830_reg/NET0131  ;
	input \g1834_reg/NET0131  ;
	input \g1840_reg/NET0131  ;
	input \g1844_reg/NET0131  ;
	input \g1848_reg/NET0131  ;
	input \g1854_reg/NET0131  ;
	input \g1858_reg/NET0131  ;
	input \g1862_reg/NET0131  ;
	input \g1870_reg/NET0131  ;
	input \g1874_reg/NET0131  ;
	input \g1878_reg/NET0131  ;
	input \g1882_reg/NET0131  ;
	input \g1886_reg/NET0131  ;
	input \g1890_reg/NET0131  ;
	input \g1894_reg/NET0131  ;
	input \g1902_reg/NET0131  ;
	input \g1906_reg/NET0131  ;
	input \g1913_reg/NET0131  ;
	input \g1917_reg/NET0131  ;
	input \g191_reg/NET0131  ;
	input \g1926_reg/NET0131  ;
	input \g1932_reg/NET0131  ;
	input \g19334_pad  ;
	input \g19357_pad  ;
	input \g1936_reg/NET0131  ;
	input \g1945_reg/NET0131  ;
	input \g1950_reg/NET0131  ;
	input \g1955_reg/NET0131  ;
	input \g1959_reg/NET0131  ;
	input \g1964_reg/NET0131  ;
	input \g1968_reg/NET0131  ;
	input \g1974_reg/NET0131  ;
	input \g1978_reg/NET0131  ;
	input \g1982_reg/NET0131  ;
	input \g1988_reg/NET0131  ;
	input \g1992_reg/NET0131  ;
	input \g1996_reg/NET0131  ;
	input \g2004_reg/NET0131  ;
	input \g2008_reg/NET0131  ;
	input \g2012_reg/NET0131  ;
	input \g2016_reg/NET0131  ;
	input \g2020_reg/NET0131  ;
	input \g2024_reg/NET0131  ;
	input \g2028_reg/NET0131  ;
	input \g2036_reg/NET0131  ;
	input \g203_reg/NET0131  ;
	input \g2040_reg/NET0131  ;
	input \g2047_reg/NET0131  ;
	input \g2051_reg/NET0131  ;
	input \g2060_reg/NET0131  ;
	input \g2066_reg/NET0131  ;
	input \g2070_reg/NET0131  ;
	input \g2079_reg/NET0131  ;
	input \g2084_reg/NET0131  ;
	input \g2089_reg/NET0131  ;
	input \g2093_reg/NET0131  ;
	input \g2098_reg/NET0131  ;
	input \g209_reg/NET0131  ;
	input \g2102_reg/NET0131  ;
	input \g2108_reg/NET0131  ;
	input \g2112_reg/NET0131  ;
	input \g2116_reg/NET0131  ;
	input \g2122_reg/NET0131  ;
	input \g2126_reg/NET0131  ;
	input \g2153_reg/NET0131  ;
	input \g2161_reg/NET0131  ;
	input \g2165_reg/NET0131  ;
	input \g2169_reg/NET0131  ;
	input \g2173_reg/NET0131  ;
	input \g2177_reg/NET0131  ;
	input \g2181_reg/NET0131  ;
	input \g2185_reg/NET0131  ;
	input \g218_reg/NET0131  ;
	input \g2193_reg/NET0131  ;
	input \g2197_reg/NET0131  ;
	input \g2204_reg/NET0131  ;
	input \g2208_reg/NET0131  ;
	input \g2217_reg/NET0131  ;
	input \g2223_reg/NET0131  ;
	input \g2227_reg/NET0131  ;
	input \g222_reg/NET0131  ;
	input \g2236_reg/NET0131  ;
	input \g2241_reg/NET0131  ;
	input \g2246_reg/NET0131  ;
	input \g2250_reg/NET0131  ;
	input \g2255_reg/NET0131  ;
	input \g2259_reg/NET0131  ;
	input \g225_reg/NET0131  ;
	input \g2265_reg/NET0131  ;
	input \g2269_reg/NET0131  ;
	input \g2273_reg/NET0131  ;
	input \g2279_reg/NET0131  ;
	input \g2283_reg/NET0131  ;
	input \g2287_reg/NET0131  ;
	input \g2295_reg/NET0131  ;
	input \g2299_reg/NET0131  ;
	input \g2303_reg/NET0131  ;
	input \g2307_reg/NET0131  ;
	input \g2311_reg/NET0131  ;
	input \g2315_reg/NET0131  ;
	input \g2319_reg/NET0131  ;
	input \g2327_reg/NET0131  ;
	input \g232_reg/NET0131  ;
	input \g2331_reg/NET0131  ;
	input \g2338_reg/NET0131  ;
	input \g2342_reg/NET0131  ;
	input \g2351_reg/NET0131  ;
	input \g2357_reg/NET0131  ;
	input \g2361_reg/NET0131  ;
	input \g2370_reg/NET0131  ;
	input \g2375_reg/NET0131  ;
	input \g2380_reg/NET0131  ;
	input \g2384_reg/NET0131  ;
	input \g2389_reg/NET0131  ;
	input \g2393_reg/NET0131  ;
	input \g2399_reg/NET0131  ;
	input \g239_reg/NET0131  ;
	input \g2403_reg/NET0131  ;
	input \g2407_reg/NET0131  ;
	input \g2413_reg/NET0131  ;
	input \g2417_reg/NET0131  ;
	input \g2421_reg/NET0131  ;
	input \g2429_reg/NET0131  ;
	input \g2433_reg/NET0131  ;
	input \g2437_reg/NET0131  ;
	input \g2441_reg/NET0131  ;
	input \g2445_reg/NET0131  ;
	input \g2449_reg/NET0131  ;
	input \g2453_reg/NET0131  ;
	input \g2461_reg/NET0131  ;
	input \g2465_reg/NET0131  ;
	input \g246_reg/NET0131  ;
	input \g2472_reg/NET0131  ;
	input \g2476_reg/NET0131  ;
	input \g2485_reg/NET0131  ;
	input \g2491_reg/NET0131  ;
	input \g2495_reg/NET0131  ;
	input \g2504_reg/NET0131  ;
	input \g2509_reg/NET0131  ;
	input \g2514_reg/NET0131  ;
	input \g2518_reg/NET0131  ;
	input \g2523_reg/NET0131  ;
	input \g2527_reg/NET0131  ;
	input \g2533_reg/NET0131  ;
	input \g2537_reg/NET0131  ;
	input \g2541_reg/NET0131  ;
	input \g2547_reg/NET0131  ;
	input \g2551_reg/NET0131  ;
	input \g2555_reg/NET0131  ;
	input \g255_reg/NET0131  ;
	input \g2563_reg/NET0131  ;
	input \g2567_reg/NET0131  ;
	input \g2571_reg/NET0131  ;
	input \g2575_reg/NET0131  ;
	input \g2579_reg/NET0131  ;
	input \g2583_reg/NET0131  ;
	input \g2587_reg/NET0131  ;
	input \g2595_reg/NET0131  ;
	input \g2599_reg/NET0131  ;
	input \g2606_reg/NET0131  ;
	input \g2610_reg/NET0131  ;
	input \g2619_reg/NET0131  ;
	input \g2625_reg/NET0131  ;
	input \g2629_reg/NET0131  ;
	input \g262_reg/NET0131  ;
	input \g2638_reg/NET0131  ;
	input \g2643_reg/NET0131  ;
	input \g2648_reg/NET0131  ;
	input \g2652_reg/NET0131  ;
	input \g2657_reg/NET0131  ;
	input \g2661_reg/NET0131  ;
	input \g2667_reg/NET0131  ;
	input \g2671_reg/NET0131  ;
	input \g2675_reg/NET0131  ;
	input \g2681_reg/NET0131  ;
	input \g2685_reg/NET0131  ;
	input \g269_reg/NET0131  ;
	input \g2715_reg/NET0131  ;
	input \g2719_reg/NET0131  ;
	input \g2724_reg/NET0131  ;
	input \g2729_reg/NET0131  ;
	input \g2735_reg/NET0131  ;
	input \g2741_reg/NET0131  ;
	input \g2748_reg/NET0131  ;
	input \g2756_reg/NET0131  ;
	input \g2759_reg/NET0131  ;
	input \g2763_reg/NET0131  ;
	input \g2767_reg/NET0131  ;
	input \g2771_reg/NET0131  ;
	input \g2775_reg/NET0131  ;
	input \g2779_reg/NET0131  ;
	input \g2783_reg/NET0131  ;
	input \g2787_reg/NET0131  ;
	input \g278_reg/NET0131  ;
	input \g2791_reg/NET0131  ;
	input \g2795_reg/NET0131  ;
	input \g2799_reg/NET0131  ;
	input \g2803_reg/NET0131  ;
	input \g2807_reg/NET0131  ;
	input \g2811_reg/NET0131  ;
	input \g2815_reg/NET0131  ;
	input \g2819_reg/NET0131  ;
	input \g2823_reg/NET0131  ;
	input \g2827_reg/NET0131  ;
	input \g2831_reg/NET0131  ;
	input \g2834_reg/NET0131  ;
	input \g283_reg/NET0131  ;
	input \g2848_reg/NET0131  ;
	input \g2856_reg/NET0131  ;
	input \g2864_reg/NET0131  ;
	input \g2873_reg/NET0131  ;
	input \g2878_reg/NET0131  ;
	input \g287_reg/NET0131  ;
	input \g2882_reg/NET0131  ;
	input \g2886_reg/NET0131  ;
	input \g2898_reg/NET0131  ;
	input \g2902_reg/NET0131  ;
	input \g2907_reg/NET0131  ;
	input \g2912_reg/NET0131  ;
	input \g2917_reg/NET0131  ;
	input \g291_reg/NET0131  ;
	input \g29211_pad  ;
	input \g29212_pad  ;
	input \g29213_pad  ;
	input \g29214_pad  ;
	input \g29215_pad  ;
	input \g29216_pad  ;
	input \g29218_pad  ;
	input \g29219_pad  ;
	input \g29220_pad  ;
	input \g29221_pad  ;
	input \g2922_reg/NET0131  ;
	input \g2927_reg/NET0131  ;
	input \g2932_reg/NET0131  ;
	input \g2936_reg/NET0131  ;
	input \g2941_reg/NET0131  ;
	input \g2946_reg/NET0131  ;
	input \g294_reg/NET0131  ;
	input \g2950_reg/NET0131  ;
	input \g2955_reg/NET0131  ;
	input \g2960_reg/NET0131  ;
	input \g2965_reg/NET0131  ;
	input \g2970_reg/NET0131  ;
	input \g2975_reg/NET0131  ;
	input \g2980_reg/NET0131  ;
	input \g2984_reg/NET0131  ;
	input \g2988_reg/NET0131  ;
	input \g298_reg/NET0131  ;
	input \g2999_reg/NET0131  ;
	input \g3003_reg/NET0131  ;
	input \g301_reg/NET0131  ;
	input \g3050_reg/NET0131  ;
	input \g305_reg/NET0131  ;
	input \g3096_reg/NET0131  ;
	input \g3100_reg/NET0131  ;
	input \g3106_reg/NET0131  ;
	input \g3111_reg/NET0131  ;
	input \g3115_reg/NET0131  ;
	input \g3119_reg/NET0131  ;
	input \g311_reg/NET0131  ;
	input \g3125_reg/NET0131  ;
	input \g3129_reg/NET0131  ;
	input \g3133_reg/NET0131  ;
	input \g3139_reg/NET0131  ;
	input \g3143_reg/NET0131  ;
	input \g3147_reg/NET0131  ;
	input \g3155_reg/NET0131  ;
	input \g3161_reg/NET0131  ;
	input \g3167_reg/NET0131  ;
	input \g316_reg/NET0131  ;
	input \g3171_reg/NET0131  ;
	input \g3179_reg/NET0131  ;
	input \g3187_reg/NET0131  ;
	input \g3191_reg/NET0131  ;
	input \g3195_reg/NET0131  ;
	input \g3199_reg/NET0131  ;
	input \g319_reg/NET0131  ;
	input \g3203_reg/NET0131  ;
	input \g3207_reg/NET0131  ;
	input \g3211_reg/NET0131  ;
	input \g3215_reg/NET0131  ;
	input \g3219_reg/NET0131  ;
	input \g3223_reg/NET0131  ;
	input \g3227_reg/NET0131  ;
	input \g3231_reg/NET0131  ;
	input \g3235_reg/NET0131  ;
	input \g3239_reg/NET0131  ;
	input \g3243_reg/NET0131  ;
	input \g3247_reg/NET0131  ;
	input \g324_reg/NET0131  ;
	input \g3251_reg/NET0131  ;
	input \g3255_reg/NET0131  ;
	input \g3259_reg/NET0131  ;
	input \g3263_reg/NET0131  ;
	input \g3288_reg/NET0131  ;
	input \g329_reg/NET0131  ;
	input \g3303_reg/NET0131  ;
	input \g3329_reg/NET0131  ;
	input \g3333_reg/NET0131  ;
	input \g3338_reg/NET0131  ;
	input \g333_reg/NET0131  ;
	input \g3343_reg/NET0131  ;
	input \g3347_reg/NET0131  ;
	input \g3352_reg/NET0131  ;
	input \g336_reg/NET0131  ;
	input \g341_reg/NET0131  ;
	input \g3457_reg/NET0131  ;
	input \g3466_reg/NET0131  ;
	input \g3470_reg/NET0131  ;
	input \g3476_reg/NET0131  ;
	input \g347_reg/NET0131  ;
	input \g3480_reg/NET0131  ;
	input \g3484_reg/NET0131  ;
	input \g3490_reg/NET0131  ;
	input \g3494_reg/NET0131  ;
	input \g34_reg/NET0131  ;
	input \g351_reg/NET0131  ;
	input \g355_reg/NET0131  ;
	input \g358_reg/NET0131  ;
	input \g35_pad  ;
	input \g3639_reg/NET0131  ;
	input \g3684_reg/NET0131  ;
	input \g3703_reg/NET0131  ;
	input \g370_reg/NET0131  ;
	input \g376_reg/NET0131  ;
	input \g37_reg/NET0131  ;
	input \g3808_reg/NET0131  ;
	input \g3817_reg/NET0131  ;
	input \g3821_reg/NET0131  ;
	input \g3827_reg/NET0131  ;
	input \g3831_reg/NET0131  ;
	input \g3835_reg/NET0131  ;
	input \g3841_reg/NET0131  ;
	input \g3845_reg/NET0131  ;
	input \g385_reg/NET0131  ;
	input \g392_reg/NET0131  ;
	input \g3990_reg/NET0131  ;
	input \g401_reg/NET0131  ;
	input \g4035_reg/NET0131  ;
	input \g4054_reg/NET0131  ;
	input \g4057_reg/NET0131  ;
	input \g405_reg/NET0131  ;
	input \g4064_reg/NET0131  ;
	input \g4072_reg/NET0131  ;
	input \g4076_reg/NET0131  ;
	input \g4082_reg/NET0131  ;
	input \g4087_reg/NET0131  ;
	input \g4093_reg/NET0131  ;
	input \g4098_reg/NET0131  ;
	input \g4104_reg/NET0131  ;
	input \g4108_reg/NET0131  ;
	input \g4112_reg/NET0131  ;
	input \g4116_reg/NET0131  ;
	input \g4119_reg/NET0131  ;
	input \g411_reg/NET0131  ;
	input \g4122_reg/NET0131  ;
	input \g4141_reg/NET0131  ;
	input \g4145_reg/NET0131  ;
	input \g4146_reg/NET0131  ;
	input \g4153_reg/NET0131  ;
	input \g4157_reg/NET0131  ;
	input \g4164_reg/NET0131  ;
	input \g4172_reg/NET0131  ;
	input \g4176_reg/NET0131  ;
	input \g417_reg/NET0131  ;
	input \g4180_reg/NET0131  ;
	input \g4235_reg/NET0131  ;
	input \g4239_reg/NET0131  ;
	input \g4242_reg/NET0131  ;
	input \g4245_reg/NET0131  ;
	input \g424_reg/NET0131  ;
	input \g4253_reg/NET0131  ;
	input \g4258_reg/NET0131  ;
	input \g4264_reg/NET0131  ;
	input \g4269_reg/NET0131  ;
	input \g4273_reg/NET0131  ;
	input \g4281_reg/NET0131  ;
	input \g4284_reg/NET0131  ;
	input \g4291_reg/NET0131  ;
	input \g4297_reg/NET0131  ;
	input \g4300_reg/NET0131  ;
	input \g4308_reg/NET0131  ;
	input \g4311_reg/NET0131  ;
	input \g4322_reg/NET0131  ;
	input \g4332_reg/NET0131  ;
	input \g433_reg/NET0131  ;
	input \g4340_reg/NET0131  ;
	input \g4349_reg/NET0131  ;
	input \g4358_reg/NET0131  ;
	input \g4366_reg/NET0131  ;
	input \g4369_reg/NET0131  ;
	input \g4372_reg/NET0131  ;
	input \g4375_reg/NET0131  ;
	input \g437_reg/NET0131  ;
	input \g4382_reg/NET0131  ;
	input \g4388_reg/NET0131  ;
	input \g4392_reg/NET0131  ;
	input \g4401_reg/NET0131  ;
	input \g4405_reg/NET0131  ;
	input \g4411_reg/NET0131  ;
	input \g4417_reg/NET0131  ;
	input \g441_reg/NET0131  ;
	input \g4420_reg/NET0131  ;
	input \g4423_reg/NET0131  ;
	input \g4427_reg/NET0131  ;
	input \g4430_reg/NET0131  ;
	input \g4434_reg/NET0131  ;
	input \g4438_reg/NET0131  ;
	input \g4443_reg/NET0131  ;
	input \g4452_reg/NET0131  ;
	input \g4455_reg/NET0131  ;
	input \g4459_reg/NET0131  ;
	input \g4462_reg/NET0131  ;
	input \g4467_reg/NET0131  ;
	input \g446_reg/NET0131  ;
	input \g4473_reg/NET0131  ;
	input \g4477_reg/NET0131  ;
	input \g4480_reg/NET0131  ;
	input \g4483_reg/NET0131  ;
	input \g4486_reg/NET0131  ;
	input \g4489_reg/NET0131  ;
	input \g4492_reg/NET0131  ;
	input \g4495_reg/NET0131  ;
	input \g4498_reg/NET0131  ;
	input \g4501_reg/NET0131  ;
	input \g4504_reg/NET0131  ;
	input \g4512_reg/NET0131  ;
	input \g4515_reg/NET0131  ;
	input \g4521_reg/NET0131  ;
	input \g4527_reg/NET0131  ;
	input \g452_reg/NET0131  ;
	input \g4531_reg/NET0131  ;
	input \g4534_reg/NET0131  ;
	input \g4540_reg/NET0131  ;
	input \g4543_reg/NET0131  ;
	input \g4546_reg/NET0131  ;
	input \g4549_reg/NET0131  ;
	input \g4552_reg/NET0131  ;
	input \g4555_reg/NET0131  ;
	input \g4558_reg/NET0131  ;
	input \g4561_reg/NET0131  ;
	input \g4564_reg/NET0131  ;
	input \g4567_reg/NET0131  ;
	input \g4572_reg/NET0131  ;
	input \g4575_reg/NET0131  ;
	input \g4581_reg/NET0131  ;
	input \g4584_reg/NET0131  ;
	input \g4593_reg/NET0131  ;
	input \g4601_reg/NET0131  ;
	input \g4608_reg/NET0131  ;
	input \g460_reg/NET0131  ;
	input \g4616_reg/NET0131  ;
	input \g4621_reg/NET0131  ;
	input \g4628_reg/NET0131  ;
	input \g4633_reg/NET0131  ;
	input \g4639_reg/NET0131  ;
	input \g4643_reg/NET0131  ;
	input \g4646_reg/NET0131  ;
	input \g4653_reg/NET0131  ;
	input \g4659_reg/NET0131  ;
	input \g4664_reg/NET0131  ;
	input \g4669_reg/NET0131  ;
	input \g4674_reg/NET0131  ;
	input \g4681_reg/NET0131  ;
	input \g4688_reg/NET0131  ;
	input \g4698_reg/NET0131  ;
	input \g4704_reg/NET0131  ;
	input \g4709_reg/NET0131  ;
	input \g4743_reg/NET0131  ;
	input \g4749_reg/NET0131  ;
	input \g4754_reg/NET0131  ;
	input \g475_reg/NET0131  ;
	input \g4760_reg/NET0131  ;
	input \g4765_reg/NET0131  ;
	input \g4771_reg/NET0131  ;
	input \g4776_reg/NET0131  ;
	input \g4785_reg/NET0131  ;
	input \g4793_reg/NET0131  ;
	input \g479_reg/NET0131  ;
	input \g4801_reg/NET0131  ;
	input \g482_reg/NET0131  ;
	input \g490_reg/NET0131  ;
	input \g496_reg/NET0131  ;
	input \g499_reg/NET0131  ;
	input \g5016_reg/NET0131  ;
	input \g5022_reg/NET0131  ;
	input \g5029_reg/NET0131  ;
	input \g5033_reg/NET0131  ;
	input \g5037_reg/NET0131  ;
	input \g5041_reg/NET0131  ;
	input \g5046_reg/NET0131  ;
	input \g504_reg/NET0131  ;
	input \g5052_reg/NET0131  ;
	input \g5057_reg/NET0131  ;
	input \g5069_reg/NET0131  ;
	input \g5073_reg/NET0131  ;
	input \g5077_reg/NET0131  ;
	input \g5080_reg/NET0131  ;
	input \g5084_reg/NET0131  ;
	input \g5092_reg/NET0131  ;
	input \g5097_reg/NET0131  ;
	input \g5101_reg/NET0131  ;
	input \g5112_reg/NET0131  ;
	input \g5115_reg/NET0131  ;
	input \g5124_reg/NET0131  ;
	input \g5128_reg/NET0131  ;
	input \g5134_reg/NET0131  ;
	input \g5138_reg/NET0131  ;
	input \g513_reg/NET0131  ;
	input \g5142_reg/NET0131  ;
	input \g5148_reg/NET0131  ;
	input \g5152_reg/NET0131  ;
	input \g518_reg/NET0131  ;
	input \g528_reg/NET0131  ;
	input \g5297_reg/NET0131  ;
	input \g534_reg/NET0131  ;
	input \g5357_reg/NET0131  ;
	input \g538_reg/NET0131  ;
	input \g542_reg/NET0131  ;
	input \g546_reg/NET0131  ;
	input \g550_reg/NET0131  ;
	input \g554_reg/NET0131  ;
	input \g645_reg/NET0131  ;
	input \g650_reg/NET0131  ;
	input \g655_reg/NET0131  ;
	input \g661_reg/NET0131  ;
	input \g667_reg/NET0131  ;
	input \g671_reg/NET0131  ;
	input \g676_reg/NET0131  ;
	input \g681_reg/NET0131  ;
	input \g686_reg/NET0131  ;
	input \g691_reg/NET0131  ;
	input \g699_reg/NET0131  ;
	input \g703_reg/NET0131  ;
	input \g714_reg/NET0131  ;
	input \g718_reg/NET0131  ;
	input \g723_reg/NET0131  ;
	input \g7243_pad  ;
	input \g7245_pad  ;
	input \g7257_pad  ;
	input \g7260_pad  ;
	input \g728_reg/NET0131  ;
	input \g732_reg/NET0131  ;
	input \g736_reg/NET0131  ;
	input \g739_reg/NET0131  ;
	input \g744_reg/NET0131  ;
	input \g749_reg/NET0131  ;
	input \g753_reg/NET0131  ;
	input \g7540_pad  ;
	input \g758_reg/NET0131  ;
	input \g763_reg/NET0131  ;
	input \g767_reg/NET0131  ;
	input \g772_reg/NET0131  ;
	input \g776_reg/NET0131  ;
	input \g781_reg/NET0131  ;
	input \g785_reg/NET0131  ;
	input \g790_reg/NET0131  ;
	input \g7916_pad  ;
	input \g7946_pad  ;
	input \g794_reg/NET0131  ;
	input \g802_reg/NET0131  ;
	input \g807_reg/NET0131  ;
	input \g812_reg/NET0131  ;
	input \g817_reg/NET0131  ;
	input \g822_reg/NET0131  ;
	input \g827_reg/NET0131  ;
	input \g8291_pad  ;
	input \g832_reg/NET0131  ;
	input \g8358_pad  ;
	input \g837_reg/NET0131  ;
	input \g8416_pad  ;
	input \g843_reg/NET0131  ;
	input \g8475_pad  ;
	input \g847_reg/NET0131  ;
	input \g854_reg/NET0131  ;
	input \g862_reg/NET0131  ;
	input \g8719_pad  ;
	input \g872_reg/NET0131  ;
	input \g8783_pad  ;
	input \g8784_pad  ;
	input \g8785_pad  ;
	input \g8786_pad  ;
	input \g8787_pad  ;
	input \g8788_pad  ;
	input \g8789_pad  ;
	input \g8839_pad  ;
	input \g8870_pad  ;
	input \g890_reg/NET0131  ;
	input \g8915_pad  ;
	input \g8916_pad  ;
	input \g8917_pad  ;
	input \g8918_pad  ;
	input \g8919_pad  ;
	input \g8920_pad  ;
	input \g896_reg/NET0131  ;
	input \g9019_pad  ;
	input \g9251_pad  ;
	input \g956_reg/NET0131  ;
	input \g962_reg/NET0131  ;
	input \g969_reg/NET0131  ;
	input \g976_reg/NET0131  ;
	input \g979_reg/NET0131  ;
	input \g990_reg/NET0131  ;
	input \g996_reg/NET0131  ;
	output \g136_reg/P0001  ;
	output \g21727_pad  ;
	output \g23190_pad  ;
	output \g26875_pad  ;
	output \g26876_pad  ;
	output \g26877_pad  ;
	output \g28041_pad  ;
	output \g28042_pad  ;
	output \g30327_pad  ;
	output \g30330_pad  ;
	output \g30331_pad  ;
	output \g31793_pad  ;
	output \g31860_pad  ;
	output \g31862_pad  ;
	output \g31863_pad  ;
	output \g32185_pad  ;
	output \g33079_pad  ;
	output \g33435_pad  ;
	output \g33959_pad  ;
	output \g34435_pad  ;
	output \g34788_pad  ;
	output \g34956_pad  ;
	output \g34_reg/P0001  ;
	output \g35_syn_2  ;
	output \g37/_0_  ;
	output \g41/_0_  ;
	output \g60853/_3_  ;
	output \g60856/_3_  ;
	output \g60879/_3_  ;
	output \g60882/_0_  ;
	output \g60888/_0_  ;
	output \g60891/_0_  ;
	output \g60896/_0_  ;
	output \g60899/_0_  ;
	output \g60900/_3_  ;
	output \g60909/_3_  ;
	output \g60911/_0_  ;
	output \g60915/_0_  ;
	output \g60918/_0_  ;
	output \g60919/_0_  ;
	output \g60928/_0_  ;
	output \g60929/_0_  ;
	output \g60936/_0_  ;
	output \g60937/_0_  ;
	output \g60939/_0_  ;
	output \g60940/_0_  ;
	output \g60941/_0_  ;
	output \g60942/_0_  ;
	output \g60943/_0_  ;
	output \g60944/_0_  ;
	output \g60952/_0_  ;
	output \g60954/_0_  ;
	output \g60958/_0_  ;
	output \g60962/_3_  ;
	output \g60972/_0_  ;
	output \g60980/_0_  ;
	output \g60984/_0_  ;
	output \g60986/_0_  ;
	output \g60989/_0_  ;
	output \g60991/_3_  ;
	output \g61006/_0_  ;
	output \g61008/_0_  ;
	output \g61013/_0_  ;
	output \g61014/_0_  ;
	output \g61015/_0_  ;
	output \g61016/_0_  ;
	output \g61017/_0_  ;
	output \g61026/_3_  ;
	output \g61027/_3_  ;
	output \g61030/_0_  ;
	output \g61031/_0_  ;
	output \g61037/_0_  ;
	output \g61038/_0_  ;
	output \g61042/_0_  ;
	output \g61044/_0_  ;
	output \g61045/_0_  ;
	output \g61046/_0_  ;
	output \g61050/_0_  ;
	output \g61051/_0_  ;
	output \g61052/_0_  ;
	output \g61078/_0_  ;
	output \g61131/_0_  ;
	output \g61137/_3_  ;
	output \g61142/_3_  ;
	output \g61143/_3_  ;
	output \g61151/_0_  ;
	output \g61152/_0_  ;
	output \g61161/_0_  ;
	output \g61168/_3_  ;
	output \g61169/_3_  ;
	output \g61170/_0_  ;
	output \g61171/_3_  ;
	output \g61172/_0_  ;
	output \g61173/_0_  ;
	output \g61174/_0_  ;
	output \g61175/_0_  ;
	output \g61176/_0_  ;
	output \g61177/_3_  ;
	output \g61178/_0_  ;
	output \g61179/_0_  ;
	output \g61180/_0_  ;
	output \g61181/_0_  ;
	output \g61182/_3_  ;
	output \g61183/_0_  ;
	output \g61184/_3_  ;
	output \g61185/_0_  ;
	output \g61186/_0_  ;
	output \g61187/_0_  ;
	output \g61188/_0_  ;
	output \g61189/_0_  ;
	output \g61190/_3_  ;
	output \g61191/_0_  ;
	output \g61192/_0_  ;
	output \g61193/_0_  ;
	output \g61194/_0_  ;
	output \g61221/_0_  ;
	output \g61222/_0_  ;
	output \g61223/_3_  ;
	output \g61224/_3_  ;
	output \g61261/_0_  ;
	output \g61295/_3_  ;
	output \g61308/_0_  ;
	output \g61316/_0_  ;
	output \g61327/_0_  ;
	output \g61329/_0_  ;
	output \g61330/_0_  ;
	output \g61331/_0_  ;
	output \g61332/_3_  ;
	output \g61333/_0_  ;
	output \g61334/_0_  ;
	output \g61335/_0_  ;
	output \g61336/_0_  ;
	output \g61337/_0_  ;
	output \g61338/_3_  ;
	output \g61339/_0_  ;
	output \g61340/_0_  ;
	output \g61341/_0_  ;
	output \g61342/_0_  ;
	output \g61343/_0_  ;
	output \g61344/_3_  ;
	output \g61345/_0_  ;
	output \g61346/_0_  ;
	output \g61347/_0_  ;
	output \g61348/_0_  ;
	output \g61349/_0_  ;
	output \g61350/_3_  ;
	output \g61351/_0_  ;
	output \g61352/_0_  ;
	output \g61353/_0_  ;
	output \g61354/_0_  ;
	output \g61367/_0_  ;
	output \g61372/_0_  ;
	output \g61373/_0_  ;
	output \g61375/_0_  ;
	output \g61382/_0_  ;
	output \g61385/_3_  ;
	output \g61386/_0_  ;
	output \g61399/_0_  ;
	output \g61400/_0_  ;
	output \g61402/_0_  ;
	output \g61405/_0_  ;
	output \g61435/_3_  ;
	output \g61449/_0_  ;
	output \g61468/_0_  ;
	output \g61475/_0_  ;
	output \g61480/_0_  ;
	output \g61482/_0_  ;
	output \g61483/_0_  ;
	output \g61484/_0_  ;
	output \g61486/_3_  ;
	output \g61494/_0_  ;
	output \g61496/_0_  ;
	output \g61497/_0_  ;
	output \g61514/_0_  ;
	output \g61517/_0_  ;
	output \g61519/_3_  ;
	output \g61520/_3_  ;
	output \g61527/_0_  ;
	output \g61541/_0_  ;
	output \g61544/_0_  ;
	output \g61550/_0_  ;
	output \g61551/_0_  ;
	output \g61554/_0_  ;
	output \g61556/_3_  ;
	output \g61567/_0_  ;
	output \g61571/_0_  ;
	output \g61574/_0_  ;
	output \g61587/_0_  ;
	output \g61592/_0_  ;
	output \g61632/_0_  ;
	output \g61634/_0_  ;
	output \g61635/_0_  ;
	output \g61639/_0_  ;
	output \g61644/_0_  ;
	output \g61652/_3_  ;
	output \g61709/_0_  ;
	output \g61714/_0_  ;
	output \g61720/_0_  ;
	output \g61721/_0_  ;
	output \g61723/_0_  ;
	output \g61725/_0_  ;
	output \g61726/_0_  ;
	output \g61734/_0_  ;
	output \g61739/_0_  ;
	output \g61744/_0_  ;
	output \g61746/_3_  ;
	output \g61747/_3_  ;
	output \g61748/_3_  ;
	output \g61750/u3_syn_7  ;
	output \g61802/_0_  ;
	output \g61804/_0_  ;
	output \g61808/_0_  ;
	output \g61811/_0_  ;
	output \g61816/_0_  ;
	output \g61818/_0_  ;
	output \g61820/_0_  ;
	output \g61823/_0_  ;
	output \g61824/_0_  ;
	output \g61841/_0_  ;
	output \g61842/_3_  ;
	output \g61844/_3_  ;
	output \g61845/_3_  ;
	output \g61846/_3_  ;
	output \g61847/u3_syn_7  ;
	output \g61848/_0_  ;
	output \g61849/_3_  ;
	output \g61850/_0_  ;
	output \g61851/u3_syn_7  ;
	output \g61852/_0_  ;
	output \g61853/_3_  ;
	output \g61854/_3_  ;
	output \g61855/_0_  ;
	output \g61856/u3_syn_7  ;
	output \g61857/_0_  ;
	output \g61858/_3_  ;
	output \g61859/_3_  ;
	output \g61860/u3_syn_7  ;
	output \g61861/_0_  ;
	output \g61862/_3_  ;
	output \g61863/_3_  ;
	output \g61864/u3_syn_7  ;
	output \g61865/_0_  ;
	output \g61866/_3_  ;
	output \g61867/_3_  ;
	output \g61868/u3_syn_7  ;
	output \g61869/_0_  ;
	output \g61870/_0_  ;
	output \g61871/_3_  ;
	output \g61872/_3_  ;
	output \g61873/u3_syn_7  ;
	output \g61874/_0_  ;
	output \g61875/_0_  ;
	output \g61877/_3_  ;
	output \g61878/_3_  ;
	output \g61879/u3_syn_7  ;
	output \g61880/_0_  ;
	output \g61881/_0_  ;
	output \g61882/_0_  ;
	output \g61883/_0_  ;
	output \g61884/_0_  ;
	output \g61914/_0_  ;
	output \g61915/_0_  ;
	output \g61917/_0_  ;
	output \g61918/_0_  ;
	output \g61922/_0_  ;
	output \g61923/_0_  ;
	output \g61924/_0_  ;
	output \g61932/_0_  ;
	output \g61936/_0_  ;
	output \g61945/_0_  ;
	output \g61947/_0_  ;
	output \g61959/_0_  ;
	output \g61960/_0_  ;
	output \g61962/_0_  ;
	output \g61973/_3_  ;
	output \g61974/u3_syn_7  ;
	output \g61975/_3_  ;
	output \g61976/u3_syn_7  ;
	output \g61977/_3_  ;
	output \g61978/_3_  ;
	output \g61979/u3_syn_7  ;
	output \g61980/_3_  ;
	output \g61981/_3_  ;
	output \g61982/_3_  ;
	output \g61983/u3_syn_7  ;
	output \g61984/_3_  ;
	output \g61985/_3_  ;
	output \g61986/u3_syn_7  ;
	output \g61987/_3_  ;
	output \g61988/_3_  ;
	output \g61989/u3_syn_7  ;
	output \g61990/_3_  ;
	output \g61991/_3_  ;
	output \g61992/u3_syn_7  ;
	output \g61993/_3_  ;
	output \g61994/u3_syn_7  ;
	output \g61995/_3_  ;
	output \g61996/_3_  ;
	output \g61997/_3_  ;
	output \g62022/_0_  ;
	output \g62028/_0_  ;
	output \g62029/_0_  ;
	output \g62031/_0_  ;
	output \g62033/_0_  ;
	output \g62038/_0_  ;
	output \g62042/_0_  ;
	output \g62046/_0_  ;
	output \g62048/_0_  ;
	output \g62049/_0_  ;
	output \g62051/_0_  ;
	output \g62053/_0_  ;
	output \g62085/_0_  ;
	output \g62101/_0_  ;
	output \g62102/_0_  ;
	output \g62103/_0_  ;
	output \g62105/_0_  ;
	output \g62108/_3_  ;
	output \g62112/_0_  ;
	output \g62137/_3_  ;
	output \g62207/_0_  ;
	output \g62239/_0_  ;
	output \g62240/_0_  ;
	output \g62267/_0_  ;
	output \g62273/_0_  ;
	output \g62284/_0_  ;
	output \g62291/_0_  ;
	output \g62293/_0_  ;
	output \g62298/_0_  ;
	output \g62303/_3_  ;
	output \g62322/_3_  ;
	output \g62323/_3_  ;
	output \g62324/_3_  ;
	output \g62325/_3_  ;
	output \g62583/_0_  ;
	output \g62598/_0_  ;
	output \g62609/_0_  ;
	output \g62636/_0_  ;
	output \g62646/_0_  ;
	output \g62649/_0_  ;
	output \g62658/_0_  ;
	output \g62663/_0_  ;
	output \g62664/_0_  ;
	output \g62667/_0_  ;
	output \g62676/_0_  ;
	output \g62677/_0_  ;
	output \g62678/_3_  ;
	output \g62679/_0_  ;
	output \g62687/u3_syn_7  ;
	output \g62688/u3_syn_7  ;
	output \g62689/_0_  ;
	output \g62690/_3_  ;
	output \g62691/_3_  ;
	output \g62693/_0_  ;
	output \g62694/_3_  ;
	output \g62695/_3_  ;
	output \g62696/_3_  ;
	output \g62697/_3_  ;
	output \g62698/_3_  ;
	output \g62699/_3_  ;
	output \g62700/_3_  ;
	output \g62701/_3_  ;
	output \g62702/_3_  ;
	output \g62703/_3_  ;
	output \g62704/u3_syn_7  ;
	output \g62705/_0_  ;
	output \g62706/_3_  ;
	output \g62707/_3_  ;
	output \g62708/u3_syn_7  ;
	output \g62709/_0_  ;
	output \g62710/_3_  ;
	output \g62711/_3_  ;
	output \g62712/u3_syn_7  ;
	output \g62713/_0_  ;
	output \g62714/_3_  ;
	output \g62715/_0_  ;
	output \g62716/u3_syn_7  ;
	output \g62717/_0_  ;
	output \g62718/_3_  ;
	output \g62719/_0_  ;
	output \g62720/u3_syn_7  ;
	output \g62721/_0_  ;
	output \g62722/_3_  ;
	output \g62723/_0_  ;
	output \g62724/u3_syn_7  ;
	output \g62725/_0_  ;
	output \g62726/_3_  ;
	output \g62728/_0_  ;
	output \g62790/_0_  ;
	output \g62791/_0_  ;
	output \g62793/_0_  ;
	output \g62794/_0_  ;
	output \g62795/_0_  ;
	output \g62796/_0_  ;
	output \g62797/_0_  ;
	output \g62807/_0_  ;
	output \g62823/_0_  ;
	output \g62824/_0_  ;
	output \g62833/_0_  ;
	output \g62846/_0_  ;
	output \g62859/_0_  ;
	output \g62860/_0_  ;
	output \g62897/_0_  ;
	output \g62898/_0_  ;
	output \g62922/_3_  ;
	output \g62923/_0_  ;
	output \g62927/_0_  ;
	output \g62938/_3_  ;
	output \g62939/_3_  ;
	output \g62940/_3_  ;
	output \g62941/u3_syn_7  ;
	output \g62942/_0_  ;
	output \g62943/_3_  ;
	output \g62987/_3_  ;
	output \g62991/_3_  ;
	output \g63015/u3_syn_7  ;
	output \g63016/_0_  ;
	output \g63017/_3_  ;
	output \g63018/_3_  ;
	output \g63019/_3_  ;
	output \g63020/_3_  ;
	output \g63021/_3_  ;
	output \g63022/_3_  ;
	output \g63025/_3_  ;
	output \g63026/_3_  ;
	output \g63027/_3_  ;
	output \g63029/_3_  ;
	output \g63030/_3_  ;
	output \g63031/_3_  ;
	output \g63033/_3_  ;
	output \g63034/_3_  ;
	output \g63043/_3_  ;
	output \g63044/_3_  ;
	output \g63051/_3_  ;
	output \g63057/_3_  ;
	output \g63068/_3_  ;
	output \g63070/_3_  ;
	output \g63073/_3_  ;
	output \g63081/_3_  ;
	output \g63082/_3_  ;
	output \g63083/u3_syn_7  ;
	output \g63084/_3_  ;
	output \g63085/_0_  ;
	output \g63086/_3_  ;
	output \g63107/_3_  ;
	output \g63108/u3_syn_7  ;
	output \g63109/u3_syn_7  ;
	output \g63110/_0_  ;
	output \g63111/_3_  ;
	output \g63132/_3_  ;
	output \g63133/_3_  ;
	output \g63134/_3_  ;
	output \g63135/_3_  ;
	output \g63136/_3_  ;
	output \g63137/_3_  ;
	output \g63138/_3_  ;
	output \g63139/u3_syn_7  ;
	output \g63140/_3_  ;
	output \g63141/_3_  ;
	output \g63142/_3_  ;
	output \g63143/_3_  ;
	output \g63144/_3_  ;
	output \g63145/_3_  ;
	output \g63146/u3_syn_7  ;
	output \g63198/_0_  ;
	output \g63205/_0_  ;
	output \g63208/_0_  ;
	output \g63212/_0_  ;
	output \g63215/_0_  ;
	output \g63219/_0_  ;
	output \g63244/_0_  ;
	output \g63246/_0_  ;
	output \g63254/_0_  ;
	output \g63255/_0_  ;
	output \g63272/_0_  ;
	output \g63276/_0_  ;
	output \g63278/_0_  ;
	output \g63279/_0_  ;
	output \g63280/_0_  ;
	output \g63327/_0_  ;
	output \g63345/_0_  ;
	output \g63346/_3_  ;
	output \g63347/_3_  ;
	output \g63354/_3_  ;
	output \g63358/_3_  ;
	output \g63359/u3_syn_7  ;
	output \g63361/_3_  ;
	output \g63365/_3_  ;
	output \g63366/_3_  ;
	output \g63367/_3_  ;
	output \g63368/_3_  ;
	output \g63370/_3_  ;
	output \g63479/_0_  ;
	output \g63484/_0_  ;
	output \g63499/_1_  ;
	output \g63520/_0_  ;
	output \g63523/_0_  ;
	output \g63526/_0_  ;
	output \g63538/_0_  ;
	output \g63539/_0_  ;
	output \g63541/_0_  ;
	output \g63555/_0_  ;
	output \g63642/_0_  ;
	output \g63645/_0_  ;
	output \g63648/_3_  ;
	output \g63777/_3_  ;
	output \g63778/_3_  ;
	output \g63781/_0_  ;
	output \g63786/u3_syn_7  ;
	output \g63787/_3_  ;
	output \g63788/_3_  ;
	output \g63790/_3_  ;
	output \g63791/_3_  ;
	output \g63792/u3_syn_7  ;
	output \g63794/_0_  ;
	output \g63795/_0_  ;
	output \g63796/_0_  ;
	output \g63798/_3_  ;
	output \g63800/_3_  ;
	output \g63804/_3_  ;
	output \g63805/_3_  ;
	output \g63806/_3_  ;
	output \g63807/_3_  ;
	output \g63808/_3_  ;
	output \g63809/_3_  ;
	output \g63870/_0_  ;
	output \g63883/_0_  ;
	output \g63934/_0_  ;
	output \g63936/_0_  ;
	output \g63938/_0_  ;
	output \g63939/_0_  ;
	output \g63966/_0_  ;
	output \g63970/_0_  ;
	output \g63999/_0_  ;
	output \g64039/_0_  ;
	output \g64040/_0_  ;
	output \g64043/_0_  ;
	output \g64062/_3_  ;
	output \g64078/_0_  ;
	output \g64091/_0_  ;
	output \g64095/_3_  ;
	output \g64096/_3_  ;
	output \g64097/u3_syn_7  ;
	output \g64098/u3_syn_7  ;
	output \g64099/u3_syn_7  ;
	output \g64100/u3_syn_7  ;
	output \g64134/_0_  ;
	output \g64135/_0_  ;
	output \g64153/_0_  ;
	output \g64155/_0_  ;
	output \g64179/_0_  ;
	output \g64229/_0_  ;
	output \g64235/_0_  ;
	output \g64236/_0_  ;
	output \g64280/_0_  ;
	output \g64315/_0_  ;
	output \g64365/_0_  ;
	output \g64426/_3_  ;
	output \g64438/_3_  ;
	output \g64442/u3_syn_7  ;
	output \g64445/_3_  ;
	output \g64447/_3_  ;
	output \g64449/_3_  ;
	output \g64451/_3_  ;
	output \g64453/_3_  ;
	output \g64454/_3_  ;
	output \g64460/_3_  ;
	output \g64461/_3_  ;
	output \g64510/_0_  ;
	output \g64527/_0_  ;
	output \g64528/_0_  ;
	output \g64544/_0_  ;
	output \g64549/_0_  ;
	output \g64566/_0_  ;
	output \g64576/_0_  ;
	output \g64602/_0_  ;
	output \g64691/_0_  ;
	output \g64697/_0_  ;
	output \g64707/_3_  ;
	output \g64778/_3_  ;
	output \g64790/_3_  ;
	output \g64791/_3_  ;
	output \g64792/_3_  ;
	output \g64793/_3_  ;
	output \g64794/_3_  ;
	output \g64795/_3_  ;
	output \g64796/_3_  ;
	output \g64797/_3_  ;
	output \g64877/_0_  ;
	output \g64912/_0_  ;
	output \g64973/_0_  ;
	output \g65047/_3_  ;
	output \g65081/_3_  ;
	output \g65088/_3_  ;
	output \g65097/_3_  ;
	output \g65100/_3_  ;
	output \g65101/_3_  ;
	output \g65104/_3_  ;
	output \g65105/_3_  ;
	output \g65107/_3_  ;
	output \g65110/_3_  ;
	output \g65111/_3_  ;
	output \g65113/_3_  ;
	output \g65114/_3_  ;
	output \g65266/_0_  ;
	output \g65267/_0_  ;
	output \g65294/_1_  ;
	output \g65328/_1_  ;
	output \g65495/_0_  ;
	output \g65499/_0_  ;
	output \g65503/_0_  ;
	output \g65529/_0_  ;
	output \g65530/_3_  ;
	output \g65531/_3_  ;
	output \g65532/_3_  ;
	output \g65533/_3_  ;
	output \g65624/_0_  ;
	output \g65625/_1_  ;
	output \g65641/_0_  ;
	output \g65701/_0_  ;
	output \g65704/_0_  ;
	output \g65853/_0_  ;
	output \g65891/_0_  ;
	output \g65901/_0_  ;
	output \g65986/_0_  ;
	output \g66029/_0_  ;
	output \g66066/_0_  ;
	output \g66067/_0_  ;
	output \g66068/_0_  ;
	output \g66154/_3_  ;
	output \g66362/_0_  ;
	output \g66369/_0_  ;
	output \g66398/_0_  ;
	output \g66409/_0_  ;
	output \g66419/_0_  ;
	output \g66439/_0_  ;
	output \g66443/_0_  ;
	output \g66464/_0_  ;
	output \g66471/_0_  ;
	output \g66512/_0_  ;
	output \g66528/_0_  ;
	output \g66541/_0_  ;
	output \g66558/_0_  ;
	output \g66644/_0_  ;
	output \g66684/_0_  ;
	output \g66697/_0_  ;
	output \g66698/_0_  ;
	output \g66701/_0_  ;
	output \g66714/_0_  ;
	output \g66715/_0_  ;
	output \g66745/_0_  ;
	output \g66750/_0_  ;
	output \g66751/_0_  ;
	output \g66810/_0_  ;
	output \g66844/_0_  ;
	output \g66853/_0_  ;
	output \g66897/_0_  ;
	output \g66905/_0_  ;
	output \g69743/_0_  ;
	output \g69750/_0_  ;
	output \g69773/_1_  ;
	output \g69792/_1_  ;
	output \g69858/_0_  ;
	output \g69938/_0_  ;
	output \g69949/_0_  ;
	output \g70167/_0_  ;
	output \g71190/_0_  ;
	output \g71198/_0_  ;
	output \g71284/_0_  ;
	output \g72369/_1_  ;
	output \g72467/_0_  ;
	output \g72476/_0_  ;
	output \g72477/_1_  ;
	output \g72648/_0_  ;
	output \g72741/_0_  ;
	output \g72772/_0_  ;
	output \g8132_pad  ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1486_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1031_ ;
	wire _w1599_ ;
	wire _w490_ ;
	wire _w2847_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w1513_ ;
	wire _w404_ ;
	wire _w2761_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w1487_ ;
	wire _w378_ ;
	wire _w2735_ ;
	wire _w917_ ;
	wire _w1485_ ;
	wire _w376_ ;
	wire _w2733_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w792_ ;
	wire _w785_ ;
	wire _w918_ ;
	wire _w1004_ ;
	wire _w871_ ;
	wire _w781_ ;
	wire _w817_ ;
	wire _w788_ ;
	wire _w884_ ;
	wire _w789_ ;
	wire _w1009_ ;
	wire _w1604_ ;
	wire _w495_ ;
	wire _w2852_ ;
	wire _w1036_ ;
	wire _w876_ ;
	wire _w790_ ;
	wire _w886_ ;
	wire _w791_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w1016_ ;
	wire _w1611_ ;
	wire _w502_ ;
	wire _w2859_ ;
	wire _w1043_ ;
	wire _w883_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w885_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2734_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\g2831_reg/NET0131 ,
		_w376_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\g2834_reg/NET0131 ,
		_w378_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\g29221_pad ,
		_w404_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\g34_reg/NET0131 ,
		_w490_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\g35_pad ,
		_w495_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\g37_reg/NET0131 ,
		_w502_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\g3003_reg/NET0131 ,
		\g35_pad ,
		_w781_
	);
	LUT4 #(
		.INIT('h0001)
	) name7 (
		\g2255_reg/NET0131 ,
		\g2389_reg/NET0131 ,
		\g2523_reg/NET0131 ,
		\g2657_reg/NET0131 ,
		_w782_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		\g1696_reg/NET0131 ,
		\g1830_reg/NET0131 ,
		\g1964_reg/NET0131 ,
		\g2098_reg/NET0131 ,
		_w783_
	);
	LUT3 #(
		.INIT('hfd)
	) name9 (
		\g35_pad ,
		_w782_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\g1978_reg/NET0131 ,
		\g1992_reg/NET0131 ,
		\g2112_reg/NET0131 ,
		\g2126_reg/NET0131 ,
		_w785_
	);
	LUT4 #(
		.INIT('h0001)
	) name11 (
		\g1710_reg/NET0131 ,
		\g1724_reg/NET0131 ,
		\g1844_reg/NET0131 ,
		\g1858_reg/NET0131 ,
		_w786_
	);
	LUT3 #(
		.INIT('h2a)
	) name12 (
		\g35_pad ,
		_w785_,
		_w786_,
		_w787_
	);
	LUT4 #(
		.INIT('h0001)
	) name13 (
		\g2537_reg/NET0131 ,
		\g2551_reg/NET0131 ,
		\g2671_reg/NET0131 ,
		\g2685_reg/NET0131 ,
		_w788_
	);
	LUT4 #(
		.INIT('h0001)
	) name14 (
		\g2269_reg/NET0131 ,
		\g2283_reg/NET0131 ,
		\g2403_reg/NET0131 ,
		\g2417_reg/NET0131 ,
		_w789_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('hd)
	) name16 (
		_w787_,
		_w790_,
		_w791_
	);
	LUT4 #(
		.INIT('h0001)
	) name17 (
		\g2472_reg/NET0131 ,
		\g2491_reg/NET0131 ,
		\g2606_reg/NET0131 ,
		\g2625_reg/NET0131 ,
		_w792_
	);
	LUT4 #(
		.INIT('h0001)
	) name18 (
		\g2204_reg/NET0131 ,
		\g2223_reg/NET0131 ,
		\g2338_reg/NET0131 ,
		\g2357_reg/NET0131 ,
		_w793_
	);
	LUT3 #(
		.INIT('h2a)
	) name19 (
		\g35_pad ,
		_w792_,
		_w793_,
		_w794_
	);
	LUT4 #(
		.INIT('h0001)
	) name20 (
		\g1913_reg/NET0131 ,
		\g1932_reg/NET0131 ,
		\g2047_reg/NET0131 ,
		\g2066_reg/NET0131 ,
		_w795_
	);
	LUT4 #(
		.INIT('h0001)
	) name21 (
		\g1644_reg/NET0131 ,
		\g1664_reg/NET0131 ,
		\g1779_reg/NET0131 ,
		\g1798_reg/NET0131 ,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('hd)
	) name23 (
		_w794_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\g1312_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w799_
	);
	LUT3 #(
		.INIT('he0)
	) name25 (
		\g1312_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\g1008_reg/NET0131 ,
		\g969_reg/NET0131 ,
		_w801_
	);
	LUT3 #(
		.INIT('hc8)
	) name27 (
		\g1008_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		\g969_reg/NET0131 ,
		_w802_
	);
	LUT4 #(
		.INIT('h3070)
	) name28 (
		\g1008_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		\g35_pad ,
		\g969_reg/NET0131 ,
		_w803_
	);
	LUT2 #(
		.INIT('hb)
	) name29 (
		_w800_,
		_w803_,
		_w804_
	);
	LUT3 #(
		.INIT('hfb)
	) name30 (
		\g1306_reg/NET0131 ,
		\g35_pad ,
		\g962_reg/NET0131 ,
		_w805_
	);
	LUT4 #(
		.INIT('h0001)
	) name31 (
		\g3115_reg/NET0131 ,
		\g3466_reg/NET0131 ,
		\g3817_reg/NET0131 ,
		\g5124_reg/NET0131 ,
		_w806_
	);
	LUT2 #(
		.INIT('hd)
	) name32 (
		\g35_pad ,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\g5297_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w808_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\g1636_reg/NET0131 ,
		\g1668_reg/NET0131 ,
		_w809_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\g1648_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\g2902_reg/NET0131 ,
		\g2907_reg/NET0131 ,
		_w811_
	);
	LUT4 #(
		.INIT('h0777)
	) name37 (
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		\g2936_reg/NET0131 ,
		\g2941_reg/NET0131 ,
		_w812_
	);
	LUT4 #(
		.INIT('h0777)
	) name38 (
		\g2960_reg/NET0131 ,
		\g2965_reg/NET0131 ,
		\g2970_reg/NET0131 ,
		\g2975_reg/NET0131 ,
		_w813_
	);
	LUT4 #(
		.INIT('h0777)
	) name39 (
		\g2922_reg/NET0131 ,
		\g2927_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		\g2955_reg/NET0131 ,
		_w814_
	);
	LUT4 #(
		.INIT('h4000)
	) name40 (
		_w811_,
		_w812_,
		_w813_,
		_w814_,
		_w815_
	);
	LUT4 #(
		.INIT('h048c)
	) name41 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2815_reg/NET0131 ,
		\g2819_reg/NET0131 ,
		_w816_
	);
	LUT4 #(
		.INIT('h0123)
	) name42 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2803_reg/NET0131 ,
		\g2807_reg/NET0131 ,
		_w817_
	);
	LUT2 #(
		.INIT('he)
	) name43 (
		_w816_,
		_w817_,
		_w818_
	);
	LUT4 #(
		.INIT('h048c)
	) name44 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		_w819_
	);
	LUT4 #(
		.INIT('h0123)
	) name45 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2771_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		_w820_
	);
	LUT2 #(
		.INIT('he)
	) name46 (
		_w819_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w822_
	);
	LUT3 #(
		.INIT('h02)
	) name48 (
		\g4698_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w823_
	);
	LUT3 #(
		.INIT('h02)
	) name49 (
		\g4776_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		\g4801_reg/NET0131 ,
		_w824_
	);
	LUT3 #(
		.INIT('h80)
	) name50 (
		\g4653_reg/NET0131 ,
		\g4659_reg/NET0131 ,
		\g4669_reg/NET0131 ,
		_w825_
	);
	LUT3 #(
		.INIT('h80)
	) name51 (
		_w823_,
		_w824_,
		_w825_,
		_w826_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name52 (
		\g4646_reg/NET0131 ,
		_w823_,
		_w824_,
		_w825_,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		_w828_
	);
	LUT4 #(
		.INIT('h1110)
	) name54 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		\g4082_reg/NET0131 ,
		\g4141_reg/NET0131 ,
		_w829_
	);
	LUT3 #(
		.INIT('h01)
	) name55 (
		\g4087_reg/NET0131 ,
		\g4093_reg/NET0131 ,
		\g4098_reg/NET0131 ,
		_w830_
	);
	LUT4 #(
		.INIT('h1000)
	) name56 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		\g4076_reg/NET0131 ,
		\g4112_reg/NET0131 ,
		_w831_
	);
	LUT3 #(
		.INIT('hea)
	) name57 (
		_w829_,
		_w830_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('h0002)
	) name58 (
		\g479_reg/NET0131 ,
		\g482_reg/NET0131 ,
		\g490_reg/NET0131 ,
		\g528_reg/NET0131 ,
		_w833_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\g890_reg/NET0131 ,
		_w833_,
		_w834_
	);
	LUT4 #(
		.INIT('h0001)
	) name60 (
		\g4311_reg/NET0131 ,
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		\g4366_reg/NET0131 ,
		_w835_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\g4369_reg/NET0131 ,
		_w835_,
		_w836_
	);
	LUT4 #(
		.INIT('h153f)
	) name62 (
		\g16624_pad ,
		\g16686_pad ,
		\g3247_reg/NET0131 ,
		\g3263_reg/NET0131 ,
		_w837_
	);
	LUT4 #(
		.INIT('h135f)
	) name63 (
		\g16874_pad ,
		\g3207_reg/NET0131 ,
		\g3223_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		_w838_
	);
	LUT3 #(
		.INIT('hd8)
	) name64 (
		\g3338_reg/NET0131 ,
		_w837_,
		_w838_,
		_w839_
	);
	LUT4 #(
		.INIT('h8008)
	) name65 (
		\g16718_pad ,
		\g3235_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w840_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\g3990_reg/NET0131 ,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w839_,
		_w841_,
		_w842_
	);
	LUT4 #(
		.INIT('h135f)
	) name68 (
		\g16874_pad ,
		\g3191_reg/NET0131 ,
		\g3215_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		_w843_
	);
	LUT4 #(
		.INIT('h135f)
	) name69 (
		\g16624_pad ,
		\g16686_pad ,
		\g3203_reg/NET0131 ,
		\g3255_reg/NET0131 ,
		_w844_
	);
	LUT3 #(
		.INIT('hd8)
	) name70 (
		\g3338_reg/NET0131 ,
		_w843_,
		_w844_,
		_w845_
	);
	LUT4 #(
		.INIT('h0880)
	) name71 (
		\g16718_pad ,
		\g3243_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w846_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\g3990_reg/NET0131 ,
		_w846_,
		_w847_
	);
	LUT3 #(
		.INIT('h2a)
	) name73 (
		\g4054_reg/NET0131 ,
		_w845_,
		_w847_,
		_w848_
	);
	LUT4 #(
		.INIT('h0770)
	) name74 (
		\g16603_pad ,
		\g3259_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w849_
	);
	LUT4 #(
		.INIT('h7007)
	) name75 (
		\g13895_pad ,
		\g3219_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w850_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w849_,
		_w850_,
		_w851_
	);
	LUT4 #(
		.INIT('h0777)
	) name77 (
		\g13039_pad ,
		\g3199_reg/NET0131 ,
		\g3211_reg/NET0131 ,
		\g3329_reg/NET0131 ,
		_w852_
	);
	LUT4 #(
		.INIT('h7f00)
	) name78 (
		\g13865_pad ,
		\g3231_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g3990_reg/NET0131 ,
		_w853_
	);
	LUT3 #(
		.INIT('he0)
	) name79 (
		\g3338_reg/NET0131 ,
		_w852_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w851_,
		_w854_,
		_w855_
	);
	LUT4 #(
		.INIT('h0770)
	) name81 (
		\g13895_pad ,
		\g3227_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w856_
	);
	LUT4 #(
		.INIT('h7007)
	) name82 (
		\g16603_pad ,
		\g3251_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w856_,
		_w857_,
		_w858_
	);
	LUT4 #(
		.INIT('h0777)
	) name84 (
		\g13039_pad ,
		\g3187_reg/NET0131 ,
		\g3195_reg/NET0131 ,
		\g3329_reg/NET0131 ,
		_w859_
	);
	LUT4 #(
		.INIT('h00f7)
	) name85 (
		\g13865_pad ,
		\g3239_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g3990_reg/NET0131 ,
		_w860_
	);
	LUT3 #(
		.INIT('hd0)
	) name86 (
		\g3338_reg/NET0131 ,
		_w859_,
		_w860_,
		_w861_
	);
	LUT3 #(
		.INIT('h45)
	) name87 (
		\g4054_reg/NET0131 ,
		_w858_,
		_w861_,
		_w862_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name88 (
		_w842_,
		_w848_,
		_w855_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w864_
	);
	LUT3 #(
		.INIT('h80)
	) name90 (
		\g4709_reg/NET0131 ,
		\g4765_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w865_
	);
	LUT3 #(
		.INIT('h80)
	) name91 (
		_w824_,
		_w825_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		\g35_pad ,
		\g4688_reg/NET0131 ,
		_w867_
	);
	LUT4 #(
		.INIT('h7f00)
	) name93 (
		_w824_,
		_w825_,
		_w865_,
		_w867_,
		_w868_
	);
	LUT4 #(
		.INIT('h8000)
	) name94 (
		\g16624_pad ,
		\g3338_reg/NET0131 ,
		\g3990_reg/NET0131 ,
		\g4054_reg/NET0131 ,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\g3808_reg/NET0131 ,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		_w868_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w868_,
		_w870_,
		_w872_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\g3111_reg/NET0131 ,
		\g35_pad ,
		_w873_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\g35_pad ,
		\g4688_reg/NET0131 ,
		_w874_
	);
	LUT4 #(
		.INIT('h8000)
	) name100 (
		\g35_pad ,
		\g4709_reg/NET0131 ,
		\g4765_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w875_
	);
	LUT4 #(
		.INIT('h070f)
	) name101 (
		_w824_,
		_w825_,
		_w874_,
		_w875_,
		_w876_
	);
	LUT3 #(
		.INIT('h31)
	) name102 (
		\g3808_reg/NET0131 ,
		_w873_,
		_w876_,
		_w877_
	);
	LUT4 #(
		.INIT('he4ff)
	) name103 (
		_w863_,
		_w871_,
		_w872_,
		_w877_,
		_w878_
	);
	LUT3 #(
		.INIT('h01)
	) name104 (
		\g482_reg/NET0131 ,
		\g490_reg/NET0131 ,
		\g528_reg/NET0131 ,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\g499_reg/NET0131 ,
		\g518_reg/NET0131 ,
		_w880_
	);
	LUT4 #(
		.INIT('h0111)
	) name106 (
		\g499_reg/NET0131 ,
		\g518_reg/NET0131 ,
		\g554_reg/NET0131 ,
		\g807_reg/NET0131 ,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w879_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		\g736_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w883_
	);
	LUT4 #(
		.INIT('h80c0)
	) name109 (
		\g736_reg/NET0131 ,
		\g749_reg/NET0131 ,
		\g758_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w884_
	);
	LUT4 #(
		.INIT('h8000)
	) name110 (
		\g739_reg/NET0131 ,
		\g744_reg/NET0131 ,
		\g763_reg/NET0131 ,
		\g767_reg/NET0131 ,
		_w885_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		_w886_
	);
	LUT4 #(
		.INIT('h8088)
	) name112 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g736_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w887_
	);
	LUT3 #(
		.INIT('h80)
	) name113 (
		_w884_,
		_w885_,
		_w887_,
		_w888_
	);
	LUT3 #(
		.INIT('h80)
	) name114 (
		\g655_reg/NET0131 ,
		\g718_reg/NET0131 ,
		\g753_reg/NET0131 ,
		_w889_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		\g370_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w890_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\g12184_pad ,
		\g802_reg/NET0131 ,
		_w891_
	);
	LUT3 #(
		.INIT('h01)
	) name117 (
		\g655_reg/NET0131 ,
		\g718_reg/NET0131 ,
		\g753_reg/NET0131 ,
		_w892_
	);
	LUT4 #(
		.INIT('h0004)
	) name118 (
		_w889_,
		_w890_,
		_w891_,
		_w892_,
		_w893_
	);
	LUT3 #(
		.INIT('h8c)
	) name119 (
		\g736_reg/NET0131 ,
		\g772_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w894_
	);
	LUT4 #(
		.INIT('h80c0)
	) name120 (
		\g736_reg/NET0131 ,
		\g772_reg/NET0131 ,
		\g776_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w895_
	);
	LUT4 #(
		.INIT('h8000)
	) name121 (
		_w882_,
		_w888_,
		_w893_,
		_w895_,
		_w896_
	);
	LUT3 #(
		.INIT('h8c)
	) name122 (
		\g736_reg/NET0131 ,
		\g785_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w897_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\g781_reg/NET0131 ,
		\g790_reg/NET0131 ,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w897_,
		_w898_,
		_w899_
	);
	LUT3 #(
		.INIT('h80)
	) name125 (
		\g794_reg/NET0131 ,
		_w897_,
		_w898_,
		_w900_
	);
	LUT4 #(
		.INIT('h8a00)
	) name126 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g802_reg/NET0131 ,
		\g807_reg/NET0131 ,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\g554_reg/NET0131 ,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w900_,
		_w902_,
		_w903_
	);
	LUT4 #(
		.INIT('h8088)
	) name129 (
		\g35_pad ,
		\g554_reg/NET0131 ,
		\g736_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w904_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		\g35_pad ,
		\g807_reg/NET0131 ,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w904_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('h8f)
	) name132 (
		_w896_,
		_w903_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\g2941_reg/NET0131 ,
		\g35_pad ,
		_w908_
	);
	LUT3 #(
		.INIT('h80)
	) name134 (
		\g35_pad ,
		_w782_,
		_w783_,
		_w909_
	);
	LUT4 #(
		.INIT('h0001)
	) name135 (
		\g2946_reg/NET0131 ,
		\g2955_reg/NET0131 ,
		\g4420_reg/NET0131 ,
		\g4427_reg/NET0131 ,
		_w910_
	);
	LUT4 #(
		.INIT('h8000)
	) name136 (
		_w785_,
		_w786_,
		_w806_,
		_w910_,
		_w911_
	);
	LUT4 #(
		.INIT('h0001)
	) name137 (
		\g3831_reg/NET0131 ,
		\g3845_reg/NET0131 ,
		\g5138_reg/NET0131 ,
		\g5152_reg/NET0131 ,
		_w912_
	);
	LUT4 #(
		.INIT('h0001)
	) name138 (
		\g3129_reg/NET0131 ,
		\g3143_reg/NET0131 ,
		\g3480_reg/NET0131 ,
		\g3494_reg/NET0131 ,
		_w913_
	);
	LUT4 #(
		.INIT('h8000)
	) name139 (
		_w788_,
		_w789_,
		_w912_,
		_w913_,
		_w914_
	);
	LUT4 #(
		.INIT('h1555)
	) name140 (
		_w908_,
		_w909_,
		_w911_,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		\g2856_reg/NET0131 ,
		\g35_pad ,
		_w916_
	);
	LUT4 #(
		.INIT('h0004)
	) name142 (
		\g2864_reg/NET0131 ,
		\g35_pad ,
		\g4420_reg/NET0131 ,
		\g4427_reg/NET0131 ,
		_w917_
	);
	LUT3 #(
		.INIT('h13)
	) name143 (
		_w806_,
		_w916_,
		_w917_,
		_w918_
	);
	LUT3 #(
		.INIT('h78)
	) name144 (
		\g10306_pad ,
		\g35_pad ,
		\g4534_reg/NET0131 ,
		_w919_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		\g35_pad ,
		\g4564_reg/NET0131 ,
		_w920_
	);
	LUT4 #(
		.INIT('h8000)
	) name146 (
		\g4555_reg/NET0131 ,
		\g4558_reg/NET0131 ,
		\g4561_reg/NET0131 ,
		\g4564_reg/NET0131 ,
		_w921_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\g2988_reg/NET0131 ,
		\g35_pad ,
		_w922_
	);
	LUT3 #(
		.INIT('hfe)
	) name148 (
		_w920_,
		_w921_,
		_w922_,
		_w923_
	);
	LUT3 #(
		.INIT('hb8)
	) name149 (
		\g18096_pad ,
		\g35_pad ,
		\g4561_reg/NET0131 ,
		_w924_
	);
	LUT3 #(
		.INIT('hb8)
	) name150 (
		\g18095_pad ,
		\g35_pad ,
		\g4558_reg/NET0131 ,
		_w925_
	);
	LUT3 #(
		.INIT('hb8)
	) name151 (
		\g18094_pad ,
		\g35_pad ,
		\g4555_reg/NET0131 ,
		_w926_
	);
	LUT4 #(
		.INIT('h8000)
	) name152 (
		\g4483_reg/NET0131 ,
		\g4486_reg/NET0131 ,
		\g4489_reg/NET0131 ,
		\g4492_reg/NET0131 ,
		_w927_
	);
	LUT4 #(
		.INIT('h4cc4)
	) name153 (
		\g35_pad ,
		\g4521_reg/NET0131 ,
		\g4527_reg/NET0131 ,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name154 (
		\g4584_reg/NET0131 ,
		\g4593_reg/NET0131 ,
		\g4601_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		_w929_
	);
	LUT4 #(
		.INIT('h1108)
	) name155 (
		\g4584_reg/NET0131 ,
		\g4593_reg/NET0131 ,
		\g4601_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		_w930_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\g35_pad ,
		\g4521_reg/NET0131 ,
		_w931_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w930_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		\g4593_reg/NET0131 ,
		\g4601_reg/NET0131 ,
		_w933_
	);
	LUT3 #(
		.INIT('h0d)
	) name159 (
		\g4584_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		\g4616_reg/NET0131 ,
		_w934_
	);
	LUT4 #(
		.INIT('h0800)
	) name160 (
		_w929_,
		_w931_,
		_w933_,
		_w934_,
		_w935_
	);
	LUT3 #(
		.INIT('hfe)
	) name161 (
		_w928_,
		_w932_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\g35_pad ,
		\g4527_reg/NET0131 ,
		_w937_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name163 (
		\g35_pad ,
		\g4515_reg/NET0131 ,
		\g4521_reg/NET0131 ,
		\g4527_reg/NET0131 ,
		_w938_
	);
	LUT4 #(
		.INIT('heb00)
	) name164 (
		\g4521_reg/NET0131 ,
		\g4527_reg/NET0131 ,
		_w927_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w937_,
		_w939_,
		_w940_
	);
	LUT3 #(
		.INIT('h80)
	) name166 (
		\g35_pad ,
		\g4572_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w941_
	);
	LUT4 #(
		.INIT('haf27)
	) name167 (
		\g35_pad ,
		\g4512_reg/NET0131 ,
		\g4515_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w942_
	);
	LUT2 #(
		.INIT('hb)
	) name168 (
		_w941_,
		_w942_,
		_w943_
	);
	LUT4 #(
		.INIT('he4cc)
	) name169 (
		\g35_pad ,
		\g4552_reg/NET0131 ,
		\g4575_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w944_
	);
	LUT4 #(
		.INIT('h4eee)
	) name170 (
		\g35_pad ,
		\g4512_reg/NET0131 ,
		\g4531_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w945_
	);
	LUT2 #(
		.INIT('h6)
	) name171 (
		\g1322_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w946_
	);
	LUT4 #(
		.INIT('h6606)
	) name172 (
		\g1322_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		\g1312_reg/NET0131 ,
		_w947_,
		_w948_
	);
	LUT3 #(
		.INIT('h80)
	) name174 (
		\g1351_reg/NET0131 ,
		\g1361_reg/NET0131 ,
		\g1373_reg/NET0131 ,
		_w949_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		\g1345_reg/NET0131 ,
		\g1361_reg/NET0131 ,
		_w950_
	);
	LUT3 #(
		.INIT('h80)
	) name176 (
		\g1345_reg/NET0131 ,
		\g1361_reg/NET0131 ,
		\g1367_reg/NET0131 ,
		_w951_
	);
	LUT3 #(
		.INIT('h0b)
	) name177 (
		_w946_,
		_w949_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\g1312_reg/NET0131 ,
		\g1373_reg/NET0131 ,
		_w954_
	);
	LUT3 #(
		.INIT('h23)
	) name180 (
		_w947_,
		_w953_,
		_w954_,
		_w955_
	);
	LUT3 #(
		.INIT('h70)
	) name181 (
		_w948_,
		_w952_,
		_w955_,
		_w956_
	);
	LUT3 #(
		.INIT('h45)
	) name182 (
		\g1379_reg/NET0131 ,
		_w946_,
		_w949_,
		_w957_
	);
	LUT3 #(
		.INIT('h2a)
	) name183 (
		\g35_pad ,
		_w948_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		\g1379_reg/NET0131 ,
		\g35_pad ,
		_w959_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\g1373_reg/NET0131 ,
		\g35_pad ,
		_w960_
	);
	LUT4 #(
		.INIT('h0027)
	) name186 (
		_w956_,
		_w958_,
		_w959_,
		_w960_,
		_w961_
	);
	LUT4 #(
		.INIT('h6aca)
	) name187 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g35_pad ,
		\g7946_pad ,
		_w962_
	);
	LUT4 #(
		.INIT('h0800)
	) name188 (
		\g1339_reg/NET0131 ,
		\g1521_reg/NET0131 ,
		\g1532_reg/NET0131 ,
		\g7946_pad ,
		_w963_
	);
	LUT3 #(
		.INIT('ha4)
	) name189 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w964_
	);
	LUT3 #(
		.INIT('h80)
	) name190 (
		\g1345_reg/NET0131 ,
		\g1367_reg/NET0131 ,
		\g1379_reg/NET0131 ,
		_w965_
	);
	LUT4 #(
		.INIT('h3bbb)
	) name191 (
		_w799_,
		_w963_,
		_w964_,
		_w965_,
		_w966_
	);
	LUT3 #(
		.INIT('hb0)
	) name192 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		_w967_
	);
	LUT4 #(
		.INIT('h4f0a)
	) name193 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		\g35_pad ,
		_w968_
	);
	LUT3 #(
		.INIT('hba)
	) name194 (
		_w962_,
		_w966_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		\g1367_reg/NET0131 ,
		\g35_pad ,
		_w970_
	);
	LUT4 #(
		.INIT('h5540)
	) name196 (
		\g1373_reg/NET0131 ,
		_w948_,
		_w952_,
		_w953_,
		_w971_
	);
	LUT4 #(
		.INIT('h80aa)
	) name197 (
		\g35_pad ,
		_w948_,
		_w952_,
		_w955_,
		_w972_
	);
	LUT3 #(
		.INIT('hba)
	) name198 (
		_w970_,
		_w971_,
		_w972_,
		_w973_
	);
	LUT4 #(
		.INIT('he4cc)
	) name199 (
		\g35_pad ,
		\g4549_reg/NET0131 ,
		\g4575_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w974_
	);
	LUT3 #(
		.INIT('h48)
	) name200 (
		\g1514_reg/NET0131 ,
		\g35_pad ,
		\g7946_pad ,
		_w975_
	);
	LUT4 #(
		.INIT('h4f00)
	) name201 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		\g35_pad ,
		_w976_
	);
	LUT3 #(
		.INIT('hdc)
	) name202 (
		_w966_,
		_w975_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('h00e0)
	) name203 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g1367_reg/NET0131 ,
		_w978_
	);
	LUT3 #(
		.INIT('hb0)
	) name204 (
		_w946_,
		_w949_,
		_w978_,
		_w979_
	);
	LUT4 #(
		.INIT('ha222)
	) name205 (
		\g1361_reg/NET0131 ,
		\g35_pad ,
		_w948_,
		_w979_,
		_w980_
	);
	LUT3 #(
		.INIT('h0b)
	) name206 (
		_w946_,
		_w949_,
		_w950_,
		_w981_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\g1367_reg/NET0131 ,
		\g35_pad ,
		_w982_
	);
	LUT4 #(
		.INIT('hec00)
	) name208 (
		_w948_,
		_w953_,
		_w981_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('he)
	) name209 (
		_w980_,
		_w983_,
		_w984_
	);
	LUT3 #(
		.INIT('h08)
	) name210 (
		\g1339_reg/NET0131 ,
		\g1521_reg/NET0131 ,
		\g1532_reg/NET0131 ,
		_w985_
	);
	LUT4 #(
		.INIT('h4000)
	) name211 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g1542_reg/NET0131 ,
		\g7946_pad ,
		_w986_
	);
	LUT3 #(
		.INIT('h8a)
	) name212 (
		\g35_pad ,
		_w985_,
		_w986_,
		_w987_
	);
	LUT4 #(
		.INIT('h8088)
	) name213 (
		\g1413_reg/NET0131 ,
		\g35_pad ,
		_w985_,
		_w986_,
		_w988_
	);
	LUT4 #(
		.INIT('h1000)
	) name214 (
		\g1413_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g7946_pad ,
		_w989_
	);
	LUT4 #(
		.INIT('h2a22)
	) name215 (
		\g1542_reg/NET0131 ,
		\g35_pad ,
		_w985_,
		_w989_,
		_w990_
	);
	LUT4 #(
		.INIT('hffe0)
	) name216 (
		_w966_,
		_w967_,
		_w988_,
		_w990_,
		_w991_
	);
	LUT3 #(
		.INIT('h08)
	) name217 (
		\g13272_pad ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		\g1442_reg/NET0131 ,
		\g1489_reg/NET0131 ,
		_w993_
	);
	LUT3 #(
		.INIT('h15)
	) name219 (
		\g1437_reg/NET0131 ,
		_w992_,
		_w993_,
		_w994_
	);
	LUT4 #(
		.INIT('h3200)
	) name220 (
		\g1312_reg/NET0131 ,
		\g1319_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		_w995_
	);
	LUT4 #(
		.INIT('h0020)
	) name221 (
		\g13272_pad ,
		\g1478_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w996_
	);
	LUT4 #(
		.INIT('h0080)
	) name222 (
		\g13272_pad ,
		\g1478_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w997_
	);
	LUT3 #(
		.INIT('h1b)
	) name223 (
		_w995_,
		_w996_,
		_w997_,
		_w998_
	);
	LUT4 #(
		.INIT('h2e22)
	) name224 (
		\g1442_reg/NET0131 ,
		\g35_pad ,
		_w994_,
		_w998_,
		_w999_
	);
	LUT3 #(
		.INIT('h20)
	) name225 (
		\g13272_pad ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1000_
	);
	LUT3 #(
		.INIT('h15)
	) name226 (
		\g1454_reg/NET0131 ,
		_w993_,
		_w1000_,
		_w1001_
	);
	LUT4 #(
		.INIT('h0200)
	) name227 (
		\g13272_pad ,
		\g1448_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1002_
	);
	LUT4 #(
		.INIT('h0800)
	) name228 (
		\g13272_pad ,
		\g1448_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1003_
	);
	LUT3 #(
		.INIT('h1b)
	) name229 (
		_w995_,
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT4 #(
		.INIT('h2e22)
	) name230 (
		\g1478_reg/NET0131 ,
		\g35_pad ,
		_w1001_,
		_w1004_,
		_w1005_
	);
	LUT3 #(
		.INIT('h80)
	) name231 (
		\g13272_pad ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1006_
	);
	LUT3 #(
		.INIT('h15)
	) name232 (
		\g1467_reg/NET0131 ,
		_w993_,
		_w1006_,
		_w1007_
	);
	LUT4 #(
		.INIT('h2000)
	) name233 (
		\g13272_pad ,
		\g1472_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1008_
	);
	LUT4 #(
		.INIT('h8000)
	) name234 (
		\g13272_pad ,
		\g1472_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1009_
	);
	LUT3 #(
		.INIT('h1b)
	) name235 (
		_w995_,
		_w1008_,
		_w1009_,
		_w1010_
	);
	LUT4 #(
		.INIT('h2e22)
	) name236 (
		\g1448_reg/NET0131 ,
		\g35_pad ,
		_w1007_,
		_w1010_,
		_w1011_
	);
	LUT3 #(
		.INIT('h02)
	) name237 (
		\g13272_pad ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1012_
	);
	LUT3 #(
		.INIT('h15)
	) name238 (
		\g1484_reg/NET0131 ,
		_w993_,
		_w1012_,
		_w1013_
	);
	LUT4 #(
		.INIT('h0004)
	) name239 (
		\g1300_reg/NET0131 ,
		\g13272_pad ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1014_
	);
	LUT4 #(
		.INIT('h0008)
	) name240 (
		\g1300_reg/NET0131 ,
		\g13272_pad ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1015_
	);
	LUT3 #(
		.INIT('h1b)
	) name241 (
		_w995_,
		_w1014_,
		_w1015_,
		_w1016_
	);
	LUT4 #(
		.INIT('h2e22)
	) name242 (
		\g1472_reg/NET0131 ,
		\g35_pad ,
		_w1013_,
		_w1016_,
		_w1017_
	);
	LUT4 #(
		.INIT('he4cc)
	) name243 (
		\g35_pad ,
		\g4504_reg/NET0131 ,
		\g4572_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1018_
	);
	LUT3 #(
		.INIT('h45)
	) name244 (
		\g1345_reg/NET0131 ,
		_w946_,
		_w949_,
		_w1019_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		\g1361_reg/NET0131 ,
		\g35_pad ,
		_w1020_
	);
	LUT4 #(
		.INIT('hec00)
	) name246 (
		_w948_,
		_w953_,
		_w1019_,
		_w1020_,
		_w1021_
	);
	LUT3 #(
		.INIT('h0e)
	) name247 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1361_reg/NET0131 ,
		_w1022_
	);
	LUT3 #(
		.INIT('hb0)
	) name248 (
		_w946_,
		_w949_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('ha222)
	) name249 (
		\g1345_reg/NET0131 ,
		\g35_pad ,
		_w948_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('he)
	) name250 (
		_w1021_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\g1532_reg/NET0131 ,
		\g35_pad ,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		\g1413_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		_w1027_
	);
	LUT4 #(
		.INIT('h2000)
	) name253 (
		\g35_pad ,
		_w985_,
		_w986_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		\g1536_reg/NET0131 ,
		\g35_pad ,
		_w1029_
	);
	LUT4 #(
		.INIT('h0103)
	) name255 (
		_w966_,
		_w1026_,
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		\g1536_reg/NET0131 ,
		\g35_pad ,
		_w1031_
	);
	LUT3 #(
		.INIT('h40)
	) name257 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g7946_pad ,
		_w1032_
	);
	LUT3 #(
		.INIT('h45)
	) name258 (
		\g1542_reg/NET0131 ,
		_w985_,
		_w1032_,
		_w1033_
	);
	LUT4 #(
		.INIT('h00e0)
	) name259 (
		_w966_,
		_w967_,
		_w987_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('he)
	) name260 (
		_w1031_,
		_w1034_,
		_w1035_
	);
	LUT4 #(
		.INIT('h040f)
	) name261 (
		\g333_reg/NET0131 ,
		\g351_reg/NET0131 ,
		\g355_reg/NET0131 ,
		\g35_pad ,
		_w1036_
	);
	LUT3 #(
		.INIT('h10)
	) name262 (
		\g29211_pad ,
		\g351_reg/NET0131 ,
		\g35_pad ,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('h2000)
	) name264 (
		\g1345_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		\g1367_reg/NET0131 ,
		\g1379_reg/NET0131 ,
		_w1039_
	);
	LUT3 #(
		.INIT('h10)
	) name265 (
		_w946_,
		_w953_,
		_w1039_,
		_w1040_
	);
	LUT3 #(
		.INIT('h60)
	) name266 (
		\g1322_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w1041_
	);
	LUT3 #(
		.INIT('h02)
	) name267 (
		_w949_,
		_w953_,
		_w1041_,
		_w1042_
	);
	LUT4 #(
		.INIT('h8a22)
	) name268 (
		\g1312_reg/NET0131 ,
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w1043_
	);
	LUT4 #(
		.INIT('haaa8)
	) name269 (
		\g35_pad ,
		_w1040_,
		_w1042_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		\g1312_reg/NET0131 ,
		\g35_pad ,
		_w1045_
	);
	LUT4 #(
		.INIT('h2088)
	) name271 (
		\g1312_reg/NET0131 ,
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w1045_,
		_w1046_,
		_w1047_
	);
	LUT4 #(
		.INIT('he000)
	) name273 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1361_reg/NET0131 ,
		\g1373_reg/NET0131 ,
		_w1048_
	);
	LUT4 #(
		.INIT('h4a00)
	) name274 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w1049_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\g1351_reg/NET0131 ,
		\g35_pad ,
		_w1050_
	);
	LUT3 #(
		.INIT('h10)
	) name276 (
		_w1048_,
		_w1049_,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('hd)
	) name277 (
		_w1047_,
		_w1051_,
		_w1052_
	);
	LUT4 #(
		.INIT('h32cc)
	) name278 (
		\g333_reg/NET0131 ,
		\g351_reg/NET0131 ,
		\g355_reg/NET0131 ,
		\g35_pad ,
		_w1053_
	);
	LUT3 #(
		.INIT('hec)
	) name279 (
		\g35_pad ,
		\g4546_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1054_
	);
	LUT4 #(
		.INIT('h0054)
	) name280 (
		\g1312_reg/NET0131 ,
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w1055_
	);
	LUT2 #(
		.INIT('h9)
	) name281 (
		\g1322_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		_w1056_
	);
	LUT3 #(
		.INIT('h08)
	) name282 (
		_w946_,
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT3 #(
		.INIT('h01)
	) name283 (
		\g1333_reg/NET0131 ,
		\g19357_pad ,
		\g7946_pad ,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		\g13272_pad ,
		\g8475_pad ,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name286 (
		\g1339_reg/NET0131 ,
		\g35_pad ,
		_w1057_,
		_w1060_,
		_w1061_
	);
	LUT3 #(
		.INIT('h60)
	) name287 (
		\g1322_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		\g35_pad ,
		_w1062_
	);
	LUT4 #(
		.INIT('h1555)
	) name288 (
		\g1333_reg/NET0131 ,
		_w946_,
		_w1055_,
		_w1062_,
		_w1063_
	);
	LUT4 #(
		.INIT('h4800)
	) name289 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		\g35_pad ,
		_w1064_
	);
	LUT3 #(
		.INIT('h80)
	) name290 (
		_w946_,
		_w1055_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w1063_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		\g1351_reg/NET0131 ,
		\g35_pad ,
		_w1067_
	);
	LUT4 #(
		.INIT('hfe00)
	) name293 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g35_pad ,
		_w1068_
	);
	LUT4 #(
		.INIT('hec00)
	) name294 (
		_w948_,
		_w953_,
		_w1019_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('he)
	) name295 (
		_w1067_,
		_w1069_,
		_w1070_
	);
	LUT3 #(
		.INIT('h01)
	) name296 (
		\g4411_reg/NET0131 ,
		\g7243_pad ,
		\g7257_pad ,
		_w1071_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		\g4375_reg/NET0131 ,
		\g4405_reg/NET0131 ,
		_w1072_
	);
	LUT4 #(
		.INIT('h0002)
	) name298 (
		\g35_pad ,
		\g4375_reg/NET0131 ,
		\g4392_reg/NET0131 ,
		\g4405_reg/NET0131 ,
		_w1073_
	);
	LUT3 #(
		.INIT('h40)
	) name299 (
		\g4417_reg/NET0131 ,
		_w1071_,
		_w1073_,
		_w1074_
	);
	LUT3 #(
		.INIT('h28)
	) name300 (
		\g35_pad ,
		\g4375_reg/NET0131 ,
		\g4382_reg/NET0131 ,
		_w1075_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		\g35_pad ,
		\g4388_reg/NET0131 ,
		_w1076_
	);
	LUT4 #(
		.INIT('h008f)
	) name302 (
		_w1071_,
		_w1072_,
		_w1075_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('hb)
	) name303 (
		_w1074_,
		_w1077_,
		_w1078_
	);
	LUT3 #(
		.INIT('h20)
	) name304 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		\g1099_reg/NET0131 ,
		\g1146_reg/NET0131 ,
		_w1080_
	);
	LUT3 #(
		.INIT('h15)
	) name306 (
		\g1094_reg/NET0131 ,
		_w1079_,
		_w1080_,
		_w1081_
	);
	LUT4 #(
		.INIT('h00c8)
	) name307 (
		\g1008_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		\g969_reg/NET0131 ,
		\g976_reg/NET0131 ,
		_w1082_
	);
	LUT4 #(
		.INIT('h0400)
	) name308 (
		\g1135_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1083_
	);
	LUT4 #(
		.INIT('h0800)
	) name309 (
		\g1135_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1084_
	);
	LUT3 #(
		.INIT('h1b)
	) name310 (
		_w1082_,
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT4 #(
		.INIT('h2e22)
	) name311 (
		\g1099_reg/NET0131 ,
		\g35_pad ,
		_w1081_,
		_w1085_,
		_w1086_
	);
	LUT3 #(
		.INIT('h40)
	) name312 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1087_
	);
	LUT3 #(
		.INIT('h15)
	) name313 (
		\g1111_reg/NET0131 ,
		_w1080_,
		_w1087_,
		_w1088_
	);
	LUT4 #(
		.INIT('h1000)
	) name314 (
		\g1105_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1089_
	);
	LUT4 #(
		.INIT('h2000)
	) name315 (
		\g1105_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1090_
	);
	LUT3 #(
		.INIT('h1b)
	) name316 (
		_w1082_,
		_w1089_,
		_w1090_,
		_w1091_
	);
	LUT4 #(
		.INIT('h2e22)
	) name317 (
		\g1135_reg/NET0131 ,
		\g35_pad ,
		_w1088_,
		_w1091_,
		_w1092_
	);
	LUT3 #(
		.INIT('h80)
	) name318 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1093_
	);
	LUT3 #(
		.INIT('h15)
	) name319 (
		\g1124_reg/NET0131 ,
		_w1080_,
		_w1093_,
		_w1094_
	);
	LUT4 #(
		.INIT('h4000)
	) name320 (
		\g1129_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1095_
	);
	LUT4 #(
		.INIT('h8000)
	) name321 (
		\g1129_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1096_
	);
	LUT3 #(
		.INIT('h1b)
	) name322 (
		_w1082_,
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT4 #(
		.INIT('h2e22)
	) name323 (
		\g1105_reg/NET0131 ,
		\g35_pad ,
		_w1094_,
		_w1097_,
		_w1098_
	);
	LUT3 #(
		.INIT('h10)
	) name324 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1099_
	);
	LUT3 #(
		.INIT('h15)
	) name325 (
		\g1141_reg/NET0131 ,
		_w1080_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('h0010)
	) name326 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		\g956_reg/NET0131 ,
		_w1101_
	);
	LUT4 #(
		.INIT('h1000)
	) name327 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		\g956_reg/NET0131 ,
		_w1102_
	);
	LUT3 #(
		.INIT('h1b)
	) name328 (
		_w1082_,
		_w1101_,
		_w1102_,
		_w1103_
	);
	LUT4 #(
		.INIT('h2e22)
	) name329 (
		\g1129_reg/NET0131 ,
		\g35_pad ,
		_w1100_,
		_w1103_,
		_w1104_
	);
	LUT3 #(
		.INIT('hec)
	) name330 (
		\g35_pad ,
		\g4501_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1105_
	);
	LUT3 #(
		.INIT('h13)
	) name331 (
		\g35_pad ,
		\g4401_reg/NET0131 ,
		\g4411_reg/NET0131 ,
		_w1106_
	);
	LUT3 #(
		.INIT('h04)
	) name332 (
		\g4375_reg/NET0131 ,
		\g4392_reg/NET0131 ,
		\g4405_reg/NET0131 ,
		_w1107_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		\g35_pad ,
		\g4411_reg/NET0131 ,
		_w1108_
	);
	LUT4 #(
		.INIT('h2033)
	) name334 (
		_w1071_,
		_w1106_,
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT4 #(
		.INIT('heccc)
	) name335 (
		\g4388_reg/NET0131 ,
		\g4405_reg/NET0131 ,
		_w1071_,
		_w1073_,
		_w1110_
	);
	LUT3 #(
		.INIT('hc4)
	) name336 (
		\g35_pad ,
		\g4375_reg/NET0131 ,
		\g4382_reg/NET0131 ,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\g35_pad ,
		\g4392_reg/NET0131 ,
		_w1112_
	);
	LUT4 #(
		.INIT('h0020)
	) name338 (
		\g35_pad ,
		\g4375_reg/NET0131 ,
		\g4392_reg/NET0131 ,
		\g4405_reg/NET0131 ,
		_w1113_
	);
	LUT3 #(
		.INIT('hec)
	) name339 (
		_w1071_,
		_w1111_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		\g35_pad ,
		\g4455_reg/NET0131 ,
		_w1115_
	);
	LUT3 #(
		.INIT('h70)
	) name341 (
		_w1071_,
		_w1072_,
		_w1112_,
		_w1116_
	);
	LUT3 #(
		.INIT('hfe)
	) name342 (
		_w1074_,
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT4 #(
		.INIT('h00e0)
	) name343 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w1118_
	);
	LUT4 #(
		.INIT('ha222)
	) name344 (
		\g1384_reg/NET0131 ,
		\g35_pad ,
		_w946_,
		_w1118_,
		_w1119_
	);
	LUT4 #(
		.INIT('hee0e)
	) name345 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		\g1384_reg/NET0131 ,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		\g1389_reg/NET0131 ,
		\g35_pad ,
		_w1121_
	);
	LUT3 #(
		.INIT('h70)
	) name347 (
		_w946_,
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT2 #(
		.INIT('he)
	) name348 (
		_w1119_,
		_w1122_,
		_w1123_
	);
	LUT4 #(
		.INIT('h8000)
	) name349 (
		\g1430_reg/NET0131 ,
		\g1548_reg/NET0131 ,
		\g1554_reg/NET0131 ,
		\g1564_reg/NET0131 ,
		_w1124_
	);
	LUT4 #(
		.INIT('h0100)
	) name350 (
		\g17320_pad ,
		\g17404_pad ,
		\g17423_pad ,
		\g35_pad ,
		_w1125_
	);
	LUT4 #(
		.INIT('h8f00)
	) name351 (
		_w946_,
		_w1055_,
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT3 #(
		.INIT('h10)
	) name352 (
		\g1478_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1127_
	);
	LUT3 #(
		.INIT('h2a)
	) name353 (
		\g35_pad ,
		_w800_,
		_w1127_,
		_w1128_
	);
	LUT4 #(
		.INIT('h0001)
	) name354 (
		\g1548_reg/NET0131 ,
		\g1554_reg/NET0131 ,
		\g1559_reg/NET0131 ,
		\g1564_reg/NET0131 ,
		_w1129_
	);
	LUT4 #(
		.INIT('h0080)
	) name355 (
		\g1322_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\g17320_pad ,
		\g35_pad ,
		_w1131_
	);
	LUT3 #(
		.INIT('h70)
	) name357 (
		_w1129_,
		_w1130_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		\g2153_reg/NET0131 ,
		\g2227_reg/NET0131 ,
		_w1133_
	);
	LUT3 #(
		.INIT('he0)
	) name359 (
		\g2153_reg/NET0131 ,
		\g2227_reg/NET0131 ,
		\g2241_reg/NET0131 ,
		_w1134_
	);
	LUT4 #(
		.INIT('h0100)
	) name360 (
		\g1478_reg/NET0131 ,
		\g1589_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1135_
	);
	LUT3 #(
		.INIT('h93)
	) name361 (
		_w800_,
		_w1134_,
		_w1135_,
		_w1136_
	);
	LUT3 #(
		.INIT('he0)
	) name362 (
		_w1128_,
		_w1132_,
		_w1136_,
		_w1137_
	);
	LUT3 #(
		.INIT('h2a)
	) name363 (
		\g17320_pad ,
		_w1129_,
		_w1130_,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\g2241_reg/NET0131 ,
		\g35_pad ,
		_w1139_
	);
	LUT3 #(
		.INIT('h80)
	) name365 (
		_w800_,
		_w1127_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		\g2227_reg/NET0131 ,
		\g35_pad ,
		_w1141_
	);
	LUT3 #(
		.INIT('h0b)
	) name367 (
		_w1138_,
		_w1140_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('hb)
	) name368 (
		_w1137_,
		_w1142_,
		_w1143_
	);
	LUT3 #(
		.INIT('h10)
	) name369 (
		\g1448_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1144_
	);
	LUT3 #(
		.INIT('h2a)
	) name370 (
		\g35_pad ,
		_w800_,
		_w1144_,
		_w1145_
	);
	LUT4 #(
		.INIT('h0800)
	) name371 (
		\g1322_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		\g17404_pad ,
		\g35_pad ,
		_w1147_
	);
	LUT3 #(
		.INIT('h70)
	) name373 (
		_w1129_,
		_w1146_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		\g2287_reg/NET0131 ,
		\g2361_reg/NET0131 ,
		_w1149_
	);
	LUT3 #(
		.INIT('he0)
	) name375 (
		\g2287_reg/NET0131 ,
		\g2361_reg/NET0131 ,
		\g2375_reg/NET0131 ,
		_w1150_
	);
	LUT4 #(
		.INIT('h0400)
	) name376 (
		\g1448_reg/NET0131 ,
		\g1589_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1151_
	);
	LUT3 #(
		.INIT('h93)
	) name377 (
		_w800_,
		_w1150_,
		_w1151_,
		_w1152_
	);
	LUT3 #(
		.INIT('he0)
	) name378 (
		_w1145_,
		_w1148_,
		_w1152_,
		_w1153_
	);
	LUT3 #(
		.INIT('h2a)
	) name379 (
		\g17404_pad ,
		_w1129_,
		_w1146_,
		_w1154_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		\g2375_reg/NET0131 ,
		\g35_pad ,
		_w1155_
	);
	LUT3 #(
		.INIT('h80)
	) name381 (
		_w800_,
		_w1144_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\g2361_reg/NET0131 ,
		\g35_pad ,
		_w1157_
	);
	LUT3 #(
		.INIT('h0b)
	) name383 (
		_w1154_,
		_w1156_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('hb)
	) name384 (
		_w1153_,
		_w1158_,
		_w1159_
	);
	LUT3 #(
		.INIT('h10)
	) name385 (
		\g1472_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1160_
	);
	LUT3 #(
		.INIT('h2a)
	) name386 (
		\g35_pad ,
		_w800_,
		_w1160_,
		_w1161_
	);
	LUT4 #(
		.INIT('h8000)
	) name387 (
		\g1322_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		\g17423_pad ,
		\g35_pad ,
		_w1163_
	);
	LUT3 #(
		.INIT('h70)
	) name389 (
		_w1129_,
		_w1162_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		\g2421_reg/NET0131 ,
		\g2495_reg/NET0131 ,
		_w1165_
	);
	LUT3 #(
		.INIT('he0)
	) name391 (
		\g2421_reg/NET0131 ,
		\g2495_reg/NET0131 ,
		\g2509_reg/NET0131 ,
		_w1166_
	);
	LUT4 #(
		.INIT('h0100)
	) name392 (
		\g1472_reg/NET0131 ,
		\g1589_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1167_
	);
	LUT3 #(
		.INIT('h93)
	) name393 (
		_w800_,
		_w1166_,
		_w1167_,
		_w1168_
	);
	LUT3 #(
		.INIT('he0)
	) name394 (
		_w1161_,
		_w1164_,
		_w1168_,
		_w1169_
	);
	LUT3 #(
		.INIT('h2a)
	) name395 (
		\g17423_pad ,
		_w1129_,
		_w1162_,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\g2509_reg/NET0131 ,
		\g35_pad ,
		_w1171_
	);
	LUT3 #(
		.INIT('h80)
	) name397 (
		_w800_,
		_w1160_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h2)
	) name398 (
		\g2495_reg/NET0131 ,
		\g35_pad ,
		_w1173_
	);
	LUT3 #(
		.INIT('h0b)
	) name399 (
		_w1170_,
		_w1172_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('hb)
	) name400 (
		_w1169_,
		_w1174_,
		_w1175_
	);
	LUT3 #(
		.INIT('h10)
	) name401 (
		\g1300_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1176_
	);
	LUT3 #(
		.INIT('h2a)
	) name402 (
		\g35_pad ,
		_w800_,
		_w1176_,
		_w1177_
	);
	LUT4 #(
		.INIT('h0008)
	) name403 (
		\g1322_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		\g1430_reg/NET0131 ,
		\g35_pad ,
		_w1179_
	);
	LUT3 #(
		.INIT('h70)
	) name405 (
		_w1129_,
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		\g2555_reg/NET0131 ,
		\g2629_reg/NET0131 ,
		_w1181_
	);
	LUT3 #(
		.INIT('he0)
	) name407 (
		\g2555_reg/NET0131 ,
		\g2629_reg/NET0131 ,
		\g2643_reg/NET0131 ,
		_w1182_
	);
	LUT4 #(
		.INIT('h0400)
	) name408 (
		\g1300_reg/NET0131 ,
		\g1589_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1183_
	);
	LUT3 #(
		.INIT('h93)
	) name409 (
		_w800_,
		_w1182_,
		_w1183_,
		_w1184_
	);
	LUT3 #(
		.INIT('he0)
	) name410 (
		_w1177_,
		_w1180_,
		_w1184_,
		_w1185_
	);
	LUT3 #(
		.INIT('h2a)
	) name411 (
		\g1430_reg/NET0131 ,
		_w1129_,
		_w1178_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		\g2643_reg/NET0131 ,
		\g35_pad ,
		_w1187_
	);
	LUT3 #(
		.INIT('h80)
	) name413 (
		_w800_,
		_w1176_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		\g2629_reg/NET0131 ,
		\g35_pad ,
		_w1189_
	);
	LUT3 #(
		.INIT('h0b)
	) name415 (
		_w1186_,
		_w1188_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('hb)
	) name416 (
		_w1185_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		\g35_pad ,
		\g4417_reg/NET0131 ,
		_w1192_
	);
	LUT3 #(
		.INIT('hfe)
	) name418 (
		_w1074_,
		_w1116_,
		_w1192_,
		_w1193_
	);
	LUT4 #(
		.INIT('ha2f7)
	) name419 (
		\g35_pad ,
		\g4375_reg/NET0131 ,
		\g4382_reg/NET0131 ,
		\g4411_reg/NET0131 ,
		_w1194_
	);
	LUT3 #(
		.INIT('h8f)
	) name420 (
		_w1071_,
		_w1073_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		\g1379_reg/NET0131 ,
		\g35_pad ,
		_w1196_
	);
	LUT4 #(
		.INIT('h00b5)
	) name422 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		\g1384_reg/NET0131 ,
		_w1197_
	);
	LUT4 #(
		.INIT('h002a)
	) name423 (
		\g35_pad ,
		_w946_,
		_w1120_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('he)
	) name424 (
		_w1196_,
		_w1198_,
		_w1199_
	);
	LUT3 #(
		.INIT('hec)
	) name425 (
		\g35_pad ,
		\g4567_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1200_
	);
	LUT3 #(
		.INIT('hec)
	) name426 (
		\g35_pad ,
		\g4498_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1201_
	);
	LUT4 #(
		.INIT('h4c00)
	) name427 (
		\g218_reg/NET0131 ,
		\g35_pad ,
		\g8291_pad ,
		\g8358_pad ,
		_w1202_
	);
	LUT4 #(
		.INIT('h4000)
	) name428 (
		\g191_reg/NET0131 ,
		\g218_reg/NET0131 ,
		\g35_pad ,
		\g8291_pad ,
		_w1203_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		\g222_reg/NET0131 ,
		\g35_pad ,
		_w1204_
	);
	LUT3 #(
		.INIT('hfe)
	) name430 (
		_w1202_,
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT3 #(
		.INIT('h62)
	) name431 (
		\g347_reg/NET0131 ,
		\g35_pad ,
		\g7540_pad ,
		_w1206_
	);
	LUT4 #(
		.INIT('hfad8)
	) name432 (
		\g35_pad ,
		\g4242_reg/NET0131 ,
		\g4297_reg/NET0131 ,
		\g4300_reg/NET0131 ,
		_w1207_
	);
	LUT3 #(
		.INIT('h10)
	) name433 (
		\g1105_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1208_
	);
	LUT3 #(
		.INIT('h2a)
	) name434 (
		\g35_pad ,
		_w802_,
		_w1208_,
		_w1209_
	);
	LUT4 #(
		.INIT('h0200)
	) name435 (
		\g1061_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		\g1221_reg/NET0131 ,
		\g979_reg/NET0131 ,
		_w1210_
	);
	LUT4 #(
		.INIT('h0004)
	) name436 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1216_reg/NET0131 ,
		_w1211_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		\g17316_pad ,
		\g35_pad ,
		_w1212_
	);
	LUT3 #(
		.INIT('h70)
	) name438 (
		_w1210_,
		_w1211_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		\g1728_reg/NET0131 ,
		\g1802_reg/NET0131 ,
		_w1214_
	);
	LUT3 #(
		.INIT('he0)
	) name440 (
		\g1728_reg/NET0131 ,
		\g1802_reg/NET0131 ,
		\g1816_reg/NET0131 ,
		_w1215_
	);
	LUT4 #(
		.INIT('h0400)
	) name441 (
		\g1105_reg/NET0131 ,
		\g1246_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1216_
	);
	LUT3 #(
		.INIT('h93)
	) name442 (
		_w802_,
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT3 #(
		.INIT('he0)
	) name443 (
		_w1209_,
		_w1213_,
		_w1217_,
		_w1218_
	);
	LUT3 #(
		.INIT('h2a)
	) name444 (
		\g17316_pad ,
		_w1210_,
		_w1211_,
		_w1219_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		\g1816_reg/NET0131 ,
		\g35_pad ,
		_w1220_
	);
	LUT3 #(
		.INIT('h80)
	) name446 (
		_w802_,
		_w1208_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		\g1802_reg/NET0131 ,
		\g35_pad ,
		_w1222_
	);
	LUT3 #(
		.INIT('h0b)
	) name448 (
		_w1219_,
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('hb)
	) name449 (
		_w1218_,
		_w1223_,
		_w1224_
	);
	LUT3 #(
		.INIT('h10)
	) name450 (
		\g1129_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1225_
	);
	LUT3 #(
		.INIT('h2a)
	) name451 (
		\g35_pad ,
		_w802_,
		_w1225_,
		_w1226_
	);
	LUT4 #(
		.INIT('h0008)
	) name452 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1216_reg/NET0131 ,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		\g17400_pad ,
		\g35_pad ,
		_w1228_
	);
	LUT3 #(
		.INIT('h70)
	) name454 (
		_w1210_,
		_w1227_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		\g1862_reg/NET0131 ,
		\g1936_reg/NET0131 ,
		_w1230_
	);
	LUT3 #(
		.INIT('he0)
	) name456 (
		\g1862_reg/NET0131 ,
		\g1936_reg/NET0131 ,
		\g1950_reg/NET0131 ,
		_w1231_
	);
	LUT4 #(
		.INIT('h0100)
	) name457 (
		\g1129_reg/NET0131 ,
		\g1246_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1232_
	);
	LUT3 #(
		.INIT('h93)
	) name458 (
		_w802_,
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT3 #(
		.INIT('he0)
	) name459 (
		_w1226_,
		_w1229_,
		_w1233_,
		_w1234_
	);
	LUT3 #(
		.INIT('h2a)
	) name460 (
		\g17400_pad ,
		_w1210_,
		_w1227_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		\g1950_reg/NET0131 ,
		\g35_pad ,
		_w1236_
	);
	LUT3 #(
		.INIT('h80)
	) name462 (
		_w802_,
		_w1225_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\g1936_reg/NET0131 ,
		\g35_pad ,
		_w1238_
	);
	LUT3 #(
		.INIT('h0b)
	) name464 (
		_w1235_,
		_w1237_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('hb)
	) name465 (
		_w1234_,
		_w1239_,
		_w1240_
	);
	LUT3 #(
		.INIT('h04)
	) name466 (
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		\g956_reg/NET0131 ,
		_w1241_
	);
	LUT3 #(
		.INIT('h2a)
	) name467 (
		\g35_pad ,
		_w802_,
		_w1241_,
		_w1242_
	);
	LUT4 #(
		.INIT('h0001)
	) name468 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1216_reg/NET0131 ,
		_w1243_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		\g1087_reg/NET0131 ,
		\g35_pad ,
		_w1244_
	);
	LUT3 #(
		.INIT('h70)
	) name470 (
		_w1210_,
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		\g1996_reg/NET0131 ,
		\g2070_reg/NET0131 ,
		_w1246_
	);
	LUT3 #(
		.INIT('he0)
	) name472 (
		\g1996_reg/NET0131 ,
		\g2070_reg/NET0131 ,
		\g2084_reg/NET0131 ,
		_w1247_
	);
	LUT4 #(
		.INIT('h0020)
	) name473 (
		\g1246_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		\g956_reg/NET0131 ,
		_w1248_
	);
	LUT3 #(
		.INIT('h93)
	) name474 (
		_w802_,
		_w1247_,
		_w1248_,
		_w1249_
	);
	LUT3 #(
		.INIT('he0)
	) name475 (
		_w1242_,
		_w1245_,
		_w1249_,
		_w1250_
	);
	LUT3 #(
		.INIT('h2a)
	) name476 (
		\g1087_reg/NET0131 ,
		_w1210_,
		_w1243_,
		_w1251_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\g2084_reg/NET0131 ,
		\g35_pad ,
		_w1252_
	);
	LUT3 #(
		.INIT('h80)
	) name478 (
		_w802_,
		_w1241_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		\g2070_reg/NET0131 ,
		\g35_pad ,
		_w1254_
	);
	LUT3 #(
		.INIT('h0b)
	) name480 (
		_w1251_,
		_w1253_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('hb)
	) name481 (
		_w1250_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		\g2970_reg/NET0131 ,
		\g35_pad ,
		_w1257_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		\g301_reg/NET0131 ,
		\g35_pad ,
		_w1258_
	);
	LUT3 #(
		.INIT('h10)
	) name484 (
		\g209_reg/NET0131 ,
		\g2902_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1259_
	);
	LUT3 #(
		.INIT('h15)
	) name485 (
		_w1257_,
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h8000)
	) name486 (
		\g1339_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g7946_pad ,
		_w1261_
	);
	LUT3 #(
		.INIT('h80)
	) name487 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g7946_pad ,
		_w1262_
	);
	LUT4 #(
		.INIT('h3f37)
	) name488 (
		\g1306_reg/NET0131 ,
		\g35_pad ,
		_w1261_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name489 (
		\g1521_reg/NET0131 ,
		\g35_pad ,
		_w1264_
	);
	LUT2 #(
		.INIT('hd)
	) name490 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT3 #(
		.INIT('h15)
	) name491 (
		\g2197_reg/NET0131 ,
		_w800_,
		_w1127_,
		_w1266_
	);
	LUT2 #(
		.INIT('h2)
	) name492 (
		\g17320_pad ,
		\g2197_reg/NET0131 ,
		_w1267_
	);
	LUT3 #(
		.INIT('h70)
	) name493 (
		_w1129_,
		_w1130_,
		_w1267_,
		_w1268_
	);
	LUT4 #(
		.INIT('h0100)
	) name494 (
		\g1478_reg/NET0131 ,
		\g1585_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1269_
	);
	LUT3 #(
		.INIT('h2a)
	) name495 (
		\g2153_reg/NET0131 ,
		_w800_,
		_w1269_,
		_w1270_
	);
	LUT4 #(
		.INIT('ha800)
	) name496 (
		\g35_pad ,
		_w1266_,
		_w1268_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		\g2161_reg/NET0131 ,
		\g35_pad ,
		_w1272_
	);
	LUT4 #(
		.INIT('h5700)
	) name498 (
		\g2153_reg/NET0131 ,
		_w1266_,
		_w1268_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h2)
	) name499 (
		\g2165_reg/NET0131 ,
		\g35_pad ,
		_w1274_
	);
	LUT3 #(
		.INIT('hfe)
	) name500 (
		_w1271_,
		_w1273_,
		_w1274_,
		_w1275_
	);
	LUT3 #(
		.INIT('h70)
	) name501 (
		_w800_,
		_w1127_,
		_w1133_,
		_w1276_
	);
	LUT3 #(
		.INIT('h02)
	) name502 (
		\g17320_pad ,
		\g2153_reg/NET0131 ,
		\g2227_reg/NET0131 ,
		_w1277_
	);
	LUT3 #(
		.INIT('h70)
	) name503 (
		_w1129_,
		_w1130_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		\g2165_reg/NET0131 ,
		\g35_pad ,
		_w1279_
	);
	LUT3 #(
		.INIT('h2a)
	) name505 (
		\g35_pad ,
		_w800_,
		_w1269_,
		_w1280_
	);
	LUT4 #(
		.INIT('h01ef)
	) name506 (
		_w1276_,
		_w1278_,
		_w1279_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h2)
	) name507 (
		\g2246_reg/NET0131 ,
		\g35_pad ,
		_w1282_
	);
	LUT2 #(
		.INIT('hd)
	) name508 (
		_w1281_,
		_w1282_,
		_w1283_
	);
	LUT3 #(
		.INIT('h2a)
	) name509 (
		\g2197_reg/NET0131 ,
		_w800_,
		_w1127_,
		_w1284_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\g17320_pad ,
		\g2197_reg/NET0131 ,
		_w1285_
	);
	LUT3 #(
		.INIT('h70)
	) name511 (
		_w1129_,
		_w1130_,
		_w1285_,
		_w1286_
	);
	LUT3 #(
		.INIT('h15)
	) name512 (
		\g2227_reg/NET0131 ,
		_w800_,
		_w1269_,
		_w1287_
	);
	LUT4 #(
		.INIT('ha800)
	) name513 (
		\g35_pad ,
		_w1284_,
		_w1286_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		\g2169_reg/NET0131 ,
		\g35_pad ,
		_w1289_
	);
	LUT4 #(
		.INIT('hab00)
	) name515 (
		\g2227_reg/NET0131 ,
		_w1284_,
		_w1286_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\g2161_reg/NET0131 ,
		\g35_pad ,
		_w1291_
	);
	LUT3 #(
		.INIT('hfe)
	) name517 (
		_w1288_,
		_w1290_,
		_w1291_,
		_w1292_
	);
	LUT3 #(
		.INIT('h2a)
	) name518 (
		\g2153_reg/NET0131 ,
		_w800_,
		_w1127_,
		_w1293_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		\g17320_pad ,
		\g2153_reg/NET0131 ,
		_w1294_
	);
	LUT3 #(
		.INIT('h70)
	) name520 (
		_w1129_,
		_w1130_,
		_w1294_,
		_w1295_
	);
	LUT3 #(
		.INIT('h2a)
	) name521 (
		\g2227_reg/NET0131 ,
		_w800_,
		_w1269_,
		_w1296_
	);
	LUT4 #(
		.INIT('ha800)
	) name522 (
		\g35_pad ,
		_w1293_,
		_w1295_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		\g2173_reg/NET0131 ,
		\g35_pad ,
		_w1298_
	);
	LUT4 #(
		.INIT('h5700)
	) name524 (
		\g2227_reg/NET0131 ,
		_w1293_,
		_w1295_,
		_w1298_,
		_w1299_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\g2177_reg/NET0131 ,
		\g35_pad ,
		_w1300_
	);
	LUT3 #(
		.INIT('hfe)
	) name526 (
		_w1297_,
		_w1299_,
		_w1300_,
		_w1301_
	);
	LUT3 #(
		.INIT('h15)
	) name527 (
		\g2153_reg/NET0131 ,
		_w800_,
		_w1269_,
		_w1302_
	);
	LUT4 #(
		.INIT('ha800)
	) name528 (
		\g35_pad ,
		_w1284_,
		_w1286_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		\g2177_reg/NET0131 ,
		\g35_pad ,
		_w1304_
	);
	LUT4 #(
		.INIT('hab00)
	) name530 (
		\g2153_reg/NET0131 ,
		_w1284_,
		_w1286_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h2)
	) name531 (
		\g2181_reg/NET0131 ,
		\g35_pad ,
		_w1306_
	);
	LUT3 #(
		.INIT('hfe)
	) name532 (
		_w1303_,
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('ha800)
	) name533 (
		\g35_pad ,
		_w1266_,
		_w1268_,
		_w1296_,
		_w1308_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		\g2181_reg/NET0131 ,
		\g35_pad ,
		_w1309_
	);
	LUT4 #(
		.INIT('h5700)
	) name535 (
		\g2227_reg/NET0131 ,
		_w1266_,
		_w1268_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		\g2169_reg/NET0131 ,
		\g35_pad ,
		_w1311_
	);
	LUT3 #(
		.INIT('hfe)
	) name537 (
		_w1308_,
		_w1310_,
		_w1311_,
		_w1312_
	);
	LUT3 #(
		.INIT('h15)
	) name538 (
		\g2331_reg/NET0131 ,
		_w800_,
		_w1144_,
		_w1313_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		\g17404_pad ,
		\g2331_reg/NET0131 ,
		_w1314_
	);
	LUT3 #(
		.INIT('h70)
	) name540 (
		_w1129_,
		_w1146_,
		_w1314_,
		_w1315_
	);
	LUT4 #(
		.INIT('h0400)
	) name541 (
		\g1448_reg/NET0131 ,
		\g1585_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1316_
	);
	LUT3 #(
		.INIT('h2a)
	) name542 (
		\g2287_reg/NET0131 ,
		_w800_,
		_w1316_,
		_w1317_
	);
	LUT4 #(
		.INIT('ha800)
	) name543 (
		\g35_pad ,
		_w1313_,
		_w1315_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		\g2295_reg/NET0131 ,
		\g35_pad ,
		_w1319_
	);
	LUT4 #(
		.INIT('h5700)
	) name545 (
		\g2287_reg/NET0131 ,
		_w1313_,
		_w1315_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h2)
	) name546 (
		\g2299_reg/NET0131 ,
		\g35_pad ,
		_w1321_
	);
	LUT3 #(
		.INIT('hfe)
	) name547 (
		_w1318_,
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT3 #(
		.INIT('h70)
	) name548 (
		_w800_,
		_w1144_,
		_w1149_,
		_w1323_
	);
	LUT3 #(
		.INIT('h02)
	) name549 (
		\g17404_pad ,
		\g2287_reg/NET0131 ,
		\g2361_reg/NET0131 ,
		_w1324_
	);
	LUT3 #(
		.INIT('h70)
	) name550 (
		_w1129_,
		_w1146_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		\g2299_reg/NET0131 ,
		\g35_pad ,
		_w1326_
	);
	LUT3 #(
		.INIT('h2a)
	) name552 (
		\g35_pad ,
		_w800_,
		_w1316_,
		_w1327_
	);
	LUT4 #(
		.INIT('h01ef)
	) name553 (
		_w1323_,
		_w1325_,
		_w1326_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		\g2380_reg/NET0131 ,
		\g35_pad ,
		_w1329_
	);
	LUT2 #(
		.INIT('hd)
	) name555 (
		_w1328_,
		_w1329_,
		_w1330_
	);
	LUT3 #(
		.INIT('h2a)
	) name556 (
		\g2331_reg/NET0131 ,
		_w800_,
		_w1144_,
		_w1331_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\g17404_pad ,
		\g2331_reg/NET0131 ,
		_w1332_
	);
	LUT3 #(
		.INIT('h70)
	) name558 (
		_w1129_,
		_w1146_,
		_w1332_,
		_w1333_
	);
	LUT3 #(
		.INIT('h15)
	) name559 (
		\g2361_reg/NET0131 ,
		_w800_,
		_w1316_,
		_w1334_
	);
	LUT4 #(
		.INIT('ha800)
	) name560 (
		\g35_pad ,
		_w1331_,
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		\g2303_reg/NET0131 ,
		\g35_pad ,
		_w1336_
	);
	LUT4 #(
		.INIT('hab00)
	) name562 (
		\g2361_reg/NET0131 ,
		_w1331_,
		_w1333_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		\g2295_reg/NET0131 ,
		\g35_pad ,
		_w1338_
	);
	LUT3 #(
		.INIT('hfe)
	) name564 (
		_w1335_,
		_w1337_,
		_w1338_,
		_w1339_
	);
	LUT3 #(
		.INIT('h2a)
	) name565 (
		\g2287_reg/NET0131 ,
		_w800_,
		_w1144_,
		_w1340_
	);
	LUT2 #(
		.INIT('h8)
	) name566 (
		\g17404_pad ,
		\g2287_reg/NET0131 ,
		_w1341_
	);
	LUT3 #(
		.INIT('h70)
	) name567 (
		_w1129_,
		_w1146_,
		_w1341_,
		_w1342_
	);
	LUT3 #(
		.INIT('h2a)
	) name568 (
		\g2361_reg/NET0131 ,
		_w800_,
		_w1316_,
		_w1343_
	);
	LUT4 #(
		.INIT('ha800)
	) name569 (
		\g35_pad ,
		_w1340_,
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		\g2307_reg/NET0131 ,
		\g35_pad ,
		_w1345_
	);
	LUT4 #(
		.INIT('h5700)
	) name571 (
		\g2361_reg/NET0131 ,
		_w1340_,
		_w1342_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		\g2311_reg/NET0131 ,
		\g35_pad ,
		_w1347_
	);
	LUT3 #(
		.INIT('hfe)
	) name573 (
		_w1344_,
		_w1346_,
		_w1347_,
		_w1348_
	);
	LUT3 #(
		.INIT('h15)
	) name574 (
		\g2287_reg/NET0131 ,
		_w800_,
		_w1316_,
		_w1349_
	);
	LUT4 #(
		.INIT('ha800)
	) name575 (
		\g35_pad ,
		_w1331_,
		_w1333_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h8)
	) name576 (
		\g2311_reg/NET0131 ,
		\g35_pad ,
		_w1351_
	);
	LUT4 #(
		.INIT('hab00)
	) name577 (
		\g2287_reg/NET0131 ,
		_w1331_,
		_w1333_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		\g2315_reg/NET0131 ,
		\g35_pad ,
		_w1353_
	);
	LUT3 #(
		.INIT('hfe)
	) name579 (
		_w1350_,
		_w1352_,
		_w1353_,
		_w1354_
	);
	LUT4 #(
		.INIT('ha800)
	) name580 (
		\g35_pad ,
		_w1313_,
		_w1315_,
		_w1343_,
		_w1355_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		\g2315_reg/NET0131 ,
		\g35_pad ,
		_w1356_
	);
	LUT4 #(
		.INIT('h5700)
	) name582 (
		\g2361_reg/NET0131 ,
		_w1313_,
		_w1315_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		\g2303_reg/NET0131 ,
		\g35_pad ,
		_w1358_
	);
	LUT3 #(
		.INIT('hfe)
	) name584 (
		_w1355_,
		_w1357_,
		_w1358_,
		_w1359_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name585 (
		\g1339_reg/NET0131 ,
		\g1521_reg/NET0131 ,
		\g35_pad ,
		\g7946_pad ,
		_w1360_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\g1526_reg/NET0131 ,
		\g35_pad ,
		_w1361_
	);
	LUT2 #(
		.INIT('he)
	) name587 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT3 #(
		.INIT('h15)
	) name588 (
		\g2465_reg/NET0131 ,
		_w800_,
		_w1160_,
		_w1363_
	);
	LUT2 #(
		.INIT('h2)
	) name589 (
		\g17423_pad ,
		\g2465_reg/NET0131 ,
		_w1364_
	);
	LUT3 #(
		.INIT('h70)
	) name590 (
		_w1129_,
		_w1162_,
		_w1364_,
		_w1365_
	);
	LUT4 #(
		.INIT('h0100)
	) name591 (
		\g1472_reg/NET0131 ,
		\g1585_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1366_
	);
	LUT3 #(
		.INIT('h2a)
	) name592 (
		\g2421_reg/NET0131 ,
		_w800_,
		_w1366_,
		_w1367_
	);
	LUT4 #(
		.INIT('ha800)
	) name593 (
		\g35_pad ,
		_w1363_,
		_w1365_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\g2429_reg/NET0131 ,
		\g35_pad ,
		_w1369_
	);
	LUT4 #(
		.INIT('h5700)
	) name595 (
		\g2421_reg/NET0131 ,
		_w1363_,
		_w1365_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		\g2433_reg/NET0131 ,
		\g35_pad ,
		_w1371_
	);
	LUT3 #(
		.INIT('hfe)
	) name597 (
		_w1368_,
		_w1370_,
		_w1371_,
		_w1372_
	);
	LUT3 #(
		.INIT('h70)
	) name598 (
		_w800_,
		_w1160_,
		_w1165_,
		_w1373_
	);
	LUT3 #(
		.INIT('h02)
	) name599 (
		\g17423_pad ,
		\g2421_reg/NET0131 ,
		\g2495_reg/NET0131 ,
		_w1374_
	);
	LUT3 #(
		.INIT('h70)
	) name600 (
		_w1129_,
		_w1162_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		\g2433_reg/NET0131 ,
		\g35_pad ,
		_w1376_
	);
	LUT3 #(
		.INIT('h2a)
	) name602 (
		\g35_pad ,
		_w800_,
		_w1366_,
		_w1377_
	);
	LUT4 #(
		.INIT('h01ef)
	) name603 (
		_w1373_,
		_w1375_,
		_w1376_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		\g2514_reg/NET0131 ,
		\g35_pad ,
		_w1379_
	);
	LUT2 #(
		.INIT('hd)
	) name605 (
		_w1378_,
		_w1379_,
		_w1380_
	);
	LUT3 #(
		.INIT('h2a)
	) name606 (
		\g2465_reg/NET0131 ,
		_w800_,
		_w1160_,
		_w1381_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		\g17423_pad ,
		\g2465_reg/NET0131 ,
		_w1382_
	);
	LUT3 #(
		.INIT('h70)
	) name608 (
		_w1129_,
		_w1162_,
		_w1382_,
		_w1383_
	);
	LUT3 #(
		.INIT('h15)
	) name609 (
		\g2495_reg/NET0131 ,
		_w800_,
		_w1366_,
		_w1384_
	);
	LUT4 #(
		.INIT('ha800)
	) name610 (
		\g35_pad ,
		_w1381_,
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		\g2437_reg/NET0131 ,
		\g35_pad ,
		_w1386_
	);
	LUT4 #(
		.INIT('hab00)
	) name612 (
		\g2495_reg/NET0131 ,
		_w1381_,
		_w1383_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		\g2429_reg/NET0131 ,
		\g35_pad ,
		_w1388_
	);
	LUT3 #(
		.INIT('hfe)
	) name614 (
		_w1385_,
		_w1387_,
		_w1388_,
		_w1389_
	);
	LUT3 #(
		.INIT('h2a)
	) name615 (
		\g2421_reg/NET0131 ,
		_w800_,
		_w1160_,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name616 (
		\g17423_pad ,
		\g2421_reg/NET0131 ,
		_w1391_
	);
	LUT3 #(
		.INIT('h70)
	) name617 (
		_w1129_,
		_w1162_,
		_w1391_,
		_w1392_
	);
	LUT3 #(
		.INIT('h2a)
	) name618 (
		\g2495_reg/NET0131 ,
		_w800_,
		_w1366_,
		_w1393_
	);
	LUT4 #(
		.INIT('ha800)
	) name619 (
		\g35_pad ,
		_w1390_,
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		\g2441_reg/NET0131 ,
		\g35_pad ,
		_w1395_
	);
	LUT4 #(
		.INIT('h5700)
	) name621 (
		\g2495_reg/NET0131 ,
		_w1390_,
		_w1392_,
		_w1395_,
		_w1396_
	);
	LUT2 #(
		.INIT('h2)
	) name622 (
		\g2445_reg/NET0131 ,
		\g35_pad ,
		_w1397_
	);
	LUT3 #(
		.INIT('hfe)
	) name623 (
		_w1394_,
		_w1396_,
		_w1397_,
		_w1398_
	);
	LUT3 #(
		.INIT('h15)
	) name624 (
		\g2421_reg/NET0131 ,
		_w800_,
		_w1366_,
		_w1399_
	);
	LUT4 #(
		.INIT('ha800)
	) name625 (
		\g35_pad ,
		_w1381_,
		_w1383_,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\g2445_reg/NET0131 ,
		\g35_pad ,
		_w1401_
	);
	LUT4 #(
		.INIT('hab00)
	) name627 (
		\g2421_reg/NET0131 ,
		_w1381_,
		_w1383_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		\g2449_reg/NET0131 ,
		\g35_pad ,
		_w1403_
	);
	LUT3 #(
		.INIT('hfe)
	) name629 (
		_w1400_,
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('ha800)
	) name630 (
		\g35_pad ,
		_w1363_,
		_w1365_,
		_w1393_,
		_w1405_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		\g2449_reg/NET0131 ,
		\g35_pad ,
		_w1406_
	);
	LUT4 #(
		.INIT('h5700)
	) name632 (
		\g2495_reg/NET0131 ,
		_w1363_,
		_w1365_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h2)
	) name633 (
		\g2437_reg/NET0131 ,
		\g35_pad ,
		_w1408_
	);
	LUT3 #(
		.INIT('hfe)
	) name634 (
		_w1405_,
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT3 #(
		.INIT('h15)
	) name635 (
		\g2599_reg/NET0131 ,
		_w800_,
		_w1176_,
		_w1410_
	);
	LUT2 #(
		.INIT('h2)
	) name636 (
		\g1430_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		_w1411_
	);
	LUT3 #(
		.INIT('h70)
	) name637 (
		_w1129_,
		_w1178_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('h0400)
	) name638 (
		\g1300_reg/NET0131 ,
		\g1585_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1413_
	);
	LUT3 #(
		.INIT('h2a)
	) name639 (
		\g2555_reg/NET0131 ,
		_w800_,
		_w1413_,
		_w1414_
	);
	LUT4 #(
		.INIT('ha800)
	) name640 (
		\g35_pad ,
		_w1410_,
		_w1412_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\g2563_reg/NET0131 ,
		\g35_pad ,
		_w1416_
	);
	LUT4 #(
		.INIT('h5700)
	) name642 (
		\g2555_reg/NET0131 ,
		_w1410_,
		_w1412_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h2)
	) name643 (
		\g2567_reg/NET0131 ,
		\g35_pad ,
		_w1418_
	);
	LUT3 #(
		.INIT('hfe)
	) name644 (
		_w1415_,
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('h70)
	) name645 (
		_w800_,
		_w1176_,
		_w1181_,
		_w1420_
	);
	LUT3 #(
		.INIT('h02)
	) name646 (
		\g1430_reg/NET0131 ,
		\g2555_reg/NET0131 ,
		\g2629_reg/NET0131 ,
		_w1421_
	);
	LUT3 #(
		.INIT('h70)
	) name647 (
		_w1129_,
		_w1178_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		\g2567_reg/NET0131 ,
		\g35_pad ,
		_w1423_
	);
	LUT3 #(
		.INIT('h2a)
	) name649 (
		\g35_pad ,
		_w800_,
		_w1413_,
		_w1424_
	);
	LUT4 #(
		.INIT('h01ef)
	) name650 (
		_w1420_,
		_w1422_,
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		\g2648_reg/NET0131 ,
		\g35_pad ,
		_w1426_
	);
	LUT2 #(
		.INIT('hd)
	) name652 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT3 #(
		.INIT('h2a)
	) name653 (
		\g2599_reg/NET0131 ,
		_w800_,
		_w1176_,
		_w1428_
	);
	LUT2 #(
		.INIT('h8)
	) name654 (
		\g1430_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		_w1429_
	);
	LUT3 #(
		.INIT('h70)
	) name655 (
		_w1129_,
		_w1178_,
		_w1429_,
		_w1430_
	);
	LUT3 #(
		.INIT('h15)
	) name656 (
		\g2629_reg/NET0131 ,
		_w800_,
		_w1413_,
		_w1431_
	);
	LUT4 #(
		.INIT('ha800)
	) name657 (
		\g35_pad ,
		_w1428_,
		_w1430_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		\g2571_reg/NET0131 ,
		\g35_pad ,
		_w1433_
	);
	LUT4 #(
		.INIT('hab00)
	) name659 (
		\g2629_reg/NET0131 ,
		_w1428_,
		_w1430_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h2)
	) name660 (
		\g2563_reg/NET0131 ,
		\g35_pad ,
		_w1435_
	);
	LUT3 #(
		.INIT('hfe)
	) name661 (
		_w1432_,
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT3 #(
		.INIT('h2a)
	) name662 (
		\g2629_reg/NET0131 ,
		_w800_,
		_w1176_,
		_w1437_
	);
	LUT2 #(
		.INIT('h8)
	) name663 (
		\g1430_reg/NET0131 ,
		\g2629_reg/NET0131 ,
		_w1438_
	);
	LUT3 #(
		.INIT('h70)
	) name664 (
		_w1129_,
		_w1178_,
		_w1438_,
		_w1439_
	);
	LUT4 #(
		.INIT('h8880)
	) name665 (
		\g35_pad ,
		_w1414_,
		_w1437_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		\g2575_reg/NET0131 ,
		\g35_pad ,
		_w1441_
	);
	LUT4 #(
		.INIT('h5700)
	) name667 (
		\g2555_reg/NET0131 ,
		_w1437_,
		_w1439_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		\g2579_reg/NET0131 ,
		\g35_pad ,
		_w1443_
	);
	LUT3 #(
		.INIT('hfe)
	) name669 (
		_w1440_,
		_w1442_,
		_w1443_,
		_w1444_
	);
	LUT3 #(
		.INIT('h15)
	) name670 (
		\g2555_reg/NET0131 ,
		_w800_,
		_w1413_,
		_w1445_
	);
	LUT4 #(
		.INIT('ha800)
	) name671 (
		\g35_pad ,
		_w1428_,
		_w1430_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h8)
	) name672 (
		\g2579_reg/NET0131 ,
		\g35_pad ,
		_w1447_
	);
	LUT4 #(
		.INIT('hab00)
	) name673 (
		\g2555_reg/NET0131 ,
		_w1428_,
		_w1430_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		\g2583_reg/NET0131 ,
		\g35_pad ,
		_w1449_
	);
	LUT3 #(
		.INIT('hfe)
	) name675 (
		_w1446_,
		_w1448_,
		_w1449_,
		_w1450_
	);
	LUT3 #(
		.INIT('h2a)
	) name676 (
		\g2629_reg/NET0131 ,
		_w800_,
		_w1413_,
		_w1451_
	);
	LUT4 #(
		.INIT('ha800)
	) name677 (
		\g35_pad ,
		_w1410_,
		_w1412_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		\g2583_reg/NET0131 ,
		\g35_pad ,
		_w1453_
	);
	LUT4 #(
		.INIT('h5700)
	) name679 (
		\g2629_reg/NET0131 ,
		_w1410_,
		_w1412_,
		_w1453_,
		_w1454_
	);
	LUT2 #(
		.INIT('h2)
	) name680 (
		\g2571_reg/NET0131 ,
		\g35_pad ,
		_w1455_
	);
	LUT3 #(
		.INIT('hfe)
	) name681 (
		_w1452_,
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT3 #(
		.INIT('hec)
	) name682 (
		\g35_pad ,
		\g4543_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1457_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		\g1395_reg/NET0131 ,
		\g35_pad ,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		\g12923_pad ,
		\g1395_reg/NET0131 ,
		_w1459_
	);
	LUT3 #(
		.INIT('h45)
	) name685 (
		\g1404_reg/NET0131 ,
		_w1058_,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		\g1322_reg/NET0131 ,
		\g35_pad ,
		_w1461_
	);
	LUT3 #(
		.INIT('h80)
	) name687 (
		\g12923_pad ,
		\g1395_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		_w1462_
	);
	LUT3 #(
		.INIT('h8c)
	) name688 (
		_w1058_,
		_w1461_,
		_w1462_,
		_w1463_
	);
	LUT3 #(
		.INIT('hba)
	) name689 (
		_w1458_,
		_w1460_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('hca00)
	) name690 (
		\g10527_pad ,
		\g12923_pad ,
		\g17423_pad ,
		\g35_pad ,
		_w1465_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		\g1589_reg/NET0131 ,
		\g35_pad ,
		_w1466_
	);
	LUT2 #(
		.INIT('he)
	) name692 (
		_w1465_,
		_w1466_,
		_w1467_
	);
	LUT4 #(
		.INIT('hfbc8)
	) name693 (
		\g301_reg/NET0131 ,
		\g35_pad ,
		\g534_reg/NET0131 ,
		\g542_reg/NET0131 ,
		_w1468_
	);
	LUT3 #(
		.INIT('hec)
	) name694 (
		\g35_pad ,
		\g4495_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		\g1404_reg/NET0131 ,
		\g35_pad ,
		_w1470_
	);
	LUT4 #(
		.INIT('h0200)
	) name696 (
		\g12923_pad ,
		\g1395_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		\g19357_pad ,
		_w1471_
	);
	LUT4 #(
		.INIT('h4000)
	) name697 (
		\g12923_pad ,
		\g1404_reg/NET0131 ,
		\g19357_pad ,
		\g35_pad ,
		_w1472_
	);
	LUT3 #(
		.INIT('h01)
	) name698 (
		_w1470_,
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT3 #(
		.INIT('h70)
	) name699 (
		_w896_,
		_w900_,
		_w901_,
		_w1474_
	);
	LUT3 #(
		.INIT('h40)
	) name700 (
		\g807_reg/NET0131 ,
		_w897_,
		_w898_,
		_w1475_
	);
	LUT4 #(
		.INIT('hc444)
	) name701 (
		\g35_pad ,
		\g794_reg/NET0131 ,
		_w896_,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('he)
	) name702 (
		_w1474_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h8)
	) name703 (
		\g35_pad ,
		\g4423_reg/NET0131 ,
		_w1478_
	);
	LUT3 #(
		.INIT('hd8)
	) name704 (
		\g35_pad ,
		\g4423_reg/NET0131 ,
		\g4427_reg/NET0131 ,
		_w1479_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		\g12923_pad ,
		\g1395_reg/NET0131 ,
		_w1480_
	);
	LUT4 #(
		.INIT('h0001)
	) name706 (
		\g1333_reg/NET0131 ,
		\g1395_reg/NET0131 ,
		\g19357_pad ,
		\g7946_pad ,
		_w1481_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w1480_,
		_w1481_,
		_w1482_
	);
	LUT3 #(
		.INIT('hb0)
	) name708 (
		_w1058_,
		_w1459_,
		_w1461_,
		_w1483_
	);
	LUT2 #(
		.INIT('h8)
	) name709 (
		_w1482_,
		_w1483_,
		_w1484_
	);
	LUT3 #(
		.INIT('h01)
	) name710 (
		\g8918_pad ,
		\g8919_pad ,
		\g8920_pad ,
		_w1485_
	);
	LUT4 #(
		.INIT('h0001)
	) name711 (
		\g11770_pad ,
		\g8915_pad ,
		\g8916_pad ,
		\g8917_pad ,
		_w1486_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w1485_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('hca)
	) name713 (
		\g4145_reg/NET0131 ,
		\g4164_reg/NET0131 ,
		\g4253_reg/NET0131 ,
		_w1488_
	);
	LUT4 #(
		.INIT('h8976)
	) name714 (
		\g4235_reg/NET0131 ,
		\g8870_pad ,
		_w1487_,
		_w1488_,
		_w1489_
	);
	LUT3 #(
		.INIT('h4e)
	) name715 (
		\g35_pad ,
		\g4235_reg/NET0131 ,
		_w1489_,
		_w1490_
	);
	LUT3 #(
		.INIT('h3a)
	) name716 (
		\g333_reg/NET0131 ,
		\g347_reg/NET0131 ,
		\g35_pad ,
		_w1491_
	);
	LUT3 #(
		.INIT('h15)
	) name717 (
		\g1772_reg/NET0131 ,
		_w802_,
		_w1208_,
		_w1492_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		\g17316_pad ,
		\g1772_reg/NET0131 ,
		_w1493_
	);
	LUT3 #(
		.INIT('h70)
	) name719 (
		_w1210_,
		_w1211_,
		_w1493_,
		_w1494_
	);
	LUT4 #(
		.INIT('h0400)
	) name720 (
		\g1105_reg/NET0131 ,
		\g1242_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1495_
	);
	LUT3 #(
		.INIT('h2a)
	) name721 (
		\g1728_reg/NET0131 ,
		_w802_,
		_w1495_,
		_w1496_
	);
	LUT4 #(
		.INIT('ha800)
	) name722 (
		\g35_pad ,
		_w1492_,
		_w1494_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h8)
	) name723 (
		\g1736_reg/NET0131 ,
		\g35_pad ,
		_w1498_
	);
	LUT4 #(
		.INIT('h5700)
	) name724 (
		\g1728_reg/NET0131 ,
		_w1492_,
		_w1494_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h2)
	) name725 (
		\g1740_reg/NET0131 ,
		\g35_pad ,
		_w1500_
	);
	LUT3 #(
		.INIT('hfe)
	) name726 (
		_w1497_,
		_w1499_,
		_w1500_,
		_w1501_
	);
	LUT3 #(
		.INIT('h70)
	) name727 (
		_w802_,
		_w1208_,
		_w1214_,
		_w1502_
	);
	LUT3 #(
		.INIT('h04)
	) name728 (
		\g1728_reg/NET0131 ,
		\g17316_pad ,
		\g1802_reg/NET0131 ,
		_w1503_
	);
	LUT3 #(
		.INIT('h70)
	) name729 (
		_w1210_,
		_w1211_,
		_w1503_,
		_w1504_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		\g1740_reg/NET0131 ,
		\g35_pad ,
		_w1505_
	);
	LUT3 #(
		.INIT('h2a)
	) name731 (
		\g35_pad ,
		_w802_,
		_w1495_,
		_w1506_
	);
	LUT4 #(
		.INIT('h01ef)
	) name732 (
		_w1502_,
		_w1504_,
		_w1505_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		\g1821_reg/NET0131 ,
		\g35_pad ,
		_w1508_
	);
	LUT2 #(
		.INIT('hd)
	) name734 (
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT3 #(
		.INIT('h2a)
	) name735 (
		\g1728_reg/NET0131 ,
		_w802_,
		_w1208_,
		_w1510_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		\g1728_reg/NET0131 ,
		\g17316_pad ,
		_w1511_
	);
	LUT3 #(
		.INIT('h70)
	) name737 (
		_w1210_,
		_w1211_,
		_w1511_,
		_w1512_
	);
	LUT3 #(
		.INIT('h2a)
	) name738 (
		\g1802_reg/NET0131 ,
		_w802_,
		_w1495_,
		_w1513_
	);
	LUT4 #(
		.INIT('ha800)
	) name739 (
		\g35_pad ,
		_w1510_,
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		\g1748_reg/NET0131 ,
		\g35_pad ,
		_w1515_
	);
	LUT4 #(
		.INIT('h5700)
	) name741 (
		\g1802_reg/NET0131 ,
		_w1510_,
		_w1512_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h2)
	) name742 (
		\g1752_reg/NET0131 ,
		\g35_pad ,
		_w1517_
	);
	LUT3 #(
		.INIT('hfe)
	) name743 (
		_w1514_,
		_w1516_,
		_w1517_,
		_w1518_
	);
	LUT3 #(
		.INIT('h2a)
	) name744 (
		\g1772_reg/NET0131 ,
		_w802_,
		_w1208_,
		_w1519_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		\g17316_pad ,
		\g1772_reg/NET0131 ,
		_w1520_
	);
	LUT3 #(
		.INIT('h70)
	) name746 (
		_w1210_,
		_w1211_,
		_w1520_,
		_w1521_
	);
	LUT3 #(
		.INIT('h15)
	) name747 (
		\g1802_reg/NET0131 ,
		_w802_,
		_w1495_,
		_w1522_
	);
	LUT4 #(
		.INIT('ha800)
	) name748 (
		\g35_pad ,
		_w1519_,
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		\g1744_reg/NET0131 ,
		\g35_pad ,
		_w1524_
	);
	LUT4 #(
		.INIT('hab00)
	) name750 (
		\g1802_reg/NET0131 ,
		_w1519_,
		_w1521_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		\g1736_reg/NET0131 ,
		\g35_pad ,
		_w1526_
	);
	LUT3 #(
		.INIT('hfe)
	) name752 (
		_w1523_,
		_w1525_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('h15)
	) name753 (
		\g1728_reg/NET0131 ,
		_w802_,
		_w1495_,
		_w1528_
	);
	LUT4 #(
		.INIT('ha800)
	) name754 (
		\g35_pad ,
		_w1519_,
		_w1521_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h8)
	) name755 (
		\g1752_reg/NET0131 ,
		\g35_pad ,
		_w1530_
	);
	LUT4 #(
		.INIT('hab00)
	) name756 (
		\g1728_reg/NET0131 ,
		_w1519_,
		_w1521_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h2)
	) name757 (
		\g1756_reg/NET0131 ,
		\g35_pad ,
		_w1532_
	);
	LUT3 #(
		.INIT('hfe)
	) name758 (
		_w1529_,
		_w1531_,
		_w1532_,
		_w1533_
	);
	LUT4 #(
		.INIT('ha800)
	) name759 (
		\g35_pad ,
		_w1492_,
		_w1494_,
		_w1513_,
		_w1534_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		\g1756_reg/NET0131 ,
		\g35_pad ,
		_w1535_
	);
	LUT4 #(
		.INIT('h5700)
	) name761 (
		\g1802_reg/NET0131 ,
		_w1492_,
		_w1494_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		\g1744_reg/NET0131 ,
		\g35_pad ,
		_w1537_
	);
	LUT3 #(
		.INIT('hfe)
	) name763 (
		_w1534_,
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('h15)
	) name764 (
		\g1906_reg/NET0131 ,
		_w802_,
		_w1225_,
		_w1539_
	);
	LUT2 #(
		.INIT('h2)
	) name765 (
		\g17400_pad ,
		\g1906_reg/NET0131 ,
		_w1540_
	);
	LUT3 #(
		.INIT('h70)
	) name766 (
		_w1210_,
		_w1227_,
		_w1540_,
		_w1541_
	);
	LUT4 #(
		.INIT('h0100)
	) name767 (
		\g1129_reg/NET0131 ,
		\g1242_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1542_
	);
	LUT3 #(
		.INIT('h2a)
	) name768 (
		\g1862_reg/NET0131 ,
		_w802_,
		_w1542_,
		_w1543_
	);
	LUT4 #(
		.INIT('ha800)
	) name769 (
		\g35_pad ,
		_w1539_,
		_w1541_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		\g1870_reg/NET0131 ,
		\g35_pad ,
		_w1545_
	);
	LUT4 #(
		.INIT('h5700)
	) name771 (
		\g1862_reg/NET0131 ,
		_w1539_,
		_w1541_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h2)
	) name772 (
		\g1874_reg/NET0131 ,
		\g35_pad ,
		_w1547_
	);
	LUT3 #(
		.INIT('hfe)
	) name773 (
		_w1544_,
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT3 #(
		.INIT('h70)
	) name774 (
		_w802_,
		_w1225_,
		_w1230_,
		_w1549_
	);
	LUT3 #(
		.INIT('h02)
	) name775 (
		\g17400_pad ,
		\g1862_reg/NET0131 ,
		\g1936_reg/NET0131 ,
		_w1550_
	);
	LUT3 #(
		.INIT('h70)
	) name776 (
		_w1210_,
		_w1227_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h8)
	) name777 (
		\g1874_reg/NET0131 ,
		\g35_pad ,
		_w1552_
	);
	LUT3 #(
		.INIT('h2a)
	) name778 (
		\g35_pad ,
		_w802_,
		_w1542_,
		_w1553_
	);
	LUT4 #(
		.INIT('h01ef)
	) name779 (
		_w1549_,
		_w1551_,
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h2)
	) name780 (
		\g1955_reg/NET0131 ,
		\g35_pad ,
		_w1555_
	);
	LUT2 #(
		.INIT('hd)
	) name781 (
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT3 #(
		.INIT('h2a)
	) name782 (
		\g1906_reg/NET0131 ,
		_w802_,
		_w1225_,
		_w1557_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		\g17400_pad ,
		\g1906_reg/NET0131 ,
		_w1558_
	);
	LUT3 #(
		.INIT('h70)
	) name784 (
		_w1210_,
		_w1227_,
		_w1558_,
		_w1559_
	);
	LUT3 #(
		.INIT('h15)
	) name785 (
		\g1936_reg/NET0131 ,
		_w802_,
		_w1542_,
		_w1560_
	);
	LUT4 #(
		.INIT('ha800)
	) name786 (
		\g35_pad ,
		_w1557_,
		_w1559_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		\g1878_reg/NET0131 ,
		\g35_pad ,
		_w1562_
	);
	LUT4 #(
		.INIT('hab00)
	) name788 (
		\g1936_reg/NET0131 ,
		_w1557_,
		_w1559_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h2)
	) name789 (
		\g1870_reg/NET0131 ,
		\g35_pad ,
		_w1564_
	);
	LUT3 #(
		.INIT('hfe)
	) name790 (
		_w1561_,
		_w1563_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('h2a)
	) name791 (
		\g1862_reg/NET0131 ,
		_w802_,
		_w1225_,
		_w1566_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		\g17400_pad ,
		\g1862_reg/NET0131 ,
		_w1567_
	);
	LUT3 #(
		.INIT('h70)
	) name793 (
		_w1210_,
		_w1227_,
		_w1567_,
		_w1568_
	);
	LUT3 #(
		.INIT('h2a)
	) name794 (
		\g1936_reg/NET0131 ,
		_w802_,
		_w1542_,
		_w1569_
	);
	LUT4 #(
		.INIT('ha800)
	) name795 (
		\g35_pad ,
		_w1566_,
		_w1568_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		\g1882_reg/NET0131 ,
		\g35_pad ,
		_w1571_
	);
	LUT4 #(
		.INIT('h5700)
	) name797 (
		\g1936_reg/NET0131 ,
		_w1566_,
		_w1568_,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		\g1886_reg/NET0131 ,
		\g35_pad ,
		_w1573_
	);
	LUT3 #(
		.INIT('hfe)
	) name799 (
		_w1570_,
		_w1572_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h15)
	) name800 (
		\g1862_reg/NET0131 ,
		_w802_,
		_w1542_,
		_w1575_
	);
	LUT4 #(
		.INIT('ha800)
	) name801 (
		\g35_pad ,
		_w1557_,
		_w1559_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\g1886_reg/NET0131 ,
		\g35_pad ,
		_w1577_
	);
	LUT4 #(
		.INIT('hab00)
	) name803 (
		\g1862_reg/NET0131 ,
		_w1557_,
		_w1559_,
		_w1577_,
		_w1578_
	);
	LUT2 #(
		.INIT('h2)
	) name804 (
		\g1890_reg/NET0131 ,
		\g35_pad ,
		_w1579_
	);
	LUT3 #(
		.INIT('hfe)
	) name805 (
		_w1576_,
		_w1578_,
		_w1579_,
		_w1580_
	);
	LUT4 #(
		.INIT('ha800)
	) name806 (
		\g35_pad ,
		_w1539_,
		_w1541_,
		_w1569_,
		_w1581_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		\g1890_reg/NET0131 ,
		\g35_pad ,
		_w1582_
	);
	LUT4 #(
		.INIT('h5700)
	) name808 (
		\g1936_reg/NET0131 ,
		_w1539_,
		_w1541_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\g1878_reg/NET0131 ,
		\g35_pad ,
		_w1584_
	);
	LUT3 #(
		.INIT('hfe)
	) name810 (
		_w1581_,
		_w1583_,
		_w1584_,
		_w1585_
	);
	LUT3 #(
		.INIT('h2a)
	) name811 (
		\g1996_reg/NET0131 ,
		_w802_,
		_w1241_,
		_w1586_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		\g1087_reg/NET0131 ,
		\g1996_reg/NET0131 ,
		_w1587_
	);
	LUT3 #(
		.INIT('h70)
	) name813 (
		_w1210_,
		_w1243_,
		_w1587_,
		_w1588_
	);
	LUT4 #(
		.INIT('h0020)
	) name814 (
		\g1242_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		\g956_reg/NET0131 ,
		_w1589_
	);
	LUT3 #(
		.INIT('h15)
	) name815 (
		\g2040_reg/NET0131 ,
		_w802_,
		_w1589_,
		_w1590_
	);
	LUT4 #(
		.INIT('ha800)
	) name816 (
		\g35_pad ,
		_w1586_,
		_w1588_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('h8)
	) name817 (
		\g2004_reg/NET0131 ,
		\g35_pad ,
		_w1592_
	);
	LUT4 #(
		.INIT('hab00)
	) name818 (
		\g2040_reg/NET0131 ,
		_w1586_,
		_w1588_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		\g2008_reg/NET0131 ,
		\g35_pad ,
		_w1594_
	);
	LUT3 #(
		.INIT('hfe)
	) name820 (
		_w1591_,
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT3 #(
		.INIT('h70)
	) name821 (
		_w802_,
		_w1241_,
		_w1246_,
		_w1596_
	);
	LUT3 #(
		.INIT('h02)
	) name822 (
		\g1087_reg/NET0131 ,
		\g1996_reg/NET0131 ,
		\g2070_reg/NET0131 ,
		_w1597_
	);
	LUT3 #(
		.INIT('h70)
	) name823 (
		_w1210_,
		_w1243_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\g2008_reg/NET0131 ,
		\g35_pad ,
		_w1599_
	);
	LUT3 #(
		.INIT('h2a)
	) name825 (
		\g35_pad ,
		_w802_,
		_w1589_,
		_w1600_
	);
	LUT4 #(
		.INIT('h01ef)
	) name826 (
		_w1596_,
		_w1598_,
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		\g2089_reg/NET0131 ,
		\g35_pad ,
		_w1602_
	);
	LUT2 #(
		.INIT('hd)
	) name828 (
		_w1601_,
		_w1602_,
		_w1603_
	);
	LUT3 #(
		.INIT('h2a)
	) name829 (
		\g2040_reg/NET0131 ,
		_w802_,
		_w1241_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		\g1087_reg/NET0131 ,
		\g2040_reg/NET0131 ,
		_w1605_
	);
	LUT3 #(
		.INIT('h70)
	) name831 (
		_w1210_,
		_w1243_,
		_w1605_,
		_w1606_
	);
	LUT3 #(
		.INIT('h15)
	) name832 (
		\g2070_reg/NET0131 ,
		_w802_,
		_w1589_,
		_w1607_
	);
	LUT4 #(
		.INIT('ha800)
	) name833 (
		\g35_pad ,
		_w1604_,
		_w1606_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		\g2012_reg/NET0131 ,
		\g35_pad ,
		_w1609_
	);
	LUT4 #(
		.INIT('hab00)
	) name835 (
		\g2070_reg/NET0131 ,
		_w1604_,
		_w1606_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h2)
	) name836 (
		\g2004_reg/NET0131 ,
		\g35_pad ,
		_w1611_
	);
	LUT3 #(
		.INIT('hfe)
	) name837 (
		_w1608_,
		_w1610_,
		_w1611_,
		_w1612_
	);
	LUT3 #(
		.INIT('h2a)
	) name838 (
		\g2070_reg/NET0131 ,
		_w802_,
		_w1589_,
		_w1613_
	);
	LUT4 #(
		.INIT('ha800)
	) name839 (
		\g35_pad ,
		_w1586_,
		_w1588_,
		_w1613_,
		_w1614_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		\g2016_reg/NET0131 ,
		\g35_pad ,
		_w1615_
	);
	LUT4 #(
		.INIT('h5700)
	) name841 (
		\g2070_reg/NET0131 ,
		_w1586_,
		_w1588_,
		_w1615_,
		_w1616_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		\g2020_reg/NET0131 ,
		\g35_pad ,
		_w1617_
	);
	LUT3 #(
		.INIT('hfe)
	) name843 (
		_w1614_,
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT3 #(
		.INIT('h15)
	) name844 (
		\g1996_reg/NET0131 ,
		_w802_,
		_w1589_,
		_w1619_
	);
	LUT4 #(
		.INIT('ha800)
	) name845 (
		\g35_pad ,
		_w1604_,
		_w1606_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		\g2020_reg/NET0131 ,
		\g35_pad ,
		_w1621_
	);
	LUT4 #(
		.INIT('hab00)
	) name847 (
		\g1996_reg/NET0131 ,
		_w1604_,
		_w1606_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h2)
	) name848 (
		\g2024_reg/NET0131 ,
		\g35_pad ,
		_w1623_
	);
	LUT3 #(
		.INIT('hfe)
	) name849 (
		_w1620_,
		_w1622_,
		_w1623_,
		_w1624_
	);
	LUT3 #(
		.INIT('h15)
	) name850 (
		\g2040_reg/NET0131 ,
		_w802_,
		_w1241_,
		_w1625_
	);
	LUT2 #(
		.INIT('h2)
	) name851 (
		\g1087_reg/NET0131 ,
		\g2040_reg/NET0131 ,
		_w1626_
	);
	LUT3 #(
		.INIT('h70)
	) name852 (
		_w1210_,
		_w1243_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('h8880)
	) name853 (
		\g35_pad ,
		_w1613_,
		_w1625_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h8)
	) name854 (
		\g2024_reg/NET0131 ,
		\g35_pad ,
		_w1629_
	);
	LUT4 #(
		.INIT('h5700)
	) name855 (
		\g2070_reg/NET0131 ,
		_w1625_,
		_w1627_,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('h2)
	) name856 (
		\g2012_reg/NET0131 ,
		\g35_pad ,
		_w1631_
	);
	LUT3 #(
		.INIT('hfe)
	) name857 (
		_w1628_,
		_w1630_,
		_w1631_,
		_w1632_
	);
	LUT3 #(
		.INIT('h10)
	) name858 (
		\g1135_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1633_
	);
	LUT3 #(
		.INIT('h2a)
	) name859 (
		\g1592_reg/NET0131 ,
		_w802_,
		_w1633_,
		_w1634_
	);
	LUT4 #(
		.INIT('h0002)
	) name860 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1216_reg/NET0131 ,
		_w1635_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		\g1592_reg/NET0131 ,
		\g17291_pad ,
		_w1636_
	);
	LUT3 #(
		.INIT('h70)
	) name862 (
		_w1210_,
		_w1635_,
		_w1636_,
		_w1637_
	);
	LUT4 #(
		.INIT('h0100)
	) name863 (
		\g1135_reg/NET0131 ,
		\g1242_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1638_
	);
	LUT3 #(
		.INIT('h15)
	) name864 (
		\g1636_reg/NET0131 ,
		_w802_,
		_w1638_,
		_w1639_
	);
	LUT4 #(
		.INIT('ha800)
	) name865 (
		\g35_pad ,
		_w1634_,
		_w1637_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\g1600_reg/NET0131 ,
		\g35_pad ,
		_w1641_
	);
	LUT4 #(
		.INIT('hab00)
	) name867 (
		\g1636_reg/NET0131 ,
		_w1634_,
		_w1637_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h2)
	) name868 (
		\g1604_reg/NET0131 ,
		\g35_pad ,
		_w1643_
	);
	LUT3 #(
		.INIT('hfe)
	) name869 (
		_w1640_,
		_w1642_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		\g1592_reg/NET0131 ,
		\g1668_reg/NET0131 ,
		_w1645_
	);
	LUT3 #(
		.INIT('h70)
	) name871 (
		_w802_,
		_w1633_,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h10)
	) name872 (
		\g1592_reg/NET0131 ,
		\g1668_reg/NET0131 ,
		\g17291_pad ,
		_w1647_
	);
	LUT3 #(
		.INIT('h70)
	) name873 (
		_w1210_,
		_w1635_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		\g1604_reg/NET0131 ,
		\g35_pad ,
		_w1649_
	);
	LUT3 #(
		.INIT('h2a)
	) name875 (
		\g35_pad ,
		_w802_,
		_w1638_,
		_w1650_
	);
	LUT4 #(
		.INIT('h01ef)
	) name876 (
		_w1646_,
		_w1648_,
		_w1649_,
		_w1650_,
		_w1651_
	);
	LUT2 #(
		.INIT('h2)
	) name877 (
		\g1687_reg/NET0131 ,
		\g35_pad ,
		_w1652_
	);
	LUT2 #(
		.INIT('hd)
	) name878 (
		_w1651_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('h2a)
	) name879 (
		\g1636_reg/NET0131 ,
		_w802_,
		_w1633_,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		\g1636_reg/NET0131 ,
		\g17291_pad ,
		_w1655_
	);
	LUT3 #(
		.INIT('h70)
	) name881 (
		_w1210_,
		_w1635_,
		_w1655_,
		_w1656_
	);
	LUT3 #(
		.INIT('h15)
	) name882 (
		\g1668_reg/NET0131 ,
		_w802_,
		_w1638_,
		_w1657_
	);
	LUT4 #(
		.INIT('ha800)
	) name883 (
		\g35_pad ,
		_w1654_,
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		\g1608_reg/NET0131 ,
		\g35_pad ,
		_w1659_
	);
	LUT4 #(
		.INIT('hab00)
	) name885 (
		\g1668_reg/NET0131 ,
		_w1654_,
		_w1656_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h2)
	) name886 (
		\g1600_reg/NET0131 ,
		\g35_pad ,
		_w1661_
	);
	LUT3 #(
		.INIT('hfe)
	) name887 (
		_w1658_,
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT3 #(
		.INIT('h2a)
	) name888 (
		\g1668_reg/NET0131 ,
		_w802_,
		_w1638_,
		_w1663_
	);
	LUT4 #(
		.INIT('ha800)
	) name889 (
		\g35_pad ,
		_w1634_,
		_w1637_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		\g1612_reg/NET0131 ,
		\g35_pad ,
		_w1665_
	);
	LUT4 #(
		.INIT('h5700)
	) name891 (
		\g1668_reg/NET0131 ,
		_w1634_,
		_w1637_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name892 (
		\g1616_reg/NET0131 ,
		\g35_pad ,
		_w1667_
	);
	LUT3 #(
		.INIT('hfe)
	) name893 (
		_w1664_,
		_w1666_,
		_w1667_,
		_w1668_
	);
	LUT3 #(
		.INIT('h15)
	) name894 (
		\g1592_reg/NET0131 ,
		_w802_,
		_w1638_,
		_w1669_
	);
	LUT4 #(
		.INIT('ha800)
	) name895 (
		\g35_pad ,
		_w1654_,
		_w1656_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		\g1616_reg/NET0131 ,
		\g35_pad ,
		_w1671_
	);
	LUT4 #(
		.INIT('hab00)
	) name897 (
		\g1592_reg/NET0131 ,
		_w1654_,
		_w1656_,
		_w1671_,
		_w1672_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		\g1620_reg/NET0131 ,
		\g35_pad ,
		_w1673_
	);
	LUT3 #(
		.INIT('hfe)
	) name899 (
		_w1670_,
		_w1672_,
		_w1673_,
		_w1674_
	);
	LUT3 #(
		.INIT('h4c)
	) name900 (
		_w802_,
		_w809_,
		_w1633_,
		_w1675_
	);
	LUT3 #(
		.INIT('h40)
	) name901 (
		\g1636_reg/NET0131 ,
		\g1668_reg/NET0131 ,
		\g17291_pad ,
		_w1676_
	);
	LUT3 #(
		.INIT('h70)
	) name902 (
		_w1210_,
		_w1635_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		\g1620_reg/NET0131 ,
		\g35_pad ,
		_w1678_
	);
	LUT4 #(
		.INIT('h5457)
	) name904 (
		_w1650_,
		_w1675_,
		_w1677_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\g1608_reg/NET0131 ,
		\g35_pad ,
		_w1680_
	);
	LUT2 #(
		.INIT('hd)
	) name906 (
		_w1679_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h4)
	) name907 (
		\g35_pad ,
		\g790_reg/NET0131 ,
		_w1682_
	);
	LUT3 #(
		.INIT('h8c)
	) name908 (
		\g736_reg/NET0131 ,
		\g794_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1683_
	);
	LUT3 #(
		.INIT('h07)
	) name909 (
		_w896_,
		_w899_,
		_w1683_,
		_w1684_
	);
	LUT3 #(
		.INIT('h2a)
	) name910 (
		\g35_pad ,
		_w896_,
		_w900_,
		_w1685_
	);
	LUT3 #(
		.INIT('hba)
	) name911 (
		_w1682_,
		_w1684_,
		_w1685_,
		_w1686_
	);
	LUT3 #(
		.INIT('hac)
	) name912 (
		\g12923_pad ,
		\g1585_reg/NET0131 ,
		\g35_pad ,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name913 (
		\g513_reg/NET0131 ,
		\g518_reg/NET0131 ,
		_w1688_
	);
	LUT3 #(
		.INIT('h20)
	) name914 (
		\g203_reg/NET0131 ,
		\g513_reg/NET0131 ,
		\g518_reg/NET0131 ,
		_w1689_
	);
	LUT3 #(
		.INIT('h01)
	) name915 (
		\g168_reg/NET0131 ,
		\g174_reg/NET0131 ,
		\g182_reg/NET0131 ,
		_w1690_
	);
	LUT3 #(
		.INIT('ha2)
	) name916 (
		\g691_reg/NET0131 ,
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h04)
	) name917 (
		_w889_,
		_w890_,
		_w892_,
		_w1692_
	);
	LUT3 #(
		.INIT('h80)
	) name918 (
		_w879_,
		_w881_,
		_w886_,
		_w1693_
	);
	LUT3 #(
		.INIT('h2a)
	) name919 (
		_w1691_,
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT4 #(
		.INIT('h0800)
	) name920 (
		\g146_reg/NET0131 ,
		\g203_reg/NET0131 ,
		\g513_reg/NET0131 ,
		\g518_reg/NET0131 ,
		_w1695_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		\g164_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1696_
	);
	LUT4 #(
		.INIT('hd000)
	) name922 (
		_w1689_,
		_w1690_,
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h8)
	) name923 (
		\g150_reg/NET0131 ,
		\g153_reg/NET0131 ,
		_w1698_
	);
	LUT3 #(
		.INIT('h40)
	) name924 (
		\g160_reg/NET0131 ,
		_w1697_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('ha222)
	) name925 (
		\g157_reg/NET0131 ,
		\g35_pad ,
		_w1694_,
		_w1699_,
		_w1700_
	);
	LUT3 #(
		.INIT('h80)
	) name926 (
		\g157_reg/NET0131 ,
		_w1697_,
		_w1698_,
		_w1701_
	);
	LUT2 #(
		.INIT('h8)
	) name927 (
		\g160_reg/NET0131 ,
		\g35_pad ,
		_w1702_
	);
	LUT4 #(
		.INIT('ha200)
	) name928 (
		\g691_reg/NET0131 ,
		_w1689_,
		_w1690_,
		_w1702_,
		_w1703_
	);
	LUT3 #(
		.INIT('h70)
	) name929 (
		_w1692_,
		_w1693_,
		_w1703_,
		_w1704_
	);
	LUT3 #(
		.INIT('h70)
	) name930 (
		_w1694_,
		_w1701_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('he)
	) name931 (
		_w1700_,
		_w1705_,
		_w1706_
	);
	LUT3 #(
		.INIT('h10)
	) name932 (
		\g225_reg/NET0131 ,
		\g232_reg/NET0131 ,
		\g255_reg/NET0131 ,
		_w1707_
	);
	LUT4 #(
		.INIT('h1000)
	) name933 (
		\g239_reg/NET0131 ,
		\g246_reg/NET0131 ,
		\g262_reg/NET0131 ,
		\g269_reg/NET0131 ,
		_w1708_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		\g278_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1709_
	);
	LUT3 #(
		.INIT('h80)
	) name935 (
		_w1707_,
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT3 #(
		.INIT('h08)
	) name936 (
		\g225_reg/NET0131 ,
		\g246_reg/NET0131 ,
		\g269_reg/NET0131 ,
		_w1711_
	);
	LUT4 #(
		.INIT('h0008)
	) name937 (
		\g232_reg/NET0131 ,
		\g239_reg/NET0131 ,
		\g255_reg/NET0131 ,
		\g262_reg/NET0131 ,
		_w1712_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		\g278_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1713_
	);
	LUT3 #(
		.INIT('h80)
	) name939 (
		_w1711_,
		_w1712_,
		_w1713_,
		_w1714_
	);
	LUT4 #(
		.INIT('h7770)
	) name940 (
		_w1692_,
		_w1693_,
		_w1710_,
		_w1714_,
		_w1715_
	);
	LUT3 #(
		.INIT('h80)
	) name941 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		\g291_reg/NET0131 ,
		_w1716_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		\g294_reg/NET0131 ,
		\g298_reg/NET0131 ,
		_w1717_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		_w1716_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		\g142_reg/NET0131 ,
		\g35_pad ,
		_w1719_
	);
	LUT3 #(
		.INIT('h20)
	) name945 (
		_w1715_,
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		\g142_reg/NET0131 ,
		\g35_pad ,
		_w1721_
	);
	LUT2 #(
		.INIT('h2)
	) name947 (
		\g298_reg/NET0131 ,
		\g35_pad ,
		_w1722_
	);
	LUT4 #(
		.INIT('h007f)
	) name948 (
		_w1715_,
		_w1718_,
		_w1721_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('hb)
	) name949 (
		_w1720_,
		_w1723_,
		_w1724_
	);
	LUT3 #(
		.INIT('hec)
	) name950 (
		\g35_pad ,
		\g4540_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1725_
	);
	LUT4 #(
		.INIT('hca00)
	) name951 (
		\g10500_pad ,
		\g12919_pad ,
		\g17400_pad ,
		\g35_pad ,
		_w1726_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		\g1246_reg/NET0131 ,
		\g35_pad ,
		_w1727_
	);
	LUT2 #(
		.INIT('he)
	) name953 (
		_w1726_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		\g1052_reg/NET0131 ,
		\g35_pad ,
		_w1729_
	);
	LUT3 #(
		.INIT('h01)
	) name955 (
		\g19334_pad ,
		\g7916_pad ,
		\g990_reg/NET0131 ,
		_w1730_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		\g1052_reg/NET0131 ,
		\g12919_pad ,
		_w1731_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		\g35_pad ,
		\g979_reg/NET0131 ,
		_w1732_
	);
	LUT4 #(
		.INIT('h9a00)
	) name958 (
		\g1061_reg/NET0131 ,
		_w1730_,
		_w1731_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('he)
	) name959 (
		_w1729_,
		_w1733_,
		_w1734_
	);
	LUT3 #(
		.INIT('hac)
	) name960 (
		\g12923_pad ,
		\g1579_reg/NET0131 ,
		\g35_pad ,
		_w1735_
	);
	LUT3 #(
		.INIT('h8c)
	) name961 (
		\g736_reg/NET0131 ,
		\g781_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1736_
	);
	LUT4 #(
		.INIT('h080c)
	) name962 (
		\g736_reg/NET0131 ,
		\g781_reg/NET0131 ,
		\g790_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1737_
	);
	LUT4 #(
		.INIT('hc444)
	) name963 (
		\g35_pad ,
		\g785_reg/NET0131 ,
		_w896_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('h80c0)
	) name964 (
		\g736_reg/NET0131 ,
		\g781_reg/NET0131 ,
		\g785_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1739_
	);
	LUT4 #(
		.INIT('h80a0)
	) name965 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g790_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1740_
	);
	LUT3 #(
		.INIT('h70)
	) name966 (
		_w896_,
		_w1739_,
		_w1740_,
		_w1741_
	);
	LUT2 #(
		.INIT('he)
	) name967 (
		_w1738_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('ha222)
	) name968 (
		\g160_reg/NET0131 ,
		\g35_pad ,
		_w1694_,
		_w1701_,
		_w1743_
	);
	LUT3 #(
		.INIT('hec)
	) name969 (
		\g35_pad ,
		\g4480_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1744_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		\g1061_reg/NET0131 ,
		\g35_pad ,
		_w1745_
	);
	LUT4 #(
		.INIT('h1000)
	) name971 (
		\g1052_reg/NET0131 ,
		\g1061_reg/NET0131 ,
		\g12919_pad ,
		\g19334_pad ,
		_w1746_
	);
	LUT4 #(
		.INIT('h2000)
	) name972 (
		\g1061_reg/NET0131 ,
		\g12919_pad ,
		\g19334_pad ,
		\g35_pad ,
		_w1747_
	);
	LUT3 #(
		.INIT('h01)
	) name973 (
		_w1745_,
		_w1746_,
		_w1747_,
		_w1748_
	);
	LUT3 #(
		.INIT('h69)
	) name974 (
		\g225_reg/NET0131 ,
		\g232_reg/NET0131 ,
		\g255_reg/NET0131 ,
		_w1749_
	);
	LUT2 #(
		.INIT('h9)
	) name975 (
		\g246_reg/NET0131 ,
		\g269_reg/NET0131 ,
		_w1750_
	);
	LUT2 #(
		.INIT('h6)
	) name976 (
		_w1749_,
		_w1750_,
		_w1751_
	);
	LUT4 #(
		.INIT('h2000)
	) name977 (
		\g358_reg/NET0131 ,
		\g370_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w1752_
	);
	LUT2 #(
		.INIT('h9)
	) name978 (
		\g239_reg/NET0131 ,
		\g262_reg/NET0131 ,
		_w1753_
	);
	LUT3 #(
		.INIT('h90)
	) name979 (
		\g239_reg/NET0131 ,
		\g262_reg/NET0131 ,
		\g732_reg/NET0131 ,
		_w1754_
	);
	LUT4 #(
		.INIT('h7f00)
	) name980 (
		_w879_,
		_w880_,
		_w1752_,
		_w1754_,
		_w1755_
	);
	LUT3 #(
		.INIT('h06)
	) name981 (
		\g239_reg/NET0131 ,
		\g262_reg/NET0131 ,
		\g732_reg/NET0131 ,
		_w1756_
	);
	LUT4 #(
		.INIT('h0080)
	) name982 (
		_w879_,
		_w880_,
		_w1752_,
		_w1753_,
		_w1757_
	);
	LUT4 #(
		.INIT('haaa8)
	) name983 (
		_w1751_,
		_w1755_,
		_w1756_,
		_w1757_,
		_w1758_
	);
	LUT4 #(
		.INIT('h0001)
	) name984 (
		_w1751_,
		_w1755_,
		_w1756_,
		_w1757_,
		_w1759_
	);
	LUT3 #(
		.INIT('h02)
	) name985 (
		\g35_pad ,
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name986 (
		\g153_reg/NET0131 ,
		\g35_pad ,
		_w1761_
	);
	LUT4 #(
		.INIT('h2a00)
	) name987 (
		\g150_reg/NET0131 ,
		_w1692_,
		_w1693_,
		_w1697_,
		_w1762_
	);
	LUT2 #(
		.INIT('h4)
	) name988 (
		\g157_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1763_
	);
	LUT4 #(
		.INIT('ha200)
	) name989 (
		\g153_reg/NET0131 ,
		_w1689_,
		_w1690_,
		_w1763_,
		_w1764_
	);
	LUT3 #(
		.INIT('h15)
	) name990 (
		_w1761_,
		_w1762_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		\g157_reg/NET0131 ,
		\g35_pad ,
		_w1766_
	);
	LUT3 #(
		.INIT('h70)
	) name992 (
		_w1697_,
		_w1698_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		_w1694_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('hd)
	) name994 (
		_w1765_,
		_w1768_,
		_w1769_
	);
	LUT3 #(
		.INIT('h80)
	) name995 (
		\g35_pad ,
		_w896_,
		_w1739_,
		_w1770_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name996 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g785_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1771_
	);
	LUT3 #(
		.INIT('h70)
	) name997 (
		_w896_,
		_w1736_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		\g35_pad ,
		\g781_reg/NET0131 ,
		_w1773_
	);
	LUT3 #(
		.INIT('h01)
	) name999 (
		_w1770_,
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		\g1052_reg/NET0131 ,
		\g12919_pad ,
		_w1775_
	);
	LUT4 #(
		.INIT('h0001)
	) name1001 (
		\g1052_reg/NET0131 ,
		\g19334_pad ,
		\g7916_pad ,
		\g990_reg/NET0131 ,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1775_,
		_w1776_,
		_w1777_
	);
	LUT3 #(
		.INIT('hb0)
	) name1003 (
		_w1730_,
		_w1731_,
		_w1732_,
		_w1778_
	);
	LUT2 #(
		.INIT('h8)
	) name1004 (
		_w1777_,
		_w1778_,
		_w1779_
	);
	LUT3 #(
		.INIT('h13)
	) name1005 (
		\g35_pad ,
		\g4434_reg/NET0131 ,
		\g4443_reg/NET0131 ,
		_w1780_
	);
	LUT3 #(
		.INIT('h01)
	) name1006 (
		\g4452_reg/NET0131 ,
		\g7245_pad ,
		\g7260_pad ,
		_w1781_
	);
	LUT3 #(
		.INIT('h02)
	) name1007 (
		\g4392_reg/NET0131 ,
		\g4438_reg/NET0131 ,
		\g4443_reg/NET0131 ,
		_w1782_
	);
	LUT2 #(
		.INIT('h2)
	) name1008 (
		\g35_pad ,
		\g4443_reg/NET0131 ,
		_w1783_
	);
	LUT4 #(
		.INIT('h4055)
	) name1009 (
		_w1780_,
		_w1781_,
		_w1782_,
		_w1783_,
		_w1784_
	);
	LUT2 #(
		.INIT('h2)
	) name1010 (
		\g329_reg/NET0131 ,
		\g35_pad ,
		_w1785_
	);
	LUT4 #(
		.INIT('h0001)
	) name1011 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		\g319_reg/NET0131 ,
		\g329_reg/NET0131 ,
		_w1786_
	);
	LUT4 #(
		.INIT('h0503)
	) name1012 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		\g319_reg/NET0131 ,
		\g336_reg/NET0131 ,
		_w1787_
	);
	LUT3 #(
		.INIT('hac)
	) name1013 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		\g324_reg/NET0131 ,
		_w1788_
	);
	LUT4 #(
		.INIT('h7577)
	) name1014 (
		\g35_pad ,
		_w1786_,
		_w1787_,
		_w1788_,
		_w1789_
	);
	LUT2 #(
		.INIT('hb)
	) name1015 (
		_w1785_,
		_w1789_,
		_w1790_
	);
	LUT3 #(
		.INIT('h08)
	) name1016 (
		\g4621_reg/NET0131 ,
		\g4628_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w1791_
	);
	LUT2 #(
		.INIT('h8)
	) name1017 (
		\g4340_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		_w1792_
	);
	LUT3 #(
		.INIT('h80)
	) name1018 (
		\g4340_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		\g4358_reg/NET0131 ,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		_w1794_
	);
	LUT4 #(
		.INIT('h8000)
	) name1020 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		\g4584_reg/NET0131 ,
		\g4593_reg/NET0131 ,
		_w1795_
	);
	LUT3 #(
		.INIT('h80)
	) name1021 (
		_w1791_,
		_w1793_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		\g4601_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		_w1797_
	);
	LUT4 #(
		.INIT('h8000)
	) name1023 (
		_w1791_,
		_w1793_,
		_w1795_,
		_w1797_,
		_w1798_
	);
	LUT3 #(
		.INIT('h80)
	) name1024 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		\g4584_reg/NET0131 ,
		_w1799_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		\g35_pad ,
		\g4616_reg/NET0131 ,
		_w1800_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1026 (
		_w1791_,
		_w1793_,
		_w1799_,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		_w1798_,
		_w1801_,
		_w1802_
	);
	LUT2 #(
		.INIT('h2)
	) name1028 (
		\g4601_reg/NET0131 ,
		\g4616_reg/NET0131 ,
		_w1803_
	);
	LUT4 #(
		.INIT('h8000)
	) name1029 (
		_w1791_,
		_w1793_,
		_w1795_,
		_w1803_,
		_w1804_
	);
	LUT3 #(
		.INIT('hc4)
	) name1030 (
		\g35_pad ,
		\g4608_reg/NET0131 ,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('he)
	) name1031 (
		_w1802_,
		_w1805_,
		_w1806_
	);
	LUT3 #(
		.INIT('h28)
	) name1032 (
		\g35_pad ,
		\g4401_reg/NET0131 ,
		\g4434_reg/NET0131 ,
		_w1807_
	);
	LUT3 #(
		.INIT('h87)
	) name1033 (
		\g35_pad ,
		\g4388_reg/NET0131 ,
		\g4430_reg/NET0131 ,
		_w1808_
	);
	LUT2 #(
		.INIT('hb)
	) name1034 (
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT3 #(
		.INIT('hca)
	) name1035 (
		\g1242_reg/NET0131 ,
		\g12919_pad ,
		\g35_pad ,
		_w1810_
	);
	LUT4 #(
		.INIT('h0080)
	) name1036 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		\g291_reg/NET0131 ,
		\g298_reg/NET0131 ,
		_w1811_
	);
	LUT4 #(
		.INIT('ha222)
	) name1037 (
		\g294_reg/NET0131 ,
		\g35_pad ,
		_w1715_,
		_w1811_,
		_w1812_
	);
	LUT4 #(
		.INIT('h8000)
	) name1038 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		\g291_reg/NET0131 ,
		\g294_reg/NET0131 ,
		_w1813_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		\g298_reg/NET0131 ,
		\g35_pad ,
		_w1814_
	);
	LUT3 #(
		.INIT('h20)
	) name1040 (
		_w1715_,
		_w1813_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('he)
	) name1041 (
		_w1812_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h080c)
	) name1042 (
		\g736_reg/NET0131 ,
		\g772_reg/NET0131 ,
		\g781_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1817_
	);
	LUT4 #(
		.INIT('h8000)
	) name1043 (
		_w882_,
		_w888_,
		_w893_,
		_w1817_,
		_w1818_
	);
	LUT3 #(
		.INIT('hc4)
	) name1044 (
		\g35_pad ,
		\g776_reg/NET0131 ,
		_w1818_,
		_w1819_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1045 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g781_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1820_
	);
	LUT2 #(
		.INIT('h4)
	) name1046 (
		_w896_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('he)
	) name1047 (
		_w1819_,
		_w1821_,
		_w1822_
	);
	LUT4 #(
		.INIT('hfad8)
	) name1048 (
		\g35_pad ,
		\g4372_reg/NET0131 ,
		\g4423_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1823_
	);
	LUT4 #(
		.INIT('h8000)
	) name1049 (
		\g358_reg/NET0131 ,
		\g370_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name1050 (
		\g817_reg/NET0131 ,
		\g832_reg/NET0131 ,
		_w1825_
	);
	LUT3 #(
		.INIT('h80)
	) name1051 (
		\g817_reg/NET0131 ,
		\g822_reg/NET0131 ,
		\g832_reg/NET0131 ,
		_w1826_
	);
	LUT2 #(
		.INIT('h8)
	) name1052 (
		_w1824_,
		_w1826_,
		_w1827_
	);
	LUT3 #(
		.INIT('hb0)
	) name1053 (
		\g812_reg/NET0131 ,
		\g837_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w1828_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1054 (
		\g35_pad ,
		\g812_reg/NET0131 ,
		\g837_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w1829_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		\g723_reg/NET0131 ,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('h1055)
	) name1056 (
		\g723_reg/NET0131 ,
		\g812_reg/NET0131 ,
		\g837_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w1831_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1057 (
		\g35_pad ,
		_w1824_,
		_w1826_,
		_w1831_,
		_w1832_
	);
	LUT4 #(
		.INIT('h70fa)
	) name1058 (
		\g827_reg/NET0131 ,
		_w1827_,
		_w1830_,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h2)
	) name1059 (
		\g3263_reg/NET0131 ,
		\g35_pad ,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		\g3333_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		_w1835_
	);
	LUT2 #(
		.INIT('h4)
	) name1061 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1836_
	);
	LUT3 #(
		.INIT('h40)
	) name1062 (
		\g4709_reg/NET0131 ,
		\g4743_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1837_
	);
	LUT4 #(
		.INIT('h1000)
	) name1063 (
		\g3333_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4743_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1838_
	);
	LUT4 #(
		.INIT('h070f)
	) name1064 (
		_w824_,
		_w825_,
		_w1835_,
		_w1838_,
		_w1839_
	);
	LUT3 #(
		.INIT('h1d)
	) name1065 (
		\g3263_reg/NET0131 ,
		\g35_pad ,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h2)
	) name1066 (
		\g3288_reg/NET0131 ,
		_w840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		_w839_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h1)
	) name1068 (
		\g3288_reg/NET0131 ,
		_w846_,
		_w1843_
	);
	LUT3 #(
		.INIT('h2a)
	) name1069 (
		\g3352_reg/NET0131 ,
		_w845_,
		_w1843_,
		_w1844_
	);
	LUT4 #(
		.INIT('h70f0)
	) name1070 (
		\g13865_pad ,
		\g3231_reg/NET0131 ,
		\g3288_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w1845_
	);
	LUT3 #(
		.INIT('he0)
	) name1071 (
		\g3338_reg/NET0131 ,
		_w852_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h4)
	) name1072 (
		_w851_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h0f07)
	) name1073 (
		\g13865_pad ,
		\g3239_reg/NET0131 ,
		\g3288_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w1848_
	);
	LUT3 #(
		.INIT('hd0)
	) name1074 (
		\g3338_reg/NET0131 ,
		_w859_,
		_w1848_,
		_w1849_
	);
	LUT3 #(
		.INIT('h45)
	) name1075 (
		\g3352_reg/NET0131 ,
		_w858_,
		_w1849_,
		_w1850_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1076 (
		_w1842_,
		_w1844_,
		_w1847_,
		_w1850_,
		_w1851_
	);
	LUT3 #(
		.INIT('h80)
	) name1077 (
		_w824_,
		_w825_,
		_w1837_,
		_w1852_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1078 (
		\g4674_reg/NET0131 ,
		_w824_,
		_w825_,
		_w1837_,
		_w1853_
	);
	LUT2 #(
		.INIT('h4)
	) name1079 (
		_w1834_,
		_w1853_,
		_w1854_
	);
	LUT3 #(
		.INIT('h15)
	) name1080 (
		_w1840_,
		_w1851_,
		_w1854_,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		\g3684_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		_w1856_
	);
	LUT2 #(
		.INIT('h2)
	) name1082 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1857_
	);
	LUT3 #(
		.INIT('h08)
	) name1083 (
		\g4709_reg/NET0131 ,
		\g4754_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1858_
	);
	LUT4 #(
		.INIT('h0040)
	) name1084 (
		\g3684_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4754_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1859_
	);
	LUT4 #(
		.INIT('h070f)
	) name1085 (
		_w824_,
		_w825_,
		_w1856_,
		_w1859_,
		_w1860_
	);
	LUT3 #(
		.INIT('h1d)
	) name1086 (
		\g3263_reg/NET0131 ,
		\g35_pad ,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		\g3703_reg/NET0131 ,
		_w840_,
		_w1862_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		_w839_,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('h007f)
	) name1089 (
		\g13865_pad ,
		\g3231_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g3703_reg/NET0131 ,
		_w1864_
	);
	LUT3 #(
		.INIT('he0)
	) name1090 (
		\g3338_reg/NET0131 ,
		_w852_,
		_w1864_,
		_w1865_
	);
	LUT3 #(
		.INIT('h8a)
	) name1091 (
		\g3639_reg/NET0131 ,
		_w851_,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h2)
	) name1092 (
		\g3703_reg/NET0131 ,
		_w846_,
		_w1867_
	);
	LUT2 #(
		.INIT('h8)
	) name1093 (
		_w845_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1094 (
		\g13865_pad ,
		\g3239_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g3703_reg/NET0131 ,
		_w1869_
	);
	LUT3 #(
		.INIT('hd0)
	) name1095 (
		\g3338_reg/NET0131 ,
		_w859_,
		_w1869_,
		_w1870_
	);
	LUT3 #(
		.INIT('h45)
	) name1096 (
		\g3639_reg/NET0131 ,
		_w858_,
		_w1870_,
		_w1871_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1097 (
		_w1863_,
		_w1866_,
		_w1868_,
		_w1871_,
		_w1872_
	);
	LUT3 #(
		.INIT('h80)
	) name1098 (
		_w824_,
		_w825_,
		_w1858_,
		_w1873_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1099 (
		\g4681_reg/NET0131 ,
		_w824_,
		_w825_,
		_w1858_,
		_w1874_
	);
	LUT2 #(
		.INIT('h4)
	) name1100 (
		_w1834_,
		_w1874_,
		_w1875_
	);
	LUT3 #(
		.INIT('h15)
	) name1101 (
		_w1861_,
		_w1872_,
		_w1875_,
		_w1876_
	);
	LUT4 #(
		.INIT('hfad8)
	) name1102 (
		\g35_pad ,
		\g4372_reg/NET0131 ,
		\g4477_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w1877_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		\g153_reg/NET0131 ,
		\g164_reg/NET0131 ,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name1104 (
		_w1695_,
		_w1878_,
		_w1879_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1105 (
		_w1691_,
		_w1692_,
		_w1693_,
		_w1879_,
		_w1880_
	);
	LUT3 #(
		.INIT('ha2)
	) name1106 (
		\g150_reg/NET0131 ,
		\g35_pad ,
		_w1880_,
		_w1881_
	);
	LUT4 #(
		.INIT('h8808)
	) name1107 (
		\g35_pad ,
		\g691_reg/NET0131 ,
		_w1689_,
		_w1690_,
		_w1882_
	);
	LUT3 #(
		.INIT('h70)
	) name1108 (
		_w1692_,
		_w1693_,
		_w1882_,
		_w1883_
	);
	LUT3 #(
		.INIT('h20)
	) name1109 (
		\g153_reg/NET0131 ,
		_w1762_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('he)
	) name1110 (
		_w1881_,
		_w1884_,
		_w1885_
	);
	LUT3 #(
		.INIT('h23)
	) name1111 (
		\g736_reg/NET0131 ,
		\g776_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1886_
	);
	LUT4 #(
		.INIT('h8000)
	) name1112 (
		_w882_,
		_w888_,
		_w893_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('hc4)
	) name1113 (
		\g35_pad ,
		\g772_reg/NET0131 ,
		_w1887_,
		_w1888_
	);
	LUT4 #(
		.INIT('h8000)
	) name1114 (
		_w882_,
		_w888_,
		_w893_,
		_w894_,
		_w1889_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1115 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g776_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1890_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w1889_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('he)
	) name1117 (
		_w1888_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('hca)
	) name1118 (
		\g1236_reg/NET0131 ,
		\g12919_pad ,
		\g35_pad ,
		_w1893_
	);
	LUT3 #(
		.INIT('he2)
	) name1119 (
		\g1554_reg/NET0131 ,
		\g35_pad ,
		\g496_reg/NET0131 ,
		_w1894_
	);
	LUT2 #(
		.INIT('h4)
	) name1120 (
		\g35_pad ,
		\g4601_reg/NET0131 ,
		_w1895_
	);
	LUT4 #(
		.INIT('h8000)
	) name1121 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		\g4584_reg/NET0131 ,
		\g4616_reg/NET0131 ,
		_w1896_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1122 (
		\g35_pad ,
		_w1791_,
		_w1793_,
		_w1896_,
		_w1897_
	);
	LUT4 #(
		.INIT('h6c00)
	) name1123 (
		\g4601_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		_w1796_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('he)
	) name1124 (
		_w1895_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1125 (
		\g4035_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w1900_
	);
	LUT4 #(
		.INIT('h4000)
	) name1126 (
		\g4035_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4765_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1901_
	);
	LUT4 #(
		.INIT('h070f)
	) name1127 (
		_w824_,
		_w825_,
		_w1900_,
		_w1901_,
		_w1902_
	);
	LUT3 #(
		.INIT('h1d)
	) name1128 (
		\g3263_reg/NET0131 ,
		\g35_pad ,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1129 (
		\g4688_reg/NET0131 ,
		_w824_,
		_w825_,
		_w865_,
		_w1904_
	);
	LUT2 #(
		.INIT('h4)
	) name1130 (
		_w1834_,
		_w1904_,
		_w1905_
	);
	LUT3 #(
		.INIT('h13)
	) name1131 (
		_w863_,
		_w1903_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h2)
	) name1132 (
		\g29219_pad ,
		\g35_pad ,
		_w1907_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1133 (
		\g2741_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		\g35_pad ,
		_w1908_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		_w1907_,
		_w1908_,
		_w1909_
	);
	LUT4 #(
		.INIT('h8000)
	) name1135 (
		\g2735_reg/NET0131 ,
		\g2741_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w1910_
	);
	LUT3 #(
		.INIT('h54)
	) name1136 (
		\g2193_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w1911_
	);
	LUT3 #(
		.INIT('h51)
	) name1137 (
		\g2799_reg/NET0131 ,
		\g29219_pad ,
		\g35_pad ,
		_w1912_
	);
	LUT3 #(
		.INIT('hb0)
	) name1138 (
		_w1910_,
		_w1911_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		_w1909_,
		_w1913_,
		_w1914_
	);
	LUT3 #(
		.INIT('h08)
	) name1140 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		\g294_reg/NET0131 ,
		_w1915_
	);
	LUT4 #(
		.INIT('ha222)
	) name1141 (
		\g291_reg/NET0131 ,
		\g35_pad ,
		_w1715_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		\g294_reg/NET0131 ,
		\g35_pad ,
		_w1917_
	);
	LUT3 #(
		.INIT('h20)
	) name1143 (
		_w1715_,
		_w1716_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('he)
	) name1144 (
		_w1916_,
		_w1918_,
		_w1919_
	);
	LUT4 #(
		.INIT('h8000)
	) name1145 (
		\g772_reg/NET0131 ,
		_w882_,
		_w888_,
		_w893_,
		_w1920_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name1146 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g772_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1921_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1147 (
		_w882_,
		_w888_,
		_w893_,
		_w1921_,
		_w1922_
	);
	LUT4 #(
		.INIT('h004e)
	) name1148 (
		\g35_pad ,
		\g767_reg/NET0131 ,
		_w1920_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h2)
	) name1149 (
		\g29211_pad ,
		\g35_pad ,
		_w1924_
	);
	LUT3 #(
		.INIT('h20)
	) name1150 (
		\g329_reg/NET0131 ,
		\g341_reg/NET0131 ,
		\g35_pad ,
		_w1925_
	);
	LUT3 #(
		.INIT('hdc)
	) name1151 (
		_w1788_,
		_w1924_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		\g35_pad ,
		\g822_reg/NET0131 ,
		_w1927_
	);
	LUT2 #(
		.INIT('h8)
	) name1153 (
		\g35_pad ,
		\g827_reg/NET0131 ,
		_w1928_
	);
	LUT4 #(
		.INIT('h0700)
	) name1154 (
		_w1824_,
		_w1826_,
		_w1828_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h2)
	) name1155 (
		\g35_pad ,
		\g827_reg/NET0131 ,
		_w1930_
	);
	LUT4 #(
		.INIT('h0800)
	) name1156 (
		_w1824_,
		_w1826_,
		_w1828_,
		_w1930_,
		_w1931_
	);
	LUT3 #(
		.INIT('hfe)
	) name1157 (
		_w1927_,
		_w1929_,
		_w1931_,
		_w1932_
	);
	LUT2 #(
		.INIT('h2)
	) name1158 (
		\g164_reg/NET0131 ,
		\g35_pad ,
		_w1933_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		\g164_reg/NET0131 ,
		\g35_pad ,
		_w1934_
	);
	LUT3 #(
		.INIT('h2a)
	) name1160 (
		\g150_reg/NET0131 ,
		\g164_reg/NET0131 ,
		_w1695_,
		_w1935_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1161 (
		_w1691_,
		_w1692_,
		_w1693_,
		_w1935_,
		_w1936_
	);
	LUT3 #(
		.INIT('h0b)
	) name1162 (
		\g150_reg/NET0131 ,
		_w1697_,
		_w1933_,
		_w1937_
	);
	LUT3 #(
		.INIT('h45)
	) name1163 (
		_w1934_,
		_w1936_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		\g35_pad ,
		\g4674_reg/NET0131 ,
		_w1939_
	);
	LUT4 #(
		.INIT('h2000)
	) name1165 (
		\g35_pad ,
		\g4709_reg/NET0131 ,
		\g4743_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w1940_
	);
	LUT4 #(
		.INIT('h070f)
	) name1166 (
		_w824_,
		_w825_,
		_w1939_,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name1167 (
		\g4749_reg/NET0131 ,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name1168 (
		\g35_pad ,
		\g4674_reg/NET0131 ,
		_w1943_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1169 (
		_w824_,
		_w825_,
		_w1837_,
		_w1943_,
		_w1944_
	);
	LUT3 #(
		.INIT('h08)
	) name1170 (
		\g4776_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		\g4801_reg/NET0131 ,
		_w1945_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		_w822_,
		_w1945_,
		_w1946_
	);
	LUT3 #(
		.INIT('h35)
	) name1172 (
		\g3343_reg/NET0131 ,
		\g3347_reg/NET0131 ,
		\g3352_reg/NET0131 ,
		_w1947_
	);
	LUT3 #(
		.INIT('hde)
	) name1173 (
		\g3288_reg/NET0131 ,
		\g4749_reg/NET0131 ,
		_w1947_,
		_w1948_
	);
	LUT3 #(
		.INIT('h80)
	) name1174 (
		_w1944_,
		_w1946_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('he)
	) name1175 (
		_w1942_,
		_w1949_,
		_w1950_
	);
	LUT2 #(
		.INIT('h2)
	) name1176 (
		\g4771_reg/NET0131 ,
		_w876_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name1177 (
		_w1857_,
		_w1945_,
		_w1952_
	);
	LUT3 #(
		.INIT('h35)
	) name1178 (
		\g3343_reg/NET0131 ,
		\g3347_reg/NET0131 ,
		\g4054_reg/NET0131 ,
		_w1953_
	);
	LUT3 #(
		.INIT('hde)
	) name1179 (
		\g3990_reg/NET0131 ,
		\g4771_reg/NET0131 ,
		_w1953_,
		_w1954_
	);
	LUT3 #(
		.INIT('h80)
	) name1180 (
		_w868_,
		_w1952_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('he)
	) name1181 (
		_w1951_,
		_w1955_,
		_w1956_
	);
	LUT3 #(
		.INIT('h8c)
	) name1182 (
		\g736_reg/NET0131 ,
		\g739_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1957_
	);
	LUT4 #(
		.INIT('h8000)
	) name1183 (
		_w879_,
		_w881_,
		_w886_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h8)
	) name1184 (
		\g744_reg/NET0131 ,
		_w884_,
		_w1959_
	);
	LUT3 #(
		.INIT('h23)
	) name1185 (
		\g736_reg/NET0131 ,
		\g767_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1960_
	);
	LUT3 #(
		.INIT('h80)
	) name1186 (
		\g744_reg/NET0131 ,
		_w884_,
		_w1960_,
		_w1961_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1187 (
		\g35_pad ,
		_w893_,
		_w1958_,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name1188 (
		\g744_reg/NET0131 ,
		\g763_reg/NET0131 ,
		_w1963_
	);
	LUT2 #(
		.INIT('h8)
	) name1189 (
		_w884_,
		_w1963_,
		_w1964_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1190 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g767_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1965_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1191 (
		_w893_,
		_w1958_,
		_w1964_,
		_w1965_,
		_w1966_
	);
	LUT3 #(
		.INIT('hf2)
	) name1192 (
		\g763_reg/NET0131 ,
		_w1962_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h0100)
	) name1193 (
		\g1099_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1968_
	);
	LUT4 #(
		.INIT('h0200)
	) name1194 (
		\g1152_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w1969_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name1195 (
		\g1146_reg/NET0131 ,
		\g35_pad ,
		_w1968_,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h9)
	) name1196 (
		\g979_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name1197 (
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w1972_
	);
	LUT4 #(
		.INIT('h1110)
	) name1198 (
		\g1008_reg/NET0131 ,
		\g969_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w1973_
	);
	LUT2 #(
		.INIT('h9)
	) name1199 (
		\g1236_reg/NET0131 ,
		\g979_reg/NET0131 ,
		_w1974_
	);
	LUT3 #(
		.INIT('h04)
	) name1200 (
		_w1971_,
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT4 #(
		.INIT('h0001)
	) name1201 (
		\g13259_pad ,
		\g19334_pad ,
		\g7916_pad ,
		\g8416_pad ,
		_w1976_
	);
	LUT4 #(
		.INIT('h7d5f)
	) name1202 (
		\g35_pad ,
		\g990_reg/NET0131 ,
		_w1975_,
		_w1976_,
		_w1977_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		\g35_pad ,
		\g996_reg/NET0131 ,
		_w1978_
	);
	LUT2 #(
		.INIT('hd)
	) name1204 (
		_w1977_,
		_w1978_,
		_w1979_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		\g35_pad ,
		\g4664_reg/NET0131 ,
		_w1980_
	);
	LUT4 #(
		.INIT('h8000)
	) name1206 (
		\g4653_reg/NET0131 ,
		\g4659_reg/NET0131 ,
		\g4669_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w1981_
	);
	LUT4 #(
		.INIT('h8000)
	) name1207 (
		\g4653_reg/NET0131 ,
		\g4659_reg/NET0131 ,
		\g4664_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w1982_
	);
	LUT4 #(
		.INIT('h0a08)
	) name1208 (
		\g35_pad ,
		\g4669_reg/NET0131 ,
		_w1981_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('he)
	) name1209 (
		_w1980_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		\g287_reg/NET0131 ,
		\g35_pad ,
		_w1985_
	);
	LUT3 #(
		.INIT('h08)
	) name1211 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		\g291_reg/NET0131 ,
		_w1986_
	);
	LUT4 #(
		.INIT('h7000)
	) name1212 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		\g291_reg/NET0131 ,
		\g35_pad ,
		_w1987_
	);
	LUT4 #(
		.INIT('heeec)
	) name1213 (
		_w1715_,
		_w1985_,
		_w1986_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('h8000)
	) name1214 (
		\g35_pad ,
		_w893_,
		_w1958_,
		_w1964_,
		_w1989_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name1215 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g763_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w1990_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1216 (
		_w893_,
		_w1958_,
		_w1959_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		\g35_pad ,
		\g758_reg/NET0131 ,
		_w1992_
	);
	LUT3 #(
		.INIT('h01)
	) name1218 (
		_w1989_,
		_w1991_,
		_w1992_,
		_w1993_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		\g35_pad ,
		\g956_reg/NET0131 ,
		_w1994_
	);
	LUT2 #(
		.INIT('h2)
	) name1220 (
		\g1141_reg/NET0131 ,
		\g35_pad ,
		_w1995_
	);
	LUT3 #(
		.INIT('h08)
	) name1221 (
		\g1099_reg/NET0131 ,
		\g1141_reg/NET0131 ,
		\g1152_reg/NET0131 ,
		_w1996_
	);
	LUT4 #(
		.INIT('h363c)
	) name1222 (
		_w1099_,
		_w1994_,
		_w1995_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h8)
	) name1223 (
		\g1105_reg/NET0131 ,
		\g35_pad ,
		_w1998_
	);
	LUT2 #(
		.INIT('h2)
	) name1224 (
		\g1111_reg/NET0131 ,
		\g35_pad ,
		_w1999_
	);
	LUT3 #(
		.INIT('h08)
	) name1225 (
		\g1099_reg/NET0131 ,
		\g1111_reg/NET0131 ,
		\g1152_reg/NET0131 ,
		_w2000_
	);
	LUT4 #(
		.INIT('h363c)
	) name1226 (
		_w1087_,
		_w1998_,
		_w1999_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		\g1129_reg/NET0131 ,
		\g35_pad ,
		_w2002_
	);
	LUT2 #(
		.INIT('h2)
	) name1228 (
		\g1124_reg/NET0131 ,
		\g35_pad ,
		_w2003_
	);
	LUT3 #(
		.INIT('h08)
	) name1229 (
		\g1099_reg/NET0131 ,
		\g1124_reg/NET0131 ,
		\g1152_reg/NET0131 ,
		_w2004_
	);
	LUT4 #(
		.INIT('h363c)
	) name1230 (
		_w1093_,
		_w2002_,
		_w2003_,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h8)
	) name1231 (
		\g1135_reg/NET0131 ,
		\g35_pad ,
		_w2006_
	);
	LUT2 #(
		.INIT('h2)
	) name1232 (
		\g1094_reg/NET0131 ,
		\g35_pad ,
		_w2007_
	);
	LUT3 #(
		.INIT('h08)
	) name1233 (
		\g1094_reg/NET0131 ,
		\g1099_reg/NET0131 ,
		\g1152_reg/NET0131 ,
		_w2008_
	);
	LUT4 #(
		.INIT('h363c)
	) name1234 (
		_w1079_,
		_w2006_,
		_w2007_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h2)
	) name1235 (
		\g35_pad ,
		\g4681_reg/NET0131 ,
		_w2010_
	);
	LUT4 #(
		.INIT('h0080)
	) name1236 (
		\g35_pad ,
		\g4709_reg/NET0131 ,
		\g4754_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w2011_
	);
	LUT4 #(
		.INIT('h070f)
	) name1237 (
		_w824_,
		_w825_,
		_w2010_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h2)
	) name1238 (
		\g4760_reg/NET0131 ,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1239 (
		\g35_pad ,
		\g4681_reg/NET0131 ,
		_w2014_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1240 (
		_w824_,
		_w825_,
		_w1858_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		_w1836_,
		_w1945_,
		_w2016_
	);
	LUT3 #(
		.INIT('h35)
	) name1242 (
		\g3343_reg/NET0131 ,
		\g3347_reg/NET0131 ,
		\g3703_reg/NET0131 ,
		_w2017_
	);
	LUT3 #(
		.INIT('hde)
	) name1243 (
		\g3639_reg/NET0131 ,
		\g4760_reg/NET0131 ,
		_w2017_,
		_w2018_
	);
	LUT3 #(
		.INIT('h80)
	) name1244 (
		_w2015_,
		_w2016_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('he)
	) name1245 (
		_w2013_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h4)
	) name1246 (
		\g35_pad ,
		\g676_reg/NET0131 ,
		_w2021_
	);
	LUT2 #(
		.INIT('h8)
	) name1247 (
		\g482_reg/NET0131 ,
		\g490_reg/NET0131 ,
		_w2022_
	);
	LUT3 #(
		.INIT('h02)
	) name1248 (
		\g499_reg/NET0131 ,
		\g504_reg/NET0131 ,
		\g528_reg/NET0131 ,
		_w2023_
	);
	LUT3 #(
		.INIT('h80)
	) name1249 (
		_w1824_,
		_w2022_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h6)
	) name1250 (
		\g655_reg/NET0131 ,
		\g718_reg/NET0131 ,
		_w2025_
	);
	LUT2 #(
		.INIT('h6)
	) name1251 (
		\g661_reg/NET0131 ,
		\g728_reg/NET0131 ,
		_w2026_
	);
	LUT4 #(
		.INIT('h1000)
	) name1252 (
		\g645_reg/NET0131 ,
		\g650_reg/NET0131 ,
		\g681_reg/NET0131 ,
		\g699_reg/NET0131 ,
		_w2027_
	);
	LUT3 #(
		.INIT('h10)
	) name1253 (
		_w2025_,
		_w2026_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h8)
	) name1254 (
		\g35_pad ,
		\g703_reg/NET0131 ,
		_w2029_
	);
	LUT3 #(
		.INIT('h70)
	) name1255 (
		_w2024_,
		_w2028_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		\g671_reg/NET0131 ,
		\g676_reg/NET0131 ,
		_w2031_
	);
	LUT4 #(
		.INIT('h8000)
	) name1257 (
		_w1824_,
		_w2022_,
		_w2023_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h6)
	) name1258 (
		\g714_reg/NET0131 ,
		_w2032_,
		_w2033_
	);
	LUT3 #(
		.INIT('hea)
	) name1259 (
		_w2021_,
		_w2030_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h4)
	) name1260 (
		\g35_pad ,
		\g4593_reg/NET0131 ,
		_w2035_
	);
	LUT4 #(
		.INIT('hff60)
	) name1261 (
		\g4601_reg/NET0131 ,
		_w1796_,
		_w1897_,
		_w2035_,
		_w2036_
	);
	LUT3 #(
		.INIT('hac)
	) name1262 (
		\g269_reg/NET0131 ,
		\g29215_pad ,
		\g35_pad ,
		_w2037_
	);
	LUT2 #(
		.INIT('h2)
	) name1263 (
		\g1146_reg/NET0131 ,
		\g35_pad ,
		_w2038_
	);
	LUT4 #(
		.INIT('h0200)
	) name1264 (
		\g1146_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		_w2039_
	);
	LUT2 #(
		.INIT('h8)
	) name1265 (
		\g1152_reg/NET0131 ,
		\g35_pad ,
		_w2040_
	);
	LUT4 #(
		.INIT('hfdfc)
	) name1266 (
		_w1099_,
		_w2038_,
		_w2039_,
		_w2040_,
		_w2041_
	);
	LUT3 #(
		.INIT('hca)
	) name1267 (
		\g1211_reg/NET0131 ,
		\g29215_pad ,
		\g35_pad ,
		_w2042_
	);
	LUT4 #(
		.INIT('h10ff)
	) name1268 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g13259_pad ,
		\g35_pad ,
		_w2043_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2044_
	);
	LUT4 #(
		.INIT('h4440)
	) name1270 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2045_
	);
	LUT4 #(
		.INIT('h0002)
	) name1271 (
		\g2735_reg/NET0131 ,
		\g2741_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w2046_
	);
	LUT3 #(
		.INIT('h04)
	) name1272 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		_w2047_
	);
	LUT3 #(
		.INIT('h15)
	) name1273 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		\g1862_reg/NET0131 ,
		\g1906_reg/NET0131 ,
		_w2049_
	);
	LUT3 #(
		.INIT('h20)
	) name1275 (
		\g1917_reg/NET0131 ,
		\g1926_reg/NET0131 ,
		\g35_pad ,
		_w2050_
	);
	LUT3 #(
		.INIT('hca)
	) name1276 (
		\g1882_reg/NET0131 ,
		\g1902_reg/NET0131 ,
		\g35_pad ,
		_w2051_
	);
	LUT4 #(
		.INIT('hbf10)
	) name1277 (
		_w2048_,
		_w2049_,
		_w2050_,
		_w2051_,
		_w2052_
	);
	LUT2 #(
		.INIT('h8)
	) name1278 (
		\g376_reg/NET0131 ,
		\g8719_pad ,
		_w2053_
	);
	LUT4 #(
		.INIT('h8000)
	) name1279 (
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		\g8719_pad ,
		\g896_reg/NET0131 ,
		_w2054_
	);
	LUT4 #(
		.INIT('h0800)
	) name1280 (
		\g370_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		\g8719_pad ,
		_w2055_
	);
	LUT3 #(
		.INIT('h1d)
	) name1281 (
		\g174_reg/NET0131 ,
		\g392_reg/NET0131 ,
		\g452_reg/NET0131 ,
		_w2056_
	);
	LUT2 #(
		.INIT('h4)
	) name1282 (
		\g392_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w2057_
	);
	LUT4 #(
		.INIT('h0013)
	) name1283 (
		\g392_reg/NET0131 ,
		\g417_reg/NET0131 ,
		\g441_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w2058_
	);
	LUT4 #(
		.INIT('h0900)
	) name1284 (
		\g182_reg/NET0131 ,
		_w2056_,
		_w2057_,
		_w2058_,
		_w2059_
	);
	LUT3 #(
		.INIT('h06)
	) name1285 (
		\g392_reg/NET0131 ,
		\g405_reg/NET0131 ,
		\g437_reg/NET0131 ,
		_w2060_
	);
	LUT4 #(
		.INIT('h2025)
	) name1286 (
		\g392_reg/NET0131 ,
		\g401_reg/NET0131 ,
		\g405_reg/NET0131 ,
		\g424_reg/NET0131 ,
		_w2061_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name1287 (
		\g417_reg/NET0131 ,
		_w2055_,
		_w2060_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		\g703_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w2063_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1289 (
		_w2055_,
		_w2059_,
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h8)
	) name1290 (
		\g35_pad ,
		\g862_reg/NET0131 ,
		_w2065_
	);
	LUT4 #(
		.INIT('h1bbb)
	) name1291 (
		\g35_pad ,
		\g446_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w2066_
	);
	LUT4 #(
		.INIT('h10ff)
	) name1292 (
		_w2054_,
		_w2064_,
		_w2065_,
		_w2066_,
		_w2067_
	);
	LUT4 #(
		.INIT('h1110)
	) name1293 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2068_
	);
	LUT3 #(
		.INIT('h01)
	) name1294 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2803_reg/NET0131 ,
		_w2069_
	);
	LUT3 #(
		.INIT('h13)
	) name1295 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h4)
	) name1296 (
		\g2153_reg/NET0131 ,
		\g2197_reg/NET0131 ,
		_w2071_
	);
	LUT3 #(
		.INIT('h20)
	) name1297 (
		\g2208_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		\g35_pad ,
		_w2072_
	);
	LUT3 #(
		.INIT('hca)
	) name1298 (
		\g2173_reg/NET0131 ,
		\g2193_reg/NET0131 ,
		\g35_pad ,
		_w2073_
	);
	LUT4 #(
		.INIT('hbf10)
	) name1299 (
		_w2070_,
		_w2071_,
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT3 #(
		.INIT('h02)
	) name1300 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2807_reg/NET0131 ,
		_w2075_
	);
	LUT4 #(
		.INIT('h2220)
	) name1301 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2076_
	);
	LUT3 #(
		.INIT('h07)
	) name1302 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		\g2287_reg/NET0131 ,
		\g2331_reg/NET0131 ,
		_w2078_
	);
	LUT3 #(
		.INIT('h20)
	) name1304 (
		\g2342_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		\g35_pad ,
		_w2079_
	);
	LUT2 #(
		.INIT('h4)
	) name1305 (
		_w2078_,
		_w2079_,
		_w2080_
	);
	LUT3 #(
		.INIT('hca)
	) name1306 (
		\g2307_reg/NET0131 ,
		\g2327_reg/NET0131 ,
		\g35_pad ,
		_w2081_
	);
	LUT2 #(
		.INIT('h4)
	) name1307 (
		_w2079_,
		_w2081_,
		_w2082_
	);
	LUT4 #(
		.INIT('h0700)
	) name1308 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2081_,
		_w2083_
	);
	LUT4 #(
		.INIT('hfff4)
	) name1309 (
		_w2077_,
		_w2080_,
		_w2082_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h2)
	) name1310 (
		\g35_pad ,
		\g4646_reg/NET0131 ,
		_w2085_
	);
	LUT4 #(
		.INIT('h0008)
	) name1311 (
		\g35_pad ,
		\g4698_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w2086_
	);
	LUT4 #(
		.INIT('h070f)
	) name1312 (
		_w824_,
		_w825_,
		_w2085_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		\g4704_reg/NET0131 ,
		_w2087_,
		_w2088_
	);
	LUT2 #(
		.INIT('h8)
	) name1314 (
		\g35_pad ,
		\g4646_reg/NET0131 ,
		_w2089_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1315 (
		_w823_,
		_w824_,
		_w825_,
		_w2089_,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		_w864_,
		_w1945_,
		_w2091_
	);
	LUT3 #(
		.INIT('h35)
	) name1317 (
		\g3343_reg/NET0131 ,
		\g3347_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w2092_
	);
	LUT3 #(
		.INIT('hbe)
	) name1318 (
		\g4704_reg/NET0131 ,
		\g5297_reg/NET0131 ,
		_w2092_,
		_w2093_
	);
	LUT3 #(
		.INIT('h80)
	) name1319 (
		_w2090_,
		_w2091_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('he)
	) name1320 (
		_w2088_,
		_w2094_,
		_w2095_
	);
	LUT3 #(
		.INIT('h04)
	) name1321 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2815_reg/NET0131 ,
		_w2096_
	);
	LUT3 #(
		.INIT('h15)
	) name1322 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h4)
	) name1323 (
		\g2421_reg/NET0131 ,
		\g2465_reg/NET0131 ,
		_w2098_
	);
	LUT3 #(
		.INIT('h20)
	) name1324 (
		\g2476_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		\g35_pad ,
		_w2099_
	);
	LUT3 #(
		.INIT('hca)
	) name1325 (
		\g2441_reg/NET0131 ,
		\g2461_reg/NET0131 ,
		\g35_pad ,
		_w2100_
	);
	LUT4 #(
		.INIT('hbf10)
	) name1326 (
		_w2097_,
		_w2098_,
		_w2099_,
		_w2100_,
		_w2101_
	);
	LUT3 #(
		.INIT('h01)
	) name1327 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2771_reg/NET0131 ,
		_w2102_
	);
	LUT4 #(
		.INIT('h00b0)
	) name1328 (
		\g1592_reg/NET0131 ,
		\g1636_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		_w2103_
	);
	LUT4 #(
		.INIT('hec00)
	) name1329 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2103_,
		_w2104_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1330 (
		_w810_,
		_w2046_,
		_w2068_,
		_w2102_,
		_w2105_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1331 (
		\g1632_reg/NET0131 ,
		\g35_pad ,
		_w2104_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h2)
	) name1332 (
		\g1612_reg/NET0131 ,
		\g35_pad ,
		_w2107_
	);
	LUT2 #(
		.INIT('hd)
	) name1333 (
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h2)
	) name1334 (
		\g146_reg/NET0131 ,
		\g35_pad ,
		_w2109_
	);
	LUT2 #(
		.INIT('h6)
	) name1335 (
		\g164_reg/NET0131 ,
		_w1695_,
		_w2110_
	);
	LUT4 #(
		.INIT('h7000)
	) name1336 (
		_w1692_,
		_w1693_,
		_w1882_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('he)
	) name1337 (
		_w2109_,
		_w2111_,
		_w2112_
	);
	LUT2 #(
		.INIT('h2)
	) name1338 (
		\g744_reg/NET0131 ,
		\g758_reg/NET0131 ,
		_w2113_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1339 (
		\g35_pad ,
		_w893_,
		_w1958_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		\g744_reg/NET0131 ,
		\g749_reg/NET0131 ,
		_w2115_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1341 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g758_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w2116_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1342 (
		_w893_,
		_w1958_,
		_w2115_,
		_w2116_,
		_w2117_
	);
	LUT3 #(
		.INIT('hf2)
	) name1343 (
		\g749_reg/NET0131 ,
		_w2114_,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h4)
	) name1344 (
		\g35_pad ,
		\g832_reg/NET0131 ,
		_w2119_
	);
	LUT4 #(
		.INIT('h6a00)
	) name1345 (
		\g822_reg/NET0131 ,
		_w1824_,
		_w1825_,
		_w1829_,
		_w2120_
	);
	LUT2 #(
		.INIT('he)
	) name1346 (
		_w2119_,
		_w2120_,
		_w2121_
	);
	LUT4 #(
		.INIT('h0002)
	) name1347 (
		\g35_pad ,
		\g4392_reg/NET0131 ,
		\g4438_reg/NET0131 ,
		\g4443_reg/NET0131 ,
		_w2122_
	);
	LUT4 #(
		.INIT('heccc)
	) name1348 (
		\g4430_reg/NET0131 ,
		\g4452_reg/NET0131 ,
		_w1781_,
		_w2122_,
		_w2123_
	);
	LUT4 #(
		.INIT('h8880)
	) name1349 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2124_
	);
	LUT3 #(
		.INIT('h08)
	) name1350 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2819_reg/NET0131 ,
		_w2125_
	);
	LUT2 #(
		.INIT('h4)
	) name1351 (
		\g2587_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		_w2126_
	);
	LUT4 #(
		.INIT('h0440)
	) name1352 (
		\g2587_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		\g2648_reg/NET0131 ,
		\g2652_reg/NET0131 ,
		_w2127_
	);
	LUT4 #(
		.INIT('hec00)
	) name1353 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2127_,
		_w2128_
	);
	LUT4 #(
		.INIT('hec00)
	) name1354 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2126_,
		_w2129_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1355 (
		\g2657_reg/NET0131 ,
		\g35_pad ,
		_w2128_,
		_w2129_,
		_w2130_
	);
	LUT2 #(
		.INIT('h2)
	) name1356 (
		\g2652_reg/NET0131 ,
		\g35_pad ,
		_w2131_
	);
	LUT2 #(
		.INIT('hd)
	) name1357 (
		_w2130_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		\g2587_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		_w2133_
	);
	LUT4 #(
		.INIT('hec00)
	) name1359 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2133_,
		_w2134_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1360 (
		\g2657_reg/NET0131 ,
		\g2661_reg/NET0131 ,
		\g35_pad ,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h4)
	) name1361 (
		\g1624_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w2136_
	);
	LUT4 #(
		.INIT('h0440)
	) name1362 (
		\g1624_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		\g1687_reg/NET0131 ,
		\g1691_reg/NET0131 ,
		_w2137_
	);
	LUT4 #(
		.INIT('hec00)
	) name1363 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2137_,
		_w2138_
	);
	LUT4 #(
		.INIT('hec00)
	) name1364 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2136_,
		_w2139_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1365 (
		\g1696_reg/NET0131 ,
		\g35_pad ,
		_w2138_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h2)
	) name1366 (
		\g1691_reg/NET0131 ,
		\g35_pad ,
		_w2141_
	);
	LUT2 #(
		.INIT('hd)
	) name1367 (
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT2 #(
		.INIT('hd)
	) name1368 (
		\g35_pad ,
		_w2134_,
		_w2143_
	);
	LUT3 #(
		.INIT('h80)
	) name1369 (
		\g2587_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		\g2675_reg/NET0131 ,
		_w2144_
	);
	LUT4 #(
		.INIT('hec00)
	) name1370 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2144_,
		_w2145_
	);
	LUT3 #(
		.INIT('h51)
	) name1371 (
		\g2681_reg/NET0131 ,
		\g35_pad ,
		_w2145_,
		_w2146_
	);
	LUT4 #(
		.INIT('h0800)
	) name1372 (
		\g2587_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		\g2675_reg/NET0131 ,
		\g2681_reg/NET0131 ,
		_w2147_
	);
	LUT4 #(
		.INIT('hec00)
	) name1373 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2147_,
		_w2148_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1374 (
		\g2685_reg/NET0131 ,
		\g35_pad ,
		_w2134_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		_w2146_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h8)
	) name1376 (
		\g1624_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		_w2151_
	);
	LUT4 #(
		.INIT('hec00)
	) name1377 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2151_,
		_w2152_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1378 (
		\g1696_reg/NET0131 ,
		\g1700_reg/NET0131 ,
		\g35_pad ,
		_w2152_,
		_w2153_
	);
	LUT3 #(
		.INIT('h80)
	) name1379 (
		\g1624_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		\g1714_reg/NET0131 ,
		_w2154_
	);
	LUT4 #(
		.INIT('hec00)
	) name1380 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2154_,
		_w2155_
	);
	LUT3 #(
		.INIT('h51)
	) name1381 (
		\g1720_reg/NET0131 ,
		\g35_pad ,
		_w2155_,
		_w2156_
	);
	LUT4 #(
		.INIT('h0800)
	) name1382 (
		\g1624_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		\g1714_reg/NET0131 ,
		\g1720_reg/NET0131 ,
		_w2157_
	);
	LUT4 #(
		.INIT('hec00)
	) name1383 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2157_,
		_w2158_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1384 (
		\g1724_reg/NET0131 ,
		\g35_pad ,
		_w2152_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h4)
	) name1385 (
		_w2156_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('hd)
	) name1386 (
		\g35_pad ,
		_w2152_,
		_w2161_
	);
	LUT3 #(
		.INIT('h02)
	) name1387 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		_w2162_
	);
	LUT3 #(
		.INIT('h13)
	) name1388 (
		_w2046_,
		_w2076_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1389 (
		\g1792_reg/NET0131 ,
		_w2046_,
		_w2076_,
		_w2162_,
		_w2164_
	);
	LUT2 #(
		.INIT('h4)
	) name1390 (
		\g1760_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w2165_
	);
	LUT4 #(
		.INIT('h0105)
	) name1391 (
		\g1760_reg/NET0131 ,
		_w2046_,
		_w2076_,
		_w2162_,
		_w2166_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1392 (
		\g35_pad ,
		_w2164_,
		_w2165_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		\g1768_reg/NET0131 ,
		\g35_pad ,
		_w2168_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('h0440)
	) name1395 (
		\g1760_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		\g1821_reg/NET0131 ,
		\g1825_reg/NET0131 ,
		_w2170_
	);
	LUT4 #(
		.INIT('hec00)
	) name1396 (
		_w2046_,
		_w2076_,
		_w2162_,
		_w2170_,
		_w2171_
	);
	LUT4 #(
		.INIT('hec00)
	) name1397 (
		_w2046_,
		_w2076_,
		_w2162_,
		_w2165_,
		_w2172_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1398 (
		\g1830_reg/NET0131 ,
		\g35_pad ,
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h2)
	) name1399 (
		\g1825_reg/NET0131 ,
		\g35_pad ,
		_w2174_
	);
	LUT2 #(
		.INIT('hd)
	) name1400 (
		_w2173_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name1401 (
		\g1760_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		_w2176_
	);
	LUT4 #(
		.INIT('hec00)
	) name1402 (
		_w2046_,
		_w2076_,
		_w2162_,
		_w2176_,
		_w2177_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1403 (
		\g1830_reg/NET0131 ,
		\g1834_reg/NET0131 ,
		\g35_pad ,
		_w2177_,
		_w2178_
	);
	LUT3 #(
		.INIT('h80)
	) name1404 (
		\g1760_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		\g1848_reg/NET0131 ,
		_w2179_
	);
	LUT4 #(
		.INIT('hec00)
	) name1405 (
		_w2046_,
		_w2076_,
		_w2162_,
		_w2179_,
		_w2180_
	);
	LUT3 #(
		.INIT('h51)
	) name1406 (
		\g1854_reg/NET0131 ,
		\g35_pad ,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h0800)
	) name1407 (
		\g1760_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		\g1848_reg/NET0131 ,
		\g1854_reg/NET0131 ,
		_w2182_
	);
	LUT4 #(
		.INIT('hec00)
	) name1408 (
		_w2046_,
		_w2076_,
		_w2162_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1409 (
		\g1858_reg/NET0131 ,
		\g35_pad ,
		_w2177_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h4)
	) name1410 (
		_w2181_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('hd)
	) name1411 (
		\g35_pad ,
		_w2177_,
		_w2186_
	);
	LUT4 #(
		.INIT('ha888)
	) name1412 (
		\g1926_reg/NET0131 ,
		_w2045_,
		_w2046_,
		_w2047_,
		_w2187_
	);
	LUT4 #(
		.INIT('h5444)
	) name1413 (
		\g1917_reg/NET0131 ,
		_w2045_,
		_w2046_,
		_w2047_,
		_w2188_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1414 (
		\g1894_reg/NET0131 ,
		\g35_pad ,
		_w2187_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		\g1902_reg/NET0131 ,
		\g35_pad ,
		_w2190_
	);
	LUT2 #(
		.INIT('h2)
	) name1416 (
		_w2189_,
		_w2190_,
		_w2191_
	);
	LUT2 #(
		.INIT('h4)
	) name1417 (
		\g1894_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w2192_
	);
	LUT4 #(
		.INIT('h0440)
	) name1418 (
		\g1894_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		\g1955_reg/NET0131 ,
		\g1959_reg/NET0131 ,
		_w2193_
	);
	LUT4 #(
		.INIT('hea00)
	) name1419 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2193_,
		_w2194_
	);
	LUT4 #(
		.INIT('hea00)
	) name1420 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2192_,
		_w2195_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1421 (
		\g1964_reg/NET0131 ,
		\g35_pad ,
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		\g1959_reg/NET0131 ,
		\g35_pad ,
		_w2197_
	);
	LUT2 #(
		.INIT('hd)
	) name1423 (
		_w2196_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h8)
	) name1424 (
		\g1894_reg/NET0131 ,
		\g1926_reg/NET0131 ,
		_w2199_
	);
	LUT4 #(
		.INIT('hea00)
	) name1425 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2199_,
		_w2200_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1426 (
		\g1964_reg/NET0131 ,
		\g1968_reg/NET0131 ,
		\g35_pad ,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('hd)
	) name1427 (
		\g35_pad ,
		_w2200_,
		_w2202_
	);
	LUT3 #(
		.INIT('h80)
	) name1428 (
		\g1894_reg/NET0131 ,
		\g1926_reg/NET0131 ,
		\g1982_reg/NET0131 ,
		_w2203_
	);
	LUT4 #(
		.INIT('hea00)
	) name1429 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('h51)
	) name1430 (
		\g1988_reg/NET0131 ,
		\g35_pad ,
		_w2204_,
		_w2205_
	);
	LUT4 #(
		.INIT('h0800)
	) name1431 (
		\g1894_reg/NET0131 ,
		\g1926_reg/NET0131 ,
		\g1982_reg/NET0131 ,
		\g1988_reg/NET0131 ,
		_w2206_
	);
	LUT4 #(
		.INIT('hea00)
	) name1432 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1433 (
		\g1992_reg/NET0131 ,
		\g35_pad ,
		_w2200_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h4)
	) name1434 (
		_w2205_,
		_w2208_,
		_w2209_
	);
	LUT3 #(
		.INIT('h08)
	) name1435 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		_w2210_
	);
	LUT2 #(
		.INIT('h4)
	) name1436 (
		\g2028_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w2211_
	);
	LUT4 #(
		.INIT('h0440)
	) name1437 (
		\g2028_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		\g2089_reg/NET0131 ,
		\g2093_reg/NET0131 ,
		_w2212_
	);
	LUT4 #(
		.INIT('hec00)
	) name1438 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2212_,
		_w2213_
	);
	LUT4 #(
		.INIT('hec00)
	) name1439 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2211_,
		_w2214_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1440 (
		\g2098_reg/NET0131 ,
		\g35_pad ,
		_w2213_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		\g2093_reg/NET0131 ,
		\g35_pad ,
		_w2216_
	);
	LUT2 #(
		.INIT('hd)
	) name1442 (
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name1443 (
		\g2028_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		_w2218_
	);
	LUT4 #(
		.INIT('hec00)
	) name1444 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2218_,
		_w2219_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1445 (
		\g2098_reg/NET0131 ,
		\g2102_reg/NET0131 ,
		\g35_pad ,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('hd)
	) name1446 (
		\g35_pad ,
		_w2219_,
		_w2221_
	);
	LUT3 #(
		.INIT('h80)
	) name1447 (
		\g2028_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		\g2116_reg/NET0131 ,
		_w2222_
	);
	LUT4 #(
		.INIT('hec00)
	) name1448 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2222_,
		_w2223_
	);
	LUT3 #(
		.INIT('h51)
	) name1449 (
		\g2122_reg/NET0131 ,
		\g35_pad ,
		_w2223_,
		_w2224_
	);
	LUT4 #(
		.INIT('h0800)
	) name1450 (
		\g2028_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		\g2116_reg/NET0131 ,
		\g2122_reg/NET0131 ,
		_w2225_
	);
	LUT4 #(
		.INIT('hec00)
	) name1451 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2225_,
		_w2226_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1452 (
		\g2126_reg/NET0131 ,
		\g35_pad ,
		_w2219_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		_w2224_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h4)
	) name1454 (
		\g2185_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		_w2229_
	);
	LUT4 #(
		.INIT('h0440)
	) name1455 (
		\g2185_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		\g2246_reg/NET0131 ,
		\g2250_reg/NET0131 ,
		_w2230_
	);
	LUT4 #(
		.INIT('hec00)
	) name1456 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2230_,
		_w2231_
	);
	LUT4 #(
		.INIT('hec00)
	) name1457 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2229_,
		_w2232_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1458 (
		\g2255_reg/NET0131 ,
		\g35_pad ,
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h2)
	) name1459 (
		\g2250_reg/NET0131 ,
		\g35_pad ,
		_w2234_
	);
	LUT2 #(
		.INIT('hd)
	) name1460 (
		_w2233_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		\g2185_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		_w2236_
	);
	LUT4 #(
		.INIT('hec00)
	) name1462 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2236_,
		_w2237_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1463 (
		\g2255_reg/NET0131 ,
		\g2259_reg/NET0131 ,
		\g35_pad ,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('hd)
	) name1464 (
		\g35_pad ,
		_w2237_,
		_w2239_
	);
	LUT3 #(
		.INIT('h80)
	) name1465 (
		\g2185_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		\g2273_reg/NET0131 ,
		_w2240_
	);
	LUT4 #(
		.INIT('hec00)
	) name1466 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2240_,
		_w2241_
	);
	LUT3 #(
		.INIT('h51)
	) name1467 (
		\g2279_reg/NET0131 ,
		\g35_pad ,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h0800)
	) name1468 (
		\g2185_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		\g2273_reg/NET0131 ,
		\g2279_reg/NET0131 ,
		_w2243_
	);
	LUT4 #(
		.INIT('hec00)
	) name1469 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2243_,
		_w2244_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1470 (
		\g2283_reg/NET0131 ,
		\g35_pad ,
		_w2237_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h4)
	) name1471 (
		_w2242_,
		_w2245_,
		_w2246_
	);
	LUT4 #(
		.INIT('haa80)
	) name1472 (
		\g2351_reg/NET0131 ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2247_
	);
	LUT2 #(
		.INIT('h4)
	) name1473 (
		\g2319_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		_w2248_
	);
	LUT4 #(
		.INIT('h0015)
	) name1474 (
		\g2319_reg/NET0131 ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2249_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1475 (
		\g35_pad ,
		_w2247_,
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT2 #(
		.INIT('h1)
	) name1476 (
		\g2327_reg/NET0131 ,
		\g35_pad ,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		_w2250_,
		_w2251_,
		_w2252_
	);
	LUT4 #(
		.INIT('h0440)
	) name1478 (
		\g2319_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		\g2380_reg/NET0131 ,
		\g2384_reg/NET0131 ,
		_w2253_
	);
	LUT4 #(
		.INIT('hf800)
	) name1479 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2253_,
		_w2254_
	);
	LUT3 #(
		.INIT('hb0)
	) name1480 (
		\g2319_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		\g2389_reg/NET0131 ,
		_w2255_
	);
	LUT4 #(
		.INIT('h002a)
	) name1481 (
		\g2389_reg/NET0131 ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2256_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1482 (
		\g35_pad ,
		_w2254_,
		_w2255_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h2)
	) name1483 (
		\g2384_reg/NET0131 ,
		\g35_pad ,
		_w2258_
	);
	LUT2 #(
		.INIT('he)
	) name1484 (
		_w2257_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h8)
	) name1485 (
		\g2319_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		_w2260_
	);
	LUT4 #(
		.INIT('hf800)
	) name1486 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2260_,
		_w2261_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1487 (
		\g2389_reg/NET0131 ,
		\g2393_reg/NET0131 ,
		\g35_pad ,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('hd)
	) name1488 (
		\g35_pad ,
		_w2261_,
		_w2263_
	);
	LUT3 #(
		.INIT('h80)
	) name1489 (
		\g2319_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		\g2407_reg/NET0131 ,
		_w2264_
	);
	LUT4 #(
		.INIT('hf800)
	) name1490 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2264_,
		_w2265_
	);
	LUT3 #(
		.INIT('h51)
	) name1491 (
		\g2413_reg/NET0131 ,
		\g35_pad ,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h0800)
	) name1492 (
		\g2319_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		\g2407_reg/NET0131 ,
		\g2413_reg/NET0131 ,
		_w2267_
	);
	LUT4 #(
		.INIT('hf800)
	) name1493 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2267_,
		_w2268_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1494 (
		\g2417_reg/NET0131 ,
		\g35_pad ,
		_w2261_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h4)
	) name1495 (
		_w2266_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('ha888)
	) name1496 (
		\g2485_reg/NET0131 ,
		_w2045_,
		_w2046_,
		_w2096_,
		_w2271_
	);
	LUT4 #(
		.INIT('h5444)
	) name1497 (
		\g2476_reg/NET0131 ,
		_w2045_,
		_w2046_,
		_w2096_,
		_w2272_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1498 (
		\g2453_reg/NET0131 ,
		\g35_pad ,
		_w2271_,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name1499 (
		\g2461_reg/NET0131 ,
		\g35_pad ,
		_w2274_
	);
	LUT2 #(
		.INIT('h2)
	) name1500 (
		_w2273_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h4)
	) name1501 (
		\g2453_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		_w2276_
	);
	LUT4 #(
		.INIT('h0440)
	) name1502 (
		\g2453_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		\g2514_reg/NET0131 ,
		\g2518_reg/NET0131 ,
		_w2277_
	);
	LUT4 #(
		.INIT('hea00)
	) name1503 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2277_,
		_w2278_
	);
	LUT4 #(
		.INIT('hea00)
	) name1504 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2276_,
		_w2279_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1505 (
		\g2523_reg/NET0131 ,
		\g35_pad ,
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT2 #(
		.INIT('h2)
	) name1506 (
		\g2518_reg/NET0131 ,
		\g35_pad ,
		_w2281_
	);
	LUT2 #(
		.INIT('hd)
	) name1507 (
		_w2280_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		\g2453_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		_w2283_
	);
	LUT4 #(
		.INIT('hea00)
	) name1509 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('h3aca)
	) name1510 (
		\g2523_reg/NET0131 ,
		\g2527_reg/NET0131 ,
		\g35_pad ,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('hd)
	) name1511 (
		\g35_pad ,
		_w2284_,
		_w2286_
	);
	LUT3 #(
		.INIT('h80)
	) name1512 (
		\g2453_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		\g2541_reg/NET0131 ,
		_w2287_
	);
	LUT4 #(
		.INIT('hea00)
	) name1513 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2287_,
		_w2288_
	);
	LUT3 #(
		.INIT('h51)
	) name1514 (
		\g2547_reg/NET0131 ,
		\g35_pad ,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('h0800)
	) name1515 (
		\g2453_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		\g2541_reg/NET0131 ,
		\g2547_reg/NET0131 ,
		_w2290_
	);
	LUT4 #(
		.INIT('hea00)
	) name1516 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('h33fb)
	) name1517 (
		\g2551_reg/NET0131 ,
		\g35_pad ,
		_w2284_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h4)
	) name1518 (
		_w2289_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1519 (
		\g2060_reg/NET0131 ,
		_w2046_,
		_w2124_,
		_w2210_,
		_w2294_
	);
	LUT4 #(
		.INIT('h5450)
	) name1520 (
		\g2051_reg/NET0131 ,
		_w2046_,
		_w2124_,
		_w2210_,
		_w2295_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1521 (
		\g2028_reg/NET0131 ,
		\g35_pad ,
		_w2294_,
		_w2295_,
		_w2296_
	);
	LUT2 #(
		.INIT('h1)
	) name1522 (
		\g2036_reg/NET0131 ,
		\g35_pad ,
		_w2297_
	);
	LUT2 #(
		.INIT('h2)
	) name1523 (
		_w2296_,
		_w2297_,
		_w2298_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1524 (
		\g2217_reg/NET0131 ,
		_w2046_,
		_w2068_,
		_w2069_,
		_w2299_
	);
	LUT4 #(
		.INIT('h5450)
	) name1525 (
		\g2208_reg/NET0131 ,
		_w2046_,
		_w2068_,
		_w2069_,
		_w2300_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1526 (
		\g2185_reg/NET0131 ,
		\g35_pad ,
		_w2299_,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1527 (
		\g2193_reg/NET0131 ,
		\g35_pad ,
		_w2302_
	);
	LUT2 #(
		.INIT('h2)
	) name1528 (
		_w2301_,
		_w2302_,
		_w2303_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1529 (
		\g1657_reg/NET0131 ,
		_w2046_,
		_w2068_,
		_w2102_,
		_w2304_
	);
	LUT4 #(
		.INIT('h5450)
	) name1530 (
		\g1648_reg/NET0131 ,
		_w2046_,
		_w2068_,
		_w2102_,
		_w2305_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1531 (
		\g1624_reg/NET0131 ,
		\g35_pad ,
		_w2304_,
		_w2305_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		\g1632_reg/NET0131 ,
		\g35_pad ,
		_w2307_
	);
	LUT2 #(
		.INIT('h2)
	) name1533 (
		_w2306_,
		_w2307_,
		_w2308_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1534 (
		\g2619_reg/NET0131 ,
		_w2046_,
		_w2124_,
		_w2125_,
		_w2309_
	);
	LUT4 #(
		.INIT('h5450)
	) name1535 (
		\g2610_reg/NET0131 ,
		_w2046_,
		_w2124_,
		_w2125_,
		_w2310_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1536 (
		\g2587_reg/NET0131 ,
		\g35_pad ,
		_w2309_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h1)
	) name1537 (
		\g2595_reg/NET0131 ,
		\g35_pad ,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		_w2311_,
		_w2312_,
		_w2313_
	);
	LUT3 #(
		.INIT('hd0)
	) name1539 (
		\g35_pad ,
		\g4382_reg/NET0131 ,
		\g4438_reg/NET0131 ,
		_w2314_
	);
	LUT4 #(
		.INIT('h0008)
	) name1540 (
		\g35_pad ,
		\g4392_reg/NET0131 ,
		\g4438_reg/NET0131 ,
		\g4443_reg/NET0131 ,
		_w2315_
	);
	LUT3 #(
		.INIT('hec)
	) name1541 (
		_w1781_,
		_w2314_,
		_w2315_,
		_w2316_
	);
	LUT3 #(
		.INIT('hc4)
	) name1542 (
		\g35_pad ,
		\g5080_reg/NET0131 ,
		\g5084_reg/NET0131 ,
		_w2317_
	);
	LUT2 #(
		.INIT('h4)
	) name1543 (
		\g5073_reg/NET0131 ,
		\g5077_reg/NET0131 ,
		_w2318_
	);
	LUT4 #(
		.INIT('h000b)
	) name1544 (
		\g5069_reg/NET0131 ,
		\g5077_reg/NET0131 ,
		\g5080_reg/NET0131 ,
		\g5084_reg/NET0131 ,
		_w2319_
	);
	LUT4 #(
		.INIT('heeec)
	) name1545 (
		\g35_pad ,
		_w2317_,
		_w2318_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name1546 (
		\g2831_reg/NET0131 ,
		\g35_pad ,
		_w2321_
	);
	LUT4 #(
		.INIT('hc840)
	) name1547 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		_w2322_
	);
	LUT4 #(
		.INIT('h3210)
	) name1548 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2771_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		_w2323_
	);
	LUT2 #(
		.INIT('h1)
	) name1549 (
		_w2322_,
		_w2323_,
		_w2324_
	);
	LUT3 #(
		.INIT('h01)
	) name1550 (
		\g2741_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w2325_
	);
	LUT3 #(
		.INIT('h01)
	) name1551 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2735_reg/NET0131 ,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name1552 (
		_w2325_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('h3500)
	) name1553 (
		\g1945_reg/NET0131 ,
		\g2079_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2328_
	);
	LUT4 #(
		.INIT('h0035)
	) name1554 (
		\g1677_reg/NET0131 ,
		\g1811_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2329_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		_w2328_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('h757f)
	) name1556 (
		\g35_pad ,
		_w2324_,
		_w2327_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('hb)
	) name1557 (
		_w2321_,
		_w2331_,
		_w2332_
	);
	LUT3 #(
		.INIT('h6a)
	) name1558 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		\g35_pad ,
		_w2333_
	);
	LUT3 #(
		.INIT('hd0)
	) name1559 (
		\g35_pad ,
		_w1715_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h4)
	) name1560 (
		\g1792_reg/NET0131 ,
		\g35_pad ,
		_w2335_
	);
	LUT3 #(
		.INIT('hb0)
	) name1561 (
		\g1728_reg/NET0131 ,
		\g1772_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w2336_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		_w2335_,
		_w2336_,
		_w2337_
	);
	LUT3 #(
		.INIT('h20)
	) name1563 (
		\g1783_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		\g35_pad ,
		_w2338_
	);
	LUT3 #(
		.INIT('hca)
	) name1564 (
		\g1748_reg/NET0131 ,
		\g1768_reg/NET0131 ,
		\g35_pad ,
		_w2339_
	);
	LUT4 #(
		.INIT('hef44)
	) name1565 (
		_w2163_,
		_w2337_,
		_w2338_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h4)
	) name1566 (
		\g35_pad ,
		\g744_reg/NET0131 ,
		_w2341_
	);
	LUT2 #(
		.INIT('h2)
	) name1567 (
		\g744_reg/NET0131 ,
		\g749_reg/NET0131 ,
		_w2342_
	);
	LUT4 #(
		.INIT('h070f)
	) name1568 (
		_w893_,
		_w1958_,
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1569 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g749_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w2344_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1570 (
		\g744_reg/NET0131 ,
		_w893_,
		_w1958_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('hd)
	) name1571 (
		_w2343_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h2)
	) name1572 (
		\g2051_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		_w2347_
	);
	LUT4 #(
		.INIT('h0040)
	) name1573 (
		\g1996_reg/NET0131 ,
		\g2040_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		_w2348_
	);
	LUT4 #(
		.INIT('hec00)
	) name1574 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2348_,
		_w2349_
	);
	LUT4 #(
		.INIT('hec00)
	) name1575 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2347_,
		_w2350_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1576 (
		\g2036_reg/NET0131 ,
		\g35_pad ,
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h1)
	) name1577 (
		\g2016_reg/NET0131 ,
		\g35_pad ,
		_w2352_
	);
	LUT2 #(
		.INIT('h2)
	) name1578 (
		_w2351_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h2)
	) name1579 (
		\g2834_reg/NET0131 ,
		\g35_pad ,
		_w2354_
	);
	LUT4 #(
		.INIT('hc840)
	) name1580 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2815_reg/NET0131 ,
		\g2819_reg/NET0131 ,
		_w2355_
	);
	LUT4 #(
		.INIT('h3210)
	) name1581 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		\g2803_reg/NET0131 ,
		\g2807_reg/NET0131 ,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		_w2355_,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('h3500)
	) name1583 (
		\g2504_reg/NET0131 ,
		\g2638_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2358_
	);
	LUT4 #(
		.INIT('h0035)
	) name1584 (
		\g2236_reg/NET0131 ,
		\g2370_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2359_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		_w2358_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1586 (
		\g35_pad ,
		_w2327_,
		_w2357_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('hb)
	) name1587 (
		_w2354_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h2)
	) name1588 (
		\g2610_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		_w2363_
	);
	LUT4 #(
		.INIT('h0040)
	) name1589 (
		\g2555_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		_w2364_
	);
	LUT4 #(
		.INIT('hec00)
	) name1590 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2364_,
		_w2365_
	);
	LUT4 #(
		.INIT('hec00)
	) name1591 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2363_,
		_w2366_
	);
	LUT4 #(
		.INIT('h3f3b)
	) name1592 (
		\g2595_reg/NET0131 ,
		\g35_pad ,
		_w2365_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h1)
	) name1593 (
		\g2575_reg/NET0131 ,
		\g35_pad ,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name1594 (
		_w2367_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h2)
	) name1595 (
		\g142_reg/NET0131 ,
		\g35_pad ,
		_w2370_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name1596 (
		\g146_reg/NET0131 ,
		\g203_reg/NET0131 ,
		\g513_reg/NET0131 ,
		\g518_reg/NET0131 ,
		_w2371_
	);
	LUT4 #(
		.INIT('h7000)
	) name1597 (
		_w1692_,
		_w1693_,
		_w1882_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('he)
	) name1598 (
		_w2370_,
		_w2372_,
		_w2373_
	);
	LUT4 #(
		.INIT('h8adf)
	) name1599 (
		\g35_pad ,
		\g4382_reg/NET0131 ,
		\g4438_reg/NET0131 ,
		\g4443_reg/NET0131 ,
		_w2374_
	);
	LUT3 #(
		.INIT('h8f)
	) name1600 (
		_w1781_,
		_w2122_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		\g35_pad ,
		\g4801_reg/NET0131 ,
		_w2376_
	);
	LUT2 #(
		.INIT('h8)
	) name1602 (
		\g4776_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		_w2377_
	);
	LUT3 #(
		.INIT('h2a)
	) name1603 (
		\g35_pad ,
		_w1981_,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h8)
	) name1604 (
		\g4793_reg/NET0131 ,
		\g4801_reg/NET0131 ,
		_w2379_
	);
	LUT3 #(
		.INIT('h15)
	) name1605 (
		\g4776_reg/NET0131 ,
		_w1981_,
		_w2379_,
		_w2380_
	);
	LUT3 #(
		.INIT('hae)
	) name1606 (
		_w2376_,
		_w2378_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h4)
	) name1607 (
		\g35_pad ,
		\g671_reg/NET0131 ,
		_w2382_
	);
	LUT4 #(
		.INIT('h8000)
	) name1608 (
		\g671_reg/NET0131 ,
		_w1824_,
		_w2022_,
		_w2023_,
		_w2383_
	);
	LUT2 #(
		.INIT('h1)
	) name1609 (
		\g676_reg/NET0131 ,
		_w2383_,
		_w2384_
	);
	LUT4 #(
		.INIT('h0070)
	) name1610 (
		_w2024_,
		_w2028_,
		_w2029_,
		_w2032_,
		_w2385_
	);
	LUT3 #(
		.INIT('hba)
	) name1611 (
		_w2382_,
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h4)
	) name1612 (
		\g35_pad ,
		\g4659_reg/NET0131 ,
		_w2387_
	);
	LUT3 #(
		.INIT('hb1)
	) name1613 (
		\g35_pad ,
		\g4659_reg/NET0131 ,
		_w1981_,
		_w2388_
	);
	LUT3 #(
		.INIT('h80)
	) name1614 (
		\g4653_reg/NET0131 ,
		\g4659_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w2389_
	);
	LUT3 #(
		.INIT('hde)
	) name1615 (
		\g4664_reg/NET0131 ,
		_w2387_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		_w2388_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		\g1798_reg/NET0131 ,
		\g35_pad ,
		_w2392_
	);
	LUT4 #(
		.INIT('h0105)
	) name1618 (
		\g1792_reg/NET0131 ,
		_w2046_,
		_w2076_,
		_w2162_,
		_w2393_
	);
	LUT2 #(
		.INIT('h8)
	) name1619 (
		\g1783_reg/NET0131 ,
		\g35_pad ,
		_w2394_
	);
	LUT4 #(
		.INIT('h020a)
	) name1620 (
		\g35_pad ,
		_w2046_,
		_w2076_,
		_w2162_,
		_w2395_
	);
	LUT4 #(
		.INIT('hfdf5)
	) name1621 (
		\g35_pad ,
		_w2046_,
		_w2076_,
		_w2162_,
		_w2396_
	);
	LUT4 #(
		.INIT('hbbba)
	) name1622 (
		_w2392_,
		_w2393_,
		_w2394_,
		_w2395_,
		_w2397_
	);
	LUT4 #(
		.INIT('h020a)
	) name1623 (
		\g1811_reg/NET0131 ,
		_w2046_,
		_w2076_,
		_w2162_,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name1624 (
		\g35_pad ,
		_w2398_,
		_w2399_
	);
	LUT4 #(
		.INIT('h51f3)
	) name1625 (
		\g1740_reg/NET0131 ,
		\g1752_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name1626 (
		\g1760_reg/NET0131 ,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('h31f5)
	) name1627 (
		\g1748_reg/NET0131 ,
		\g1756_reg/NET0131 ,
		\g1760_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w2402_
	);
	LUT3 #(
		.INIT('h20)
	) name1628 (
		\g1736_reg/NET0131 ,
		\g1760_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w2403_
	);
	LUT2 #(
		.INIT('h2)
	) name1629 (
		\g1744_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w2404_
	);
	LUT4 #(
		.INIT('h040e)
	) name1630 (
		\g1792_reg/NET0131 ,
		_w2402_,
		_w2403_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1631 (
		\g35_pad ,
		_w2046_,
		_w2076_,
		_w2162_,
		_w2406_
	);
	LUT3 #(
		.INIT('hb0)
	) name1632 (
		_w2401_,
		_w2405_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		\g1792_reg/NET0131 ,
		\g35_pad ,
		_w2408_
	);
	LUT3 #(
		.INIT('hfe)
	) name1634 (
		_w2399_,
		_w2407_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('h0222)
	) name1635 (
		\g35_pad ,
		_w2045_,
		_w2046_,
		_w2047_,
		_w2410_
	);
	LUT4 #(
		.INIT('hfddd)
	) name1636 (
		\g35_pad ,
		_w2045_,
		_w2046_,
		_w2047_,
		_w2411_
	);
	LUT2 #(
		.INIT('h4)
	) name1637 (
		\g1926_reg/NET0131 ,
		\g35_pad ,
		_w2412_
	);
	LUT4 #(
		.INIT('h1500)
	) name1638 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h4)
	) name1639 (
		\g1917_reg/NET0131 ,
		\g35_pad ,
		_w2414_
	);
	LUT4 #(
		.INIT('hea00)
	) name1640 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		\g1932_reg/NET0131 ,
		\g35_pad ,
		_w2416_
	);
	LUT3 #(
		.INIT('h01)
	) name1642 (
		_w2413_,
		_w2415_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('h0222)
	) name1643 (
		\g1945_reg/NET0131 ,
		_w2045_,
		_w2046_,
		_w2047_,
		_w2418_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		\g35_pad ,
		_w2418_,
		_w2419_
	);
	LUT4 #(
		.INIT('h51f3)
	) name1645 (
		\g1874_reg/NET0131 ,
		\g1886_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		\g1926_reg/NET0131 ,
		_w2420_
	);
	LUT2 #(
		.INIT('h2)
	) name1646 (
		\g1894_reg/NET0131 ,
		_w2420_,
		_w2421_
	);
	LUT4 #(
		.INIT('h31f5)
	) name1647 (
		\g1882_reg/NET0131 ,
		\g1890_reg/NET0131 ,
		\g1894_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w2422_
	);
	LUT3 #(
		.INIT('h20)
	) name1648 (
		\g1870_reg/NET0131 ,
		\g1894_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name1649 (
		\g1878_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w2424_
	);
	LUT4 #(
		.INIT('h040e)
	) name1650 (
		\g1926_reg/NET0131 ,
		_w2422_,
		_w2423_,
		_w2424_,
		_w2425_
	);
	LUT4 #(
		.INIT('ha888)
	) name1651 (
		\g35_pad ,
		_w2045_,
		_w2046_,
		_w2047_,
		_w2426_
	);
	LUT3 #(
		.INIT('hb0)
	) name1652 (
		_w2421_,
		_w2425_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		\g1926_reg/NET0131 ,
		\g35_pad ,
		_w2428_
	);
	LUT3 #(
		.INIT('hfe)
	) name1654 (
		_w2419_,
		_w2427_,
		_w2428_,
		_w2429_
	);
	LUT4 #(
		.INIT('h020a)
	) name1655 (
		\g35_pad ,
		_w2046_,
		_w2124_,
		_w2210_,
		_w2430_
	);
	LUT4 #(
		.INIT('hfdf5)
	) name1656 (
		\g35_pad ,
		_w2046_,
		_w2124_,
		_w2210_,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name1657 (
		\g2066_reg/NET0131 ,
		\g35_pad ,
		_w2432_
	);
	LUT2 #(
		.INIT('h8)
	) name1658 (
		\g2060_reg/NET0131 ,
		\g35_pad ,
		_w2433_
	);
	LUT4 #(
		.INIT('h1300)
	) name1659 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		\g2051_reg/NET0131 ,
		\g35_pad ,
		_w2435_
	);
	LUT4 #(
		.INIT('hec00)
	) name1661 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('hfe)
	) name1662 (
		_w2432_,
		_w2434_,
		_w2436_,
		_w2437_
	);
	LUT4 #(
		.INIT('h020a)
	) name1663 (
		\g2079_reg/NET0131 ,
		_w2046_,
		_w2124_,
		_w2210_,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		\g35_pad ,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('h51f3)
	) name1665 (
		\g2008_reg/NET0131 ,
		\g2020_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		\g2028_reg/NET0131 ,
		_w2440_,
		_w2441_
	);
	LUT4 #(
		.INIT('h31f5)
	) name1667 (
		\g2016_reg/NET0131 ,
		\g2024_reg/NET0131 ,
		\g2028_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w2442_
	);
	LUT3 #(
		.INIT('h20)
	) name1668 (
		\g2004_reg/NET0131 ,
		\g2028_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w2443_
	);
	LUT2 #(
		.INIT('h2)
	) name1669 (
		\g2012_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w2444_
	);
	LUT4 #(
		.INIT('h040e)
	) name1670 (
		\g2060_reg/NET0131 ,
		_w2442_,
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1671 (
		\g35_pad ,
		_w2046_,
		_w2124_,
		_w2210_,
		_w2446_
	);
	LUT3 #(
		.INIT('hb0)
	) name1672 (
		_w2441_,
		_w2445_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h2)
	) name1673 (
		\g2060_reg/NET0131 ,
		\g35_pad ,
		_w2448_
	);
	LUT3 #(
		.INIT('hfe)
	) name1674 (
		_w2439_,
		_w2447_,
		_w2448_,
		_w2449_
	);
	LUT3 #(
		.INIT('h08)
	) name1675 (
		\g35_pad ,
		\g411_reg/NET0131 ,
		_w1824_,
		_w2450_
	);
	LUT4 #(
		.INIT('h8880)
	) name1676 (
		\g35_pad ,
		_w1824_,
		_w2060_,
		_w2061_,
		_w2451_
	);
	LUT2 #(
		.INIT('h4)
	) name1677 (
		\g35_pad ,
		\g417_reg/NET0131 ,
		_w2452_
	);
	LUT3 #(
		.INIT('hfe)
	) name1678 (
		_w2450_,
		_w2451_,
		_w2452_,
		_w2453_
	);
	LUT4 #(
		.INIT('h020a)
	) name1679 (
		\g35_pad ,
		_w2046_,
		_w2068_,
		_w2069_,
		_w2454_
	);
	LUT4 #(
		.INIT('hfdf5)
	) name1680 (
		\g35_pad ,
		_w2046_,
		_w2068_,
		_w2069_,
		_w2455_
	);
	LUT2 #(
		.INIT('h4)
	) name1681 (
		\g2217_reg/NET0131 ,
		\g35_pad ,
		_w2456_
	);
	LUT4 #(
		.INIT('h1300)
	) name1682 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h4)
	) name1683 (
		\g2208_reg/NET0131 ,
		\g35_pad ,
		_w2458_
	);
	LUT4 #(
		.INIT('hec00)
	) name1684 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		\g2223_reg/NET0131 ,
		\g35_pad ,
		_w2460_
	);
	LUT3 #(
		.INIT('h01)
	) name1686 (
		_w2457_,
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT4 #(
		.INIT('h020a)
	) name1687 (
		\g2236_reg/NET0131 ,
		_w2046_,
		_w2068_,
		_w2069_,
		_w2462_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		\g35_pad ,
		_w2462_,
		_w2463_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1689 (
		\g2165_reg/NET0131 ,
		\g2169_reg/NET0131 ,
		\g2185_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		_w2464_
	);
	LUT2 #(
		.INIT('h2)
	) name1690 (
		\g2217_reg/NET0131 ,
		_w2464_,
		_w2465_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1691 (
		\g2161_reg/NET0131 ,
		\g2173_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		_w2466_
	);
	LUT3 #(
		.INIT('h08)
	) name1692 (
		\g2181_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		_w2467_
	);
	LUT3 #(
		.INIT('h08)
	) name1693 (
		\g2177_reg/NET0131 ,
		\g2185_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		_w2468_
	);
	LUT4 #(
		.INIT('h000e)
	) name1694 (
		\g2185_reg/NET0131 ,
		_w2466_,
		_w2467_,
		_w2468_,
		_w2469_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1695 (
		\g35_pad ,
		_w2046_,
		_w2068_,
		_w2069_,
		_w2470_
	);
	LUT3 #(
		.INIT('hb0)
	) name1696 (
		_w2465_,
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h2)
	) name1697 (
		\g2217_reg/NET0131 ,
		\g35_pad ,
		_w2472_
	);
	LUT3 #(
		.INIT('hfe)
	) name1698 (
		_w2463_,
		_w2471_,
		_w2472_,
		_w2473_
	);
	LUT4 #(
		.INIT('h002a)
	) name1699 (
		\g35_pad ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2474_
	);
	LUT4 #(
		.INIT('hffd5)
	) name1700 (
		\g35_pad ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2475_
	);
	LUT4 #(
		.INIT('h0015)
	) name1701 (
		\g2351_reg/NET0131 ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2476_
	);
	LUT2 #(
		.INIT('h4)
	) name1702 (
		\g2342_reg/NET0131 ,
		\g35_pad ,
		_w2477_
	);
	LUT4 #(
		.INIT('hf800)
	) name1703 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('h002e)
	) name1704 (
		\g2357_reg/NET0131 ,
		\g35_pad ,
		_w2476_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('h002a)
	) name1705 (
		\g2370_reg/NET0131 ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2480_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		\g35_pad ,
		_w2480_,
		_w2481_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1707 (
		\g2299_reg/NET0131 ,
		\g2303_reg/NET0131 ,
		\g2319_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		_w2482_
	);
	LUT2 #(
		.INIT('h2)
	) name1708 (
		\g2351_reg/NET0131 ,
		_w2482_,
		_w2483_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1709 (
		\g2295_reg/NET0131 ,
		\g2307_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		_w2484_
	);
	LUT3 #(
		.INIT('h08)
	) name1710 (
		\g2315_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		_w2485_
	);
	LUT3 #(
		.INIT('h08)
	) name1711 (
		\g2311_reg/NET0131 ,
		\g2319_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		_w2486_
	);
	LUT4 #(
		.INIT('h000e)
	) name1712 (
		\g2319_reg/NET0131 ,
		_w2484_,
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('haa80)
	) name1713 (
		\g35_pad ,
		_w2046_,
		_w2075_,
		_w2076_,
		_w2488_
	);
	LUT3 #(
		.INIT('hb0)
	) name1714 (
		_w2483_,
		_w2487_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h2)
	) name1715 (
		\g2351_reg/NET0131 ,
		\g35_pad ,
		_w2490_
	);
	LUT3 #(
		.INIT('hfe)
	) name1716 (
		_w2481_,
		_w2489_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('h0222)
	) name1717 (
		\g35_pad ,
		_w2045_,
		_w2046_,
		_w2096_,
		_w2492_
	);
	LUT4 #(
		.INIT('hfddd)
	) name1718 (
		\g35_pad ,
		_w2045_,
		_w2046_,
		_w2096_,
		_w2493_
	);
	LUT2 #(
		.INIT('h4)
	) name1719 (
		\g2485_reg/NET0131 ,
		\g35_pad ,
		_w2494_
	);
	LUT4 #(
		.INIT('h1500)
	) name1720 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h4)
	) name1721 (
		\g2476_reg/NET0131 ,
		\g35_pad ,
		_w2496_
	);
	LUT4 #(
		.INIT('hea00)
	) name1722 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		\g2491_reg/NET0131 ,
		\g35_pad ,
		_w2498_
	);
	LUT3 #(
		.INIT('h01)
	) name1724 (
		_w2495_,
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('h0222)
	) name1725 (
		\g2504_reg/NET0131 ,
		_w2045_,
		_w2046_,
		_w2096_,
		_w2500_
	);
	LUT2 #(
		.INIT('h8)
	) name1726 (
		\g35_pad ,
		_w2500_,
		_w2501_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1727 (
		\g2433_reg/NET0131 ,
		\g2437_reg/NET0131 ,
		\g2453_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		_w2502_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		\g2485_reg/NET0131 ,
		_w2502_,
		_w2503_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1729 (
		\g2429_reg/NET0131 ,
		\g2441_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		_w2504_
	);
	LUT3 #(
		.INIT('h08)
	) name1730 (
		\g2449_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		_w2505_
	);
	LUT3 #(
		.INIT('h08)
	) name1731 (
		\g2445_reg/NET0131 ,
		\g2453_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		_w2506_
	);
	LUT4 #(
		.INIT('h000e)
	) name1732 (
		\g2453_reg/NET0131 ,
		_w2504_,
		_w2505_,
		_w2506_,
		_w2507_
	);
	LUT4 #(
		.INIT('ha888)
	) name1733 (
		\g35_pad ,
		_w2045_,
		_w2046_,
		_w2096_,
		_w2508_
	);
	LUT3 #(
		.INIT('hb0)
	) name1734 (
		_w2503_,
		_w2507_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h2)
	) name1735 (
		\g2485_reg/NET0131 ,
		\g35_pad ,
		_w2510_
	);
	LUT3 #(
		.INIT('hfe)
	) name1736 (
		_w2501_,
		_w2509_,
		_w2510_,
		_w2511_
	);
	LUT4 #(
		.INIT('h020a)
	) name1737 (
		\g35_pad ,
		_w2046_,
		_w2068_,
		_w2102_,
		_w2512_
	);
	LUT4 #(
		.INIT('hfdf5)
	) name1738 (
		\g35_pad ,
		_w2046_,
		_w2068_,
		_w2102_,
		_w2513_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		\g1657_reg/NET0131 ,
		\g35_pad ,
		_w2514_
	);
	LUT4 #(
		.INIT('h1300)
	) name1740 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2514_,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1741 (
		\g1648_reg/NET0131 ,
		\g35_pad ,
		_w2516_
	);
	LUT4 #(
		.INIT('hec00)
	) name1742 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		\g1664_reg/NET0131 ,
		\g35_pad ,
		_w2518_
	);
	LUT3 #(
		.INIT('h01)
	) name1744 (
		_w2515_,
		_w2517_,
		_w2518_,
		_w2519_
	);
	LUT4 #(
		.INIT('h020a)
	) name1745 (
		\g35_pad ,
		_w2046_,
		_w2124_,
		_w2125_,
		_w2520_
	);
	LUT4 #(
		.INIT('hfdf5)
	) name1746 (
		\g35_pad ,
		_w2046_,
		_w2124_,
		_w2125_,
		_w2521_
	);
	LUT4 #(
		.INIT('h020a)
	) name1747 (
		\g1677_reg/NET0131 ,
		_w2046_,
		_w2068_,
		_w2102_,
		_w2522_
	);
	LUT2 #(
		.INIT('h8)
	) name1748 (
		\g35_pad ,
		_w2522_,
		_w2523_
	);
	LUT4 #(
		.INIT('h51f3)
	) name1749 (
		\g1604_reg/NET0131 ,
		\g1616_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name1750 (
		\g1624_reg/NET0131 ,
		_w2524_,
		_w2525_
	);
	LUT4 #(
		.INIT('h31f5)
	) name1751 (
		\g1612_reg/NET0131 ,
		\g1620_reg/NET0131 ,
		\g1624_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w2526_
	);
	LUT3 #(
		.INIT('h20)
	) name1752 (
		\g1600_reg/NET0131 ,
		\g1624_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w2527_
	);
	LUT2 #(
		.INIT('h2)
	) name1753 (
		\g1608_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w2528_
	);
	LUT4 #(
		.INIT('h040e)
	) name1754 (
		\g1657_reg/NET0131 ,
		_w2526_,
		_w2527_,
		_w2528_,
		_w2529_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1755 (
		\g35_pad ,
		_w2046_,
		_w2068_,
		_w2102_,
		_w2530_
	);
	LUT3 #(
		.INIT('hb0)
	) name1756 (
		_w2525_,
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h2)
	) name1757 (
		\g1657_reg/NET0131 ,
		\g35_pad ,
		_w2532_
	);
	LUT3 #(
		.INIT('hfe)
	) name1758 (
		_w2523_,
		_w2531_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		\g2625_reg/NET0131 ,
		\g35_pad ,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		\g2619_reg/NET0131 ,
		\g35_pad ,
		_w2535_
	);
	LUT4 #(
		.INIT('h1300)
	) name1761 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		\g2610_reg/NET0131 ,
		\g35_pad ,
		_w2537_
	);
	LUT4 #(
		.INIT('hec00)
	) name1763 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2537_,
		_w2538_
	);
	LUT3 #(
		.INIT('hfe)
	) name1764 (
		_w2534_,
		_w2536_,
		_w2538_,
		_w2539_
	);
	LUT4 #(
		.INIT('h020a)
	) name1765 (
		\g2638_reg/NET0131 ,
		_w2046_,
		_w2124_,
		_w2125_,
		_w2540_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		\g35_pad ,
		_w2540_,
		_w2541_
	);
	LUT4 #(
		.INIT('h153f)
	) name1767 (
		\g2571_reg/NET0131 ,
		\g2579_reg/NET0131 ,
		\g2587_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		_w2542_
	);
	LUT2 #(
		.INIT('h1)
	) name1768 (
		\g2610_reg/NET0131 ,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('h31f5)
	) name1769 (
		\g2575_reg/NET0131 ,
		\g2583_reg/NET0131 ,
		\g2587_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		_w2544_
	);
	LUT3 #(
		.INIT('h20)
	) name1770 (
		\g2563_reg/NET0131 ,
		\g2587_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		_w2545_
	);
	LUT2 #(
		.INIT('h8)
	) name1771 (
		\g2567_reg/NET0131 ,
		\g2587_reg/NET0131 ,
		_w2546_
	);
	LUT4 #(
		.INIT('h040e)
	) name1772 (
		\g2619_reg/NET0131 ,
		_w2544_,
		_w2545_,
		_w2546_,
		_w2547_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1773 (
		\g35_pad ,
		_w2046_,
		_w2124_,
		_w2125_,
		_w2548_
	);
	LUT3 #(
		.INIT('hb0)
	) name1774 (
		_w2543_,
		_w2547_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h2)
	) name1775 (
		\g2619_reg/NET0131 ,
		\g35_pad ,
		_w2550_
	);
	LUT3 #(
		.INIT('hfe)
	) name1776 (
		_w2541_,
		_w2549_,
		_w2550_,
		_w2551_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		\g1691_reg/NET0131 ,
		\g35_pad ,
		_w2552_
	);
	LUT4 #(
		.INIT('h1300)
	) name1778 (
		_w2046_,
		_w2068_,
		_w2102_,
		_w2552_,
		_w2553_
	);
	LUT4 #(
		.INIT('hb000)
	) name1779 (
		\g1624_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		\g1691_reg/NET0131 ,
		\g35_pad ,
		_w2554_
	);
	LUT2 #(
		.INIT('h6)
	) name1780 (
		\g1677_reg/NET0131 ,
		_w2554_,
		_w2555_
	);
	LUT3 #(
		.INIT('hdc)
	) name1781 (
		_w2512_,
		_w2553_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h8)
	) name1782 (
		\g1825_reg/NET0131 ,
		\g35_pad ,
		_w2557_
	);
	LUT4 #(
		.INIT('h1300)
	) name1783 (
		_w2046_,
		_w2076_,
		_w2162_,
		_w2557_,
		_w2558_
	);
	LUT4 #(
		.INIT('hb000)
	) name1784 (
		\g1760_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		\g1825_reg/NET0131 ,
		\g35_pad ,
		_w2559_
	);
	LUT2 #(
		.INIT('h6)
	) name1785 (
		\g1811_reg/NET0131 ,
		_w2559_,
		_w2560_
	);
	LUT3 #(
		.INIT('hdc)
	) name1786 (
		_w2395_,
		_w2558_,
		_w2560_,
		_w2561_
	);
	LUT4 #(
		.INIT('heef0)
	) name1787 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		\g316_reg/NET0131 ,
		\g35_pad ,
		_w2562_
	);
	LUT4 #(
		.INIT('h0dd0)
	) name1788 (
		\g1008_reg/NET0131 ,
		\g1046_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w2563_
	);
	LUT2 #(
		.INIT('h1)
	) name1789 (
		\g969_reg/NET0131 ,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h80)
	) name1790 (
		\g1008_reg/NET0131 ,
		\g1018_reg/NET0131 ,
		\g1030_reg/NET0131 ,
		_w2565_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		\g1002_reg/NET0131 ,
		\g1018_reg/NET0131 ,
		_w2566_
	);
	LUT3 #(
		.INIT('h07)
	) name1792 (
		_w1971_,
		_w2565_,
		_w2566_,
		_w2567_
	);
	LUT3 #(
		.INIT('h15)
	) name1793 (
		_w1972_,
		_w2564_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('h15)
	) name1794 (
		\g1024_reg/NET0131 ,
		_w1971_,
		_w2565_,
		_w2569_
	);
	LUT2 #(
		.INIT('h1)
	) name1795 (
		\g1030_reg/NET0131 ,
		\g969_reg/NET0131 ,
		_w2570_
	);
	LUT2 #(
		.INIT('h4)
	) name1796 (
		_w2563_,
		_w2570_,
		_w2571_
	);
	LUT3 #(
		.INIT('h07)
	) name1797 (
		_w2564_,
		_w2569_,
		_w2571_,
		_w2572_
	);
	LUT3 #(
		.INIT('h15)
	) name1798 (
		\g1036_reg/NET0131 ,
		_w1971_,
		_w2565_,
		_w2573_
	);
	LUT3 #(
		.INIT('h2a)
	) name1799 (
		\g35_pad ,
		_w2564_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		\g1036_reg/NET0131 ,
		\g35_pad ,
		_w2575_
	);
	LUT4 #(
		.INIT('h087f)
	) name1801 (
		_w2568_,
		_w2572_,
		_w2574_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		\g1030_reg/NET0131 ,
		\g35_pad ,
		_w2577_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		_w2576_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		\g1959_reg/NET0131 ,
		\g35_pad ,
		_w2579_
	);
	LUT4 #(
		.INIT('h1500)
	) name1805 (
		_w2045_,
		_w2046_,
		_w2047_,
		_w2579_,
		_w2580_
	);
	LUT4 #(
		.INIT('hb000)
	) name1806 (
		\g1894_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		\g1959_reg/NET0131 ,
		\g35_pad ,
		_w2581_
	);
	LUT2 #(
		.INIT('h6)
	) name1807 (
		\g1945_reg/NET0131 ,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('hdc)
	) name1808 (
		_w2410_,
		_w2580_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		\g2250_reg/NET0131 ,
		\g35_pad ,
		_w2584_
	);
	LUT4 #(
		.INIT('h1300)
	) name1810 (
		_w2046_,
		_w2068_,
		_w2069_,
		_w2584_,
		_w2585_
	);
	LUT4 #(
		.INIT('hb000)
	) name1811 (
		\g2185_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		\g2250_reg/NET0131 ,
		\g35_pad ,
		_w2586_
	);
	LUT2 #(
		.INIT('h6)
	) name1812 (
		\g2236_reg/NET0131 ,
		_w2586_,
		_w2587_
	);
	LUT3 #(
		.INIT('hdc)
	) name1813 (
		_w2454_,
		_w2585_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		\g2384_reg/NET0131 ,
		\g35_pad ,
		_w2589_
	);
	LUT4 #(
		.INIT('h0700)
	) name1815 (
		_w2046_,
		_w2075_,
		_w2076_,
		_w2589_,
		_w2590_
	);
	LUT4 #(
		.INIT('hb000)
	) name1816 (
		\g2319_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		\g2384_reg/NET0131 ,
		\g35_pad ,
		_w2591_
	);
	LUT2 #(
		.INIT('h6)
	) name1817 (
		\g2370_reg/NET0131 ,
		_w2591_,
		_w2592_
	);
	LUT3 #(
		.INIT('hdc)
	) name1818 (
		_w2474_,
		_w2590_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h8)
	) name1819 (
		\g2518_reg/NET0131 ,
		\g35_pad ,
		_w2594_
	);
	LUT4 #(
		.INIT('h1500)
	) name1820 (
		_w2045_,
		_w2046_,
		_w2096_,
		_w2594_,
		_w2595_
	);
	LUT4 #(
		.INIT('hb000)
	) name1821 (
		\g2453_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		\g2518_reg/NET0131 ,
		\g35_pad ,
		_w2596_
	);
	LUT2 #(
		.INIT('h6)
	) name1822 (
		\g2504_reg/NET0131 ,
		_w2596_,
		_w2597_
	);
	LUT3 #(
		.INIT('hdc)
	) name1823 (
		_w2492_,
		_w2595_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h4)
	) name1824 (
		\g35_pad ,
		\g739_reg/NET0131 ,
		_w2599_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1825 (
		\g35_pad ,
		\g744_reg/NET0131 ,
		_w893_,
		_w1958_,
		_w2600_
	);
	LUT3 #(
		.INIT('h80)
	) name1826 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g739_reg/NET0131 ,
		_w2601_
	);
	LUT3 #(
		.INIT('h80)
	) name1827 (
		_w879_,
		_w881_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('h3222)
	) name1828 (
		\g744_reg/NET0131 ,
		_w883_,
		_w893_,
		_w2602_,
		_w2603_
	);
	LUT3 #(
		.INIT('hea)
	) name1829 (
		_w2599_,
		_w2600_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h8)
	) name1830 (
		\g2093_reg/NET0131 ,
		\g35_pad ,
		_w2605_
	);
	LUT4 #(
		.INIT('h1300)
	) name1831 (
		_w2046_,
		_w2124_,
		_w2210_,
		_w2605_,
		_w2606_
	);
	LUT4 #(
		.INIT('hb000)
	) name1832 (
		\g2028_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		\g2093_reg/NET0131 ,
		\g35_pad ,
		_w2607_
	);
	LUT2 #(
		.INIT('h6)
	) name1833 (
		\g2079_reg/NET0131 ,
		_w2607_,
		_w2608_
	);
	LUT3 #(
		.INIT('hdc)
	) name1834 (
		_w2430_,
		_w2606_,
		_w2608_,
		_w2609_
	);
	LUT2 #(
		.INIT('h8)
	) name1835 (
		\g2652_reg/NET0131 ,
		\g35_pad ,
		_w2610_
	);
	LUT4 #(
		.INIT('h1300)
	) name1836 (
		_w2046_,
		_w2124_,
		_w2125_,
		_w2610_,
		_w2611_
	);
	LUT4 #(
		.INIT('hb000)
	) name1837 (
		\g2587_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		\g2652_reg/NET0131 ,
		\g35_pad ,
		_w2612_
	);
	LUT2 #(
		.INIT('h6)
	) name1838 (
		\g2638_reg/NET0131 ,
		_w2612_,
		_w2613_
	);
	LUT3 #(
		.INIT('hdc)
	) name1839 (
		_w2520_,
		_w2611_,
		_w2613_,
		_w2614_
	);
	LUT3 #(
		.INIT('h20)
	) name1840 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w2615_
	);
	LUT3 #(
		.INIT('h07)
	) name1841 (
		\g482_reg/NET0131 ,
		\g490_reg/NET0131 ,
		\g528_reg/NET0131 ,
		_w2616_
	);
	LUT3 #(
		.INIT('ha2)
	) name1842 (
		\g490_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w2617_
	);
	LUT4 #(
		.INIT('h0008)
	) name1843 (
		_w1688_,
		_w2615_,
		_w2616_,
		_w2617_,
		_w2618_
	);
	LUT3 #(
		.INIT('ha8)
	) name1844 (
		\g482_reg/NET0131 ,
		\g490_reg/NET0131 ,
		\g528_reg/NET0131 ,
		_w2619_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1845 (
		\g35_pad ,
		\g490_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w2620_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1846 (
		_w1688_,
		_w2615_,
		_w2619_,
		_w2620_,
		_w2621_
	);
	LUT4 #(
		.INIT('hffc4)
	) name1847 (
		\g35_pad ,
		\g482_reg/NET0131 ,
		_w2618_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h4)
	) name1848 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		_w2623_
	);
	LUT3 #(
		.INIT('h15)
	) name1849 (
		\g739_reg/NET0131 ,
		_w893_,
		_w1693_,
		_w2624_
	);
	LUT3 #(
		.INIT('h8a)
	) name1850 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w2625_
	);
	LUT3 #(
		.INIT('h70)
	) name1851 (
		_w893_,
		_w2602_,
		_w2625_,
		_w2626_
	);
	LUT3 #(
		.INIT('hba)
	) name1852 (
		_w2623_,
		_w2624_,
		_w2626_,
		_w2627_
	);
	LUT3 #(
		.INIT('h80)
	) name1853 (
		\g1087_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		\g1221_reg/NET0131 ,
		_w2628_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		\g1211_reg/NET0131 ,
		\g35_pad ,
		_w2629_
	);
	LUT2 #(
		.INIT('h4)
	) name1855 (
		_w2628_,
		_w2629_,
		_w2630_
	);
	LUT4 #(
		.INIT('h0800)
	) name1856 (
		\g1087_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1221_reg/NET0131 ,
		_w2631_
	);
	LUT3 #(
		.INIT('ha2)
	) name1857 (
		\g1216_reg/NET0131 ,
		\g35_pad ,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('he)
	) name1858 (
		_w2630_,
		_w2632_,
		_w2633_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1859 (
		\g35_pad ,
		_w1791_,
		_w1793_,
		_w1794_,
		_w2634_
	);
	LUT4 #(
		.INIT('h0080)
	) name1860 (
		\g4311_reg/NET0131 ,
		\g4621_reg/NET0131 ,
		\g4628_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w2635_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name1861 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		_w1793_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name1862 (
		\g35_pad ,
		\g4322_reg/NET0131 ,
		_w2637_
	);
	LUT2 #(
		.INIT('h2)
	) name1863 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		_w2638_
	);
	LUT4 #(
		.INIT('h070f)
	) name1864 (
		_w1793_,
		_w2635_,
		_w2637_,
		_w2638_,
		_w2639_
	);
	LUT3 #(
		.INIT('h8f)
	) name1865 (
		_w2634_,
		_w2636_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h2)
	) name1866 (
		\g1559_reg/NET0131 ,
		\g35_pad ,
		_w2641_
	);
	LUT4 #(
		.INIT('h8000)
	) name1867 (
		\g1430_reg/NET0131 ,
		\g1548_reg/NET0131 ,
		\g1559_reg/NET0131 ,
		\g1564_reg/NET0131 ,
		_w2642_
	);
	LUT4 #(
		.INIT('h0c08)
	) name1868 (
		\g1554_reg/NET0131 ,
		\g35_pad ,
		_w1124_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('he)
	) name1869 (
		_w2641_,
		_w2643_,
		_w2644_
	);
	LUT4 #(
		.INIT('h88a0)
	) name1870 (
		\g35_pad ,
		\g5069_reg/NET0131 ,
		\g5073_reg/NET0131 ,
		\g5084_reg/NET0131 ,
		_w2645_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		\g5077_reg/NET0131 ,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name1872 (
		\g246_reg/NET0131 ,
		\g35_pad ,
		_w2647_
	);
	LUT3 #(
		.INIT('hb8)
	) name1873 (
		\g246_reg/NET0131 ,
		\g35_pad ,
		\g479_reg/NET0131 ,
		_w2648_
	);
	LUT2 #(
		.INIT('h4)
	) name1874 (
		\g35_pad ,
		\g4584_reg/NET0131 ,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		\g35_pad ,
		\g4593_reg/NET0131 ,
		_w2650_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1876 (
		_w1791_,
		_w1793_,
		_w1799_,
		_w2650_,
		_w2651_
	);
	LUT3 #(
		.INIT('h02)
	) name1877 (
		\g35_pad ,
		\g4593_reg/NET0131 ,
		\g4616_reg/NET0131 ,
		_w2652_
	);
	LUT4 #(
		.INIT('h8000)
	) name1878 (
		_w1791_,
		_w1793_,
		_w1799_,
		_w2652_,
		_w2653_
	);
	LUT3 #(
		.INIT('hfe)
	) name1879 (
		_w2649_,
		_w2651_,
		_w2653_,
		_w2654_
	);
	LUT4 #(
		.INIT('h0040)
	) name1880 (
		\g862_reg/NET0131 ,
		\g872_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w2655_
	);
	LUT3 #(
		.INIT('h04)
	) name1881 (
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name1882 (
		\g35_pad ,
		\g446_reg/NET0131 ,
		_w2657_
	);
	LUT4 #(
		.INIT('h5f57)
	) name1883 (
		\g35_pad ,
		\g446_reg/NET0131 ,
		_w2655_,
		_w2656_,
		_w2658_
	);
	LUT2 #(
		.INIT('h2)
	) name1884 (
		\g246_reg/NET0131 ,
		\g35_pad ,
		_w2659_
	);
	LUT2 #(
		.INIT('hd)
	) name1885 (
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT4 #(
		.INIT('h1d00)
	) name1886 (
		\g854_reg/NET0131 ,
		_w2055_,
		_w2059_,
		_w2062_,
		_w2661_
	);
	LUT2 #(
		.INIT('h2)
	) name1887 (
		\g35_pad ,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h4)
	) name1888 (
		\g4340_reg/NET0131 ,
		_w930_,
		_w2663_
	);
	LUT4 #(
		.INIT('h0400)
	) name1889 (
		\g4340_reg/NET0131 ,
		_w929_,
		_w933_,
		_w934_,
		_w2664_
	);
	LUT3 #(
		.INIT('h20)
	) name1890 (
		\g4311_reg/NET0131 ,
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		_w2665_
	);
	LUT3 #(
		.INIT('h02)
	) name1891 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		\g4515_reg/NET0131 ,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name1892 (
		\g4340_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		_w2667_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		\g35_pad ,
		\g4358_reg/NET0131 ,
		_w2668_
	);
	LUT4 #(
		.INIT('hef00)
	) name1894 (
		_w2665_,
		_w2666_,
		_w2667_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1895 (
		\g4349_reg/NET0131 ,
		_w2663_,
		_w2664_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h8)
	) name1896 (
		\g35_pad ,
		\g4358_reg/NET0131 ,
		_w2671_
	);
	LUT3 #(
		.INIT('h27)
	) name1897 (
		\g35_pad ,
		\g4358_reg/NET0131 ,
		\g4366_reg/NET0131 ,
		_w2672_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name1898 (
		\g35_pad ,
		\g4340_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		\g4366_reg/NET0131 ,
		_w2673_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1899 (
		_w2663_,
		_w2664_,
		_w2672_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('he)
	) name1900 (
		_w2670_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		\g1024_reg/NET0131 ,
		\g35_pad ,
		_w2676_
	);
	LUT4 #(
		.INIT('h1115)
	) name1902 (
		_w1972_,
		_w2564_,
		_w2567_,
		_w2569_,
		_w2677_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		\g1030_reg/NET0131 ,
		_w2677_,
		_w2678_
	);
	LUT3 #(
		.INIT('h2a)
	) name1904 (
		\g35_pad ,
		_w2568_,
		_w2572_,
		_w2679_
	);
	LUT3 #(
		.INIT('hba)
	) name1905 (
		_w2676_,
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT3 #(
		.INIT('h80)
	) name1906 (
		\g4776_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		_w2681_
	);
	LUT2 #(
		.INIT('h8)
	) name1907 (
		\g35_pad ,
		\g4709_reg/NET0131 ,
		_w2682_
	);
	LUT3 #(
		.INIT('h70)
	) name1908 (
		_w1981_,
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT3 #(
		.INIT('h70)
	) name1909 (
		\g35_pad ,
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w2684_
	);
	LUT4 #(
		.INIT('hd500)
	) name1910 (
		\g35_pad ,
		_w1981_,
		_w2377_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('he)
	) name1911 (
		_w2683_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h8)
	) name1912 (
		\g843_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w2687_
	);
	LUT3 #(
		.INIT('h15)
	) name1913 (
		\g812_reg/NET0131 ,
		_w1824_,
		_w2687_,
		_w2688_
	);
	LUT3 #(
		.INIT('h80)
	) name1914 (
		\g812_reg/NET0131 ,
		\g843_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w2689_
	);
	LUT3 #(
		.INIT('h2a)
	) name1915 (
		\g837_reg/NET0131 ,
		_w1824_,
		_w2689_,
		_w2690_
	);
	LUT4 #(
		.INIT('h4e44)
	) name1916 (
		\g35_pad ,
		\g843_reg/NET0131 ,
		_w2688_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h4)
	) name1917 (
		\g35_pad ,
		\g667_reg/NET0131 ,
		_w2692_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1918 (
		\g671_reg/NET0131 ,
		_w1824_,
		_w2022_,
		_w2023_,
		_w2693_
	);
	LUT4 #(
		.INIT('h7000)
	) name1919 (
		_w2024_,
		_w2028_,
		_w2029_,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('he)
	) name1920 (
		_w2692_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h4)
	) name1921 (
		\g283_reg/NET0131 ,
		\g35_pad ,
		_w2696_
	);
	LUT2 #(
		.INIT('h2)
	) name1922 (
		\g278_reg/NET0131 ,
		\g35_pad ,
		_w2697_
	);
	LUT3 #(
		.INIT('hf8)
	) name1923 (
		_w1715_,
		_w2696_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		\g35_pad ,
		\g817_reg/NET0131 ,
		_w2699_
	);
	LUT4 #(
		.INIT('h6c00)
	) name1925 (
		\g817_reg/NET0131 ,
		\g832_reg/NET0131 ,
		_w1824_,
		_w1829_,
		_w2700_
	);
	LUT2 #(
		.INIT('he)
	) name1926 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		\g35_pad ,
		\g4793_reg/NET0131 ,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		\g35_pad ,
		\g4801_reg/NET0131 ,
		_w2703_
	);
	LUT3 #(
		.INIT('h02)
	) name1929 (
		\g35_pad ,
		\g4776_reg/NET0131 ,
		\g4801_reg/NET0131 ,
		_w2704_
	);
	LUT4 #(
		.INIT('h078f)
	) name1930 (
		\g4793_reg/NET0131 ,
		_w1981_,
		_w2703_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('hb)
	) name1931 (
		_w2702_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h0004)
	) name1932 (
		\g5016_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		\g5029_reg/NET0131 ,
		\g5033_reg/NET0131 ,
		_w2707_
	);
	LUT3 #(
		.INIT('h01)
	) name1933 (
		\g5037_reg/NET0131 ,
		\g5041_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		_w2708_
	);
	LUT4 #(
		.INIT('h8000)
	) name1934 (
		\g3050_reg/NET0131 ,
		\g5016_reg/NET0131 ,
		\g5029_reg/NET0131 ,
		\g5033_reg/NET0131 ,
		_w2709_
	);
	LUT3 #(
		.INIT('h80)
	) name1935 (
		\g5037_reg/NET0131 ,
		\g5041_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		_w2710_
	);
	LUT4 #(
		.INIT('h0777)
	) name1936 (
		_w2707_,
		_w2708_,
		_w2709_,
		_w2710_,
		_w2711_
	);
	LUT4 #(
		.INIT('h0080)
	) name1937 (
		\g3050_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w2712_
	);
	LUT4 #(
		.INIT('hf070)
	) name1938 (
		\g3050_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name1939 (
		\g35_pad ,
		_w2713_,
		_w2714_
	);
	LUT2 #(
		.INIT('h2)
	) name1940 (
		\g35_pad ,
		\g5052_reg/NET0131 ,
		_w2715_
	);
	LUT2 #(
		.INIT('h4)
	) name1941 (
		\g35_pad ,
		\g5046_reg/NET0131 ,
		_w2716_
	);
	LUT4 #(
		.INIT('hffd8)
	) name1942 (
		_w2711_,
		_w2714_,
		_w2715_,
		_w2716_,
		_w2717_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1943 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w2718_
	);
	LUT2 #(
		.INIT('h8)
	) name1944 (
		\g35_pad ,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('h2010)
	) name1945 (
		\g655_reg/NET0131 ,
		\g691_reg/NET0131 ,
		\g703_reg/NET0131 ,
		\g718_reg/NET0131 ,
		_w2720_
	);
	LUT4 #(
		.INIT('h0800)
	) name1946 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w2721_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1947 (
		_w2026_,
		_w2027_,
		_w2720_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name1948 (
		\g35_pad ,
		\g691_reg/NET0131 ,
		_w2723_
	);
	LUT3 #(
		.INIT('hfe)
	) name1949 (
		_w2719_,
		_w2722_,
		_w2723_,
		_w2724_
	);
	LUT3 #(
		.INIT('hca)
	) name1950 (
		\g29216_pad ,
		\g316_reg/NET0131 ,
		\g35_pad ,
		_w2725_
	);
	LUT2 #(
		.INIT('h4)
	) name1951 (
		\g35_pad ,
		\g4776_reg/NET0131 ,
		_w2726_
	);
	LUT4 #(
		.INIT('h2888)
	) name1952 (
		\g35_pad ,
		\g4785_reg/NET0131 ,
		_w1981_,
		_w2377_,
		_w2727_
	);
	LUT2 #(
		.INIT('he)
	) name1953 (
		_w2726_,
		_w2727_,
		_w2728_
	);
	LUT4 #(
		.INIT('h0020)
	) name1954 (
		\g14167_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w2729_
	);
	LUT4 #(
		.INIT('h33f7)
	) name1955 (
		\g246_reg/NET0131 ,
		\g35_pad ,
		_w2656_,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h2)
	) name1956 (
		\g269_reg/NET0131 ,
		\g35_pad ,
		_w2731_
	);
	LUT2 #(
		.INIT('hd)
	) name1957 (
		_w2730_,
		_w2731_,
		_w2732_
	);
	LUT3 #(
		.INIT('h48)
	) name1958 (
		\g1171_reg/NET0131 ,
		\g35_pad ,
		\g7916_pad ,
		_w2733_
	);
	LUT4 #(
		.INIT('h2000)
	) name1959 (
		\g1178_reg/NET0131 ,
		\g1189_reg/NET0131 ,
		\g7916_pad ,
		\g996_reg/NET0131 ,
		_w2734_
	);
	LUT3 #(
		.INIT('ha4)
	) name1960 (
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w2735_
	);
	LUT3 #(
		.INIT('h80)
	) name1961 (
		\g1002_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1036_reg/NET0131 ,
		_w2736_
	);
	LUT4 #(
		.INIT('h3bbb)
	) name1962 (
		_w801_,
		_w2734_,
		_w2735_,
		_w2736_,
		_w2737_
	);
	LUT3 #(
		.INIT('hb0)
	) name1963 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		_w2738_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1964 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		\g35_pad ,
		_w2739_
	);
	LUT3 #(
		.INIT('hba)
	) name1965 (
		_w2733_,
		_w2737_,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h2)
	) name1966 (
		\g1018_reg/NET0131 ,
		\g35_pad ,
		_w2741_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		\g1024_reg/NET0131 ,
		\g35_pad ,
		_w2742_
	);
	LUT3 #(
		.INIT('h80)
	) name1968 (
		\g35_pad ,
		_w2564_,
		_w2569_,
		_w2743_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1969 (
		_w2568_,
		_w2741_,
		_w2742_,
		_w2743_,
		_w2744_
	);
	LUT3 #(
		.INIT('h20)
	) name1970 (
		\g1178_reg/NET0131 ,
		\g1189_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w2745_
	);
	LUT4 #(
		.INIT('h4000)
	) name1971 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1199_reg/NET0131 ,
		\g7916_pad ,
		_w2746_
	);
	LUT3 #(
		.INIT('h8a)
	) name1972 (
		\g35_pad ,
		_w2745_,
		_w2746_,
		_w2747_
	);
	LUT4 #(
		.INIT('h8088)
	) name1973 (
		\g1070_reg/NET0131 ,
		\g35_pad ,
		_w2745_,
		_w2746_,
		_w2748_
	);
	LUT4 #(
		.INIT('h1000)
	) name1974 (
		\g1070_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g7916_pad ,
		_w2749_
	);
	LUT4 #(
		.INIT('h2a22)
	) name1975 (
		\g1199_reg/NET0131 ,
		\g35_pad ,
		_w2745_,
		_w2749_,
		_w2750_
	);
	LUT4 #(
		.INIT('hffe0)
	) name1976 (
		_w2737_,
		_w2738_,
		_w2748_,
		_w2750_,
		_w2751_
	);
	LUT3 #(
		.INIT('h40)
	) name1977 (
		\g5052_reg/NET0131 ,
		_w2707_,
		_w2708_,
		_w2752_
	);
	LUT3 #(
		.INIT('h80)
	) name1978 (
		\g5052_reg/NET0131 ,
		_w2709_,
		_w2710_,
		_w2753_
	);
	LUT4 #(
		.INIT('h0200)
	) name1979 (
		\g5022_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w2754_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1980 (
		\g5022_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w2755_
	);
	LUT3 #(
		.INIT('h20)
	) name1981 (
		\g35_pad ,
		_w2712_,
		_w2755_,
		_w2756_
	);
	LUT3 #(
		.INIT('h10)
	) name1982 (
		_w2752_,
		_w2753_,
		_w2756_,
		_w2757_
	);
	LUT2 #(
		.INIT('h4)
	) name1983 (
		\g35_pad ,
		\g5052_reg/NET0131 ,
		_w2758_
	);
	LUT3 #(
		.INIT('h08)
	) name1984 (
		\g35_pad ,
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w2759_
	);
	LUT3 #(
		.INIT('h80)
	) name1985 (
		_w2709_,
		_w2710_,
		_w2759_,
		_w2760_
	);
	LUT3 #(
		.INIT('h02)
	) name1986 (
		\g35_pad ,
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w2761_
	);
	LUT3 #(
		.INIT('h80)
	) name1987 (
		_w2707_,
		_w2708_,
		_w2761_,
		_w2762_
	);
	LUT3 #(
		.INIT('h01)
	) name1988 (
		_w2758_,
		_w2760_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('hb)
	) name1989 (
		_w2757_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name1990 (
		\g1216_reg/NET0131 ,
		\g35_pad ,
		_w2765_
	);
	LUT3 #(
		.INIT('he0)
	) name1991 (
		\g1211_reg/NET0131 ,
		\g1216_reg/NET0131 ,
		\g35_pad ,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name1992 (
		\g1221_reg/NET0131 ,
		\g35_pad ,
		_w2767_
	);
	LUT4 #(
		.INIT('h001b)
	) name1993 (
		_w2628_,
		_w2765_,
		_w2766_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h8)
	) name1994 (
		\g3338_reg/NET0131 ,
		\g35_pad ,
		_w2769_
	);
	LUT4 #(
		.INIT('h8000)
	) name1995 (
		\g13895_pad ,
		\g16603_pad ,
		\g16718_pad ,
		\g3303_reg/NET0131 ,
		_w2770_
	);
	LUT3 #(
		.INIT('h2a)
	) name1996 (
		\g3343_reg/NET0131 ,
		_w2769_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name1997 (
		\g1564_reg/NET0131 ,
		\g35_pad ,
		_w2772_
	);
	LUT3 #(
		.INIT('h80)
	) name1998 (
		\g1430_reg/NET0131 ,
		\g1548_reg/NET0131 ,
		\g1564_reg/NET0131 ,
		_w2773_
	);
	LUT2 #(
		.INIT('h8)
	) name1999 (
		\g1559_reg/NET0131 ,
		\g35_pad ,
		_w2774_
	);
	LUT3 #(
		.INIT('h10)
	) name2000 (
		\g1554_reg/NET0131 ,
		\g1559_reg/NET0131 ,
		\g35_pad ,
		_w2775_
	);
	LUT4 #(
		.INIT('hfeba)
	) name2001 (
		_w2772_,
		_w2773_,
		_w2774_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h2)
	) name2002 (
		\g2771_reg/NET0131 ,
		\g35_pad ,
		_w2777_
	);
	LUT2 #(
		.INIT('hd)
	) name2003 (
		_w2331_,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		\g2803_reg/NET0131 ,
		\g35_pad ,
		_w2779_
	);
	LUT2 #(
		.INIT('hd)
	) name2005 (
		_w2361_,
		_w2779_,
		_w2780_
	);
	LUT3 #(
		.INIT('h70)
	) name2006 (
		_w1791_,
		_w1792_,
		_w2671_,
		_w2781_
	);
	LUT4 #(
		.INIT('h0080)
	) name2007 (
		\g4340_reg/NET0131 ,
		\g4621_reg/NET0131 ,
		\g4628_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w2782_
	);
	LUT3 #(
		.INIT('h4c)
	) name2008 (
		\g35_pad ,
		\g4349_reg/NET0131 ,
		\g4358_reg/NET0131 ,
		_w2783_
	);
	LUT3 #(
		.INIT('hd0)
	) name2009 (
		\g35_pad ,
		_w2782_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('he)
	) name2010 (
		_w2781_,
		_w2784_,
		_w2785_
	);
	LUT4 #(
		.INIT('ha800)
	) name2011 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		\g324_reg/NET0131 ,
		\g35_pad ,
		_w2786_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		\g336_reg/NET0131 ,
		\g35_pad ,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2013 (
		\g311_reg/NET0131 ,
		\g35_pad ,
		_w2788_
	);
	LUT4 #(
		.INIT('hffdc)
	) name2014 (
		_w1788_,
		_w2786_,
		_w2787_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h4)
	) name2015 (
		\g35_pad ,
		\g4311_reg/NET0131 ,
		_w2790_
	);
	LUT3 #(
		.INIT('h6a)
	) name2016 (
		\g4322_reg/NET0131 ,
		_w1793_,
		_w2635_,
		_w2791_
	);
	LUT3 #(
		.INIT('hec)
	) name2017 (
		_w2634_,
		_w2790_,
		_w2791_,
		_w2792_
	);
	LUT4 #(
		.INIT('h0020)
	) name2018 (
		\g14189_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w2793_
	);
	LUT4 #(
		.INIT('h33f7)
	) name2019 (
		\g225_reg/NET0131 ,
		\g35_pad ,
		_w2656_,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h4)
	) name2020 (
		\g35_pad ,
		\g872_reg/NET0131 ,
		_w2795_
	);
	LUT2 #(
		.INIT('hd)
	) name2021 (
		_w2794_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('h6ce4)
	) name2022 (
		\g35_pad ,
		\g4653_reg/NET0131 ,
		\g4659_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w2797_
	);
	LUT3 #(
		.INIT('hfd)
	) name2023 (
		\g35_pad ,
		_w1646_,
		_w1648_,
		_w2798_
	);
	LUT3 #(
		.INIT('hfd)
	) name2024 (
		\g35_pad ,
		_w1420_,
		_w1422_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name2025 (
		\g2667_reg/NET0131 ,
		\g35_pad ,
		_w2800_
	);
	LUT2 #(
		.INIT('h2)
	) name2026 (
		\g2661_reg/NET0131 ,
		\g2667_reg/NET0131 ,
		_w2801_
	);
	LUT4 #(
		.INIT('h010f)
	) name2027 (
		_w1420_,
		_w1422_,
		_w2800_,
		_w2801_,
		_w2802_
	);
	LUT3 #(
		.INIT('h40)
	) name2028 (
		\g2661_reg/NET0131 ,
		\g2667_reg/NET0131 ,
		\g35_pad ,
		_w2803_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		\g2671_reg/NET0131 ,
		\g35_pad ,
		_w2804_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2030 (
		_w1420_,
		_w1422_,
		_w2803_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		_w2802_,
		_w2805_,
		_w2806_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2032 (
		\g2675_reg/NET0131 ,
		\g35_pad ,
		_w1420_,
		_w1422_,
		_w2807_
	);
	LUT2 #(
		.INIT('h2)
	) name2033 (
		\g2671_reg/NET0131 ,
		\g35_pad ,
		_w2808_
	);
	LUT2 #(
		.INIT('hd)
	) name2034 (
		_w2807_,
		_w2808_,
		_w2809_
	);
	LUT4 #(
		.INIT('h0020)
	) name2035 (
		\g14147_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w2810_
	);
	LUT2 #(
		.INIT('h8)
	) name2036 (
		\g269_reg/NET0131 ,
		\g35_pad ,
		_w2811_
	);
	LUT4 #(
		.INIT('h33f7)
	) name2037 (
		\g269_reg/NET0131 ,
		\g35_pad ,
		_w2656_,
		_w2810_,
		_w2812_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		\g239_reg/NET0131 ,
		\g35_pad ,
		_w2813_
	);
	LUT2 #(
		.INIT('hd)
	) name2039 (
		_w2812_,
		_w2813_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name2040 (
		\g1706_reg/NET0131 ,
		\g35_pad ,
		_w2815_
	);
	LUT2 #(
		.INIT('h2)
	) name2041 (
		\g1700_reg/NET0131 ,
		\g1706_reg/NET0131 ,
		_w2816_
	);
	LUT4 #(
		.INIT('h010f)
	) name2042 (
		_w1646_,
		_w1648_,
		_w2815_,
		_w2816_,
		_w2817_
	);
	LUT3 #(
		.INIT('h40)
	) name2043 (
		\g1700_reg/NET0131 ,
		\g1706_reg/NET0131 ,
		\g35_pad ,
		_w2818_
	);
	LUT2 #(
		.INIT('h4)
	) name2044 (
		\g1710_reg/NET0131 ,
		\g35_pad ,
		_w2819_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2045 (
		_w1646_,
		_w1648_,
		_w2818_,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h8)
	) name2046 (
		_w2817_,
		_w2820_,
		_w2821_
	);
	LUT3 #(
		.INIT('h01)
	) name2047 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2767_reg/NET0131 ,
		_w2822_
	);
	LUT3 #(
		.INIT('h80)
	) name2048 (
		\g35_pad ,
		_w1910_,
		_w2822_,
		_w2823_
	);
	LUT2 #(
		.INIT('h8)
	) name2049 (
		\g2771_reg/NET0131 ,
		\g35_pad ,
		_w2824_
	);
	LUT3 #(
		.INIT('h70)
	) name2050 (
		_w1910_,
		_w2044_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		\g2775_reg/NET0131 ,
		\g35_pad ,
		_w2826_
	);
	LUT3 #(
		.INIT('hfe)
	) name2052 (
		_w2823_,
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name2053 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2828_
	);
	LUT3 #(
		.INIT('h02)
	) name2054 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2779_reg/NET0131 ,
		_w2829_
	);
	LUT3 #(
		.INIT('h80)
	) name2055 (
		\g35_pad ,
		_w1910_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		\g2775_reg/NET0131 ,
		\g35_pad ,
		_w2831_
	);
	LUT3 #(
		.INIT('h70)
	) name2057 (
		_w1910_,
		_w2828_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h2)
	) name2058 (
		\g2783_reg/NET0131 ,
		\g35_pad ,
		_w2833_
	);
	LUT3 #(
		.INIT('hfe)
	) name2059 (
		_w2830_,
		_w2832_,
		_w2833_,
		_w2834_
	);
	LUT3 #(
		.INIT('h04)
	) name2060 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2791_reg/NET0131 ,
		_w2835_
	);
	LUT3 #(
		.INIT('h80)
	) name2061 (
		\g35_pad ,
		_w1910_,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h4)
	) name2062 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2837_
	);
	LUT2 #(
		.INIT('h8)
	) name2063 (
		\g2783_reg/NET0131 ,
		\g35_pad ,
		_w2838_
	);
	LUT3 #(
		.INIT('h70)
	) name2064 (
		_w1910_,
		_w2837_,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('h2)
	) name2065 (
		\g2787_reg/NET0131 ,
		\g35_pad ,
		_w2840_
	);
	LUT3 #(
		.INIT('hfe)
	) name2066 (
		_w2836_,
		_w2839_,
		_w2840_,
		_w2841_
	);
	LUT3 #(
		.INIT('h08)
	) name2067 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2795_reg/NET0131 ,
		_w2842_
	);
	LUT3 #(
		.INIT('h80)
	) name2068 (
		\g35_pad ,
		_w1910_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2844_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		\g2787_reg/NET0131 ,
		\g35_pad ,
		_w2845_
	);
	LUT3 #(
		.INIT('h70)
	) name2071 (
		_w1910_,
		_w2844_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name2072 (
		\g2795_reg/NET0131 ,
		\g35_pad ,
		_w2847_
	);
	LUT3 #(
		.INIT('hfe)
	) name2073 (
		_w2843_,
		_w2846_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2074 (
		\g1714_reg/NET0131 ,
		\g35_pad ,
		_w1646_,
		_w1648_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2075 (
		\g1710_reg/NET0131 ,
		\g35_pad ,
		_w2850_
	);
	LUT2 #(
		.INIT('hd)
	) name2076 (
		_w2849_,
		_w2850_,
		_w2851_
	);
	LUT3 #(
		.INIT('h01)
	) name2077 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2799_reg/NET0131 ,
		_w2852_
	);
	LUT3 #(
		.INIT('h80)
	) name2078 (
		\g35_pad ,
		_w1910_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h8)
	) name2079 (
		\g2803_reg/NET0131 ,
		\g35_pad ,
		_w2854_
	);
	LUT3 #(
		.INIT('h70)
	) name2080 (
		_w1910_,
		_w2044_,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h2)
	) name2081 (
		\g2807_reg/NET0131 ,
		\g35_pad ,
		_w2856_
	);
	LUT3 #(
		.INIT('hfe)
	) name2082 (
		_w2853_,
		_w2855_,
		_w2856_,
		_w2857_
	);
	LUT3 #(
		.INIT('h02)
	) name2083 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2811_reg/NET0131 ,
		_w2858_
	);
	LUT3 #(
		.INIT('h80)
	) name2084 (
		\g35_pad ,
		_w1910_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		\g2807_reg/NET0131 ,
		\g35_pad ,
		_w2860_
	);
	LUT3 #(
		.INIT('h70)
	) name2086 (
		_w1910_,
		_w2828_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h2)
	) name2087 (
		\g2815_reg/NET0131 ,
		\g35_pad ,
		_w2862_
	);
	LUT3 #(
		.INIT('hfe)
	) name2088 (
		_w2859_,
		_w2861_,
		_w2862_,
		_w2863_
	);
	LUT3 #(
		.INIT('h04)
	) name2089 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2823_reg/NET0131 ,
		_w2864_
	);
	LUT3 #(
		.INIT('h80)
	) name2090 (
		\g35_pad ,
		_w1910_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h8)
	) name2091 (
		\g2815_reg/NET0131 ,
		\g35_pad ,
		_w2866_
	);
	LUT3 #(
		.INIT('h70)
	) name2092 (
		_w1910_,
		_w2837_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h2)
	) name2093 (
		\g2819_reg/NET0131 ,
		\g35_pad ,
		_w2868_
	);
	LUT3 #(
		.INIT('hfe)
	) name2094 (
		_w2865_,
		_w2867_,
		_w2868_,
		_w2869_
	);
	LUT3 #(
		.INIT('h08)
	) name2095 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		\g2827_reg/NET0131 ,
		_w2870_
	);
	LUT3 #(
		.INIT('h80)
	) name2096 (
		\g35_pad ,
		_w1910_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		\g2819_reg/NET0131 ,
		\g35_pad ,
		_w2872_
	);
	LUT3 #(
		.INIT('h70)
	) name2098 (
		_w1910_,
		_w2844_,
		_w2872_,
		_w2873_
	);
	LUT2 #(
		.INIT('h2)
	) name2099 (
		\g2827_reg/NET0131 ,
		\g35_pad ,
		_w2874_
	);
	LUT3 #(
		.INIT('hfe)
	) name2100 (
		_w2871_,
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT3 #(
		.INIT('hfd)
	) name2101 (
		\g35_pad ,
		_w1502_,
		_w1504_,
		_w2876_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2102 (
		\g1816_reg/NET0131 ,
		\g35_pad ,
		_w1502_,
		_w1504_,
		_w2877_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		\g1821_reg/NET0131 ,
		\g35_pad ,
		_w2878_
	);
	LUT3 #(
		.INIT('h10)
	) name2104 (
		_w1502_,
		_w1504_,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('he)
	) name2105 (
		_w2877_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h1)
	) name2106 (
		\g1840_reg/NET0131 ,
		\g35_pad ,
		_w2881_
	);
	LUT2 #(
		.INIT('h2)
	) name2107 (
		\g1834_reg/NET0131 ,
		\g1840_reg/NET0131 ,
		_w2882_
	);
	LUT4 #(
		.INIT('h010f)
	) name2108 (
		_w1502_,
		_w1504_,
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT3 #(
		.INIT('h40)
	) name2109 (
		\g1834_reg/NET0131 ,
		\g1840_reg/NET0131 ,
		\g35_pad ,
		_w2884_
	);
	LUT2 #(
		.INIT('h4)
	) name2110 (
		\g1844_reg/NET0131 ,
		\g35_pad ,
		_w2885_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2111 (
		_w1502_,
		_w1504_,
		_w2884_,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name2112 (
		_w2883_,
		_w2886_,
		_w2887_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2113 (
		\g1848_reg/NET0131 ,
		\g35_pad ,
		_w1502_,
		_w1504_,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name2114 (
		\g1844_reg/NET0131 ,
		\g35_pad ,
		_w2889_
	);
	LUT2 #(
		.INIT('hd)
	) name2115 (
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT3 #(
		.INIT('hfd)
	) name2116 (
		\g35_pad ,
		_w1549_,
		_w1551_,
		_w2891_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2117 (
		\g1950_reg/NET0131 ,
		\g35_pad ,
		_w1549_,
		_w1551_,
		_w2892_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		\g1955_reg/NET0131 ,
		\g35_pad ,
		_w2893_
	);
	LUT3 #(
		.INIT('h10)
	) name2119 (
		_w1549_,
		_w1551_,
		_w2893_,
		_w2894_
	);
	LUT2 #(
		.INIT('he)
	) name2120 (
		_w2892_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name2121 (
		\g1974_reg/NET0131 ,
		\g35_pad ,
		_w2896_
	);
	LUT2 #(
		.INIT('h2)
	) name2122 (
		\g1968_reg/NET0131 ,
		\g1974_reg/NET0131 ,
		_w2897_
	);
	LUT4 #(
		.INIT('h010f)
	) name2123 (
		_w1549_,
		_w1551_,
		_w2896_,
		_w2897_,
		_w2898_
	);
	LUT3 #(
		.INIT('h40)
	) name2124 (
		\g1968_reg/NET0131 ,
		\g1974_reg/NET0131 ,
		\g35_pad ,
		_w2899_
	);
	LUT2 #(
		.INIT('h4)
	) name2125 (
		\g1978_reg/NET0131 ,
		\g35_pad ,
		_w2900_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2126 (
		_w1549_,
		_w1551_,
		_w2899_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		_w2898_,
		_w2901_,
		_w2902_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2128 (
		\g1982_reg/NET0131 ,
		\g35_pad ,
		_w1549_,
		_w1551_,
		_w2903_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		\g1978_reg/NET0131 ,
		\g35_pad ,
		_w2904_
	);
	LUT2 #(
		.INIT('hd)
	) name2130 (
		_w2903_,
		_w2904_,
		_w2905_
	);
	LUT3 #(
		.INIT('hfd)
	) name2131 (
		\g35_pad ,
		_w1596_,
		_w1598_,
		_w2906_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2132 (
		\g2084_reg/NET0131 ,
		\g35_pad ,
		_w1596_,
		_w1598_,
		_w2907_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		\g2089_reg/NET0131 ,
		\g35_pad ,
		_w2908_
	);
	LUT3 #(
		.INIT('h10)
	) name2134 (
		_w1596_,
		_w1598_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('he)
	) name2135 (
		_w2907_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		\g2108_reg/NET0131 ,
		\g35_pad ,
		_w2911_
	);
	LUT2 #(
		.INIT('h2)
	) name2137 (
		\g2102_reg/NET0131 ,
		\g2108_reg/NET0131 ,
		_w2912_
	);
	LUT4 #(
		.INIT('h010f)
	) name2138 (
		_w1596_,
		_w1598_,
		_w2911_,
		_w2912_,
		_w2913_
	);
	LUT3 #(
		.INIT('h40)
	) name2139 (
		\g2102_reg/NET0131 ,
		\g2108_reg/NET0131 ,
		\g35_pad ,
		_w2914_
	);
	LUT2 #(
		.INIT('h4)
	) name2140 (
		\g2112_reg/NET0131 ,
		\g35_pad ,
		_w2915_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2141 (
		_w1596_,
		_w1598_,
		_w2914_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		_w2913_,
		_w2916_,
		_w2917_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2143 (
		\g2116_reg/NET0131 ,
		\g35_pad ,
		_w1596_,
		_w1598_,
		_w2918_
	);
	LUT2 #(
		.INIT('h2)
	) name2144 (
		\g2112_reg/NET0131 ,
		\g35_pad ,
		_w2919_
	);
	LUT2 #(
		.INIT('hd)
	) name2145 (
		_w2918_,
		_w2919_,
		_w2920_
	);
	LUT3 #(
		.INIT('hfd)
	) name2146 (
		\g35_pad ,
		_w1276_,
		_w1278_,
		_w2921_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2147 (
		\g2241_reg/NET0131 ,
		\g35_pad ,
		_w1276_,
		_w1278_,
		_w2922_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		\g2246_reg/NET0131 ,
		\g35_pad ,
		_w2923_
	);
	LUT3 #(
		.INIT('h10)
	) name2149 (
		_w1276_,
		_w1278_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('he)
	) name2150 (
		_w2922_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		\g2265_reg/NET0131 ,
		\g35_pad ,
		_w2926_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		\g2259_reg/NET0131 ,
		\g2265_reg/NET0131 ,
		_w2927_
	);
	LUT4 #(
		.INIT('h010f)
	) name2153 (
		_w1276_,
		_w1278_,
		_w2926_,
		_w2927_,
		_w2928_
	);
	LUT3 #(
		.INIT('h40)
	) name2154 (
		\g2259_reg/NET0131 ,
		\g2265_reg/NET0131 ,
		\g35_pad ,
		_w2929_
	);
	LUT2 #(
		.INIT('h4)
	) name2155 (
		\g2269_reg/NET0131 ,
		\g35_pad ,
		_w2930_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2156 (
		_w1276_,
		_w1278_,
		_w2929_,
		_w2930_,
		_w2931_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		_w2928_,
		_w2931_,
		_w2932_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2158 (
		\g2273_reg/NET0131 ,
		\g35_pad ,
		_w1276_,
		_w1278_,
		_w2933_
	);
	LUT2 #(
		.INIT('h2)
	) name2159 (
		\g2269_reg/NET0131 ,
		\g35_pad ,
		_w2934_
	);
	LUT2 #(
		.INIT('hd)
	) name2160 (
		_w2933_,
		_w2934_,
		_w2935_
	);
	LUT3 #(
		.INIT('hfd)
	) name2161 (
		\g35_pad ,
		_w1323_,
		_w1325_,
		_w2936_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2162 (
		\g2375_reg/NET0131 ,
		\g35_pad ,
		_w1323_,
		_w1325_,
		_w2937_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		\g2380_reg/NET0131 ,
		\g35_pad ,
		_w2938_
	);
	LUT3 #(
		.INIT('h10)
	) name2164 (
		_w1323_,
		_w1325_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('he)
	) name2165 (
		_w2937_,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h1)
	) name2166 (
		\g2399_reg/NET0131 ,
		\g35_pad ,
		_w2941_
	);
	LUT2 #(
		.INIT('h2)
	) name2167 (
		\g2393_reg/NET0131 ,
		\g2399_reg/NET0131 ,
		_w2942_
	);
	LUT4 #(
		.INIT('h010f)
	) name2168 (
		_w1323_,
		_w1325_,
		_w2941_,
		_w2942_,
		_w2943_
	);
	LUT3 #(
		.INIT('h40)
	) name2169 (
		\g2393_reg/NET0131 ,
		\g2399_reg/NET0131 ,
		\g35_pad ,
		_w2944_
	);
	LUT2 #(
		.INIT('h4)
	) name2170 (
		\g2403_reg/NET0131 ,
		\g35_pad ,
		_w2945_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2171 (
		_w1323_,
		_w1325_,
		_w2944_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h8)
	) name2172 (
		_w2943_,
		_w2946_,
		_w2947_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2173 (
		\g2407_reg/NET0131 ,
		\g35_pad ,
		_w1323_,
		_w1325_,
		_w2948_
	);
	LUT2 #(
		.INIT('h2)
	) name2174 (
		\g2403_reg/NET0131 ,
		\g35_pad ,
		_w2949_
	);
	LUT2 #(
		.INIT('hd)
	) name2175 (
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT3 #(
		.INIT('hfd)
	) name2176 (
		\g35_pad ,
		_w1373_,
		_w1375_,
		_w2951_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2177 (
		\g2509_reg/NET0131 ,
		\g35_pad ,
		_w1373_,
		_w1375_,
		_w2952_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		\g2514_reg/NET0131 ,
		\g35_pad ,
		_w2953_
	);
	LUT3 #(
		.INIT('h10)
	) name2179 (
		_w1373_,
		_w1375_,
		_w2953_,
		_w2954_
	);
	LUT2 #(
		.INIT('he)
	) name2180 (
		_w2952_,
		_w2954_,
		_w2955_
	);
	LUT2 #(
		.INIT('h1)
	) name2181 (
		\g2533_reg/NET0131 ,
		\g35_pad ,
		_w2956_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		\g2527_reg/NET0131 ,
		\g2533_reg/NET0131 ,
		_w2957_
	);
	LUT4 #(
		.INIT('h010f)
	) name2183 (
		_w1373_,
		_w1375_,
		_w2956_,
		_w2957_,
		_w2958_
	);
	LUT3 #(
		.INIT('h40)
	) name2184 (
		\g2527_reg/NET0131 ,
		\g2533_reg/NET0131 ,
		\g35_pad ,
		_w2959_
	);
	LUT2 #(
		.INIT('h4)
	) name2185 (
		\g2537_reg/NET0131 ,
		\g35_pad ,
		_w2960_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2186 (
		_w1373_,
		_w1375_,
		_w2959_,
		_w2960_,
		_w2961_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		_w2958_,
		_w2961_,
		_w2962_
	);
	LUT4 #(
		.INIT('hbbb7)
	) name2188 (
		\g2541_reg/NET0131 ,
		\g35_pad ,
		_w1373_,
		_w1375_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name2189 (
		\g2537_reg/NET0131 ,
		\g35_pad ,
		_w2964_
	);
	LUT2 #(
		.INIT('hd)
	) name2190 (
		_w2963_,
		_w2964_,
		_w2965_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2191 (
		\g2643_reg/NET0131 ,
		\g35_pad ,
		_w1420_,
		_w1422_,
		_w2966_
	);
	LUT2 #(
		.INIT('h8)
	) name2192 (
		\g2648_reg/NET0131 ,
		\g35_pad ,
		_w2967_
	);
	LUT3 #(
		.INIT('h10)
	) name2193 (
		_w1420_,
		_w1422_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('he)
	) name2194 (
		_w2966_,
		_w2968_,
		_w2969_
	);
	LUT3 #(
		.INIT('h15)
	) name2195 (
		\g1636_reg/NET0131 ,
		_w802_,
		_w1633_,
		_w2970_
	);
	LUT2 #(
		.INIT('h4)
	) name2196 (
		\g1636_reg/NET0131 ,
		\g17291_pad ,
		_w2971_
	);
	LUT3 #(
		.INIT('h70)
	) name2197 (
		_w1210_,
		_w1635_,
		_w2971_,
		_w2972_
	);
	LUT3 #(
		.INIT('h01)
	) name2198 (
		\g1592_reg/NET0131 ,
		_w2970_,
		_w2972_,
		_w2973_
	);
	LUT3 #(
		.INIT('h2a)
	) name2199 (
		\g1668_reg/NET0131 ,
		_w802_,
		_w1633_,
		_w2974_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		\g1668_reg/NET0131 ,
		\g17291_pad ,
		_w2975_
	);
	LUT3 #(
		.INIT('h70)
	) name2201 (
		_w1210_,
		_w1635_,
		_w2975_,
		_w2976_
	);
	LUT3 #(
		.INIT('h02)
	) name2202 (
		\g35_pad ,
		_w2974_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h4)
	) name2203 (
		_w2973_,
		_w2977_,
		_w2978_
	);
	LUT4 #(
		.INIT('h2000)
	) name2204 (
		\g1002_reg/NET0131 ,
		\g1008_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1036_reg/NET0131 ,
		_w2979_
	);
	LUT3 #(
		.INIT('h20)
	) name2205 (
		_w1971_,
		_w1972_,
		_w2979_,
		_w2980_
	);
	LUT3 #(
		.INIT('h28)
	) name2206 (
		\g1046_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w2981_
	);
	LUT3 #(
		.INIT('h04)
	) name2207 (
		_w1972_,
		_w2565_,
		_w2981_,
		_w2982_
	);
	LUT4 #(
		.INIT('h8a22)
	) name2208 (
		\g969_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w2983_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2209 (
		\g35_pad ,
		_w2980_,
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h2)
	) name2210 (
		\g2763_reg/NET0131 ,
		\g35_pad ,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w1908_,
		_w2985_,
		_w2986_
	);
	LUT3 #(
		.INIT('h54)
	) name2212 (
		\g1632_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w2987_
	);
	LUT3 #(
		.INIT('h31)
	) name2213 (
		\g2763_reg/NET0131 ,
		\g2767_reg/NET0131 ,
		\g35_pad ,
		_w2988_
	);
	LUT3 #(
		.INIT('hb0)
	) name2214 (
		_w1910_,
		_w2987_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		_w2986_,
		_w2989_,
		_w2990_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		\g2767_reg/NET0131 ,
		\g35_pad ,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name2217 (
		_w1908_,
		_w2991_,
		_w2992_
	);
	LUT3 #(
		.INIT('h54)
	) name2218 (
		\g1768_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w2993_
	);
	LUT3 #(
		.INIT('h31)
	) name2219 (
		\g2767_reg/NET0131 ,
		\g2779_reg/NET0131 ,
		\g35_pad ,
		_w2994_
	);
	LUT3 #(
		.INIT('hb0)
	) name2220 (
		_w1910_,
		_w2993_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h1)
	) name2221 (
		_w2992_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('h2)
	) name2222 (
		\g2779_reg/NET0131 ,
		\g35_pad ,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name2223 (
		_w1908_,
		_w2997_,
		_w2998_
	);
	LUT3 #(
		.INIT('h54)
	) name2224 (
		\g1902_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w2999_
	);
	LUT3 #(
		.INIT('h31)
	) name2225 (
		\g2779_reg/NET0131 ,
		\g2791_reg/NET0131 ,
		\g35_pad ,
		_w3000_
	);
	LUT3 #(
		.INIT('hb0)
	) name2226 (
		_w1910_,
		_w2999_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		_w2998_,
		_w3001_,
		_w3002_
	);
	LUT2 #(
		.INIT('h2)
	) name2228 (
		\g2791_reg/NET0131 ,
		\g35_pad ,
		_w3003_
	);
	LUT2 #(
		.INIT('h1)
	) name2229 (
		_w1908_,
		_w3003_,
		_w3004_
	);
	LUT3 #(
		.INIT('h54)
	) name2230 (
		\g2036_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w3005_
	);
	LUT3 #(
		.INIT('h31)
	) name2231 (
		\g2791_reg/NET0131 ,
		\g2795_reg/NET0131 ,
		\g35_pad ,
		_w3006_
	);
	LUT3 #(
		.INIT('hb0)
	) name2232 (
		_w1910_,
		_w3005_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w3004_,
		_w3007_,
		_w3008_
	);
	LUT2 #(
		.INIT('h2)
	) name2234 (
		\g2799_reg/NET0131 ,
		\g35_pad ,
		_w3009_
	);
	LUT2 #(
		.INIT('h1)
	) name2235 (
		_w1908_,
		_w3009_,
		_w3010_
	);
	LUT3 #(
		.INIT('h54)
	) name2236 (
		\g2327_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w3011_
	);
	LUT3 #(
		.INIT('h31)
	) name2237 (
		\g2799_reg/NET0131 ,
		\g2811_reg/NET0131 ,
		\g35_pad ,
		_w3012_
	);
	LUT3 #(
		.INIT('hb0)
	) name2238 (
		_w1910_,
		_w3011_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w3010_,
		_w3013_,
		_w3014_
	);
	LUT3 #(
		.INIT('h15)
	) name2240 (
		\g1002_reg/NET0131 ,
		_w1971_,
		_w2565_,
		_w3015_
	);
	LUT2 #(
		.INIT('h8)
	) name2241 (
		\g1018_reg/NET0131 ,
		\g35_pad ,
		_w3016_
	);
	LUT4 #(
		.INIT('hea00)
	) name2242 (
		_w1972_,
		_w2564_,
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT3 #(
		.INIT('h54)
	) name2243 (
		\g1018_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w3018_
	);
	LUT3 #(
		.INIT('h70)
	) name2244 (
		_w1971_,
		_w2565_,
		_w3018_,
		_w3019_
	);
	LUT4 #(
		.INIT('ha222)
	) name2245 (
		\g1002_reg/NET0131 ,
		\g35_pad ,
		_w2564_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('he)
	) name2246 (
		_w3017_,
		_w3020_,
		_w3021_
	);
	LUT3 #(
		.INIT('h28)
	) name2247 (
		\g35_pad ,
		\g4793_reg/NET0131 ,
		_w1981_,
		_w3022_
	);
	LUT3 #(
		.INIT('h15)
	) name2248 (
		\g168_reg/NET0131 ,
		\g174_reg/NET0131 ,
		\g182_reg/NET0131 ,
		_w3023_
	);
	LUT3 #(
		.INIT('he0)
	) name2249 (
		\g174_reg/NET0131 ,
		\g182_reg/NET0131 ,
		\g35_pad ,
		_w3024_
	);
	LUT3 #(
		.INIT('h20)
	) name2250 (
		_w1689_,
		_w3023_,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h2)
	) name2251 (
		\g1189_reg/NET0131 ,
		\g35_pad ,
		_w3026_
	);
	LUT3 #(
		.INIT('h20)
	) name2252 (
		\g1070_reg/NET0131 ,
		_w2745_,
		_w2746_,
		_w3027_
	);
	LUT4 #(
		.INIT('hfb73)
	) name2253 (
		\g1193_reg/NET0131 ,
		\g35_pad ,
		_w2737_,
		_w3027_,
		_w3028_
	);
	LUT2 #(
		.INIT('hb)
	) name2254 (
		_w3026_,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('h2)
	) name2255 (
		\g29218_pad ,
		\g35_pad ,
		_w3030_
	);
	LUT4 #(
		.INIT('h0001)
	) name2256 (
		\g4311_reg/NET0131 ,
		\g4322_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		\g4358_reg/NET0131 ,
		_w3031_
	);
	LUT4 #(
		.INIT('h0200)
	) name2257 (
		\g35_pad ,
		\g4332_reg/NET0131 ,
		\g4340_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3032_
	);
	LUT3 #(
		.INIT('hea)
	) name2258 (
		_w3030_,
		_w3031_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h2)
	) name2259 (
		\g2811_reg/NET0131 ,
		\g35_pad ,
		_w3034_
	);
	LUT2 #(
		.INIT('h1)
	) name2260 (
		_w1908_,
		_w3034_,
		_w3035_
	);
	LUT3 #(
		.INIT('h54)
	) name2261 (
		\g2461_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w3036_
	);
	LUT3 #(
		.INIT('h31)
	) name2262 (
		\g2811_reg/NET0131 ,
		\g2823_reg/NET0131 ,
		\g35_pad ,
		_w3037_
	);
	LUT3 #(
		.INIT('hb0)
	) name2263 (
		_w1910_,
		_w3036_,
		_w3037_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name2264 (
		_w3035_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h2)
	) name2265 (
		\g2823_reg/NET0131 ,
		\g35_pad ,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		_w1908_,
		_w3040_,
		_w3041_
	);
	LUT3 #(
		.INIT('h54)
	) name2267 (
		\g2595_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w3042_
	);
	LUT3 #(
		.INIT('h31)
	) name2268 (
		\g2823_reg/NET0131 ,
		\g2827_reg/NET0131 ,
		\g35_pad ,
		_w3043_
	);
	LUT3 #(
		.INIT('hb0)
	) name2269 (
		_w1910_,
		_w3042_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name2270 (
		_w3041_,
		_w3044_,
		_w3045_
	);
	LUT2 #(
		.INIT('h1)
	) name2271 (
		\g2927_reg/NET0131 ,
		\g35_pad ,
		_w3046_
	);
	LUT4 #(
		.INIT('h0004)
	) name2272 (
		\g2941_reg/NET0131 ,
		\g35_pad ,
		\g4072_reg/NET0131 ,
		\g4153_reg/NET0131 ,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w3046_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h2)
	) name2274 (
		\g1193_reg/NET0131 ,
		\g35_pad ,
		_w3049_
	);
	LUT3 #(
		.INIT('h40)
	) name2275 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g7916_pad ,
		_w3050_
	);
	LUT3 #(
		.INIT('h45)
	) name2276 (
		\g1199_reg/NET0131 ,
		_w2745_,
		_w3050_,
		_w3051_
	);
	LUT4 #(
		.INIT('h00e0)
	) name2277 (
		_w2737_,
		_w2738_,
		_w2747_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('he)
	) name2278 (
		_w3049_,
		_w3052_,
		_w3053_
	);
	LUT4 #(
		.INIT('h3aca)
	) name2279 (
		\g3329_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g35_pad ,
		_w2770_,
		_w3054_
	);
	LUT4 #(
		.INIT('h7ddd)
	) name2280 (
		\g35_pad ,
		\g843_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w1824_,
		_w3055_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		\g837_reg/NET0131 ,
		_w3055_,
		_w3056_
	);
	LUT4 #(
		.INIT('h1555)
	) name2282 (
		\g4584_reg/NET0131 ,
		_w1791_,
		_w1793_,
		_w1794_,
		_w3057_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2283 (
		\g35_pad ,
		_w1791_,
		_w1793_,
		_w1799_,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name2284 (
		\g35_pad ,
		\g4332_reg/NET0131 ,
		_w3059_
	);
	LUT3 #(
		.INIT('hf4)
	) name2285 (
		_w3057_,
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2286 (
		\g2856_reg/NET0131 ,
		\g35_pad ,
		_w788_,
		_w789_,
		_w3061_
	);
	LUT4 #(
		.INIT('hd111)
	) name2287 (
		\g2848_reg/NET0131 ,
		\g35_pad ,
		_w785_,
		_w786_,
		_w3062_
	);
	LUT2 #(
		.INIT('hb)
	) name2288 (
		_w3061_,
		_w3062_,
		_w3063_
	);
	LUT3 #(
		.INIT('h1b)
	) name2289 (
		\g5037_reg/NET0131 ,
		_w2707_,
		_w2709_,
		_w3064_
	);
	LUT2 #(
		.INIT('h2)
	) name2290 (
		\g35_pad ,
		\g5041_reg/NET0131 ,
		_w3065_
	);
	LUT2 #(
		.INIT('h8)
	) name2291 (
		\g35_pad ,
		\g5041_reg/NET0131 ,
		_w3066_
	);
	LUT3 #(
		.INIT('h10)
	) name2292 (
		_w2712_,
		_w2754_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h4)
	) name2293 (
		\g35_pad ,
		\g5037_reg/NET0131 ,
		_w3068_
	);
	LUT4 #(
		.INIT('hffe4)
	) name2294 (
		_w3064_,
		_w3065_,
		_w3067_,
		_w3068_,
		_w3069_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2295 (
		\g2882_reg/NET0131 ,
		\g35_pad ,
		_w795_,
		_w796_,
		_w3070_
	);
	LUT4 #(
		.INIT('hd111)
	) name2296 (
		\g2898_reg/NET0131 ,
		\g35_pad ,
		_w792_,
		_w793_,
		_w3071_
	);
	LUT2 #(
		.INIT('hb)
	) name2297 (
		_w3070_,
		_w3071_,
		_w3072_
	);
	LUT4 #(
		.INIT('h8000)
	) name2298 (
		\g16624_pad ,
		\g3338_reg/NET0131 ,
		\g5297_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w3073_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		\g4646_reg/NET0131 ,
		_w3073_,
		_w3074_
	);
	LUT3 #(
		.INIT('h75)
	) name2300 (
		\g35_pad ,
		_w826_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		\g4646_reg/NET0131 ,
		\g5128_reg/NET0131 ,
		_w3076_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		_w3073_,
		_w3076_,
		_w3077_
	);
	LUT4 #(
		.INIT('h1311)
	) name2303 (
		\g35_pad ,
		\g5134_reg/NET0131 ,
		_w826_,
		_w3077_,
		_w3078_
	);
	LUT3 #(
		.INIT('h20)
	) name2304 (
		\g4646_reg/NET0131 ,
		\g5128_reg/NET0131 ,
		\g5134_reg/NET0131 ,
		_w3079_
	);
	LUT2 #(
		.INIT('h8)
	) name2305 (
		_w3073_,
		_w3079_,
		_w3080_
	);
	LUT3 #(
		.INIT('h20)
	) name2306 (
		\g35_pad ,
		_w826_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h2)
	) name2307 (
		\g35_pad ,
		\g5138_reg/NET0131 ,
		_w3082_
	);
	LUT3 #(
		.INIT('hb0)
	) name2308 (
		_w826_,
		_w3074_,
		_w3082_,
		_w3083_
	);
	LUT3 #(
		.INIT('h01)
	) name2309 (
		_w3078_,
		_w3081_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('h7d77)
	) name2310 (
		\g35_pad ,
		\g5142_reg/NET0131 ,
		_w826_,
		_w3074_,
		_w3085_
	);
	LUT2 #(
		.INIT('h4)
	) name2311 (
		\g35_pad ,
		\g5138_reg/NET0131 ,
		_w3086_
	);
	LUT2 #(
		.INIT('hd)
	) name2312 (
		_w3085_,
		_w3086_,
		_w3087_
	);
	LUT3 #(
		.INIT('h80)
	) name2313 (
		\g1772_reg/NET0131 ,
		_w802_,
		_w1208_,
		_w3088_
	);
	LUT4 #(
		.INIT('h0203)
	) name2314 (
		_w1219_,
		_w1510_,
		_w1512_,
		_w3088_,
		_w3089_
	);
	LUT3 #(
		.INIT('h2e)
	) name2315 (
		\g1779_reg/NET0131 ,
		\g35_pad ,
		_w3089_,
		_w3090_
	);
	LUT3 #(
		.INIT('h80)
	) name2316 (
		\g35_pad ,
		_w802_,
		_w1208_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name2317 (
		\g1802_reg/NET0131 ,
		\g35_pad ,
		_w3092_
	);
	LUT3 #(
		.INIT('h80)
	) name2318 (
		_w802_,
		_w1208_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name2319 (
		\g1772_reg/NET0131 ,
		_w1219_,
		_w3091_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		\g3352_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		_w3095_
	);
	LUT3 #(
		.INIT('h80)
	) name2321 (
		\g16624_pad ,
		\g3288_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w3096_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT3 #(
		.INIT('h75)
	) name2323 (
		\g35_pad ,
		_w1852_,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		\g3125_reg/NET0131 ,
		\g35_pad ,
		_w3099_
	);
	LUT2 #(
		.INIT('h2)
	) name2325 (
		\g3119_reg/NET0131 ,
		\g3125_reg/NET0131 ,
		_w3100_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2326 (
		_w1852_,
		_w3097_,
		_w3099_,
		_w3100_,
		_w3101_
	);
	LUT3 #(
		.INIT('h40)
	) name2327 (
		\g3119_reg/NET0131 ,
		\g3125_reg/NET0131 ,
		\g35_pad ,
		_w3102_
	);
	LUT2 #(
		.INIT('h4)
	) name2328 (
		\g3129_reg/NET0131 ,
		\g35_pad ,
		_w3103_
	);
	LUT4 #(
		.INIT('h04bf)
	) name2329 (
		_w1852_,
		_w3097_,
		_w3102_,
		_w3103_,
		_w3104_
	);
	LUT2 #(
		.INIT('h8)
	) name2330 (
		_w3101_,
		_w3104_,
		_w3105_
	);
	LUT3 #(
		.INIT('h01)
	) name2331 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3167_reg/NET0131 ,
		_w3106_
	);
	LUT2 #(
		.INIT('h1)
	) name2332 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name2333 (
		\g4180_reg/NET0131 ,
		\g4284_reg/NET0131 ,
		_w3108_
	);
	LUT4 #(
		.INIT('h1101)
	) name2334 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		\g4180_reg/NET0131 ,
		\g4284_reg/NET0131 ,
		_w3109_
	);
	LUT3 #(
		.INIT('h80)
	) name2335 (
		\g35_pad ,
		_w3106_,
		_w3109_,
		_w3110_
	);
	LUT2 #(
		.INIT('h8)
	) name2336 (
		\g3187_reg/NET0131 ,
		\g35_pad ,
		_w3111_
	);
	LUT3 #(
		.INIT('h70)
	) name2337 (
		_w3106_,
		_w3107_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		\g3179_reg/NET0131 ,
		\g35_pad ,
		_w3113_
	);
	LUT3 #(
		.INIT('hfe)
	) name2339 (
		_w3110_,
		_w3112_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3115_
	);
	LUT4 #(
		.INIT('h2202)
	) name2341 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		\g4180_reg/NET0131 ,
		\g4284_reg/NET0131 ,
		_w3116_
	);
	LUT3 #(
		.INIT('h80)
	) name2342 (
		\g35_pad ,
		_w3106_,
		_w3116_,
		_w3117_
	);
	LUT2 #(
		.INIT('h8)
	) name2343 (
		\g3191_reg/NET0131 ,
		\g35_pad ,
		_w3118_
	);
	LUT3 #(
		.INIT('h70)
	) name2344 (
		_w3106_,
		_w3115_,
		_w3118_,
		_w3119_
	);
	LUT2 #(
		.INIT('h2)
	) name2345 (
		\g3195_reg/NET0131 ,
		\g35_pad ,
		_w3120_
	);
	LUT3 #(
		.INIT('hfe)
	) name2346 (
		_w3117_,
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT4 #(
		.INIT('h7b77)
	) name2347 (
		\g3133_reg/NET0131 ,
		\g35_pad ,
		_w1852_,
		_w3097_,
		_w3122_
	);
	LUT2 #(
		.INIT('h2)
	) name2348 (
		\g3129_reg/NET0131 ,
		\g35_pad ,
		_w3123_
	);
	LUT2 #(
		.INIT('hd)
	) name2349 (
		_w3122_,
		_w3123_,
		_w3124_
	);
	LUT3 #(
		.INIT('h02)
	) name2350 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3125_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		\g3195_reg/NET0131 ,
		\g35_pad ,
		_w3126_
	);
	LUT3 #(
		.INIT('ha2)
	) name2352 (
		\g35_pad ,
		\g4180_reg/NET0131 ,
		\g4284_reg/NET0131 ,
		_w3127_
	);
	LUT2 #(
		.INIT('h2)
	) name2353 (
		\g3247_reg/NET0131 ,
		\g35_pad ,
		_w3128_
	);
	LUT4 #(
		.INIT('hffe4)
	) name2354 (
		_w3125_,
		_w3126_,
		_w3127_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h4)
	) name2355 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3130_
	);
	LUT4 #(
		.INIT('h4404)
	) name2356 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		\g4180_reg/NET0131 ,
		\g4284_reg/NET0131 ,
		_w3131_
	);
	LUT3 #(
		.INIT('h80)
	) name2357 (
		\g35_pad ,
		_w3106_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		\g3199_reg/NET0131 ,
		\g35_pad ,
		_w3133_
	);
	LUT3 #(
		.INIT('h70)
	) name2359 (
		_w3106_,
		_w3130_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h2)
	) name2360 (
		\g3203_reg/NET0131 ,
		\g35_pad ,
		_w3135_
	);
	LUT3 #(
		.INIT('hfe)
	) name2361 (
		_w3132_,
		_w3134_,
		_w3135_,
		_w3136_
	);
	LUT3 #(
		.INIT('h08)
	) name2362 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3137_
	);
	LUT2 #(
		.INIT('h8)
	) name2363 (
		\g3203_reg/NET0131 ,
		\g35_pad ,
		_w3138_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		\g3251_reg/NET0131 ,
		\g35_pad ,
		_w3139_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2365 (
		_w3127_,
		_w3137_,
		_w3138_,
		_w3139_,
		_w3140_
	);
	LUT4 #(
		.INIT('h0002)
	) name2366 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3141_
	);
	LUT2 #(
		.INIT('h8)
	) name2367 (
		\g3215_reg/NET0131 ,
		\g35_pad ,
		_w3142_
	);
	LUT2 #(
		.INIT('h2)
	) name2368 (
		\g3187_reg/NET0131 ,
		\g35_pad ,
		_w3143_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2369 (
		_w3127_,
		_w3141_,
		_w3142_,
		_w3143_,
		_w3144_
	);
	LUT4 #(
		.INIT('h0020)
	) name2370 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3145_
	);
	LUT2 #(
		.INIT('h8)
	) name2371 (
		\g3219_reg/NET0131 ,
		\g35_pad ,
		_w3146_
	);
	LUT2 #(
		.INIT('h2)
	) name2372 (
		\g3191_reg/NET0131 ,
		\g35_pad ,
		_w3147_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2373 (
		_w3127_,
		_w3145_,
		_w3146_,
		_w3147_,
		_w3148_
	);
	LUT4 #(
		.INIT('h0200)
	) name2374 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3149_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		\g3223_reg/NET0131 ,
		\g35_pad ,
		_w3150_
	);
	LUT2 #(
		.INIT('h2)
	) name2376 (
		\g3199_reg/NET0131 ,
		\g35_pad ,
		_w3151_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2377 (
		_w3127_,
		_w3149_,
		_w3150_,
		_w3151_,
		_w3152_
	);
	LUT4 #(
		.INIT('h0004)
	) name2378 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3153_
	);
	LUT2 #(
		.INIT('h8)
	) name2379 (
		\g3231_reg/NET0131 ,
		\g35_pad ,
		_w3154_
	);
	LUT2 #(
		.INIT('h2)
	) name2380 (
		\g3215_reg/NET0131 ,
		\g35_pad ,
		_w3155_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2381 (
		_w3127_,
		_w3153_,
		_w3154_,
		_w3155_,
		_w3156_
	);
	LUT4 #(
		.INIT('h0040)
	) name2382 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name2383 (
		\g3235_reg/NET0131 ,
		\g35_pad ,
		_w3158_
	);
	LUT2 #(
		.INIT('h2)
	) name2384 (
		\g3219_reg/NET0131 ,
		\g35_pad ,
		_w3159_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2385 (
		_w3127_,
		_w3157_,
		_w3158_,
		_w3159_,
		_w3160_
	);
	LUT4 #(
		.INIT('h0400)
	) name2386 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3161_
	);
	LUT2 #(
		.INIT('h8)
	) name2387 (
		\g3239_reg/NET0131 ,
		\g35_pad ,
		_w3162_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		\g3223_reg/NET0131 ,
		\g35_pad ,
		_w3163_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2389 (
		_w3127_,
		_w3161_,
		_w3162_,
		_w3163_,
		_w3164_
	);
	LUT4 #(
		.INIT('h0008)
	) name2390 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3165_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		\g3247_reg/NET0131 ,
		\g35_pad ,
		_w3166_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		\g3231_reg/NET0131 ,
		\g35_pad ,
		_w3167_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2393 (
		_w3127_,
		_w3165_,
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h0080)
	) name2394 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3169_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		\g3251_reg/NET0131 ,
		\g35_pad ,
		_w3170_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		\g3235_reg/NET0131 ,
		\g35_pad ,
		_w3171_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2397 (
		_w3127_,
		_w3169_,
		_w3170_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3173_
	);
	LUT4 #(
		.INIT('h8808)
	) name2399 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		\g4180_reg/NET0131 ,
		\g4284_reg/NET0131 ,
		_w3174_
	);
	LUT3 #(
		.INIT('h80)
	) name2400 (
		\g35_pad ,
		_w3106_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		\g3207_reg/NET0131 ,
		\g35_pad ,
		_w3176_
	);
	LUT3 #(
		.INIT('h70)
	) name2402 (
		_w3106_,
		_w3173_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h2)
	) name2403 (
		\g3211_reg/NET0131 ,
		\g35_pad ,
		_w3178_
	);
	LUT3 #(
		.INIT('hfe)
	) name2404 (
		_w3175_,
		_w3177_,
		_w3178_,
		_w3179_
	);
	LUT3 #(
		.INIT('h20)
	) name2405 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3180_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		\g3211_reg/NET0131 ,
		\g35_pad ,
		_w3181_
	);
	LUT2 #(
		.INIT('h2)
	) name2407 (
		\g3255_reg/NET0131 ,
		\g35_pad ,
		_w3182_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2408 (
		_w3127_,
		_w3180_,
		_w3181_,
		_w3182_,
		_w3183_
	);
	LUT4 #(
		.INIT('h2000)
	) name2409 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3184_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		\g3227_reg/NET0131 ,
		\g35_pad ,
		_w3185_
	);
	LUT2 #(
		.INIT('h2)
	) name2411 (
		\g3207_reg/NET0131 ,
		\g35_pad ,
		_w3186_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2412 (
		_w3127_,
		_w3184_,
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT4 #(
		.INIT('h4000)
	) name2413 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3188_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		\g3243_reg/NET0131 ,
		\g35_pad ,
		_w3189_
	);
	LUT2 #(
		.INIT('h2)
	) name2415 (
		\g3227_reg/NET0131 ,
		\g35_pad ,
		_w3190_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2416 (
		_w3127_,
		_w3188_,
		_w3189_,
		_w3190_,
		_w3191_
	);
	LUT4 #(
		.INIT('h0800)
	) name2417 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3192_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		\g3255_reg/NET0131 ,
		\g35_pad ,
		_w3193_
	);
	LUT2 #(
		.INIT('h2)
	) name2419 (
		\g3239_reg/NET0131 ,
		\g35_pad ,
		_w3194_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2420 (
		_w3127_,
		_w3192_,
		_w3193_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h8000)
	) name2421 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3196_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		\g3259_reg/NET0131 ,
		\g35_pad ,
		_w3197_
	);
	LUT2 #(
		.INIT('h2)
	) name2423 (
		\g3243_reg/NET0131 ,
		\g35_pad ,
		_w3198_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2424 (
		_w3127_,
		_w3196_,
		_w3197_,
		_w3198_,
		_w3199_
	);
	LUT3 #(
		.INIT('h80)
	) name2425 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w3200_
	);
	LUT2 #(
		.INIT('h8)
	) name2426 (
		\g3263_reg/NET0131 ,
		\g35_pad ,
		_w3201_
	);
	LUT2 #(
		.INIT('h2)
	) name2427 (
		\g3259_reg/NET0131 ,
		\g35_pad ,
		_w3202_
	);
	LUT4 #(
		.INIT('hffb8)
	) name2428 (
		_w3127_,
		_w3200_,
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT3 #(
		.INIT('h80)
	) name2429 (
		\g1906_reg/NET0131 ,
		_w802_,
		_w1225_,
		_w3204_
	);
	LUT4 #(
		.INIT('h0203)
	) name2430 (
		_w1235_,
		_w1566_,
		_w1568_,
		_w3204_,
		_w3205_
	);
	LUT3 #(
		.INIT('h2e)
	) name2431 (
		\g1913_reg/NET0131 ,
		\g35_pad ,
		_w3205_,
		_w3206_
	);
	LUT3 #(
		.INIT('h80)
	) name2432 (
		\g35_pad ,
		_w802_,
		_w1225_,
		_w3207_
	);
	LUT2 #(
		.INIT('h8)
	) name2433 (
		\g1936_reg/NET0131 ,
		\g35_pad ,
		_w3208_
	);
	LUT3 #(
		.INIT('h80)
	) name2434 (
		_w802_,
		_w1225_,
		_w3208_,
		_w3209_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name2435 (
		\g1906_reg/NET0131 ,
		_w1235_,
		_w3207_,
		_w3209_,
		_w3210_
	);
	LUT4 #(
		.INIT('hd555)
	) name2436 (
		\g35_pad ,
		_w879_,
		_w880_,
		_w1752_,
		_w3211_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		\g29213_pad ,
		\g35_pad ,
		_w3212_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		\g5084_reg/NET0131 ,
		\g5092_reg/NET0131 ,
		_w3213_
	);
	LUT4 #(
		.INIT('h3cf4)
	) name2439 (
		\g35_pad ,
		\g5097_reg/NET0131 ,
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT4 #(
		.INIT('h8000)
	) name2440 (
		\g16624_pad ,
		\g3338_reg/NET0131 ,
		\g3639_reg/NET0131 ,
		\g3703_reg/NET0131 ,
		_w3215_
	);
	LUT2 #(
		.INIT('h8)
	) name2441 (
		\g3470_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name2442 (
		_w3215_,
		_w3216_,
		_w3217_
	);
	LUT4 #(
		.INIT('h1511)
	) name2443 (
		\g3476_reg/NET0131 ,
		\g35_pad ,
		_w1873_,
		_w3217_,
		_w3218_
	);
	LUT3 #(
		.INIT('h40)
	) name2444 (
		\g3470_reg/NET0131 ,
		\g3476_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		_w3219_
	);
	LUT2 #(
		.INIT('h8)
	) name2445 (
		_w3215_,
		_w3219_,
		_w3220_
	);
	LUT3 #(
		.INIT('h20)
	) name2446 (
		\g35_pad ,
		_w1873_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h8)
	) name2447 (
		\g4681_reg/NET0131 ,
		_w3215_,
		_w3222_
	);
	LUT2 #(
		.INIT('h4)
	) name2448 (
		\g3480_reg/NET0131 ,
		\g35_pad ,
		_w3223_
	);
	LUT3 #(
		.INIT('hb0)
	) name2449 (
		_w1873_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT3 #(
		.INIT('h01)
	) name2450 (
		_w3218_,
		_w3221_,
		_w3224_,
		_w3225_
	);
	LUT4 #(
		.INIT('h7b77)
	) name2451 (
		\g3484_reg/NET0131 ,
		\g35_pad ,
		_w1873_,
		_w3222_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name2452 (
		\g3480_reg/NET0131 ,
		\g35_pad ,
		_w3227_
	);
	LUT2 #(
		.INIT('hd)
	) name2453 (
		_w3226_,
		_w3227_,
		_w3228_
	);
	LUT3 #(
		.INIT('h80)
	) name2454 (
		\g2040_reg/NET0131 ,
		_w802_,
		_w1241_,
		_w3229_
	);
	LUT4 #(
		.INIT('h0203)
	) name2455 (
		_w1251_,
		_w1586_,
		_w1588_,
		_w3229_,
		_w3230_
	);
	LUT3 #(
		.INIT('h2e)
	) name2456 (
		\g2047_reg/NET0131 ,
		\g35_pad ,
		_w3230_,
		_w3231_
	);
	LUT3 #(
		.INIT('h80)
	) name2457 (
		\g35_pad ,
		_w802_,
		_w1241_,
		_w3232_
	);
	LUT2 #(
		.INIT('hb)
	) name2458 (
		_w1251_,
		_w3232_,
		_w3233_
	);
	LUT3 #(
		.INIT('h80)
	) name2459 (
		\g16624_pad ,
		\g3338_reg/NET0131 ,
		\g3990_reg/NET0131 ,
		_w3234_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		\g4054_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w3235_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		_w3234_,
		_w3235_,
		_w3236_
	);
	LUT3 #(
		.INIT('h75)
	) name2462 (
		\g35_pad ,
		_w866_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		\g35_pad ,
		\g3827_reg/NET0131 ,
		_w3238_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		\g3821_reg/NET0131 ,
		\g3827_reg/NET0131 ,
		_w3239_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2465 (
		_w866_,
		_w3236_,
		_w3238_,
		_w3239_,
		_w3240_
	);
	LUT3 #(
		.INIT('h20)
	) name2466 (
		\g35_pad ,
		\g3821_reg/NET0131 ,
		\g3827_reg/NET0131 ,
		_w3241_
	);
	LUT2 #(
		.INIT('h2)
	) name2467 (
		\g35_pad ,
		\g3831_reg/NET0131 ,
		_w3242_
	);
	LUT4 #(
		.INIT('h04bf)
	) name2468 (
		_w866_,
		_w3236_,
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		_w3240_,
		_w3243_,
		_w3244_
	);
	LUT4 #(
		.INIT('h7d77)
	) name2470 (
		\g35_pad ,
		\g3835_reg/NET0131 ,
		_w866_,
		_w3236_,
		_w3245_
	);
	LUT2 #(
		.INIT('h4)
	) name2471 (
		\g35_pad ,
		\g3831_reg/NET0131 ,
		_w3246_
	);
	LUT2 #(
		.INIT('hd)
	) name2472 (
		_w3245_,
		_w3246_,
		_w3247_
	);
	LUT3 #(
		.INIT('h80)
	) name2473 (
		\g2197_reg/NET0131 ,
		_w800_,
		_w1127_,
		_w3248_
	);
	LUT4 #(
		.INIT('h0203)
	) name2474 (
		_w1138_,
		_w1293_,
		_w1295_,
		_w3248_,
		_w3249_
	);
	LUT3 #(
		.INIT('h2e)
	) name2475 (
		\g2204_reg/NET0131 ,
		\g35_pad ,
		_w3249_,
		_w3250_
	);
	LUT3 #(
		.INIT('h80)
	) name2476 (
		\g35_pad ,
		_w800_,
		_w1127_,
		_w3251_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		\g2227_reg/NET0131 ,
		\g35_pad ,
		_w3252_
	);
	LUT3 #(
		.INIT('h80)
	) name2478 (
		_w800_,
		_w1127_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name2479 (
		\g2197_reg/NET0131 ,
		_w1138_,
		_w3251_,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h8)
	) name2480 (
		\g4258_reg/NET0131 ,
		\g4264_reg/NET0131 ,
		_w3255_
	);
	LUT4 #(
		.INIT('h6ce4)
	) name2481 (
		\g35_pad ,
		\g4269_reg/NET0131 ,
		\g4273_reg/NET0131 ,
		_w3255_,
		_w3256_
	);
	LUT4 #(
		.INIT('h6ce4)
	) name2482 (
		\g35_pad ,
		\g4340_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		_w1791_,
		_w3257_
	);
	LUT3 #(
		.INIT('h80)
	) name2483 (
		\g2331_reg/NET0131 ,
		_w800_,
		_w1144_,
		_w3258_
	);
	LUT4 #(
		.INIT('h0203)
	) name2484 (
		_w1154_,
		_w1340_,
		_w1342_,
		_w3258_,
		_w3259_
	);
	LUT3 #(
		.INIT('h2e)
	) name2485 (
		\g2338_reg/NET0131 ,
		\g35_pad ,
		_w3259_,
		_w3260_
	);
	LUT3 #(
		.INIT('h80)
	) name2486 (
		\g35_pad ,
		_w800_,
		_w1144_,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		\g2361_reg/NET0131 ,
		\g35_pad ,
		_w3262_
	);
	LUT3 #(
		.INIT('h80)
	) name2488 (
		_w800_,
		_w1144_,
		_w3262_,
		_w3263_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name2489 (
		\g2331_reg/NET0131 ,
		_w1154_,
		_w3261_,
		_w3263_,
		_w3264_
	);
	LUT4 #(
		.INIT('h0020)
	) name2490 (
		\g14125_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w3265_
	);
	LUT4 #(
		.INIT('h33f7)
	) name2491 (
		\g239_reg/NET0131 ,
		\g35_pad ,
		_w2656_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h2)
	) name2492 (
		\g262_reg/NET0131 ,
		\g35_pad ,
		_w3267_
	);
	LUT2 #(
		.INIT('hd)
	) name2493 (
		_w3266_,
		_w3267_,
		_w3268_
	);
	LUT3 #(
		.INIT('h75)
	) name2494 (
		\g35_pad ,
		_w1873_,
		_w3222_,
		_w3269_
	);
	LUT3 #(
		.INIT('h80)
	) name2495 (
		\g2465_reg/NET0131 ,
		_w800_,
		_w1160_,
		_w3270_
	);
	LUT4 #(
		.INIT('h0203)
	) name2496 (
		_w1170_,
		_w1390_,
		_w1392_,
		_w3270_,
		_w3271_
	);
	LUT3 #(
		.INIT('h2e)
	) name2497 (
		\g2472_reg/NET0131 ,
		\g35_pad ,
		_w3271_,
		_w3272_
	);
	LUT3 #(
		.INIT('h80)
	) name2498 (
		\g35_pad ,
		_w800_,
		_w1160_,
		_w3273_
	);
	LUT2 #(
		.INIT('h8)
	) name2499 (
		\g2495_reg/NET0131 ,
		\g35_pad ,
		_w3274_
	);
	LUT3 #(
		.INIT('h80)
	) name2500 (
		_w800_,
		_w1160_,
		_w3274_,
		_w3275_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name2501 (
		\g2465_reg/NET0131 ,
		_w1170_,
		_w3273_,
		_w3275_,
		_w3276_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		\g35_pad ,
		\g528_reg/NET0131 ,
		_w3277_
	);
	LUT3 #(
		.INIT('ha2)
	) name2503 (
		\g35_pad ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3278_
	);
	LUT4 #(
		.INIT('h2202)
	) name2504 (
		\g35_pad ,
		\g482_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3279_
	);
	LUT4 #(
		.INIT('hf700)
	) name2505 (
		_w1688_,
		_w2615_,
		_w2616_,
		_w3279_,
		_w3280_
	);
	LUT4 #(
		.INIT('h8808)
	) name2506 (
		\g35_pad ,
		\g482_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3281_
	);
	LUT4 #(
		.INIT('h0800)
	) name2507 (
		_w1688_,
		_w2615_,
		_w2616_,
		_w3281_,
		_w3282_
	);
	LUT3 #(
		.INIT('h01)
	) name2508 (
		_w3277_,
		_w3280_,
		_w3282_,
		_w3283_
	);
	LUT3 #(
		.INIT('h2a)
	) name2509 (
		\g17291_pad ,
		_w1210_,
		_w1635_,
		_w3284_
	);
	LUT3 #(
		.INIT('h80)
	) name2510 (
		\g1636_reg/NET0131 ,
		_w802_,
		_w1633_,
		_w3285_
	);
	LUT4 #(
		.INIT('h1011)
	) name2511 (
		_w1634_,
		_w1637_,
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT3 #(
		.INIT('h2e)
	) name2512 (
		\g1644_reg/NET0131 ,
		\g35_pad ,
		_w3286_,
		_w3287_
	);
	LUT3 #(
		.INIT('h15)
	) name2513 (
		\g2555_reg/NET0131 ,
		_w800_,
		_w1176_,
		_w3288_
	);
	LUT2 #(
		.INIT('h2)
	) name2514 (
		\g1430_reg/NET0131 ,
		\g2555_reg/NET0131 ,
		_w3289_
	);
	LUT3 #(
		.INIT('h70)
	) name2515 (
		_w1129_,
		_w1178_,
		_w3289_,
		_w3290_
	);
	LUT3 #(
		.INIT('h40)
	) name2516 (
		\g2599_reg/NET0131 ,
		_w800_,
		_w1176_,
		_w3291_
	);
	LUT4 #(
		.INIT('h0203)
	) name2517 (
		_w1186_,
		_w3288_,
		_w3290_,
		_w3291_,
		_w3292_
	);
	LUT3 #(
		.INIT('he2)
	) name2518 (
		\g2606_reg/NET0131 ,
		\g35_pad ,
		_w3292_,
		_w3293_
	);
	LUT3 #(
		.INIT('h80)
	) name2519 (
		\g35_pad ,
		_w802_,
		_w1633_,
		_w3294_
	);
	LUT2 #(
		.INIT('h8)
	) name2520 (
		\g1668_reg/NET0131 ,
		\g35_pad ,
		_w3295_
	);
	LUT3 #(
		.INIT('h80)
	) name2521 (
		_w802_,
		_w1633_,
		_w3295_,
		_w3296_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name2522 (
		\g1636_reg/NET0131 ,
		_w3284_,
		_w3294_,
		_w3296_,
		_w3297_
	);
	LUT3 #(
		.INIT('h80)
	) name2523 (
		\g35_pad ,
		_w800_,
		_w1176_,
		_w3298_
	);
	LUT2 #(
		.INIT('hb)
	) name2524 (
		_w1186_,
		_w3298_,
		_w3299_
	);
	LUT3 #(
		.INIT('h78)
	) name2525 (
		\g3111_reg/NET0131 ,
		\g35_pad ,
		\g5115_reg/NET0131 ,
		_w3300_
	);
	LUT4 #(
		.INIT('h0075)
	) name2526 (
		\g35_pad ,
		_w826_,
		_w3074_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h2)
	) name2527 (
		\g35_pad ,
		\g5124_reg/NET0131 ,
		_w3302_
	);
	LUT3 #(
		.INIT('hb0)
	) name2528 (
		_w826_,
		_w3074_,
		_w3302_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		_w3301_,
		_w3303_,
		_w3304_
	);
	LUT3 #(
		.INIT('h6a)
	) name2530 (
		\g3106_reg/NET0131 ,
		\g3111_reg/NET0131 ,
		\g35_pad ,
		_w3305_
	);
	LUT4 #(
		.INIT('h0075)
	) name2531 (
		\g35_pad ,
		_w1852_,
		_w3097_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h4)
	) name2532 (
		\g3115_reg/NET0131 ,
		\g35_pad ,
		_w3307_
	);
	LUT3 #(
		.INIT('hb0)
	) name2533 (
		_w1852_,
		_w3097_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w3306_,
		_w3308_,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name2535 (
		\g336_reg/NET0131 ,
		\g35_pad ,
		_w3310_
	);
	LUT4 #(
		.INIT('h4500)
	) name2536 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		\g324_reg/NET0131 ,
		\g35_pad ,
		_w3311_
	);
	LUT2 #(
		.INIT('h1)
	) name2537 (
		_w3310_,
		_w3311_,
		_w3312_
	);
	LUT4 #(
		.INIT('h4000)
	) name2538 (
		\g661_reg/NET0131 ,
		_w1824_,
		_w2022_,
		_w2023_,
		_w3313_
	);
	LUT2 #(
		.INIT('h4)
	) name2539 (
		\g29212_pad ,
		\g35_pad ,
		_w3314_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2540 (
		_w1824_,
		_w2022_,
		_w2023_,
		_w3314_,
		_w3315_
	);
	LUT4 #(
		.INIT('h00ce)
	) name2541 (
		\g35_pad ,
		\g728_reg/NET0131 ,
		_w3313_,
		_w3315_,
		_w3316_
	);
	LUT3 #(
		.INIT('h6c)
	) name2542 (
		\g3111_reg/NET0131 ,
		\g3457_reg/NET0131 ,
		\g35_pad ,
		_w3317_
	);
	LUT4 #(
		.INIT('h0075)
	) name2543 (
		\g35_pad ,
		_w1873_,
		_w3222_,
		_w3317_,
		_w3318_
	);
	LUT2 #(
		.INIT('h4)
	) name2544 (
		\g3466_reg/NET0131 ,
		\g35_pad ,
		_w3319_
	);
	LUT3 #(
		.INIT('hb0)
	) name2545 (
		_w1873_,
		_w3222_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h1)
	) name2546 (
		_w3318_,
		_w3320_,
		_w3321_
	);
	LUT3 #(
		.INIT('h78)
	) name2547 (
		\g3111_reg/NET0131 ,
		\g35_pad ,
		\g3808_reg/NET0131 ,
		_w3322_
	);
	LUT4 #(
		.INIT('h0075)
	) name2548 (
		\g35_pad ,
		_w866_,
		_w3236_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h2)
	) name2549 (
		\g35_pad ,
		\g3817_reg/NET0131 ,
		_w3324_
	);
	LUT3 #(
		.INIT('hb0)
	) name2550 (
		_w866_,
		_w3236_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h1)
	) name2551 (
		_w3323_,
		_w3325_,
		_w3326_
	);
	LUT4 #(
		.INIT('h67ef)
	) name2552 (
		\g5037_reg/NET0131 ,
		\g5041_reg/NET0131 ,
		_w2707_,
		_w2709_,
		_w3327_
	);
	LUT2 #(
		.INIT('h4)
	) name2553 (
		\g35_pad ,
		\g5041_reg/NET0131 ,
		_w3328_
	);
	LUT3 #(
		.INIT('hb1)
	) name2554 (
		\g35_pad ,
		\g5041_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		_w3329_
	);
	LUT2 #(
		.INIT('h8)
	) name2555 (
		\g35_pad ,
		\g5046_reg/NET0131 ,
		_w3330_
	);
	LUT3 #(
		.INIT('h23)
	) name2556 (
		_w2712_,
		_w3328_,
		_w3330_,
		_w3331_
	);
	LUT3 #(
		.INIT('h1b)
	) name2557 (
		_w3327_,
		_w3329_,
		_w3331_,
		_w3332_
	);
	LUT3 #(
		.INIT('hd0)
	) name2558 (
		\g35_pad ,
		\g5069_reg/NET0131 ,
		\g5073_reg/NET0131 ,
		_w3333_
	);
	LUT4 #(
		.INIT('h0c84)
	) name2559 (
		\g3147_reg/NET0131 ,
		\g35_pad ,
		_w3108_,
		_w3200_,
		_w3334_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		\g35_pad ,
		\g969_reg/NET0131 ,
		_w3335_
	);
	LUT4 #(
		.INIT('h2088)
	) name2561 (
		\g969_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w3336_
	);
	LUT2 #(
		.INIT('h1)
	) name2562 (
		_w3335_,
		_w3336_,
		_w3337_
	);
	LUT4 #(
		.INIT('h8880)
	) name2563 (
		\g1018_reg/NET0131 ,
		\g1030_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w3338_
	);
	LUT4 #(
		.INIT('h2088)
	) name2564 (
		\g1046_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w3339_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		\g1008_reg/NET0131 ,
		\g35_pad ,
		_w3340_
	);
	LUT3 #(
		.INIT('h10)
	) name2566 (
		_w3338_,
		_w3339_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('hd)
	) name2567 (
		_w3337_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		\g4646_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w3343_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2569 (
		_w823_,
		_w824_,
		_w825_,
		_w3343_,
		_w3344_
	);
	LUT2 #(
		.INIT('h8)
	) name2570 (
		\g35_pad ,
		\g5297_reg/NET0131 ,
		_w3345_
	);
	LUT4 #(
		.INIT('h0f88)
	) name2571 (
		\g5357_reg/NET0131 ,
		_w2087_,
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		\g3288_reg/NET0131 ,
		\g35_pad ,
		_w3347_
	);
	LUT3 #(
		.INIT('h78)
	) name2573 (
		\g3352_reg/NET0131 ,
		_w1941_,
		_w3347_,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name2574 (
		\g3703_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		_w3349_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2575 (
		_w824_,
		_w825_,
		_w1858_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h8)
	) name2576 (
		\g35_pad ,
		\g3639_reg/NET0131 ,
		_w3351_
	);
	LUT4 #(
		.INIT('h0f88)
	) name2577 (
		\g3703_reg/NET0131 ,
		_w2012_,
		_w3350_,
		_w3351_,
		_w3352_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2578 (
		_w824_,
		_w825_,
		_w865_,
		_w3235_,
		_w3353_
	);
	LUT2 #(
		.INIT('h8)
	) name2579 (
		\g35_pad ,
		\g3990_reg/NET0131 ,
		_w3354_
	);
	LUT4 #(
		.INIT('h0f88)
	) name2580 (
		\g4054_reg/NET0131 ,
		_w876_,
		_w3353_,
		_w3354_,
		_w3355_
	);
	LUT3 #(
		.INIT('h3a)
	) name2581 (
		\g3338_reg/NET0131 ,
		\g3347_reg/NET0131 ,
		\g35_pad ,
		_w3356_
	);
	LUT3 #(
		.INIT('h70)
	) name2582 (
		_w2769_,
		_w2770_,
		_w3356_,
		_w3357_
	);
	LUT2 #(
		.INIT('h4)
	) name2583 (
		\g35_pad ,
		\g812_reg/NET0131 ,
		_w3358_
	);
	LUT4 #(
		.INIT('h9b11)
	) name2584 (
		\g35_pad ,
		\g812_reg/NET0131 ,
		\g837_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w3359_
	);
	LUT4 #(
		.INIT('h00f6)
	) name2585 (
		\g817_reg/NET0131 ,
		_w1824_,
		_w3358_,
		_w3359_,
		_w3360_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		\g2864_reg/NET0131 ,
		\g35_pad ,
		_w3361_
	);
	LUT2 #(
		.INIT('h4)
	) name2587 (
		\g2898_reg/NET0131 ,
		\g35_pad ,
		_w3362_
	);
	LUT4 #(
		.INIT('h070f)
	) name2588 (
		_w912_,
		_w913_,
		_w3361_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('hfad8)
	) name2589 (
		\g35_pad ,
		\g4072_reg/NET0131 ,
		\g4172_reg/NET0131 ,
		\g4176_reg/NET0131 ,
		_w3364_
	);
	LUT4 #(
		.INIT('h0080)
	) name2590 (
		\g3050_reg/NET0131 ,
		\g5016_reg/NET0131 ,
		\g5029_reg/NET0131 ,
		\g5033_reg/NET0131 ,
		_w3365_
	);
	LUT3 #(
		.INIT('ha8)
	) name2591 (
		\g35_pad ,
		_w3365_,
		_w2707_,
		_w3366_
	);
	LUT3 #(
		.INIT('h02)
	) name2592 (
		\g5033_reg/NET0131 ,
		_w2712_,
		_w2754_,
		_w3367_
	);
	LUT4 #(
		.INIT('h77cf)
	) name2593 (
		\g3050_reg/NET0131 ,
		\g5016_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		\g5029_reg/NET0131 ,
		_w3368_
	);
	LUT2 #(
		.INIT('h8)
	) name2594 (
		\g35_pad ,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('h4)
	) name2595 (
		\g35_pad ,
		\g5029_reg/NET0131 ,
		_w3370_
	);
	LUT4 #(
		.INIT('hffea)
	) name2596 (
		_w3366_,
		_w3367_,
		_w3369_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h1)
	) name2597 (
		\g4646_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w3372_
	);
	LUT4 #(
		.INIT('h0002)
	) name2598 (
		\g4698_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w3373_
	);
	LUT4 #(
		.INIT('h070f)
	) name2599 (
		_w824_,
		_w825_,
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT4 #(
		.INIT('h2e22)
	) name2600 (
		\g3347_reg/NET0131 ,
		\g35_pad ,
		_w3344_,
		_w3374_,
		_w3375_
	);
	LUT3 #(
		.INIT('h10)
	) name2601 (
		\g499_reg/NET0131 ,
		\g518_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w3376_
	);
	LUT4 #(
		.INIT('h0004)
	) name2602 (
		\g411_reg/NET0131 ,
		\g417_reg/NET0131 ,
		\g424_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w3377_
	);
	LUT4 #(
		.INIT('h8880)
	) name2603 (
		\g681_reg/NET0131 ,
		_w1752_,
		_w3376_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h8)
	) name2604 (
		\g35_pad ,
		\g650_reg/NET0131 ,
		_w3379_
	);
	LUT4 #(
		.INIT('h5700)
	) name2605 (
		_w1752_,
		_w3376_,
		_w3377_,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('hffe4)
	) name2606 (
		\g35_pad ,
		\g699_reg/NET0131 ,
		_w3378_,
		_w3380_,
		_w3381_
	);
	LUT4 #(
		.INIT('hddd5)
	) name2607 (
		\g35_pad ,
		_w1752_,
		_w3376_,
		_w3377_,
		_w3382_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		\g3352_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		_w3383_
	);
	LUT4 #(
		.INIT('h1000)
	) name2609 (
		\g3352_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4743_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w3384_
	);
	LUT4 #(
		.INIT('h070f)
	) name2610 (
		_w824_,
		_w825_,
		_w3383_,
		_w3384_,
		_w3385_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2611 (
		_w824_,
		_w825_,
		_w1837_,
		_w3095_,
		_w3386_
	);
	LUT4 #(
		.INIT('h22e2)
	) name2612 (
		\g3347_reg/NET0131 ,
		\g35_pad ,
		_w3385_,
		_w3386_,
		_w3387_
	);
	LUT4 #(
		.INIT('hff48)
	) name2613 (
		\g1236_reg/NET0131 ,
		\g35_pad ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w3388_
	);
	LUT4 #(
		.INIT('h4800)
	) name2614 (
		\g1236_reg/NET0131 ,
		\g35_pad ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w3389_
	);
	LUT4 #(
		.INIT('h8aba)
	) name2615 (
		\g990_reg/NET0131 ,
		_w1971_,
		_w1973_,
		_w3389_,
		_w3390_
	);
	LUT2 #(
		.INIT('h8)
	) name2616 (
		_w3388_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h1)
	) name2617 (
		\g3703_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		_w3392_
	);
	LUT4 #(
		.INIT('h0040)
	) name2618 (
		\g3703_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4754_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w3393_
	);
	LUT4 #(
		.INIT('h070f)
	) name2619 (
		_w824_,
		_w825_,
		_w3392_,
		_w3393_,
		_w3394_
	);
	LUT4 #(
		.INIT('h2e22)
	) name2620 (
		\g3347_reg/NET0131 ,
		\g35_pad ,
		_w3350_,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		\g4054_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w3396_
	);
	LUT4 #(
		.INIT('h4000)
	) name2622 (
		\g4054_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4765_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w3397_
	);
	LUT4 #(
		.INIT('h070f)
	) name2623 (
		_w824_,
		_w825_,
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT4 #(
		.INIT('h2e22)
	) name2624 (
		\g3347_reg/NET0131 ,
		\g35_pad ,
		_w3353_,
		_w3398_,
		_w3399_
	);
	LUT4 #(
		.INIT('hacf0)
	) name2625 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		\g324_reg/NET0131 ,
		\g35_pad ,
		_w3400_
	);
	LUT4 #(
		.INIT('h0020)
	) name2626 (
		\g14096_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w3401_
	);
	LUT4 #(
		.INIT('h33f7)
	) name2627 (
		\g262_reg/NET0131 ,
		\g35_pad ,
		_w2656_,
		_w3401_,
		_w3402_
	);
	LUT2 #(
		.INIT('h2)
	) name2628 (
		\g232_reg/NET0131 ,
		\g35_pad ,
		_w3403_
	);
	LUT2 #(
		.INIT('hd)
	) name2629 (
		_w3402_,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h2)
	) name2630 (
		\g1008_reg/NET0131 ,
		\g35_pad ,
		_w3405_
	);
	LUT4 #(
		.INIT('hccc8)
	) name2631 (
		\g1002_reg/NET0131 ,
		\g35_pad ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w3406_
	);
	LUT4 #(
		.INIT('hea00)
	) name2632 (
		_w1972_,
		_w2564_,
		_w3015_,
		_w3406_,
		_w3407_
	);
	LUT2 #(
		.INIT('he)
	) name2633 (
		_w3405_,
		_w3407_,
		_w3408_
	);
	LUT4 #(
		.INIT('h4440)
	) name2634 (
		\g446_reg/NET0131 ,
		_w1752_,
		_w3376_,
		_w3377_,
		_w3409_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		\g35_pad ,
		\g645_reg/NET0131 ,
		_w3410_
	);
	LUT4 #(
		.INIT('h8880)
	) name2636 (
		\g35_pad ,
		_w1752_,
		_w3376_,
		_w3377_,
		_w3411_
	);
	LUT3 #(
		.INIT('h54)
	) name2637 (
		_w3409_,
		_w3410_,
		_w3411_,
		_w3412_
	);
	LUT2 #(
		.INIT('h4)
	) name2638 (
		\g35_pad ,
		\g546_reg/NET0131 ,
		_w3413_
	);
	LUT2 #(
		.INIT('h4)
	) name2639 (
		\g542_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w3414_
	);
	LUT3 #(
		.INIT('hce)
	) name2640 (
		_w2625_,
		_w3413_,
		_w3414_,
		_w3415_
	);
	LUT3 #(
		.INIT('h4e)
	) name2641 (
		\g13895_pad ,
		\g16718_pad ,
		\g3303_reg/NET0131 ,
		_w3416_
	);
	LUT4 #(
		.INIT('h0100)
	) name2642 (
		\g13039_pad ,
		\g16603_pad ,
		\g16624_pad ,
		\g35_pad ,
		_w3417_
	);
	LUT2 #(
		.INIT('h4)
	) name2643 (
		_w3416_,
		_w3417_,
		_w3418_
	);
	LUT3 #(
		.INIT('h08)
	) name2644 (
		\g4621_reg/NET0131 ,
		\g4633_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w3419_
	);
	LUT3 #(
		.INIT('h2a)
	) name2645 (
		\g35_pad ,
		_w1793_,
		_w3419_,
		_w3420_
	);
	LUT3 #(
		.INIT('h20)
	) name2646 (
		_w929_,
		_w933_,
		_w934_,
		_w3421_
	);
	LUT2 #(
		.INIT('h2)
	) name2647 (
		\g35_pad ,
		_w930_,
		_w3422_
	);
	LUT3 #(
		.INIT('hba)
	) name2648 (
		_w3420_,
		_w3421_,
		_w3422_,
		_w3423_
	);
	LUT3 #(
		.INIT('h78)
	) name2649 (
		\g35_pad ,
		\g4653_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w3424_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		\g4621_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w3425_
	);
	LUT3 #(
		.INIT('h80)
	) name2651 (
		\g4621_reg/NET0131 ,
		\g4628_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w3426_
	);
	LUT2 #(
		.INIT('h2)
	) name2652 (
		\g35_pad ,
		\g4643_reg/NET0131 ,
		_w3427_
	);
	LUT3 #(
		.INIT('h08)
	) name2653 (
		\g35_pad ,
		\g4633_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name2654 (
		_w3426_,
		_w3428_,
		_w3429_
	);
	LUT4 #(
		.INIT('h0020)
	) name2655 (
		\g4621_reg/NET0131 ,
		\g4633_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3430_
	);
	LUT3 #(
		.INIT('hc4)
	) name2656 (
		\g35_pad ,
		\g4628_reg/NET0131 ,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('he)
	) name2657 (
		_w3429_,
		_w3431_,
		_w3432_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name2658 (
		\g2878_reg/NET0131 ,
		\g2886_reg/NET0131 ,
		\g2946_reg/NET0131 ,
		\g35_pad ,
		_w3433_
	);
	LUT3 #(
		.INIT('h80)
	) name2659 (
		\g35_pad ,
		\g4180_reg/NET0131 ,
		\g8786_pad ,
		_w3434_
	);
	LUT3 #(
		.INIT('h01)
	) name2660 (
		\g8787_pad ,
		\g8788_pad ,
		\g8789_pad ,
		_w3435_
	);
	LUT4 #(
		.INIT('h0001)
	) name2661 (
		\g11447_pad ,
		\g8783_pad ,
		\g8784_pad ,
		\g8785_pad ,
		_w3436_
	);
	LUT3 #(
		.INIT('h02)
	) name2662 (
		\g35_pad ,
		\g4180_reg/NET0131 ,
		\g8786_pad ,
		_w3437_
	);
	LUT4 #(
		.INIT('h4055)
	) name2663 (
		_w3434_,
		_w3435_,
		_w3436_,
		_w3437_,
		_w3438_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		\g2946_reg/NET0131 ,
		\g35_pad ,
		_w3439_
	);
	LUT2 #(
		.INIT('h2)
	) name2665 (
		_w3438_,
		_w3439_,
		_w3440_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		\g35_pad ,
		\g4145_reg/NET0131 ,
		_w3441_
	);
	LUT3 #(
		.INIT('h01)
	) name2667 (
		\g4076_reg/NET0131 ,
		\g4082_reg/NET0131 ,
		\g4141_reg/NET0131 ,
		_w3442_
	);
	LUT3 #(
		.INIT('h10)
	) name2668 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		\g4145_reg/NET0131 ,
		_w3443_
	);
	LUT4 #(
		.INIT('h1333)
	) name2669 (
		_w830_,
		_w3441_,
		_w3442_,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h8)
	) name2670 (
		\g35_pad ,
		\g4112_reg/NET0131 ,
		_w3445_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2671 (
		_w828_,
		_w830_,
		_w3442_,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('hd)
	) name2672 (
		_w3444_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		\g35_pad ,
		\g4369_reg/NET0131 ,
		_w3448_
	);
	LUT4 #(
		.INIT('h2022)
	) name2674 (
		\g35_pad ,
		\g4459_reg/NET0131 ,
		\g4462_reg/NET0131 ,
		\g4473_reg/NET0131 ,
		_w3449_
	);
	LUT2 #(
		.INIT('h1)
	) name2675 (
		_w3448_,
		_w3449_,
		_w3450_
	);
	LUT2 #(
		.INIT('h4)
	) name2676 (
		\g35_pad ,
		\g518_reg/NET0131 ,
		_w3451_
	);
	LUT4 #(
		.INIT('h8808)
	) name2677 (
		\g35_pad ,
		\g528_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3452_
	);
	LUT3 #(
		.INIT('h70)
	) name2678 (
		_w1688_,
		_w2615_,
		_w3452_,
		_w3453_
	);
	LUT4 #(
		.INIT('h8000)
	) name2679 (
		_w1688_,
		_w2615_,
		_w2616_,
		_w3278_,
		_w3454_
	);
	LUT3 #(
		.INIT('hfe)
	) name2680 (
		_w3451_,
		_w3453_,
		_w3454_,
		_w3455_
	);
	LUT3 #(
		.INIT('h08)
	) name2681 (
		\g35_pad ,
		\g699_reg/NET0131 ,
		_w1824_,
		_w3456_
	);
	LUT2 #(
		.INIT('h4)
	) name2682 (
		\g35_pad ,
		\g681_reg/NET0131 ,
		_w3457_
	);
	LUT3 #(
		.INIT('hfe)
	) name2683 (
		_w3411_,
		_w3456_,
		_w3457_,
		_w3458_
	);
	LUT4 #(
		.INIT('h0080)
	) name2684 (
		\g723_reg/NET0131 ,
		\g817_reg/NET0131 ,
		\g822_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w3459_
	);
	LUT3 #(
		.INIT('h80)
	) name2685 (
		\g35_pad ,
		_w1824_,
		_w3459_,
		_w3460_
	);
	LUT3 #(
		.INIT('h80)
	) name2686 (
		\g812_reg/NET0131 ,
		\g837_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w3461_
	);
	LUT3 #(
		.INIT('h4c)
	) name2687 (
		_w1824_,
		_w2029_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h4)
	) name2688 (
		\g35_pad ,
		\g847_reg/NET0131 ,
		_w3463_
	);
	LUT3 #(
		.INIT('hfe)
	) name2689 (
		_w3460_,
		_w3462_,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('hd)
	) name2690 (
		\g35_pad ,
		_w1824_,
		_w3465_
	);
	LUT4 #(
		.INIT('hf0d8)
	) name2691 (
		\g35_pad ,
		\g847_reg/NET0131 ,
		\g854_reg/NET0131 ,
		_w1824_,
		_w3466_
	);
	LUT2 #(
		.INIT('hd)
	) name2692 (
		\g35_pad ,
		_w1752_,
		_w3467_
	);
	LUT4 #(
		.INIT('h7ad0)
	) name2693 (
		\g35_pad ,
		\g5084_reg/NET0131 ,
		\g5092_reg/NET0131 ,
		\g5097_reg/NET0131 ,
		_w3468_
	);
	LUT4 #(
		.INIT('h78cc)
	) name2694 (
		\g1087_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		\g1221_reg/NET0131 ,
		\g35_pad ,
		_w3469_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		\g182_reg/NET0131 ,
		\g35_pad ,
		_w3470_
	);
	LUT2 #(
		.INIT('h4)
	) name2696 (
		\g35_pad ,
		\g405_reg/NET0131 ,
		_w3471_
	);
	LUT4 #(
		.INIT('hffd8)
	) name2697 (
		_w1752_,
		_w2657_,
		_w3470_,
		_w3471_,
		_w3472_
	);
	LUT2 #(
		.INIT('h4)
	) name2698 (
		\g837_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w3473_
	);
	LUT4 #(
		.INIT('hc444)
	) name2699 (
		\g35_pad ,
		\g703_reg/NET0131 ,
		_w1824_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('h153f)
	) name2700 (
		\g812_reg/NET0131 ,
		\g827_reg/NET0131 ,
		\g832_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w3475_
	);
	LUT2 #(
		.INIT('h8)
	) name2701 (
		\g35_pad ,
		\g837_reg/NET0131 ,
		_w3476_
	);
	LUT3 #(
		.INIT('hd0)
	) name2702 (
		_w1824_,
		_w3475_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('he)
	) name2703 (
		_w3474_,
		_w3477_,
		_w3478_
	);
	LUT4 #(
		.INIT('h0002)
	) name2704 (
		\g4064_reg/NET0131 ,
		\g4087_reg/NET0131 ,
		\g4093_reg/NET0131 ,
		\g4098_reg/NET0131 ,
		_w3479_
	);
	LUT2 #(
		.INIT('h4)
	) name2705 (
		\g4057_reg/NET0131 ,
		\g4145_reg/NET0131 ,
		_w3480_
	);
	LUT4 #(
		.INIT('h8000)
	) name2706 (
		\g35_pad ,
		_w3442_,
		_w3479_,
		_w3480_,
		_w3481_
	);
	LUT2 #(
		.INIT('h8)
	) name2707 (
		\g35_pad ,
		\g4116_reg/NET0131 ,
		_w3482_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2708 (
		\g4057_reg/NET0131 ,
		_w3442_,
		_w3479_,
		_w3482_,
		_w3483_
	);
	LUT2 #(
		.INIT('h4)
	) name2709 (
		\g35_pad ,
		\g4112_reg/NET0131 ,
		_w3484_
	);
	LUT3 #(
		.INIT('hfe)
	) name2710 (
		_w3481_,
		_w3483_,
		_w3484_,
		_w3485_
	);
	LUT2 #(
		.INIT('h2)
	) name2711 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		_w3486_
	);
	LUT3 #(
		.INIT('h20)
	) name2712 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		\g4145_reg/NET0131 ,
		_w3487_
	);
	LUT4 #(
		.INIT('h8000)
	) name2713 (
		\g35_pad ,
		_w830_,
		_w3442_,
		_w3487_,
		_w3488_
	);
	LUT2 #(
		.INIT('h8)
	) name2714 (
		\g35_pad ,
		\g4119_reg/NET0131 ,
		_w3489_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2715 (
		_w830_,
		_w3442_,
		_w3486_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h4)
	) name2716 (
		\g35_pad ,
		\g4116_reg/NET0131 ,
		_w3491_
	);
	LUT3 #(
		.INIT('hfe)
	) name2717 (
		_w3488_,
		_w3490_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h8)
	) name2718 (
		\g4057_reg/NET0131 ,
		\g4145_reg/NET0131 ,
		_w3493_
	);
	LUT4 #(
		.INIT('h8000)
	) name2719 (
		\g35_pad ,
		_w3442_,
		_w3479_,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h8)
	) name2720 (
		\g35_pad ,
		\g4122_reg/NET0131 ,
		_w3495_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2721 (
		\g4057_reg/NET0131 ,
		_w3442_,
		_w3479_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name2722 (
		\g35_pad ,
		\g4119_reg/NET0131 ,
		_w3497_
	);
	LUT3 #(
		.INIT('hfe)
	) name2723 (
		_w3494_,
		_w3496_,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h2)
	) name2724 (
		\g35_pad ,
		\g4258_reg/NET0131 ,
		_w3499_
	);
	LUT4 #(
		.INIT('h7ad0)
	) name2725 (
		\g35_pad ,
		\g4258_reg/NET0131 ,
		\g4264_reg/NET0131 ,
		\g4269_reg/NET0131 ,
		_w3500_
	);
	LUT2 #(
		.INIT('h8)
	) name2726 (
		\g35_pad ,
		\g433_reg/NET0131 ,
		_w3501_
	);
	LUT2 #(
		.INIT('h4)
	) name2727 (
		\g35_pad ,
		\g437_reg/NET0131 ,
		_w3502_
	);
	LUT4 #(
		.INIT('hffd8)
	) name2728 (
		_w1824_,
		_w2811_,
		_w3501_,
		_w3502_,
		_w3503_
	);
	LUT4 #(
		.INIT('h0020)
	) name2729 (
		\g14217_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w3504_
	);
	LUT4 #(
		.INIT('h33f7)
	) name2730 (
		\g232_reg/NET0131 ,
		\g35_pad ,
		_w2656_,
		_w3504_,
		_w3505_
	);
	LUT2 #(
		.INIT('h2)
	) name2731 (
		\g255_reg/NET0131 ,
		\g35_pad ,
		_w3506_
	);
	LUT2 #(
		.INIT('hd)
	) name2732 (
		_w3505_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h8)
	) name2733 (
		\g35_pad ,
		\g460_reg/NET0131 ,
		_w3508_
	);
	LUT2 #(
		.INIT('h2)
	) name2734 (
		\g168_reg/NET0131 ,
		\g35_pad ,
		_w3509_
	);
	LUT4 #(
		.INIT('hffd8)
	) name2735 (
		_w1752_,
		_w2647_,
		_w3508_,
		_w3509_,
		_w3510_
	);
	LUT4 #(
		.INIT('h78cc)
	) name2736 (
		\g1430_reg/NET0131 ,
		\g1548_reg/NET0131 ,
		\g1564_reg/NET0131 ,
		\g35_pad ,
		_w3511_
	);
	LUT2 #(
		.INIT('h8)
	) name2737 (
		\g35_pad ,
		\g475_reg/NET0131 ,
		_w3512_
	);
	LUT2 #(
		.INIT('h4)
	) name2738 (
		\g35_pad ,
		\g424_reg/NET0131 ,
		_w3513_
	);
	LUT4 #(
		.INIT('hffd8)
	) name2739 (
		_w1824_,
		_w2647_,
		_w3512_,
		_w3513_,
		_w3514_
	);
	LUT4 #(
		.INIT('h0020)
	) name2740 (
		\g14201_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w3515_
	);
	LUT4 #(
		.INIT('h33f7)
	) name2741 (
		\g255_reg/NET0131 ,
		\g35_pad ,
		_w2656_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h2)
	) name2742 (
		\g225_reg/NET0131 ,
		\g35_pad ,
		_w3517_
	);
	LUT2 #(
		.INIT('hd)
	) name2743 (
		_w3516_,
		_w3517_,
		_w3518_
	);
	LUT4 #(
		.INIT('h0040)
	) name2744 (
		\g3050_reg/NET0131 ,
		\g35_pad ,
		\g5016_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		_w3519_
	);
	LUT4 #(
		.INIT('h0c08)
	) name2745 (
		\g3050_reg/NET0131 ,
		\g35_pad ,
		\g5016_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		_w3520_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2746 (
		_w2712_,
		_w2754_,
		_w3519_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h4)
	) name2747 (
		\g35_pad ,
		\g5022_reg/NET0131 ,
		_w3522_
	);
	LUT2 #(
		.INIT('hd)
	) name2748 (
		_w3521_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h2)
	) name2749 (
		\g3100_reg/NET0131 ,
		\g35_pad ,
		_w3524_
	);
	LUT3 #(
		.INIT('h45)
	) name2750 (
		\g3050_reg/NET0131 ,
		\g3100_reg/NET0131 ,
		\g5101_reg/NET0131 ,
		_w3525_
	);
	LUT2 #(
		.INIT('h4)
	) name2751 (
		\g3096_reg/NET0131 ,
		\g35_pad ,
		_w3526_
	);
	LUT3 #(
		.INIT('hba)
	) name2752 (
		_w3524_,
		_w3525_,
		_w3526_,
		_w3527_
	);
	LUT3 #(
		.INIT('he0)
	) name2753 (
		\g2932_reg/NET0131 ,
		\g2999_reg/NET0131 ,
		\g35_pad ,
		_w3528_
	);
	LUT4 #(
		.INIT('h8000)
	) name2754 (
		\g1087_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1221_reg/NET0131 ,
		_w3529_
	);
	LUT4 #(
		.INIT('h0100)
	) name2755 (
		\g17291_pad ,
		\g17316_pad ,
		\g17400_pad ,
		\g35_pad ,
		_w3530_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2756 (
		_w1971_,
		_w1973_,
		_w3529_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('he)
	) name2757 (
		\g35_pad ,
		\g4072_reg/NET0131 ,
		_w3532_
	);
	LUT2 #(
		.INIT('h8)
	) name2758 (
		\g35_pad ,
		\g417_reg/NET0131 ,
		_w3533_
	);
	LUT3 #(
		.INIT('hd8)
	) name2759 (
		_w1824_,
		_w2657_,
		_w3533_,
		_w3534_
	);
	LUT4 #(
		.INIT('h0222)
	) name2760 (
		\g35_pad ,
		\g4311_reg/NET0131 ,
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		_w3535_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		\g35_pad ,
		\g4311_reg/NET0131 ,
		_w3536_
	);
	LUT4 #(
		.INIT('hf780)
	) name2762 (
		_w1791_,
		_w1793_,
		_w3535_,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w2707_,
		_w2709_,
		_w3538_
	);
	LUT4 #(
		.INIT('h0008)
	) name2764 (
		\g35_pad ,
		\g5037_reg/NET0131 ,
		_w2712_,
		_w2754_,
		_w3539_
	);
	LUT2 #(
		.INIT('h4)
	) name2765 (
		\g35_pad ,
		\g5033_reg/NET0131 ,
		_w3540_
	);
	LUT2 #(
		.INIT('h2)
	) name2766 (
		\g35_pad ,
		\g5037_reg/NET0131 ,
		_w3541_
	);
	LUT4 #(
		.INIT('h010f)
	) name2767 (
		_w2707_,
		_w2709_,
		_w3540_,
		_w3541_,
		_w3542_
	);
	LUT3 #(
		.INIT('h8f)
	) name2768 (
		_w3538_,
		_w3539_,
		_w3542_,
		_w3543_
	);
	LUT4 #(
		.INIT('h2220)
	) name2769 (
		\g1008_reg/NET0131 ,
		\g1046_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w3544_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2770 (
		\g1041_reg/NET0131 ,
		\g35_pad ,
		_w1971_,
		_w3544_,
		_w3545_
	);
	LUT4 #(
		.INIT('hddd0)
	) name2771 (
		\g1008_reg/NET0131 ,
		\g1041_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w3546_
	);
	LUT2 #(
		.INIT('h8)
	) name2772 (
		\g1046_reg/NET0131 ,
		\g35_pad ,
		_w3547_
	);
	LUT3 #(
		.INIT('hb0)
	) name2773 (
		_w1971_,
		_w3546_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('he)
	) name2774 (
		_w3545_,
		_w3548_,
		_w3549_
	);
	LUT3 #(
		.INIT('h8a)
	) name2775 (
		\g35_pad ,
		\g703_reg/NET0131 ,
		\g854_reg/NET0131 ,
		_w3550_
	);
	LUT2 #(
		.INIT('h2)
	) name2776 (
		\g35_pad ,
		\g392_reg/NET0131 ,
		_w3551_
	);
	LUT2 #(
		.INIT('h1)
	) name2777 (
		\g35_pad ,
		\g401_reg/NET0131 ,
		_w3552_
	);
	LUT4 #(
		.INIT('h0027)
	) name2778 (
		_w1824_,
		_w3550_,
		_w3551_,
		_w3552_,
		_w3553_
	);
	LUT2 #(
		.INIT('h2)
	) name2779 (
		\g1036_reg/NET0131 ,
		\g35_pad ,
		_w3554_
	);
	LUT4 #(
		.INIT('h4511)
	) name2780 (
		\g1041_reg/NET0131 ,
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w3555_
	);
	LUT4 #(
		.INIT('h008a)
	) name2781 (
		\g35_pad ,
		_w1971_,
		_w3546_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('he)
	) name2782 (
		_w3554_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h4)
	) name2783 (
		\g35_pad ,
		\g4358_reg/NET0131 ,
		_w3558_
	);
	LUT4 #(
		.INIT('h0001)
	) name2784 (
		\g4593_reg/NET0131 ,
		\g4601_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		\g4616_reg/NET0131 ,
		_w3559_
	);
	LUT4 #(
		.INIT('h0020)
	) name2785 (
		\g35_pad ,
		\g4332_reg/NET0131 ,
		\g4340_reg/NET0131 ,
		\g4584_reg/NET0131 ,
		_w3560_
	);
	LUT4 #(
		.INIT('h8000)
	) name2786 (
		_w3031_,
		_w3419_,
		_w3559_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('he)
	) name2787 (
		_w3558_,
		_w3561_,
		_w3562_
	);
	LUT4 #(
		.INIT('h7cb0)
	) name2788 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w3563_
	);
	LUT3 #(
		.INIT('h4e)
	) name2789 (
		\g35_pad ,
		\g5069_reg/NET0131 ,
		_w2712_,
		_w3564_
	);
	LUT3 #(
		.INIT('h4e)
	) name2790 (
		\g35_pad ,
		\g4284_reg/NET0131 ,
		\g4291_reg/NET0131 ,
		_w3565_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		\g2902_reg/NET0131 ,
		\g35_pad ,
		_w3566_
	);
	LUT2 #(
		.INIT('h4)
	) name2792 (
		\g2917_reg/NET0131 ,
		\g35_pad ,
		_w3567_
	);
	LUT4 #(
		.INIT('h070f)
	) name2793 (
		_w800_,
		_w802_,
		_w3566_,
		_w3567_,
		_w3568_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		\g29214_pad ,
		\g35_pad ,
		_w3569_
	);
	LUT4 #(
		.INIT('h4000)
	) name2795 (
		\g2848_reg/NET0131 ,
		\g35_pad ,
		_w782_,
		_w783_,
		_w3570_
	);
	LUT2 #(
		.INIT('h1)
	) name2796 (
		_w3569_,
		_w3570_,
		_w3571_
	);
	LUT4 #(
		.INIT('h5515)
	) name2797 (
		\g4340_reg/NET0131 ,
		\g4621_reg/NET0131 ,
		\g4628_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w3572_
	);
	LUT4 #(
		.INIT('h444e)
	) name2798 (
		\g35_pad ,
		\g4643_reg/NET0131 ,
		_w2782_,
		_w3572_,
		_w3573_
	);
	LUT3 #(
		.INIT('hd5)
	) name2799 (
		\g35_pad ,
		_w864_,
		_w1945_,
		_w3574_
	);
	LUT3 #(
		.INIT('hd5)
	) name2800 (
		\g35_pad ,
		_w822_,
		_w1945_,
		_w3575_
	);
	LUT3 #(
		.INIT('hd5)
	) name2801 (
		\g35_pad ,
		_w1836_,
		_w1945_,
		_w3576_
	);
	LUT3 #(
		.INIT('hd5)
	) name2802 (
		\g35_pad ,
		_w1857_,
		_w1945_,
		_w3577_
	);
	LUT4 #(
		.INIT('h2000)
	) name2803 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		\g513_reg/NET0131 ,
		_w3578_
	);
	LUT3 #(
		.INIT('ha2)
	) name2804 (
		\g518_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3579_
	);
	LUT4 #(
		.INIT('hf531)
	) name2805 (
		\g499_reg/NET0131 ,
		_w2615_,
		_w3578_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('h2)
	) name2806 (
		\g35_pad ,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h4)
	) name2807 (
		\g35_pad ,
		\g5112_reg/NET0131 ,
		_w3582_
	);
	LUT3 #(
		.INIT('h31)
	) name2808 (
		\g3096_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		\g5112_reg/NET0131 ,
		_w3583_
	);
	LUT2 #(
		.INIT('h2)
	) name2809 (
		\g35_pad ,
		\g5101_reg/NET0131 ,
		_w3584_
	);
	LUT3 #(
		.INIT('hba)
	) name2810 (
		_w3582_,
		_w3583_,
		_w3584_,
		_w3585_
	);
	LUT4 #(
		.INIT('h80ff)
	) name2811 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		\g35_pad ,
		_w3586_
	);
	LUT3 #(
		.INIT('hd2)
	) name2812 (
		\g35_pad ,
		\g5142_reg/NET0131 ,
		\g5148_reg/NET0131 ,
		_w3587_
	);
	LUT4 #(
		.INIT('hfd08)
	) name2813 (
		\g35_pad ,
		\g5152_reg/NET0131 ,
		_w3200_,
		_w3587_,
		_w3588_
	);
	LUT3 #(
		.INIT('h15)
	) name2814 (
		\g278_reg/NET0131 ,
		_w1707_,
		_w1708_,
		_w3589_
	);
	LUT3 #(
		.INIT('h2a)
	) name2815 (
		\g35_pad ,
		_w1711_,
		_w1712_,
		_w3590_
	);
	LUT2 #(
		.INIT('h4)
	) name2816 (
		_w3589_,
		_w3590_,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name2817 (
		\g1300_reg/NET0131 ,
		\g35_pad ,
		_w3592_
	);
	LUT2 #(
		.INIT('h2)
	) name2818 (
		\g1484_reg/NET0131 ,
		\g35_pad ,
		_w3593_
	);
	LUT3 #(
		.INIT('h08)
	) name2819 (
		\g1442_reg/NET0131 ,
		\g1484_reg/NET0131 ,
		\g1495_reg/NET0131 ,
		_w3594_
	);
	LUT4 #(
		.INIT('h363c)
	) name2820 (
		_w1012_,
		_w3592_,
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h8)
	) name2821 (
		\g1448_reg/NET0131 ,
		\g35_pad ,
		_w3596_
	);
	LUT2 #(
		.INIT('h2)
	) name2822 (
		\g1454_reg/NET0131 ,
		\g35_pad ,
		_w3597_
	);
	LUT3 #(
		.INIT('h08)
	) name2823 (
		\g1442_reg/NET0131 ,
		\g1454_reg/NET0131 ,
		\g1495_reg/NET0131 ,
		_w3598_
	);
	LUT4 #(
		.INIT('h363c)
	) name2824 (
		_w1000_,
		_w3596_,
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('h8)
	) name2825 (
		\g1472_reg/NET0131 ,
		\g35_pad ,
		_w3600_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		\g1467_reg/NET0131 ,
		\g35_pad ,
		_w3601_
	);
	LUT3 #(
		.INIT('h08)
	) name2827 (
		\g1442_reg/NET0131 ,
		\g1467_reg/NET0131 ,
		\g1495_reg/NET0131 ,
		_w3602_
	);
	LUT4 #(
		.INIT('h363c)
	) name2828 (
		_w1006_,
		_w3600_,
		_w3601_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name2829 (
		\g1478_reg/NET0131 ,
		\g35_pad ,
		_w3604_
	);
	LUT2 #(
		.INIT('h2)
	) name2830 (
		\g1437_reg/NET0131 ,
		\g35_pad ,
		_w3605_
	);
	LUT3 #(
		.INIT('h08)
	) name2831 (
		\g1437_reg/NET0131 ,
		\g1442_reg/NET0131 ,
		\g1495_reg/NET0131 ,
		_w3606_
	);
	LUT4 #(
		.INIT('h363c)
	) name2832 (
		_w992_,
		_w3604_,
		_w3605_,
		_w3606_,
		_w3607_
	);
	LUT3 #(
		.INIT('h47)
	) name2833 (
		\g3050_reg/NET0131 ,
		\g5016_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		_w3608_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		\g35_pad ,
		\g5029_reg/NET0131 ,
		_w3609_
	);
	LUT4 #(
		.INIT('h1000)
	) name2835 (
		_w2712_,
		_w2754_,
		_w3608_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h4)
	) name2836 (
		\g35_pad ,
		\g5016_reg/NET0131 ,
		_w3611_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		\g35_pad ,
		\g5029_reg/NET0131 ,
		_w3612_
	);
	LUT3 #(
		.INIT('h23)
	) name2838 (
		_w3608_,
		_w3611_,
		_w3612_,
		_w3613_
	);
	LUT2 #(
		.INIT('hb)
	) name2839 (
		_w3610_,
		_w3613_,
		_w3614_
	);
	LUT4 #(
		.INIT('h0002)
	) name2840 (
		\g35_pad ,
		\g4646_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		_w3615_
	);
	LUT2 #(
		.INIT('h4)
	) name2841 (
		_w1981_,
		_w3615_,
		_w3616_
	);
	LUT2 #(
		.INIT('h4)
	) name2842 (
		\g35_pad ,
		\g4621_reg/NET0131 ,
		_w3617_
	);
	LUT4 #(
		.INIT('hff60)
	) name2843 (
		\g4628_reg/NET0131 ,
		_w3425_,
		_w3427_,
		_w3617_,
		_w3618_
	);
	LUT4 #(
		.INIT('h4ee4)
	) name2844 (
		\g35_pad ,
		\g5124_reg/NET0131 ,
		\g5128_reg/NET0131 ,
		_w3200_,
		_w3619_
	);
	LUT4 #(
		.INIT('h3aca)
	) name2845 (
		\g3115_reg/NET0131 ,
		\g3119_reg/NET0131 ,
		\g35_pad ,
		_w3200_,
		_w3620_
	);
	LUT4 #(
		.INIT('h3b33)
	) name2846 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w3621_
	);
	LUT4 #(
		.INIT('h3aca)
	) name2847 (
		\g3466_reg/NET0131 ,
		\g3470_reg/NET0131 ,
		\g35_pad ,
		_w3200_,
		_w3622_
	);
	LUT4 #(
		.INIT('hd777)
	) name2848 (
		\g35_pad ,
		\g370_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w2053_,
		_w3623_
	);
	LUT2 #(
		.INIT('h2)
	) name2849 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		_w3624_
	);
	LUT2 #(
		.INIT('hd)
	) name2850 (
		_w3623_,
		_w3624_,
		_w3625_
	);
	LUT4 #(
		.INIT('h4ee4)
	) name2851 (
		\g35_pad ,
		\g3817_reg/NET0131 ,
		\g3821_reg/NET0131 ,
		_w3200_,
		_w3626_
	);
	LUT3 #(
		.INIT('h2a)
	) name2852 (
		\g209_reg/NET0131 ,
		\g218_reg/NET0131 ,
		\g8291_pad ,
		_w3627_
	);
	LUT4 #(
		.INIT('h4000)
	) name2853 (
		\g191_reg/NET0131 ,
		\g218_reg/NET0131 ,
		\g8291_pad ,
		\g8358_pad ,
		_w3628_
	);
	LUT3 #(
		.INIT('ha8)
	) name2854 (
		\g35_pad ,
		_w3627_,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		\g191_reg/NET0131 ,
		\g35_pad ,
		_w3630_
	);
	LUT4 #(
		.INIT('h0080)
	) name2856 (
		\g191_reg/NET0131 ,
		\g218_reg/NET0131 ,
		\g8291_pad ,
		\g8358_pad ,
		_w3631_
	);
	LUT2 #(
		.INIT('h1)
	) name2857 (
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT2 #(
		.INIT('hb)
	) name2858 (
		_w3629_,
		_w3632_,
		_w3633_
	);
	LUT2 #(
		.INIT('h4)
	) name2859 (
		\g35_pad ,
		\g4180_reg/NET0131 ,
		_w3634_
	);
	LUT4 #(
		.INIT('h0a22)
	) name2860 (
		\g35_pad ,
		\g4145_reg/NET0131 ,
		\g4164_reg/NET0131 ,
		\g4253_reg/NET0131 ,
		_w3635_
	);
	LUT2 #(
		.INIT('he)
	) name2861 (
		_w3634_,
		_w3635_,
		_w3636_
	);
	LUT3 #(
		.INIT('h4e)
	) name2862 (
		\g35_pad ,
		\g4245_reg/NET0131 ,
		\g4281_reg/NET0131 ,
		_w3637_
	);
	LUT4 #(
		.INIT('h8000)
	) name2863 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g7916_pad ,
		\g996_reg/NET0131 ,
		_w3638_
	);
	LUT3 #(
		.INIT('h80)
	) name2864 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g7916_pad ,
		_w3639_
	);
	LUT4 #(
		.INIT('h5f57)
	) name2865 (
		\g35_pad ,
		\g962_reg/NET0131 ,
		_w3638_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h2)
	) name2866 (
		\g1178_reg/NET0131 ,
		\g35_pad ,
		_w3641_
	);
	LUT2 #(
		.INIT('hd)
	) name2867 (
		_w3640_,
		_w3641_,
		_w3642_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		\g35_pad ,
		\g499_reg/NET0131 ,
		_w3643_
	);
	LUT3 #(
		.INIT('h51)
	) name2869 (
		\g499_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3644_
	);
	LUT2 #(
		.INIT('h2)
	) name2870 (
		\g35_pad ,
		\g504_reg/NET0131 ,
		_w3645_
	);
	LUT4 #(
		.INIT('h0213)
	) name2871 (
		_w2615_,
		_w3643_,
		_w3644_,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h2)
	) name2872 (
		\g35_pad ,
		\g4308_reg/NET0131 ,
		_w3647_
	);
	LUT2 #(
		.INIT('h4)
	) name2873 (
		\g35_pad ,
		\g504_reg/NET0131 ,
		_w3648_
	);
	LUT3 #(
		.INIT('ha2)
	) name2874 (
		\g504_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3649_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		\g35_pad ,
		\g513_reg/NET0131 ,
		_w3650_
	);
	LUT4 #(
		.INIT('hfdec)
	) name2876 (
		_w2615_,
		_w3648_,
		_w3649_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('he)
	) name2877 (
		\g2748_reg/NET0131 ,
		\g35_pad ,
		_w3652_
	);
	LUT3 #(
		.INIT('h9c)
	) name2878 (
		\g3133_reg/NET0131 ,
		\g3139_reg/NET0131 ,
		\g35_pad ,
		_w3653_
	);
	LUT4 #(
		.INIT('hfb08)
	) name2879 (
		\g3143_reg/NET0131 ,
		\g35_pad ,
		_w3200_,
		_w3653_,
		_w3654_
	);
	LUT3 #(
		.INIT('h9c)
	) name2880 (
		\g3484_reg/NET0131 ,
		\g3490_reg/NET0131 ,
		\g35_pad ,
		_w3655_
	);
	LUT4 #(
		.INIT('hfb08)
	) name2881 (
		\g3494_reg/NET0131 ,
		\g35_pad ,
		_w3200_,
		_w3655_,
		_w3656_
	);
	LUT3 #(
		.INIT('hd2)
	) name2882 (
		\g35_pad ,
		\g3835_reg/NET0131 ,
		\g3841_reg/NET0131 ,
		_w3657_
	);
	LUT4 #(
		.INIT('hfd08)
	) name2883 (
		\g35_pad ,
		\g3845_reg/NET0131 ,
		_w3200_,
		_w3657_,
		_w3658_
	);
	LUT4 #(
		.INIT('h0800)
	) name2884 (
		\g4076_reg/NET0131 ,
		\g4087_reg/NET0131 ,
		\g4093_reg/NET0131 ,
		\g4098_reg/NET0131 ,
		_w3659_
	);
	LUT4 #(
		.INIT('h0001)
	) name2885 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		\g4082_reg/NET0131 ,
		\g4141_reg/NET0131 ,
		_w3660_
	);
	LUT3 #(
		.INIT('h2a)
	) name2886 (
		\g35_pad ,
		_w3659_,
		_w3660_,
		_w3661_
	);
	LUT4 #(
		.INIT('h5078)
	) name2887 (
		\g35_pad ,
		\g4621_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3662_
	);
	LUT2 #(
		.INIT('h1)
	) name2888 (
		\g2965_reg/NET0131 ,
		\g35_pad ,
		_w3663_
	);
	LUT4 #(
		.INIT('h2000)
	) name2889 (
		\g1306_reg/NET0131 ,
		\g2975_reg/NET0131 ,
		\g35_pad ,
		\g962_reg/NET0131 ,
		_w3664_
	);
	LUT2 #(
		.INIT('h1)
	) name2890 (
		_w3663_,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		\g35_pad ,
		\g518_reg/NET0131 ,
		_w3666_
	);
	LUT2 #(
		.INIT('h4)
	) name2892 (
		\g35_pad ,
		\g513_reg/NET0131 ,
		_w3667_
	);
	LUT3 #(
		.INIT('ha2)
	) name2893 (
		\g513_reg/NET0131 ,
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3668_
	);
	LUT4 #(
		.INIT('hfef4)
	) name2894 (
		_w2615_,
		_w3666_,
		_w3667_,
		_w3668_,
		_w3669_
	);
	LUT4 #(
		.INIT('h0002)
	) name2895 (
		\g13272_pad ,
		\g1442_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w3670_
	);
	LUT4 #(
		.INIT('h0008)
	) name2896 (
		\g13272_pad ,
		\g1495_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w3671_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name2897 (
		\g1489_reg/NET0131 ,
		\g35_pad ,
		_w3670_,
		_w3671_,
		_w3672_
	);
	LUT3 #(
		.INIT('he4)
	) name2898 (
		\g35_pad ,
		\g4459_reg/NET0131 ,
		\g4473_reg/NET0131 ,
		_w3673_
	);
	LUT2 #(
		.INIT('h1)
	) name2899 (
		\g35_pad ,
		\g4492_reg/NET0131 ,
		_w3674_
	);
	LUT2 #(
		.INIT('h4)
	) name2900 (
		\g2988_reg/NET0131 ,
		\g35_pad ,
		_w3675_
	);
	LUT3 #(
		.INIT('h23)
	) name2901 (
		_w927_,
		_w3674_,
		_w3675_,
		_w3676_
	);
	LUT4 #(
		.INIT('h0800)
	) name2902 (
		\g35_pad ,
		\g4462_reg/NET0131 ,
		\g4467_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3677_
	);
	LUT2 #(
		.INIT('h2)
	) name2903 (
		\g4473_reg/NET0131 ,
		_w3677_,
		_w3678_
	);
	LUT3 #(
		.INIT('h6c)
	) name2904 (
		\g35_pad ,
		\g5084_reg/NET0131 ,
		\g5092_reg/NET0131 ,
		_w3679_
	);
	LUT3 #(
		.INIT('h6a)
	) name2905 (
		\g1087_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		\g35_pad ,
		_w3680_
	);
	LUT4 #(
		.INIT('h74b8)
	) name2906 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		\g370_reg/NET0131 ,
		\g376_reg/NET0131 ,
		_w3681_
	);
	LUT3 #(
		.INIT('h6c)
	) name2907 (
		\g35_pad ,
		\g4258_reg/NET0131 ,
		\g4264_reg/NET0131 ,
		_w3682_
	);
	LUT3 #(
		.INIT('hc6)
	) name2908 (
		\g35_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		_w3683_
	);
	LUT3 #(
		.INIT('h6a)
	) name2909 (
		\g1430_reg/NET0131 ,
		\g1548_reg/NET0131 ,
		\g35_pad ,
		_w3684_
	);
	LUT3 #(
		.INIT('hd5)
	) name2910 (
		\g35_pad ,
		_w912_,
		_w913_,
		_w3685_
	);
	LUT2 #(
		.INIT('h4)
	) name2911 (
		\g35_pad ,
		\g4633_reg/NET0131 ,
		_w3686_
	);
	LUT4 #(
		.INIT('h0008)
	) name2912 (
		\g4621_reg/NET0131 ,
		\g4633_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3687_
	);
	LUT2 #(
		.INIT('he)
	) name2913 (
		_w3686_,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h8)
	) name2914 (
		\g3179_reg/NET0131 ,
		\g35_pad ,
		_w3689_
	);
	LUT4 #(
		.INIT('h78cc)
	) name2915 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		\g35_pad ,
		_w3690_
	);
	LUT3 #(
		.INIT('hac)
	) name2916 (
		\g18098_pad ,
		\g305_reg/NET0131 ,
		\g35_pad ,
		_w3691_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name2917 (
		\g2886_reg/NET0131 ,
		\g2980_reg/NET0131 ,
		\g34_reg/NET0131 ,
		\g35_pad ,
		_w3692_
	);
	LUT3 #(
		.INIT('h6a)
	) name2918 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g35_pad ,
		_w3693_
	);
	LUT3 #(
		.INIT('h4e)
	) name2919 (
		\g35_pad ,
		\g5057_reg/NET0131 ,
		_w2754_,
		_w3694_
	);
	LUT3 #(
		.INIT('h6c)
	) name2920 (
		\g35_pad ,
		\g4308_reg/NET0131 ,
		\g9251_pad ,
		_w3695_
	);
	LUT3 #(
		.INIT('h6a)
	) name2921 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		\g35_pad ,
		_w3696_
	);
	LUT4 #(
		.INIT('h5ad8)
	) name2922 (
		\g35_pad ,
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		\g896_reg/NET0131 ,
		_w3697_
	);
	LUT3 #(
		.INIT('h6c)
	) name2923 (
		\g35_pad ,
		\g4291_reg/NET0131 ,
		\g9019_pad ,
		_w3698_
	);
	LUT4 #(
		.INIT('hd050)
	) name2924 (
		\g35_pad ,
		\g376_reg/NET0131 ,
		\g385_reg/NET0131 ,
		\g8719_pad ,
		_w3699_
	);
	LUT3 #(
		.INIT('h6c)
	) name2925 (
		\g35_pad ,
		\g4281_reg/NET0131 ,
		\g8839_pad ,
		_w3700_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name2926 (
		\g1521_reg/NET0131 ,
		\g1532_reg/NET0131 ,
		\g35_pad ,
		\g7946_pad ,
		_w3701_
	);
	LUT2 #(
		.INIT('h2)
	) name2927 (
		\g1306_reg/NET0131 ,
		\g35_pad ,
		_w3702_
	);
	LUT2 #(
		.INIT('he)
	) name2928 (
		_w3701_,
		_w3702_,
		_w3703_
	);
	LUT4 #(
		.INIT('hc808)
	) name2929 (
		\g1178_reg/NET0131 ,
		\g35_pad ,
		\g7916_pad ,
		\g996_reg/NET0131 ,
		_w3704_
	);
	LUT2 #(
		.INIT('h2)
	) name2930 (
		\g1183_reg/NET0131 ,
		\g35_pad ,
		_w3705_
	);
	LUT2 #(
		.INIT('he)
	) name2931 (
		_w3704_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name2932 (
		\g1178_reg/NET0131 ,
		\g1189_reg/NET0131 ,
		\g35_pad ,
		\g7916_pad ,
		_w3707_
	);
	LUT2 #(
		.INIT('h4)
	) name2933 (
		\g35_pad ,
		\g962_reg/NET0131 ,
		_w3708_
	);
	LUT2 #(
		.INIT('he)
	) name2934 (
		_w3707_,
		_w3708_,
		_w3709_
	);
	LUT2 #(
		.INIT('he)
	) name2935 (
		\g2724_reg/NET0131 ,
		\g35_pad ,
		_w3710_
	);
	LUT2 #(
		.INIT('h2)
	) name2936 (
		\g2741_reg/NET0131 ,
		\g35_pad ,
		_w3711_
	);
	LUT4 #(
		.INIT('h02ff)
	) name2937 (
		\g13272_pad ,
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g35_pad ,
		_w3712_
	);
	LUT4 #(
		.INIT('h08cc)
	) name2938 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		\g3167_reg/NET0131 ,
		\g35_pad ,
		_w3713_
	);
	LUT4 #(
		.INIT('h3074)
	) name2939 (
		\g10122_pad ,
		\g35_pad ,
		\g4239_reg/NET0131 ,
		\g4297_reg/NET0131 ,
		_w3714_
	);
	LUT4 #(
		.INIT('h444e)
	) name2940 (
		\g35_pad ,
		\g4462_reg/NET0131 ,
		\g4467_reg/NET0131 ,
		\g4473_reg/NET0131 ,
		_w3715_
	);
	LUT4 #(
		.INIT('hfc74)
	) name2941 (
		\g29212_pad ,
		\g35_pad ,
		\g534_reg/NET0131 ,
		\g550_reg/NET0131 ,
		_w3716_
	);
	LUT4 #(
		.INIT('hcfaa)
	) name2942 (
		\g2980_reg/NET0131 ,
		\g2984_reg/NET0131 ,
		\g34_reg/NET0131 ,
		\g35_pad ,
		_w3717_
	);
	LUT4 #(
		.INIT('he4ee)
	) name2943 (
		\g35_pad ,
		\g538_reg/NET0131 ,
		\g546_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w3718_
	);
	LUT3 #(
		.INIT('h3a)
	) name2944 (
		\g209_reg/NET0131 ,
		\g218_reg/NET0131 ,
		\g35_pad ,
		_w3719_
	);
	LUT4 #(
		.INIT('h4eee)
	) name2945 (
		\g35_pad ,
		\g4122_reg/NET0131 ,
		\g4146_reg/NET0131 ,
		\g4157_reg/NET0131 ,
		_w3720_
	);
	LUT3 #(
		.INIT('hc8)
	) name2946 (
		\g209_reg/NET0131 ,
		\g35_pad ,
		\g538_reg/NET0131 ,
		_w3721_
	);
	LUT3 #(
		.INIT('ha8)
	) name2947 (
		\g35_pad ,
		\g4153_reg/NET0131 ,
		\g4172_reg/NET0131 ,
		_w3722_
	);
	LUT4 #(
		.INIT('hfddd)
	) name2948 (
		\g35_pad ,
		\g4462_reg/NET0131 ,
		\g4467_reg/NET0131 ,
		\g4473_reg/NET0131 ,
		_w3723_
	);
	LUT3 #(
		.INIT('h10)
	) name2949 (
		\g3155_reg/NET0131 ,
		\g3167_reg/NET0131 ,
		\g35_pad ,
		_w3724_
	);
	LUT2 #(
		.INIT('he)
	) name2950 (
		\g2715_reg/NET0131 ,
		\g35_pad ,
		_w3725_
	);
	LUT3 #(
		.INIT('h02)
	) name2951 (
		\g35_pad ,
		\g4639_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3726_
	);
	LUT3 #(
		.INIT('h04)
	) name2952 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		\g8719_pad ,
		_w3727_
	);
	LUT3 #(
		.INIT('h2a)
	) name2953 (
		\g35_pad ,
		\g4462_reg/NET0131 ,
		\g4467_reg/NET0131 ,
		_w3728_
	);
	LUT3 #(
		.INIT('hca)
	) name2954 (
		\g3050_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g35_pad ,
		_w3729_
	);
	LUT3 #(
		.INIT('hb8)
	) name2955 (
		\g18094_pad ,
		\g35_pad ,
		\g4483_reg/NET0131 ,
		_w3730_
	);
	LUT3 #(
		.INIT('hb8)
	) name2956 (
		\g18095_pad ,
		\g35_pad ,
		\g4486_reg/NET0131 ,
		_w3731_
	);
	LUT3 #(
		.INIT('hb8)
	) name2957 (
		\g18096_pad ,
		\g35_pad ,
		\g4489_reg/NET0131 ,
		_w3732_
	);
	LUT3 #(
		.INIT('h72)
	) name2958 (
		\g35_pad ,
		\g4239_reg/NET0131 ,
		\g4273_reg/NET0131 ,
		_w3733_
	);
	LUT2 #(
		.INIT('h2)
	) name2959 (
		\g2735_reg/NET0131 ,
		\g35_pad ,
		_w3734_
	);
	LUT2 #(
		.INIT('h4)
	) name2960 (
		\g35_pad ,
		\g4382_reg/NET0131 ,
		_w3735_
	);
	LUT2 #(
		.INIT('h2)
	) name2961 (
		\g2719_reg/NET0131 ,
		\g35_pad ,
		_w3736_
	);
	LUT2 #(
		.INIT('h4)
	) name2962 (
		\g35_pad ,
		\g4392_reg/NET0131 ,
		_w3737_
	);
	LUT2 #(
		.INIT('h4)
	) name2963 (
		\g35_pad ,
		\g4153_reg/NET0131 ,
		_w3738_
	);
	LUT2 #(
		.INIT('h2)
	) name2964 (
		\g2975_reg/NET0131 ,
		\g35_pad ,
		_w3739_
	);
	LUT2 #(
		.INIT('h4)
	) name2965 (
		\g35_pad ,
		\g4104_reg/NET0131 ,
		_w3740_
	);
	LUT2 #(
		.INIT('h4)
	) name2966 (
		\g35_pad ,
		\g4087_reg/NET0131 ,
		_w3741_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		\g35_pad ,
		\g4057_reg/NET0131 ,
		_w3742_
	);
	LUT2 #(
		.INIT('h4)
	) name2968 (
		\g35_pad ,
		\g4076_reg/NET0131 ,
		_w3743_
	);
	LUT2 #(
		.INIT('h4)
	) name2969 (
		\g35_pad ,
		\g4064_reg/NET0131 ,
		_w3744_
	);
	LUT2 #(
		.INIT('h4)
	) name2970 (
		\g35_pad ,
		\g753_reg/NET0131 ,
		_w3745_
	);
	LUT2 #(
		.INIT('he)
	) name2971 (
		\g2759_reg/NET0131 ,
		\g35_pad ,
		_w3746_
	);
	LUT2 #(
		.INIT('he)
	) name2972 (
		\g35_pad ,
		\g4108_reg/NET0131 ,
		_w3747_
	);
	LUT2 #(
		.INIT('he)
	) name2973 (
		\g2756_reg/NET0131 ,
		\g35_pad ,
		_w3748_
	);
	LUT2 #(
		.INIT('he)
	) name2974 (
		\g2917_reg/NET0131 ,
		\g35_pad ,
		_w3749_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		\g18099_pad ,
		\g35_pad ,
		_w3750_
	);
	LUT2 #(
		.INIT('he)
	) name2976 (
		\g2882_reg/NET0131 ,
		\g35_pad ,
		_w3751_
	);
	LUT2 #(
		.INIT('he)
	) name2977 (
		\g35_pad ,
		\g4141_reg/NET0131 ,
		_w3752_
	);
	LUT2 #(
		.INIT('he)
	) name2978 (
		\g35_pad ,
		\g4082_reg/NET0131 ,
		_w3753_
	);
	LUT2 #(
		.INIT('h8)
	) name2979 (
		\g29216_pad ,
		\g35_pad ,
		_w3754_
	);
	LUT2 #(
		.INIT('he)
	) name2980 (
		\g2955_reg/NET0131 ,
		\g35_pad ,
		_w3755_
	);
	LUT2 #(
		.INIT('he)
	) name2981 (
		\g35_pad ,
		\g4098_reg/NET0131 ,
		_w3756_
	);
	LUT2 #(
		.INIT('he)
	) name2982 (
		\g35_pad ,
		\g4093_reg/NET0131 ,
		_w3757_
	);
	LUT2 #(
		.INIT('he)
	) name2983 (
		\g2873_reg/NET0131 ,
		\g35_pad ,
		_w3758_
	);
	LUT2 #(
		.INIT('he)
	) name2984 (
		\g2729_reg/NET0131 ,
		\g35_pad ,
		_w3759_
	);
	LUT3 #(
		.INIT('h01)
	) name2985 (
		\g2421_reg/NET0131 ,
		_w1363_,
		_w1365_,
		_w3760_
	);
	LUT3 #(
		.INIT('h2a)
	) name2986 (
		\g2495_reg/NET0131 ,
		_w800_,
		_w1160_,
		_w3761_
	);
	LUT2 #(
		.INIT('h8)
	) name2987 (
		\g17423_pad ,
		\g2495_reg/NET0131 ,
		_w3762_
	);
	LUT3 #(
		.INIT('h70)
	) name2988 (
		_w1129_,
		_w1162_,
		_w3762_,
		_w3763_
	);
	LUT3 #(
		.INIT('h02)
	) name2989 (
		\g35_pad ,
		_w3761_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h4)
	) name2990 (
		_w3760_,
		_w3764_,
		_w3765_
	);
	LUT3 #(
		.INIT('h01)
	) name2991 (
		\g2287_reg/NET0131 ,
		_w1313_,
		_w1315_,
		_w3766_
	);
	LUT3 #(
		.INIT('h2a)
	) name2992 (
		\g2361_reg/NET0131 ,
		_w800_,
		_w1144_,
		_w3767_
	);
	LUT2 #(
		.INIT('h8)
	) name2993 (
		\g17404_pad ,
		\g2361_reg/NET0131 ,
		_w3768_
	);
	LUT3 #(
		.INIT('h70)
	) name2994 (
		_w1129_,
		_w1146_,
		_w3768_,
		_w3769_
	);
	LUT3 #(
		.INIT('h02)
	) name2995 (
		\g35_pad ,
		_w3767_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h4)
	) name2996 (
		_w3766_,
		_w3770_,
		_w3771_
	);
	LUT3 #(
		.INIT('h01)
	) name2997 (
		\g2555_reg/NET0131 ,
		_w1410_,
		_w1412_,
		_w3772_
	);
	LUT3 #(
		.INIT('h02)
	) name2998 (
		\g35_pad ,
		_w1437_,
		_w1439_,
		_w3773_
	);
	LUT2 #(
		.INIT('h4)
	) name2999 (
		_w3772_,
		_w3773_,
		_w3774_
	);
	LUT3 #(
		.INIT('h01)
	) name3000 (
		\g1862_reg/NET0131 ,
		_w1539_,
		_w1541_,
		_w3775_
	);
	LUT3 #(
		.INIT('h2a)
	) name3001 (
		\g1936_reg/NET0131 ,
		_w802_,
		_w1225_,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name3002 (
		\g17400_pad ,
		\g1936_reg/NET0131 ,
		_w3777_
	);
	LUT3 #(
		.INIT('h70)
	) name3003 (
		_w1210_,
		_w1227_,
		_w3777_,
		_w3778_
	);
	LUT3 #(
		.INIT('h02)
	) name3004 (
		\g35_pad ,
		_w3776_,
		_w3778_,
		_w3779_
	);
	LUT2 #(
		.INIT('h4)
	) name3005 (
		_w3775_,
		_w3779_,
		_w3780_
	);
	LUT3 #(
		.INIT('h01)
	) name3006 (
		\g1996_reg/NET0131 ,
		_w1625_,
		_w1627_,
		_w3781_
	);
	LUT3 #(
		.INIT('h2a)
	) name3007 (
		\g2070_reg/NET0131 ,
		_w802_,
		_w1241_,
		_w3782_
	);
	LUT2 #(
		.INIT('h8)
	) name3008 (
		\g1087_reg/NET0131 ,
		\g2070_reg/NET0131 ,
		_w3783_
	);
	LUT3 #(
		.INIT('h70)
	) name3009 (
		_w1210_,
		_w1243_,
		_w3783_,
		_w3784_
	);
	LUT3 #(
		.INIT('h02)
	) name3010 (
		\g35_pad ,
		_w3782_,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('h4)
	) name3011 (
		_w3781_,
		_w3785_,
		_w3786_
	);
	LUT3 #(
		.INIT('h2a)
	) name3012 (
		\g35_pad ,
		_w802_,
		_w1633_,
		_w3787_
	);
	LUT2 #(
		.INIT('h8)
	) name3013 (
		\g17291_pad ,
		\g35_pad ,
		_w3788_
	);
	LUT3 #(
		.INIT('h70)
	) name3014 (
		_w1210_,
		_w1635_,
		_w3788_,
		_w3789_
	);
	LUT3 #(
		.INIT('he0)
	) name3015 (
		\g1592_reg/NET0131 ,
		\g1668_reg/NET0131 ,
		\g1682_reg/NET0131 ,
		_w3790_
	);
	LUT4 #(
		.INIT('h0100)
	) name3016 (
		\g1135_reg/NET0131 ,
		\g1246_reg/NET0131 ,
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w3791_
	);
	LUT3 #(
		.INIT('h93)
	) name3017 (
		_w802_,
		_w3790_,
		_w3791_,
		_w3792_
	);
	LUT3 #(
		.INIT('he0)
	) name3018 (
		_w3787_,
		_w3789_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h8)
	) name3019 (
		\g1682_reg/NET0131 ,
		\g35_pad ,
		_w3794_
	);
	LUT3 #(
		.INIT('h80)
	) name3020 (
		_w802_,
		_w1633_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('h2)
	) name3021 (
		\g1668_reg/NET0131 ,
		\g35_pad ,
		_w3796_
	);
	LUT3 #(
		.INIT('h0b)
	) name3022 (
		_w3284_,
		_w3795_,
		_w3796_,
		_w3797_
	);
	LUT2 #(
		.INIT('hb)
	) name3023 (
		_w3793_,
		_w3797_,
		_w3798_
	);
	LUT3 #(
		.INIT('h01)
	) name3024 (
		\g1728_reg/NET0131 ,
		_w1492_,
		_w1494_,
		_w3799_
	);
	LUT3 #(
		.INIT('h2a)
	) name3025 (
		\g1802_reg/NET0131 ,
		_w802_,
		_w1208_,
		_w3800_
	);
	LUT2 #(
		.INIT('h8)
	) name3026 (
		\g17316_pad ,
		\g1802_reg/NET0131 ,
		_w3801_
	);
	LUT3 #(
		.INIT('h70)
	) name3027 (
		_w1210_,
		_w1211_,
		_w3801_,
		_w3802_
	);
	LUT3 #(
		.INIT('h02)
	) name3028 (
		\g35_pad ,
		_w3800_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h4)
	) name3029 (
		_w3799_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('h2)
	) name3030 (
		\g3457_reg/NET0131 ,
		_w3215_,
		_w3805_
	);
	LUT2 #(
		.INIT('h2)
	) name3031 (
		_w2015_,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h8)
	) name3032 (
		_w2015_,
		_w3805_,
		_w3807_
	);
	LUT3 #(
		.INIT('h31)
	) name3033 (
		\g3457_reg/NET0131 ,
		_w873_,
		_w2012_,
		_w3808_
	);
	LUT4 #(
		.INIT('he4ff)
	) name3034 (
		_w1872_,
		_w3806_,
		_w3807_,
		_w3808_,
		_w3809_
	);
	LUT4 #(
		.INIT('h8000)
	) name3035 (
		\g16624_pad ,
		\g3288_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g3352_reg/NET0131 ,
		_w3810_
	);
	LUT2 #(
		.INIT('h2)
	) name3036 (
		\g3106_reg/NET0131 ,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h2)
	) name3037 (
		_w1944_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h8)
	) name3038 (
		_w1944_,
		_w3811_,
		_w3813_
	);
	LUT3 #(
		.INIT('h31)
	) name3039 (
		\g3106_reg/NET0131 ,
		_w873_,
		_w1941_,
		_w3814_
	);
	LUT4 #(
		.INIT('he4ff)
	) name3040 (
		_w1851_,
		_w3812_,
		_w3813_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('h2)
	) name3041 (
		\g1171_reg/NET0131 ,
		\g35_pad ,
		_w3816_
	);
	LUT2 #(
		.INIT('h2)
	) name3042 (
		\g1171_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		_w3817_
	);
	LUT3 #(
		.INIT('h23)
	) name3043 (
		_w2737_,
		_w3816_,
		_w3817_,
		_w3818_
	);
	LUT3 #(
		.INIT('h45)
	) name3044 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		_w3819_
	);
	LUT3 #(
		.INIT('h6c)
	) name3045 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g7916_pad ,
		_w3820_
	);
	LUT4 #(
		.INIT('haa20)
	) name3046 (
		\g35_pad ,
		_w2737_,
		_w3819_,
		_w3820_,
		_w3821_
	);
	LUT2 #(
		.INIT('hd)
	) name3047 (
		_w3818_,
		_w3821_,
		_w3822_
	);
	LUT2 #(
		.INIT('h2)
	) name3048 (
		\g5297_reg/NET0131 ,
		_w840_,
		_w3823_
	);
	LUT2 #(
		.INIT('h8)
	) name3049 (
		_w839_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name3050 (
		\g5297_reg/NET0131 ,
		_w846_,
		_w3825_
	);
	LUT3 #(
		.INIT('h2a)
	) name3051 (
		\g5357_reg/NET0131 ,
		_w845_,
		_w3825_,
		_w3826_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3052 (
		\g13865_pad ,
		\g3231_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g5297_reg/NET0131 ,
		_w3827_
	);
	LUT3 #(
		.INIT('he0)
	) name3053 (
		\g3338_reg/NET0131 ,
		_w852_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h4)
	) name3054 (
		_w851_,
		_w3828_,
		_w3829_
	);
	LUT4 #(
		.INIT('h00f7)
	) name3055 (
		\g13865_pad ,
		\g3239_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		\g5297_reg/NET0131 ,
		_w3830_
	);
	LUT3 #(
		.INIT('hd0)
	) name3056 (
		\g3338_reg/NET0131 ,
		_w859_,
		_w3830_,
		_w3831_
	);
	LUT3 #(
		.INIT('h45)
	) name3057 (
		\g5357_reg/NET0131 ,
		_w858_,
		_w3831_,
		_w3832_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3058 (
		_w3824_,
		_w3826_,
		_w3829_,
		_w3832_,
		_w3833_
	);
	LUT2 #(
		.INIT('h2)
	) name3059 (
		\g5115_reg/NET0131 ,
		_w3073_,
		_w3834_
	);
	LUT2 #(
		.INIT('h2)
	) name3060 (
		_w2090_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h8)
	) name3061 (
		_w2090_,
		_w3834_,
		_w3836_
	);
	LUT3 #(
		.INIT('h31)
	) name3062 (
		\g5115_reg/NET0131 ,
		_w873_,
		_w2087_,
		_w3837_
	);
	LUT4 #(
		.INIT('he4ff)
	) name3063 (
		_w3833_,
		_w3835_,
		_w3836_,
		_w3837_,
		_w3838_
	);
	LUT3 #(
		.INIT('h01)
	) name3064 (
		\g2153_reg/NET0131 ,
		_w1266_,
		_w1268_,
		_w3839_
	);
	LUT3 #(
		.INIT('h2a)
	) name3065 (
		\g2227_reg/NET0131 ,
		_w800_,
		_w1127_,
		_w3840_
	);
	LUT2 #(
		.INIT('h8)
	) name3066 (
		\g17320_pad ,
		\g2227_reg/NET0131 ,
		_w3841_
	);
	LUT3 #(
		.INIT('h70)
	) name3067 (
		_w1129_,
		_w1130_,
		_w3841_,
		_w3842_
	);
	LUT3 #(
		.INIT('h02)
	) name3068 (
		\g35_pad ,
		_w3840_,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name3069 (
		_w3839_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h4)
	) name3070 (
		\g35_pad ,
		\g4572_reg/NET0131 ,
		_w3845_
	);
	LUT2 #(
		.INIT('h1)
	) name3071 (
		\g35_pad ,
		\g4572_reg/NET0131 ,
		_w3846_
	);
	LUT3 #(
		.INIT('h01)
	) name3072 (
		\g4776_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		\g4801_reg/NET0131 ,
		_w3847_
	);
	LUT4 #(
		.INIT('h0001)
	) name3073 (
		\g4646_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w3848_
	);
	LUT4 #(
		.INIT('hdc00)
	) name3074 (
		_w822_,
		_w1945_,
		_w3847_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('h3fdd)
	) name3075 (
		\g4698_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4765_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w3850_
	);
	LUT4 #(
		.INIT('hbb5f)
	) name3076 (
		\g4709_reg/NET0131 ,
		\g4743_reg/NET0131 ,
		\g4754_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w3851_
	);
	LUT3 #(
		.INIT('hb9)
	) name3077 (
		\g4776_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		\g4801_reg/NET0131 ,
		_w3852_
	);
	LUT4 #(
		.INIT('h002a)
	) name3078 (
		_w3848_,
		_w3850_,
		_w3851_,
		_w3852_,
		_w3853_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3079 (
		\g3684_reg/NET0131 ,
		\g4035_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w3854_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3080 (
		\g29220_pad ,
		\g3333_reg/NET0131 ,
		\g4646_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		_w3855_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT3 #(
		.INIT('h40)
	) name3082 (
		_w3845_,
		_w3854_,
		_w3855_,
		_w3857_
	);
	LUT4 #(
		.INIT('h5455)
	) name3083 (
		_w3846_,
		_w3849_,
		_w3853_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3084 (
		\g35_pad ,
		_w3849_,
		_w3853_,
		_w3856_,
		_w3859_
	);
	LUT3 #(
		.INIT('h08)
	) name3085 (
		\g691_reg/NET0131 ,
		\g703_reg/NET0131 ,
		\g714_reg/NET0131 ,
		_w3860_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3086 (
		_w2026_,
		_w2027_,
		_w2720_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h8)
	) name3087 (
		\g35_pad ,
		\g691_reg/NET0131 ,
		_w3862_
	);
	LUT2 #(
		.INIT('h2)
	) name3088 (
		\g29212_pad ,
		\g35_pad ,
		_w3863_
	);
	LUT3 #(
		.INIT('h0b)
	) name3089 (
		_w2615_,
		_w3862_,
		_w3863_,
		_w3864_
	);
	LUT3 #(
		.INIT('h4f)
	) name3090 (
		_w3861_,
		_w2721_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h1)
	) name3091 (
		\g29220_pad ,
		\g4646_reg/NET0131 ,
		_w3866_
	);
	LUT4 #(
		.INIT('h0004)
	) name3092 (
		\g29220_pad ,
		\g4698_reg/NET0131 ,
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w3867_
	);
	LUT4 #(
		.INIT('h070f)
	) name3093 (
		_w824_,
		_w825_,
		_w3866_,
		_w3867_,
		_w3868_
	);
	LUT3 #(
		.INIT('h1d)
	) name3094 (
		\g3263_reg/NET0131 ,
		\g35_pad ,
		_w3868_,
		_w3869_
	);
	LUT2 #(
		.INIT('h2)
	) name3095 (
		_w827_,
		_w1834_,
		_w3870_
	);
	LUT3 #(
		.INIT('h13)
	) name3096 (
		_w3833_,
		_w3869_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h2)
	) name3097 (
		\g301_reg/NET0131 ,
		\g35_pad ,
		_w3872_
	);
	LUT4 #(
		.INIT('hff80)
	) name3098 (
		_w1715_,
		_w1718_,
		_w1719_,
		_w3872_,
		_w3873_
	);
	assign \g136_reg/P0001  = _w404_ ;
	assign \g21727_pad  = _w781_ ;
	assign \g23190_pad  = 1'b1;
	assign \g26875_pad  = _w784_ ;
	assign \g26876_pad  = _w791_ ;
	assign \g26877_pad  = _w798_ ;
	assign \g28041_pad  = _w804_ ;
	assign \g28042_pad  = _w805_ ;
	assign \g30327_pad  = _w502_ ;
	assign \g30330_pad  = _w378_ ;
	assign \g30331_pad  = _w376_ ;
	assign \g31793_pad  = _w807_ ;
	assign \g31860_pad  = _w808_ ;
	assign \g31862_pad  = _w809_ ;
	assign \g31863_pad  = _w810_ ;
	assign \g32185_pad  = _w815_ ;
	assign \g33079_pad  = _w818_ ;
	assign \g33435_pad  = _w821_ ;
	assign \g33959_pad  = _w827_ ;
	assign \g34435_pad  = _w832_ ;
	assign \g34788_pad  = _w834_ ;
	assign \g34956_pad  = _w836_ ;
	assign \g34_reg/P0001  = _w490_ ;
	assign \g35_syn_2  = _w495_ ;
	assign \g37/_0_  = _w878_ ;
	assign \g41/_0_  = _w907_ ;
	assign \g60853/_3_  = _w915_ ;
	assign \g60856/_3_  = _w918_ ;
	assign \g60879/_3_  = _w919_ ;
	assign \g60882/_0_  = _w923_ ;
	assign \g60888/_0_  = _w924_ ;
	assign \g60891/_0_  = _w925_ ;
	assign \g60896/_0_  = _w926_ ;
	assign \g60899/_0_  = _w936_ ;
	assign \g60900/_3_  = _w940_ ;
	assign \g60909/_3_  = _w943_ ;
	assign \g60911/_0_  = _w944_ ;
	assign \g60915/_0_  = _w945_ ;
	assign \g60918/_0_  = _w961_ ;
	assign \g60919/_0_  = _w969_ ;
	assign \g60928/_0_  = _w973_ ;
	assign \g60929/_0_  = _w974_ ;
	assign \g60936/_0_  = _w977_ ;
	assign \g60937/_0_  = _w984_ ;
	assign \g60939/_0_  = _w991_ ;
	assign \g60940/_0_  = _w999_ ;
	assign \g60941/_0_  = _w1005_ ;
	assign \g60942/_0_  = _w1011_ ;
	assign \g60943/_0_  = _w1017_ ;
	assign \g60944/_0_  = _w1018_ ;
	assign \g60952/_0_  = _w1025_ ;
	assign \g60954/_0_  = _w1030_ ;
	assign \g60958/_0_  = _w1035_ ;
	assign \g60962/_3_  = _w1038_ ;
	assign \g60972/_0_  = _w1044_ ;
	assign \g60980/_0_  = _w1052_ ;
	assign \g60984/_0_  = _w1053_ ;
	assign \g60986/_0_  = _w1054_ ;
	assign \g60989/_0_  = _w1061_ ;
	assign \g60991/_3_  = _w1066_ ;
	assign \g61006/_0_  = _w1070_ ;
	assign \g61008/_0_  = _w1078_ ;
	assign \g61013/_0_  = _w1086_ ;
	assign \g61014/_0_  = _w1092_ ;
	assign \g61015/_0_  = _w1098_ ;
	assign \g61016/_0_  = _w1104_ ;
	assign \g61017/_0_  = _w1105_ ;
	assign \g61026/_3_  = _w1109_ ;
	assign \g61027/_3_  = _w1110_ ;
	assign \g61030/_0_  = _w1114_ ;
	assign \g61031/_0_  = _w1117_ ;
	assign \g61037/_0_  = _w1123_ ;
	assign \g61038/_0_  = _w1126_ ;
	assign \g61042/_0_  = _w1143_ ;
	assign \g61044/_0_  = _w1159_ ;
	assign \g61045/_0_  = _w1175_ ;
	assign \g61046/_0_  = _w1191_ ;
	assign \g61050/_0_  = _w1193_ ;
	assign \g61051/_0_  = _w1195_ ;
	assign \g61052/_0_  = _w1199_ ;
	assign \g61078/_0_  = _w1200_ ;
	assign \g61131/_0_  = _w1201_ ;
	assign \g61137/_3_  = _w1205_ ;
	assign \g61142/_3_  = _w1206_ ;
	assign \g61143/_3_  = _w1207_ ;
	assign \g61151/_0_  = _w1224_ ;
	assign \g61152/_0_  = _w1240_ ;
	assign \g61161/_0_  = _w1256_ ;
	assign \g61168/_3_  = _w1260_ ;
	assign \g61169/_3_  = _w1265_ ;
	assign \g61170/_0_  = _w1275_ ;
	assign \g61171/_3_  = _w1283_ ;
	assign \g61172/_0_  = _w1292_ ;
	assign \g61173/_0_  = _w1301_ ;
	assign \g61174/_0_  = _w1307_ ;
	assign \g61175/_0_  = _w1312_ ;
	assign \g61176/_0_  = _w1322_ ;
	assign \g61177/_3_  = _w1330_ ;
	assign \g61178/_0_  = _w1339_ ;
	assign \g61179/_0_  = _w1348_ ;
	assign \g61180/_0_  = _w1354_ ;
	assign \g61181/_0_  = _w1359_ ;
	assign \g61182/_3_  = _w1362_ ;
	assign \g61183/_0_  = _w1372_ ;
	assign \g61184/_3_  = _w1380_ ;
	assign \g61185/_0_  = _w1389_ ;
	assign \g61186/_0_  = _w1398_ ;
	assign \g61187/_0_  = _w1404_ ;
	assign \g61188/_0_  = _w1409_ ;
	assign \g61189/_0_  = _w1419_ ;
	assign \g61190/_3_  = _w1427_ ;
	assign \g61191/_0_  = _w1436_ ;
	assign \g61192/_0_  = _w1444_ ;
	assign \g61193/_0_  = _w1450_ ;
	assign \g61194/_0_  = _w1456_ ;
	assign \g61221/_0_  = _w1457_ ;
	assign \g61222/_0_  = _w1464_ ;
	assign \g61223/_3_  = _w1467_ ;
	assign \g61224/_3_  = _w1468_ ;
	assign \g61261/_0_  = _w1469_ ;
	assign \g61295/_3_  = _w1473_ ;
	assign \g61308/_0_  = _w1477_ ;
	assign \g61316/_0_  = _w1479_ ;
	assign \g61327/_0_  = _w1484_ ;
	assign \g61329/_0_  = _w1490_ ;
	assign \g61330/_0_  = _w1491_ ;
	assign \g61331/_0_  = _w1501_ ;
	assign \g61332/_3_  = _w1509_ ;
	assign \g61333/_0_  = _w1518_ ;
	assign \g61334/_0_  = _w1527_ ;
	assign \g61335/_0_  = _w1533_ ;
	assign \g61336/_0_  = _w1538_ ;
	assign \g61337/_0_  = _w1548_ ;
	assign \g61338/_3_  = _w1556_ ;
	assign \g61339/_0_  = _w1565_ ;
	assign \g61340/_0_  = _w1574_ ;
	assign \g61341/_0_  = _w1580_ ;
	assign \g61342/_0_  = _w1585_ ;
	assign \g61343/_0_  = _w1595_ ;
	assign \g61344/_3_  = _w1603_ ;
	assign \g61345/_0_  = _w1612_ ;
	assign \g61346/_0_  = _w1618_ ;
	assign \g61347/_0_  = _w1624_ ;
	assign \g61348/_0_  = _w1632_ ;
	assign \g61349/_0_  = _w1644_ ;
	assign \g61350/_3_  = _w1653_ ;
	assign \g61351/_0_  = _w1662_ ;
	assign \g61352/_0_  = _w1668_ ;
	assign \g61353/_0_  = _w1674_ ;
	assign \g61354/_0_  = _w1681_ ;
	assign \g61367/_0_  = _w1686_ ;
	assign \g61372/_0_  = _w1687_ ;
	assign \g61373/_0_  = _w1706_ ;
	assign \g61375/_0_  = _w1724_ ;
	assign \g61382/_0_  = _w1725_ ;
	assign \g61385/_3_  = _w1728_ ;
	assign \g61386/_0_  = _w1734_ ;
	assign \g61399/_0_  = _w1735_ ;
	assign \g61400/_0_  = _w1742_ ;
	assign \g61402/_0_  = _w1743_ ;
	assign \g61405/_0_  = _w1744_ ;
	assign \g61435/_3_  = _w1748_ ;
	assign \g61449/_0_  = _w1760_ ;
	assign \g61468/_0_  = _w1769_ ;
	assign \g61475/_0_  = _w1774_ ;
	assign \g61480/_0_  = _w1779_ ;
	assign \g61482/_0_  = _w1784_ ;
	assign \g61483/_0_  = _w1790_ ;
	assign \g61484/_0_  = _w1806_ ;
	assign \g61486/_3_  = _w1809_ ;
	assign \g61494/_0_  = _w1810_ ;
	assign \g61496/_0_  = _w1816_ ;
	assign \g61497/_0_  = _w1822_ ;
	assign \g61514/_0_  = _w1823_ ;
	assign \g61517/_0_  = _w1833_ ;
	assign \g61519/_3_  = _w1855_ ;
	assign \g61520/_3_  = _w1876_ ;
	assign \g61527/_0_  = _w1877_ ;
	assign \g61541/_0_  = _w1885_ ;
	assign \g61544/_0_  = _w1892_ ;
	assign \g61550/_0_  = _w1893_ ;
	assign \g61551/_0_  = _w1894_ ;
	assign \g61554/_0_  = _w1899_ ;
	assign \g61556/_3_  = _w1906_ ;
	assign \g61567/_0_  = _w1914_ ;
	assign \g61571/_0_  = _w1919_ ;
	assign \g61574/_0_  = _w1923_ ;
	assign \g61587/_0_  = _w1926_ ;
	assign \g61592/_0_  = _w1932_ ;
	assign \g61632/_0_  = _w1938_ ;
	assign \g61634/_0_  = _w1950_ ;
	assign \g61635/_0_  = _w1956_ ;
	assign \g61639/_0_  = _w1967_ ;
	assign \g61644/_0_  = _w1970_ ;
	assign \g61652/_3_  = _w1979_ ;
	assign \g61709/_0_  = _w1984_ ;
	assign \g61714/_0_  = _w1988_ ;
	assign \g61720/_0_  = _w1993_ ;
	assign \g61721/_0_  = _w1997_ ;
	assign \g61723/_0_  = _w2001_ ;
	assign \g61725/_0_  = _w2005_ ;
	assign \g61726/_0_  = _w2009_ ;
	assign \g61734/_0_  = _w2020_ ;
	assign \g61739/_0_  = _w2034_ ;
	assign \g61744/_0_  = _w2036_ ;
	assign \g61746/_3_  = _w2037_ ;
	assign \g61747/_3_  = _w2041_ ;
	assign \g61748/_3_  = _w2042_ ;
	assign \g61750/u3_syn_7  = _w2043_ ;
	assign \g61802/_0_  = _w2052_ ;
	assign \g61804/_0_  = _w2067_ ;
	assign \g61808/_0_  = _w2074_ ;
	assign \g61811/_0_  = _w2084_ ;
	assign \g61816/_0_  = _w2095_ ;
	assign \g61818/_0_  = _w2101_ ;
	assign \g61820/_0_  = _w2108_ ;
	assign \g61823/_0_  = _w2112_ ;
	assign \g61824/_0_  = _w2118_ ;
	assign \g61841/_0_  = _w2121_ ;
	assign \g61842/_3_  = _w2123_ ;
	assign \g61844/_3_  = _w2132_ ;
	assign \g61845/_3_  = _w2135_ ;
	assign \g61846/_3_  = _w2142_ ;
	assign \g61847/u3_syn_7  = _w2143_ ;
	assign \g61848/_0_  = _w2150_ ;
	assign \g61849/_3_  = _w2153_ ;
	assign \g61850/_0_  = _w2160_ ;
	assign \g61851/u3_syn_7  = _w2161_ ;
	assign \g61852/_0_  = _w2169_ ;
	assign \g61853/_3_  = _w2175_ ;
	assign \g61854/_3_  = _w2178_ ;
	assign \g61855/_0_  = _w2185_ ;
	assign \g61856/u3_syn_7  = _w2186_ ;
	assign \g61857/_0_  = _w2191_ ;
	assign \g61858/_3_  = _w2198_ ;
	assign \g61859/_3_  = _w2201_ ;
	assign \g61860/u3_syn_7  = _w2202_ ;
	assign \g61861/_0_  = _w2209_ ;
	assign \g61862/_3_  = _w2217_ ;
	assign \g61863/_3_  = _w2220_ ;
	assign \g61864/u3_syn_7  = _w2221_ ;
	assign \g61865/_0_  = _w2228_ ;
	assign \g61866/_3_  = _w2235_ ;
	assign \g61867/_3_  = _w2238_ ;
	assign \g61868/u3_syn_7  = _w2239_ ;
	assign \g61869/_0_  = _w2246_ ;
	assign \g61870/_0_  = _w2252_ ;
	assign \g61871/_3_  = _w2259_ ;
	assign \g61872/_3_  = _w2262_ ;
	assign \g61873/u3_syn_7  = _w2263_ ;
	assign \g61874/_0_  = _w2270_ ;
	assign \g61875/_0_  = _w2275_ ;
	assign \g61877/_3_  = _w2282_ ;
	assign \g61878/_3_  = _w2285_ ;
	assign \g61879/u3_syn_7  = _w2286_ ;
	assign \g61880/_0_  = _w2293_ ;
	assign \g61881/_0_  = _w2298_ ;
	assign \g61882/_0_  = _w2303_ ;
	assign \g61883/_0_  = _w2308_ ;
	assign \g61884/_0_  = _w2313_ ;
	assign \g61914/_0_  = _w2316_ ;
	assign \g61915/_0_  = _w2320_ ;
	assign \g61917/_0_  = _w2332_ ;
	assign \g61918/_0_  = _w2334_ ;
	assign \g61922/_0_  = _w2340_ ;
	assign \g61923/_0_  = _w2346_ ;
	assign \g61924/_0_  = _w2353_ ;
	assign \g61932/_0_  = _w2362_ ;
	assign \g61936/_0_  = _w2369_ ;
	assign \g61945/_0_  = _w2373_ ;
	assign \g61947/_0_  = _w2375_ ;
	assign \g61959/_0_  = _w2381_ ;
	assign \g61960/_0_  = _w2386_ ;
	assign \g61962/_0_  = _w2391_ ;
	assign \g61973/_3_  = _w2397_ ;
	assign \g61974/u3_syn_7  = _w2396_ ;
	assign \g61975/_3_  = _w2409_ ;
	assign \g61976/u3_syn_7  = _w2411_ ;
	assign \g61977/_3_  = _w2417_ ;
	assign \g61978/_3_  = _w2429_ ;
	assign \g61979/u3_syn_7  = _w2431_ ;
	assign \g61980/_3_  = _w2437_ ;
	assign \g61981/_3_  = _w2449_ ;
	assign \g61982/_3_  = _w2453_ ;
	assign \g61983/u3_syn_7  = _w2455_ ;
	assign \g61984/_3_  = _w2461_ ;
	assign \g61985/_3_  = _w2473_ ;
	assign \g61986/u3_syn_7  = _w2475_ ;
	assign \g61987/_3_  = _w2479_ ;
	assign \g61988/_3_  = _w2491_ ;
	assign \g61989/u3_syn_7  = _w2493_ ;
	assign \g61990/_3_  = _w2499_ ;
	assign \g61991/_3_  = _w2511_ ;
	assign \g61992/u3_syn_7  = _w2513_ ;
	assign \g61993/_3_  = _w2519_ ;
	assign \g61994/u3_syn_7  = _w2521_ ;
	assign \g61995/_3_  = _w2533_ ;
	assign \g61996/_3_  = _w2539_ ;
	assign \g61997/_3_  = _w2551_ ;
	assign \g62022/_0_  = _w2556_ ;
	assign \g62028/_0_  = _w2561_ ;
	assign \g62029/_0_  = _w2562_ ;
	assign \g62031/_0_  = _w2578_ ;
	assign \g62033/_0_  = _w2583_ ;
	assign \g62038/_0_  = _w2588_ ;
	assign \g62042/_0_  = _w2593_ ;
	assign \g62046/_0_  = _w2598_ ;
	assign \g62048/_0_  = _w2604_ ;
	assign \g62049/_0_  = _w2609_ ;
	assign \g62051/_0_  = _w2614_ ;
	assign \g62053/_0_  = _w2622_ ;
	assign \g62085/_0_  = _w2627_ ;
	assign \g62101/_0_  = _w2633_ ;
	assign \g62102/_0_  = _w2640_ ;
	assign \g62103/_0_  = _w2644_ ;
	assign \g62105/_0_  = _w2646_ ;
	assign \g62108/_3_  = _w2648_ ;
	assign \g62112/_0_  = _w2654_ ;
	assign \g62137/_3_  = _w2660_ ;
	assign \g62207/_0_  = _w2662_ ;
	assign \g62239/_0_  = _w2675_ ;
	assign \g62240/_0_  = _w2680_ ;
	assign \g62267/_0_  = _w2686_ ;
	assign \g62273/_0_  = _w2691_ ;
	assign \g62284/_0_  = _w2695_ ;
	assign \g62291/_0_  = _w2698_ ;
	assign \g62293/_0_  = _w2701_ ;
	assign \g62298/_0_  = _w2706_ ;
	assign \g62303/_3_  = _w2717_ ;
	assign \g62322/_3_  = _w2724_ ;
	assign \g62323/_3_  = _w2725_ ;
	assign \g62324/_3_  = _w2728_ ;
	assign \g62325/_3_  = _w2732_ ;
	assign \g62583/_0_  = _w2740_ ;
	assign \g62598/_0_  = _w2744_ ;
	assign \g62609/_0_  = _w2751_ ;
	assign \g62636/_0_  = _w2764_ ;
	assign \g62646/_0_  = _w2768_ ;
	assign \g62649/_0_  = _w2771_ ;
	assign \g62658/_0_  = _w2776_ ;
	assign \g62663/_0_  = _w2778_ ;
	assign \g62664/_0_  = _w2780_ ;
	assign \g62667/_0_  = _w2785_ ;
	assign \g62676/_0_  = _w2789_ ;
	assign \g62677/_0_  = _w2792_ ;
	assign \g62678/_3_  = _w2796_ ;
	assign \g62679/_0_  = _w2797_ ;
	assign \g62687/u3_syn_7  = _w2798_ ;
	assign \g62688/u3_syn_7  = _w2799_ ;
	assign \g62689/_0_  = _w2806_ ;
	assign \g62690/_3_  = _w2809_ ;
	assign \g62691/_3_  = _w2814_ ;
	assign \g62693/_0_  = _w2821_ ;
	assign \g62694/_3_  = _w2827_ ;
	assign \g62695/_3_  = _w2834_ ;
	assign \g62696/_3_  = _w2841_ ;
	assign \g62697/_3_  = _w2848_ ;
	assign \g62698/_3_  = _w2851_ ;
	assign \g62699/_3_  = _w2857_ ;
	assign \g62700/_3_  = _w2863_ ;
	assign \g62701/_3_  = _w2869_ ;
	assign \g62702/_3_  = _w2875_ ;
	assign \g62703/_3_  = _w2880_ ;
	assign \g62704/u3_syn_7  = _w2876_ ;
	assign \g62705/_0_  = _w2887_ ;
	assign \g62706/_3_  = _w2890_ ;
	assign \g62707/_3_  = _w2895_ ;
	assign \g62708/u3_syn_7  = _w2891_ ;
	assign \g62709/_0_  = _w2902_ ;
	assign \g62710/_3_  = _w2905_ ;
	assign \g62711/_3_  = _w2910_ ;
	assign \g62712/u3_syn_7  = _w2906_ ;
	assign \g62713/_0_  = _w2917_ ;
	assign \g62714/_3_  = _w2920_ ;
	assign \g62715/_0_  = _w2925_ ;
	assign \g62716/u3_syn_7  = _w2921_ ;
	assign \g62717/_0_  = _w2932_ ;
	assign \g62718/_3_  = _w2935_ ;
	assign \g62719/_0_  = _w2940_ ;
	assign \g62720/u3_syn_7  = _w2936_ ;
	assign \g62721/_0_  = _w2947_ ;
	assign \g62722/_3_  = _w2950_ ;
	assign \g62723/_0_  = _w2955_ ;
	assign \g62724/u3_syn_7  = _w2951_ ;
	assign \g62725/_0_  = _w2962_ ;
	assign \g62726/_3_  = _w2965_ ;
	assign \g62728/_0_  = _w2969_ ;
	assign \g62790/_0_  = _w2978_ ;
	assign \g62791/_0_  = _w2984_ ;
	assign \g62793/_0_  = _w2990_ ;
	assign \g62794/_0_  = _w2996_ ;
	assign \g62795/_0_  = _w3002_ ;
	assign \g62796/_0_  = _w3008_ ;
	assign \g62797/_0_  = _w3014_ ;
	assign \g62807/_0_  = _w3021_ ;
	assign \g62823/_0_  = _w3022_ ;
	assign \g62824/_0_  = _w3025_ ;
	assign \g62833/_0_  = _w3029_ ;
	assign \g62846/_0_  = _w3033_ ;
	assign \g62859/_0_  = _w3039_ ;
	assign \g62860/_0_  = _w3045_ ;
	assign \g62897/_0_  = _w3048_ ;
	assign \g62898/_0_  = _w3053_ ;
	assign \g62922/_3_  = _w3054_ ;
	assign \g62923/_0_  = _w3056_ ;
	assign \g62927/_0_  = _w3060_ ;
	assign \g62938/_3_  = _w3063_ ;
	assign \g62939/_3_  = _w3069_ ;
	assign \g62940/_3_  = _w3072_ ;
	assign \g62941/u3_syn_7  = _w3075_ ;
	assign \g62942/_0_  = _w3084_ ;
	assign \g62943/_3_  = _w3087_ ;
	assign \g62987/_3_  = _w3090_ ;
	assign \g62991/_3_  = _w3094_ ;
	assign \g63015/u3_syn_7  = _w3098_ ;
	assign \g63016/_0_  = _w3105_ ;
	assign \g63017/_3_  = _w3114_ ;
	assign \g63018/_3_  = _w3121_ ;
	assign \g63019/_3_  = _w3124_ ;
	assign \g63020/_3_  = _w3129_ ;
	assign \g63021/_3_  = _w3136_ ;
	assign \g63022/_3_  = _w3140_ ;
	assign \g63025/_3_  = _w3144_ ;
	assign \g63026/_3_  = _w3148_ ;
	assign \g63027/_3_  = _w3152_ ;
	assign \g63029/_3_  = _w3156_ ;
	assign \g63030/_3_  = _w3160_ ;
	assign \g63031/_3_  = _w3164_ ;
	assign \g63033/_3_  = _w3168_ ;
	assign \g63034/_3_  = _w3172_ ;
	assign \g63043/_3_  = _w3179_ ;
	assign \g63044/_3_  = _w3183_ ;
	assign \g63051/_3_  = _w3187_ ;
	assign \g63057/_3_  = _w3191_ ;
	assign \g63068/_3_  = _w3195_ ;
	assign \g63070/_3_  = _w3199_ ;
	assign \g63073/_3_  = _w3203_ ;
	assign \g63081/_3_  = _w3206_ ;
	assign \g63082/_3_  = _w3210_ ;
	assign \g63083/u3_syn_7  = _w3211_ ;
	assign \g63084/_3_  = _w3214_ ;
	assign \g63085/_0_  = _w3225_ ;
	assign \g63086/_3_  = _w3228_ ;
	assign \g63107/_3_  = _w3231_ ;
	assign \g63108/u3_syn_7  = _w3233_ ;
	assign \g63109/u3_syn_7  = _w3237_ ;
	assign \g63110/_0_  = _w3244_ ;
	assign \g63111/_3_  = _w3247_ ;
	assign \g63132/_3_  = _w3250_ ;
	assign \g63133/_3_  = _w3254_ ;
	assign \g63134/_3_  = _w3256_ ;
	assign \g63135/_3_  = _w3257_ ;
	assign \g63136/_3_  = _w3260_ ;
	assign \g63137/_3_  = _w3264_ ;
	assign \g63138/_3_  = _w3268_ ;
	assign \g63139/u3_syn_7  = _w3269_ ;
	assign \g63140/_3_  = _w3272_ ;
	assign \g63141/_3_  = _w3276_ ;
	assign \g63142/_3_  = _w3283_ ;
	assign \g63143/_3_  = _w3287_ ;
	assign \g63144/_3_  = _w3293_ ;
	assign \g63145/_3_  = _w3297_ ;
	assign \g63146/u3_syn_7  = _w3299_ ;
	assign \g63198/_0_  = _w3304_ ;
	assign \g63205/_0_  = _w3309_ ;
	assign \g63208/_0_  = _w3312_ ;
	assign \g63212/_0_  = _w3316_ ;
	assign \g63215/_0_  = _w3321_ ;
	assign \g63219/_0_  = _w3326_ ;
	assign \g63244/_0_  = _w3332_ ;
	assign \g63246/_0_  = _w3333_ ;
	assign \g63254/_0_  = _w3334_ ;
	assign \g63255/_0_  = _w3342_ ;
	assign \g63272/_0_  = _w3346_ ;
	assign \g63276/_0_  = _w3348_ ;
	assign \g63278/_0_  = _w3352_ ;
	assign \g63279/_0_  = _w3355_ ;
	assign \g63280/_0_  = _w3357_ ;
	assign \g63327/_0_  = _w3360_ ;
	assign \g63345/_0_  = _w3363_ ;
	assign \g63346/_3_  = _w3364_ ;
	assign \g63347/_3_  = _w3371_ ;
	assign \g63354/_3_  = _w3375_ ;
	assign \g63358/_3_  = _w3381_ ;
	assign \g63359/u3_syn_7  = _w3382_ ;
	assign \g63361/_3_  = _w3387_ ;
	assign \g63365/_3_  = _w3391_ ;
	assign \g63366/_3_  = _w3395_ ;
	assign \g63367/_3_  = _w3399_ ;
	assign \g63368/_3_  = _w3400_ ;
	assign \g63370/_3_  = _w3404_ ;
	assign \g63479/_0_  = _w3408_ ;
	assign \g63484/_0_  = _w3412_ ;
	assign \g63499/_1_  = _w1478_ ;
	assign \g63520/_0_  = _w3415_ ;
	assign \g63523/_0_  = _w3418_ ;
	assign \g63526/_0_  = _w3423_ ;
	assign \g63538/_0_  = _w3424_ ;
	assign \g63539/_0_  = _w3432_ ;
	assign \g63541/_0_  = _w3433_ ;
	assign \g63555/_0_  = _w3440_ ;
	assign \g63642/_0_  = _w3447_ ;
	assign \g63645/_0_  = _w3450_ ;
	assign \g63648/_3_  = _w3455_ ;
	assign \g63777/_3_  = _w3458_ ;
	assign \g63778/_3_  = _w3464_ ;
	assign \g63781/_0_  = _w3466_ ;
	assign \g63786/u3_syn_7  = _w3467_ ;
	assign \g63787/_3_  = _w3468_ ;
	assign \g63788/_3_  = _w3469_ ;
	assign \g63790/_3_  = _w3472_ ;
	assign \g63791/_3_  = _w3478_ ;
	assign \g63792/u3_syn_7  = _w3465_ ;
	assign \g63794/_0_  = _w3485_ ;
	assign \g63795/_0_  = _w3492_ ;
	assign \g63796/_0_  = _w3498_ ;
	assign \g63798/_3_  = _w3500_ ;
	assign \g63800/_3_  = _w3503_ ;
	assign \g63804/_3_  = _w3507_ ;
	assign \g63805/_3_  = _w3510_ ;
	assign \g63806/_3_  = _w3511_ ;
	assign \g63807/_3_  = _w3514_ ;
	assign \g63808/_3_  = _w3518_ ;
	assign \g63809/_3_  = _w3523_ ;
	assign \g63870/_0_  = _w3527_ ;
	assign \g63883/_0_  = _w3528_ ;
	assign \g63934/_0_  = _w3531_ ;
	assign \g63936/_0_  = _w3532_ ;
	assign \g63938/_0_  = _w3534_ ;
	assign \g63939/_0_  = _w3537_ ;
	assign \g63966/_0_  = _w3543_ ;
	assign \g63970/_0_  = _w3549_ ;
	assign \g63999/_0_  = _w3553_ ;
	assign \g64039/_0_  = _w3557_ ;
	assign \g64040/_0_  = _w3562_ ;
	assign \g64043/_0_  = _w3563_ ;
	assign \g64062/_3_  = _w3564_ ;
	assign \g64078/_0_  = _w3565_ ;
	assign \g64091/_0_  = _w3568_ ;
	assign \g64095/_3_  = _w3571_ ;
	assign \g64096/_3_  = _w3573_ ;
	assign \g64097/u3_syn_7  = _w3574_ ;
	assign \g64098/u3_syn_7  = _w3575_ ;
	assign \g64099/u3_syn_7  = _w3576_ ;
	assign \g64100/u3_syn_7  = _w3577_ ;
	assign \g64134/_0_  = _w3581_ ;
	assign \g64135/_0_  = _w3585_ ;
	assign \g64153/_0_  = _w3588_ ;
	assign \g64155/_0_  = _w3591_ ;
	assign \g64179/_0_  = _w3595_ ;
	assign \g64229/_0_  = _w3599_ ;
	assign \g64235/_0_  = _w3603_ ;
	assign \g64236/_0_  = _w3607_ ;
	assign \g64280/_0_  = _w3614_ ;
	assign \g64315/_0_  = _w3616_ ;
	assign \g64365/_0_  = _w3618_ ;
	assign \g64426/_3_  = _w3619_ ;
	assign \g64438/_3_  = _w3620_ ;
	assign \g64442/u3_syn_7  = _w3621_ ;
	assign \g64445/_3_  = _w3622_ ;
	assign \g64447/_3_  = _w3625_ ;
	assign \g64449/_3_  = _w3626_ ;
	assign \g64451/_3_  = _w3633_ ;
	assign \g64453/_3_  = _w3636_ ;
	assign \g64454/_3_  = _w3637_ ;
	assign \g64460/_3_  = _w3642_ ;
	assign \g64461/_3_  = _w3646_ ;
	assign \g64510/_0_  = _w3647_ ;
	assign \g64527/_0_  = _w3651_ ;
	assign \g64528/_0_  = _w3652_ ;
	assign \g64544/_0_  = _w3654_ ;
	assign \g64549/_0_  = _w3656_ ;
	assign \g64566/_0_  = _w3658_ ;
	assign \g64576/_0_  = _w3661_ ;
	assign \g64602/_0_  = _w3662_ ;
	assign \g64691/_0_  = _w3665_ ;
	assign \g64697/_0_  = _w3669_ ;
	assign \g64707/_3_  = _w3672_ ;
	assign \g64778/_3_  = _w3673_ ;
	assign \g64790/_3_  = _w3676_ ;
	assign \g64791/_3_  = _w3678_ ;
	assign \g64792/_3_  = _w3679_ ;
	assign \g64793/_3_  = _w3680_ ;
	assign \g64794/_3_  = _w3681_ ;
	assign \g64795/_3_  = _w3682_ ;
	assign \g64796/_3_  = _w3683_ ;
	assign \g64797/_3_  = _w3684_ ;
	assign \g64877/_0_  = _w3685_ ;
	assign \g64912/_0_  = _w3688_ ;
	assign \g64973/_0_  = _w3690_ ;
	assign \g65047/_3_  = _w3691_ ;
	assign \g65081/_3_  = _w3692_ ;
	assign \g65088/_3_  = _w3693_ ;
	assign \g65097/_3_  = _w3694_ ;
	assign \g65100/_3_  = _w3695_ ;
	assign \g65101/_3_  = _w3696_ ;
	assign \g65104/_3_  = _w3697_ ;
	assign \g65105/_3_  = _w3698_ ;
	assign \g65107/_3_  = _w3699_ ;
	assign \g65110/_3_  = _w3700_ ;
	assign \g65111/_3_  = _w3703_ ;
	assign \g65113/_3_  = _w3706_ ;
	assign \g65114/_3_  = _w3709_ ;
	assign \g65266/_0_  = _w3710_ ;
	assign \g65267/_0_  = _w3711_ ;
	assign \g65294/_1_  = _w3586_ ;
	assign \g65328/_1_  = _w3712_ ;
	assign \g65495/_0_  = _w3713_ ;
	assign \g65499/_0_  = _w3714_ ;
	assign \g65503/_0_  = _w3715_ ;
	assign \g65529/_0_  = _w3716_ ;
	assign \g65530/_3_  = _w3717_ ;
	assign \g65531/_3_  = _w3718_ ;
	assign \g65532/_3_  = _w3719_ ;
	assign \g65533/_3_  = _w3720_ ;
	assign \g65624/_0_  = _w3721_ ;
	assign \g65625/_1_  = _w3200_ ;
	assign \g65641/_0_  = _w3722_ ;
	assign \g65701/_0_  = _w3723_ ;
	assign \g65704/_0_  = _w3724_ ;
	assign \g65853/_0_  = _w3725_ ;
	assign \g65891/_0_  = _w3726_ ;
	assign \g65901/_0_  = _w3727_ ;
	assign \g65986/_0_  = _w3728_ ;
	assign \g66029/_0_  = _w3729_ ;
	assign \g66066/_0_  = _w3730_ ;
	assign \g66067/_0_  = _w3731_ ;
	assign \g66068/_0_  = _w3732_ ;
	assign \g66154/_3_  = _w3733_ ;
	assign \g66362/_0_  = _w3734_ ;
	assign \g66369/_0_  = _w3735_ ;
	assign \g66398/_0_  = _w3736_ ;
	assign \g66409/_0_  = _w3737_ ;
	assign \g66419/_0_  = _w3738_ ;
	assign \g66439/_0_  = _w3739_ ;
	assign \g66443/_0_  = _w3740_ ;
	assign \g66464/_0_  = _w3741_ ;
	assign \g66471/_0_  = _w3742_ ;
	assign \g66512/_0_  = _w3743_ ;
	assign \g66528/_0_  = _w3744_ ;
	assign \g66541/_0_  = _w3499_ ;
	assign \g66558/_0_  = _w3745_ ;
	assign \g66644/_0_  = _w3746_ ;
	assign \g66684/_0_  = _w3747_ ;
	assign \g66697/_0_  = _w3748_ ;
	assign \g66698/_0_  = _w3689_ ;
	assign \g66701/_0_  = _w3749_ ;
	assign \g66714/_0_  = _w3750_ ;
	assign \g66715/_0_  = _w3751_ ;
	assign \g66745/_0_  = _w3752_ ;
	assign \g66750/_0_  = _w3753_ ;
	assign \g66751/_0_  = _w3754_ ;
	assign \g66810/_0_  = _w3755_ ;
	assign \g66844/_0_  = _w3756_ ;
	assign \g66853/_0_  = _w3757_ ;
	assign \g66897/_0_  = _w3758_ ;
	assign \g66905/_0_  = _w3759_ ;
	assign \g69743/_0_  = _w3765_ ;
	assign \g69750/_0_  = _w3771_ ;
	assign \g69773/_1_  = _w3774_ ;
	assign \g69792/_1_  = _w3780_ ;
	assign \g69858/_0_  = _w3786_ ;
	assign \g69938/_0_  = _w3798_ ;
	assign \g69949/_0_  = _w3804_ ;
	assign \g70167/_0_  = _w3809_ ;
	assign \g71190/_0_  = _w3815_ ;
	assign \g71198/_0_  = _w3822_ ;
	assign \g71284/_0_  = _w3838_ ;
	assign \g72369/_1_  = _w3284_ ;
	assign \g72467/_0_  = _w3844_ ;
	assign \g72476/_0_  = _w3858_ ;
	assign \g72477/_1_  = _w3859_ ;
	assign \g72648/_0_  = _w3865_ ;
	assign \g72741/_0_  = _w3871_ ;
	assign \g72772/_0_  = _w3873_ ;
	assign \g8132_pad  = 1'b0;
endmodule;