module top (\a0_pad , \a1_pad , \a2_pad , a_pad, \b0_pad , \b1_pad , \b2_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \d0_pad , \d1_pad , \d2_pad , \e0_pad , \e1_pad , \e2_pad , \f0_pad , \f1_pad , \f2_pad , \g0_pad , \g1_pad , \g2_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , h_pad, \i0_pad , \i1_pad , \i2_pad , i_pad, \j1_pad , \j2_pad , \k0_pad , \k1_pad , \k2_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , o_pad, \p0_pad , \p1_pad , \p2_pad , p_pad, \q0_pad , \q1_pad , \q2_pad , q_pad, \r0_pad , \r1_pad , \r2_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , v_pad, \w0_pad , \w1_pad , w_pad, \x0_pad , \x1_pad , x_pad, \y0_pad , \y1_pad , y_pad, \z0_pad , \z1_pad , z_pad, \a3_pad , \a4_pad , \a5_pad , \b3_pad , \b4_pad , \b5_pad , \c3_pad , \c4_pad , \c5_pad , \d3_pad , \d4_pad , \d5_pad , \e3_pad , \e4_pad , \e5_pad , \f3_pad , \f4_pad , \f5_pad , \g3_pad , \g4_pad , \g5_pad , \h3_pad , \h4_pad , \h5_pad , \i3_pad , \i4_pad , \i5_pad , \j3_pad , \j4_pad , \j5_pad , \k3_pad , \k4_pad , \k5_pad , \l3_pad , \l4_pad , \l5_pad , \m3_pad , \m4_pad , \m5_pad , \n3_pad , \n4_pad , \n5_pad , \o3_pad , \o4_pad , \o5_pad , \p3_pad , \p4_pad , \q3_pad , \q4_pad , \r3_pad , \r4_pad , \s3_pad , \s4_pad , \t3_pad , \t4_pad , \u3_pad , \u4_pad , \v3_pad , \v4_pad , \w2_pad , \w3_pad , \w4_pad , \x2_pad , \x3_pad , \x4_pad , \y2_pad , \y3_pad , \y4_pad , \z2_pad , \z3_pad , \z4_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \e0_pad  ;
	input \e1_pad  ;
	input \e2_pad  ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input i_pad ;
	input \j1_pad  ;
	input \j2_pad  ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input \p1_pad  ;
	input \p2_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input \q1_pad  ;
	input \q2_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input \r1_pad  ;
	input \r2_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input x_pad ;
	input \y0_pad  ;
	input \y1_pad  ;
	input y_pad ;
	input \z0_pad  ;
	input \z1_pad  ;
	input z_pad ;
	output \a3_pad  ;
	output \a4_pad  ;
	output \a5_pad  ;
	output \b3_pad  ;
	output \b4_pad  ;
	output \b5_pad  ;
	output \c3_pad  ;
	output \c4_pad  ;
	output \c5_pad  ;
	output \d3_pad  ;
	output \d4_pad  ;
	output \d5_pad  ;
	output \e3_pad  ;
	output \e4_pad  ;
	output \e5_pad  ;
	output \f3_pad  ;
	output \f4_pad  ;
	output \f5_pad  ;
	output \g3_pad  ;
	output \g4_pad  ;
	output \g5_pad  ;
	output \h3_pad  ;
	output \h4_pad  ;
	output \h5_pad  ;
	output \i3_pad  ;
	output \i4_pad  ;
	output \i5_pad  ;
	output \j3_pad  ;
	output \j4_pad  ;
	output \j5_pad  ;
	output \k3_pad  ;
	output \k4_pad  ;
	output \k5_pad  ;
	output \l3_pad  ;
	output \l4_pad  ;
	output \l5_pad  ;
	output \m3_pad  ;
	output \m4_pad  ;
	output \m5_pad  ;
	output \n3_pad  ;
	output \n4_pad  ;
	output \n5_pad  ;
	output \o3_pad  ;
	output \o4_pad  ;
	output \o5_pad  ;
	output \p3_pad  ;
	output \p4_pad  ;
	output \q3_pad  ;
	output \q4_pad  ;
	output \r3_pad  ;
	output \r4_pad  ;
	output \s3_pad  ;
	output \s4_pad  ;
	output \t3_pad  ;
	output \t4_pad  ;
	output \u3_pad  ;
	output \u4_pad  ;
	output \v3_pad  ;
	output \v4_pad  ;
	output \w2_pad  ;
	output \w3_pad  ;
	output \w4_pad  ;
	output \x2_pad  ;
	output \x3_pad  ;
	output \x4_pad  ;
	output \y2_pad  ;
	output \y3_pad  ;
	output \y4_pad  ;
	output \z2_pad  ;
	output \z3_pad  ;
	output \z4_pad  ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w154_ ;
	wire _w152_ ;
	wire _w282_ ;
	wire _w25_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w296_ ;
	wire _w39_ ;
	wire _w166_ ;
	wire _w153_ ;
	wire _w292_ ;
	wire _w35_ ;
	wire _w162_ ;
	wire _w122_ ;
	wire _w108_ ;
	wire _w139_ ;
	wire _w278_ ;
	wire _w21_ ;
	wire _w148_ ;
	wire _w102_ ;
	wire _w300_ ;
	wire _w43_ ;
	wire _w170_ ;
	wire _w287_ ;
	wire _w30_ ;
	wire _w157_ ;
	wire _w117_ ;
	wire _w103_ ;
	wire _w143_ ;
	wire _w112_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\f1_pad ,
		_w21_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\g1_pad ,
		_w25_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\h1_pad ,
		_w30_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\i1_pad ,
		_w35_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\j1_pad ,
		_w39_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\k1_pad ,
		_w43_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		\p2_pad ,
		\q2_pad ,
		\r2_pad ,
		_w102_
	);
	LUT3 #(
		.INIT('h20)
	) name7 (
		\e1_pad ,
		\n2_pad ,
		\o2_pad ,
		_w103_
	);
	LUT3 #(
		.INIT('h15)
	) name8 (
		\h1_pad ,
		_w102_,
		_w103_,
		_w104_
	);
	LUT4 #(
		.INIT('h0001)
	) name9 (
		\p2_pad ,
		\q0_pad ,
		\q2_pad ,
		\r2_pad ,
		_w105_
	);
	LUT3 #(
		.INIT('h15)
	) name10 (
		\c1_pad ,
		_w103_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w104_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		g_pad,
		h_pad,
		_w108_
	);
	LUT4 #(
		.INIT('h0004)
	) name13 (
		g_pad,
		\h0_pad ,
		h_pad,
		i_pad,
		_w109_
	);
	LUT4 #(
		.INIT('h8000)
	) name14 (
		\c0_pad ,
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		_w110_
	);
	LUT3 #(
		.INIT('h80)
	) name15 (
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		_w111_
	);
	LUT4 #(
		.INIT('hcce4)
	) name16 (
		\e1_pad ,
		\h2_pad ,
		\i2_pad ,
		\m0_pad ,
		_w112_
	);
	LUT4 #(
		.INIT('h10bb)
	) name17 (
		_w109_,
		_w110_,
		_w111_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\i0_pad ,
		_w113_,
		_w114_
	);
	LUT3 #(
		.INIT('h15)
	) name19 (
		\i1_pad ,
		_w102_,
		_w103_,
		_w115_
	);
	LUT4 #(
		.INIT('h0001)
	) name20 (
		\p2_pad ,
		\q2_pad ,
		\r0_pad ,
		\r2_pad ,
		_w116_
	);
	LUT3 #(
		.INIT('h15)
	) name21 (
		\c1_pad ,
		_w103_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w115_,
		_w117_,
		_w118_
	);
	LUT4 #(
		.INIT('h8000)
	) name23 (
		\d0_pad ,
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		_w119_
	);
	LUT4 #(
		.INIT('hcce4)
	) name24 (
		\e1_pad ,
		\i2_pad ,
		\j2_pad ,
		\m0_pad ,
		_w120_
	);
	LUT4 #(
		.INIT('h04af)
	) name25 (
		_w109_,
		_w111_,
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\i0_pad ,
		_w121_,
		_w122_
	);
	LUT3 #(
		.INIT('h08)
	) name27 (
		\e1_pad ,
		\n2_pad ,
		\o2_pad ,
		_w123_
	);
	LUT4 #(
		.INIT('h3200)
	) name28 (
		i_pad,
		\p2_pad ,
		\q2_pad ,
		\r2_pad ,
		_w124_
	);
	LUT3 #(
		.INIT('h21)
	) name29 (
		\h0_pad ,
		\i0_pad ,
		\t2_pad ,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		\i0_pad ,
		\s2_pad ,
		_w126_
	);
	LUT4 #(
		.INIT('hf780)
	) name31 (
		_w123_,
		_w124_,
		_w125_,
		_w126_,
		_w127_
	);
	LUT3 #(
		.INIT('h15)
	) name32 (
		\j1_pad ,
		_w102_,
		_w103_,
		_w128_
	);
	LUT4 #(
		.INIT('h0001)
	) name33 (
		\p2_pad ,
		\q2_pad ,
		\r2_pad ,
		\s0_pad ,
		_w129_
	);
	LUT3 #(
		.INIT('h15)
	) name34 (
		\c1_pad ,
		_w103_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w128_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		\i0_pad ,
		\m1_pad ,
		_w132_
	);
	LUT4 #(
		.INIT('h2000)
	) name37 (
		\g0_pad ,
		\i0_pad ,
		\m1_pad ,
		\v2_pad ,
		_w133_
	);
	LUT3 #(
		.INIT('h20)
	) name38 (
		\e0_pad ,
		_w109_,
		_w133_,
		_w134_
	);
	LUT4 #(
		.INIT('h3010)
	) name39 (
		\e1_pad ,
		\i0_pad ,
		\j2_pad ,
		\m0_pad ,
		_w135_
	);
	LUT3 #(
		.INIT('hb0)
	) name40 (
		_w109_,
		_w111_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('he)
	) name41 (
		_w134_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\f0_pad ,
		\v2_pad ,
		_w138_
	);
	LUT4 #(
		.INIT('h5450)
	) name43 (
		\c1_pad ,
		\f0_pad ,
		\k0_pad ,
		\v2_pad ,
		_w139_
	);
	LUT3 #(
		.INIT('h40)
	) name44 (
		\c1_pad ,
		\g0_pad ,
		\v2_pad ,
		_w140_
	);
	LUT4 #(
		.INIT('hfdf0)
	) name45 (
		\m1_pad ,
		_w109_,
		_w139_,
		_w140_,
		_w141_
	);
	LUT3 #(
		.INIT('h15)
	) name46 (
		\k1_pad ,
		_w102_,
		_w103_,
		_w142_
	);
	LUT4 #(
		.INIT('h0001)
	) name47 (
		\p2_pad ,
		\q2_pad ,
		\r2_pad ,
		\t0_pad ,
		_w143_
	);
	LUT3 #(
		.INIT('h15)
	) name48 (
		\c1_pad ,
		_w103_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w142_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		b_pad,
		\u0_pad ,
		_w146_
	);
	LUT4 #(
		.INIT('h0031)
	) name51 (
		b_pad,
		\k2_pad ,
		\u0_pad ,
		\u2_pad ,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\c1_pad ,
		\k2_pad ,
		_w148_
	);
	LUT4 #(
		.INIT('h0031)
	) name53 (
		b_pad,
		\c1_pad ,
		\u0_pad ,
		\u2_pad ,
		_w149_
	);
	LUT3 #(
		.INIT('h54)
	) name54 (
		_w147_,
		_w148_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h5444)
	) name55 (
		\c1_pad ,
		\l0_pad ,
		_w102_,
		_w123_,
		_w151_
	);
	LUT4 #(
		.INIT('h5444)
	) name56 (
		\c1_pad ,
		\l1_pad ,
		_w102_,
		_w123_,
		_w152_
	);
	LUT3 #(
		.INIT('h0d)
	) name57 (
		b_pad,
		\u0_pad ,
		\u2_pad ,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\k2_pad ,
		\l2_pad ,
		_w154_
	);
	LUT4 #(
		.INIT('h4050)
	) name59 (
		\c1_pad ,
		\k2_pad ,
		\l2_pad ,
		\m2_pad ,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		\c1_pad ,
		\k2_pad ,
		_w156_
	);
	LUT4 #(
		.INIT('hb1b0)
	) name61 (
		_w153_,
		_w154_,
		_w155_,
		_w156_,
		_w157_
	);
	LUT3 #(
		.INIT('h13)
	) name62 (
		\g0_pad ,
		\i0_pad ,
		\v2_pad ,
		_w158_
	);
	LUT3 #(
		.INIT('h0b)
	) name63 (
		_w109_,
		_w132_,
		_w158_,
		_w159_
	);
	LUT3 #(
		.INIT('h4c)
	) name64 (
		\g0_pad ,
		\m0_pad ,
		\v2_pad ,
		_w160_
	);
	LUT4 #(
		.INIT('hff0b)
	) name65 (
		_w109_,
		_w132_,
		_w158_,
		_w160_,
		_w161_
	);
	LUT3 #(
		.INIT('h40)
	) name66 (
		\k2_pad ,
		\l2_pad ,
		\m2_pad ,
		_w162_
	);
	LUT4 #(
		.INIT('he0a0)
	) name67 (
		\m1_pad ,
		_w108_,
		_w158_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\l2_pad ,
		\m2_pad ,
		_w164_
	);
	LUT4 #(
		.INIT('h0031)
	) name69 (
		b_pad,
		\m2_pad ,
		\u0_pad ,
		\u2_pad ,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w164_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\l2_pad ,
		\m2_pad ,
		_w167_
	);
	LUT3 #(
		.INIT('h45)
	) name72 (
		\c1_pad ,
		\k2_pad ,
		\l2_pad ,
		_w168_
	);
	LUT3 #(
		.INIT('hb0)
	) name73 (
		_w153_,
		_w167_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w166_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\c1_pad ,
		\i0_pad ,
		_w171_
	);
	LUT4 #(
		.INIT('hea00)
	) name76 (
		\n0_pad ,
		_w102_,
		_w123_,
		_w171_,
		_w172_
	);
	LUT4 #(
		.INIT('h8000)
	) name77 (
		\g0_pad ,
		i_pad,
		\m1_pad ,
		\v2_pad ,
		_w173_
	);
	LUT3 #(
		.INIT('h04)
	) name78 (
		g_pad,
		\h0_pad ,
		h_pad,
		_w174_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name79 (
		\e1_pad ,
		\m0_pad ,
		\n1_pad ,
		\o1_pad ,
		_w175_
	);
	LUT4 #(
		.INIT('h0233)
	) name80 (
		_w111_,
		_w173_,
		_w174_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\i0_pad ,
		_w176_,
		_w177_
	);
	LUT3 #(
		.INIT('h01)
	) name82 (
		\d1_pad ,
		\e1_pad ,
		\n2_pad ,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w162_,
		_w178_,
		_w179_
	);
	LUT3 #(
		.INIT('he0)
	) name84 (
		\d1_pad ,
		\e1_pad ,
		\n2_pad ,
		_w180_
	);
	LUT4 #(
		.INIT('h4000)
	) name85 (
		\k2_pad ,
		\l2_pad ,
		\m2_pad ,
		\n2_pad ,
		_w181_
	);
	LUT3 #(
		.INIT('h01)
	) name86 (
		\c1_pad ,
		_w180_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w179_,
		_w182_,
		_w183_
	);
	LUT3 #(
		.INIT('h10)
	) name88 (
		\c1_pad ,
		\i0_pad ,
		\o0_pad ,
		_w184_
	);
	LUT4 #(
		.INIT('h2f0d)
	) name89 (
		\e1_pad ,
		\m0_pad ,
		\o1_pad ,
		\p1_pad ,
		_w185_
	);
	LUT4 #(
		.INIT('hbaff)
	) name90 (
		\i0_pad ,
		_w109_,
		_w111_,
		_w185_,
		_w186_
	);
	LUT4 #(
		.INIT('h1114)
	) name91 (
		\c1_pad ,
		\o2_pad ,
		_w180_,
		_w181_,
		_w187_
	);
	LUT3 #(
		.INIT('h10)
	) name92 (
		\c1_pad ,
		\i0_pad ,
		\p0_pad ,
		_w188_
	);
	LUT3 #(
		.INIT('h20)
	) name93 (
		k_pad,
		_w109_,
		_w133_,
		_w189_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name94 (
		\e1_pad ,
		\m0_pad ,
		\p1_pad ,
		\q1_pad ,
		_w190_
	);
	LUT4 #(
		.INIT('h4500)
	) name95 (
		\i0_pad ,
		_w109_,
		_w111_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('he)
	) name96 (
		_w189_,
		_w191_,
		_w192_
	);
	LUT4 #(
		.INIT('h1113)
	) name97 (
		\o2_pad ,
		\p2_pad ,
		_w180_,
		_w181_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\o2_pad ,
		\p2_pad ,
		_w194_
	);
	LUT4 #(
		.INIT('h0155)
	) name99 (
		\c1_pad ,
		_w180_,
		_w181_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		_w193_,
		_w195_,
		_w196_
	);
	LUT3 #(
		.INIT('h10)
	) name101 (
		\c1_pad ,
		\i0_pad ,
		\q0_pad ,
		_w197_
	);
	LUT4 #(
		.INIT('h8000)
	) name102 (
		\g0_pad ,
		l_pad,
		\m1_pad ,
		\v2_pad ,
		_w198_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name103 (
		\e1_pad ,
		\m0_pad ,
		\q1_pad ,
		\r1_pad ,
		_w199_
	);
	LUT4 #(
		.INIT('h04af)
	) name104 (
		_w109_,
		_w111_,
		_w198_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\i0_pad ,
		_w200_,
		_w201_
	);
	LUT4 #(
		.INIT('h0155)
	) name106 (
		\q2_pad ,
		_w180_,
		_w181_,
		_w194_,
		_w202_
	);
	LUT3 #(
		.INIT('h80)
	) name107 (
		\o2_pad ,
		\p2_pad ,
		\q2_pad ,
		_w203_
	);
	LUT4 #(
		.INIT('h0155)
	) name108 (
		\c1_pad ,
		_w180_,
		_w181_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w202_,
		_w204_,
		_w205_
	);
	LUT3 #(
		.INIT('h10)
	) name110 (
		\c1_pad ,
		\i0_pad ,
		\r0_pad ,
		_w206_
	);
	LUT4 #(
		.INIT('h8000)
	) name111 (
		\g0_pad ,
		\m1_pad ,
		m_pad,
		\v2_pad ,
		_w207_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name112 (
		\e1_pad ,
		\m0_pad ,
		\r1_pad ,
		\s1_pad ,
		_w208_
	);
	LUT4 #(
		.INIT('h04af)
	) name113 (
		_w109_,
		_w111_,
		_w207_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\i0_pad ,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		\c1_pad ,
		\r2_pad ,
		_w211_
	);
	LUT4 #(
		.INIT('h1f00)
	) name116 (
		_w180_,
		_w181_,
		_w203_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\c1_pad ,
		\r2_pad ,
		_w213_
	);
	LUT4 #(
		.INIT('he000)
	) name118 (
		_w180_,
		_w181_,
		_w203_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('he)
	) name119 (
		_w212_,
		_w214_,
		_w215_
	);
	LUT3 #(
		.INIT('h10)
	) name120 (
		\c1_pad ,
		\i0_pad ,
		\s0_pad ,
		_w216_
	);
	LUT4 #(
		.INIT('h8000)
	) name121 (
		\g0_pad ,
		\m1_pad ,
		n_pad,
		\v2_pad ,
		_w217_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name122 (
		\e1_pad ,
		\m0_pad ,
		\s1_pad ,
		\t1_pad ,
		_w218_
	);
	LUT4 #(
		.INIT('h04af)
	) name123 (
		_w109_,
		_w111_,
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\i0_pad ,
		_w219_,
		_w220_
	);
	LUT4 #(
		.INIT('h0a02)
	) name125 (
		\b1_pad ,
		\e1_pad ,
		\i0_pad ,
		\m0_pad ,
		_w221_
	);
	LUT4 #(
		.INIT('h0200)
	) name126 (
		\e1_pad ,
		\i0_pad ,
		\m0_pad ,
		\n1_pad ,
		_w222_
	);
	LUT2 #(
		.INIT('he)
	) name127 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT3 #(
		.INIT('h10)
	) name128 (
		\c1_pad ,
		\i0_pad ,
		\t0_pad ,
		_w224_
	);
	LUT4 #(
		.INIT('h8000)
	) name129 (
		\g0_pad ,
		\m1_pad ,
		o_pad,
		\v2_pad ,
		_w225_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name130 (
		\e1_pad ,
		\m0_pad ,
		\t1_pad ,
		\u1_pad ,
		_w226_
	);
	LUT4 #(
		.INIT('h04af)
	) name131 (
		_w109_,
		_w111_,
		_w225_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		\i0_pad ,
		_w227_,
		_w228_
	);
	LUT4 #(
		.INIT('h1540)
	) name133 (
		\c1_pad ,
		\l1_pad ,
		\s2_pad ,
		\t2_pad ,
		_w229_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		b_pad,
		\i0_pad ,
		_w230_
	);
	LUT4 #(
		.INIT('h8000)
	) name135 (
		\g0_pad ,
		\m1_pad ,
		p_pad,
		\v2_pad ,
		_w231_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name136 (
		\e1_pad ,
		\m0_pad ,
		\u1_pad ,
		\v1_pad ,
		_w232_
	);
	LUT4 #(
		.INIT('h04af)
	) name137 (
		_w109_,
		_w111_,
		_w231_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\i0_pad ,
		_w233_,
		_w234_
	);
	LUT4 #(
		.INIT('h3302)
	) name139 (
		b_pad,
		\i0_pad ,
		\u0_pad ,
		\u2_pad ,
		_w235_
	);
	LUT3 #(
		.INIT('hb0)
	) name140 (
		_w146_,
		_w162_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		a_pad,
		\i0_pad ,
		_w237_
	);
	LUT4 #(
		.INIT('h8000)
	) name142 (
		\g0_pad ,
		\m1_pad ,
		q_pad,
		\v2_pad ,
		_w238_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name143 (
		\e1_pad ,
		\m0_pad ,
		\v1_pad ,
		\w1_pad ,
		_w239_
	);
	LUT4 #(
		.INIT('h04af)
	) name144 (
		_w109_,
		_w111_,
		_w238_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\i0_pad ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		\f0_pad ,
		\v2_pad ,
		_w242_
	);
	LUT4 #(
		.INIT('hf080)
	) name147 (
		_w123_,
		_w124_,
		_w158_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\i0_pad ,
		\v0_pad ,
		_w244_
	);
	LUT4 #(
		.INIT('h8000)
	) name149 (
		\g0_pad ,
		\m1_pad ,
		r_pad,
		\v2_pad ,
		_w245_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name150 (
		\e1_pad ,
		\m0_pad ,
		\w1_pad ,
		\x1_pad ,
		_w246_
	);
	LUT4 #(
		.INIT('h04af)
	) name151 (
		_w109_,
		_w111_,
		_w245_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\i0_pad ,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\i0_pad ,
		\w0_pad ,
		_w249_
	);
	LUT4 #(
		.INIT('h8000)
	) name154 (
		\g0_pad ,
		\m1_pad ,
		s_pad,
		\v2_pad ,
		_w250_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name155 (
		\e1_pad ,
		\m0_pad ,
		\x1_pad ,
		\y1_pad ,
		_w251_
	);
	LUT4 #(
		.INIT('h04af)
	) name156 (
		_w109_,
		_w111_,
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\i0_pad ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		\i0_pad ,
		\x0_pad ,
		_w254_
	);
	LUT4 #(
		.INIT('h8000)
	) name159 (
		\g0_pad ,
		\m1_pad ,
		t_pad,
		\v2_pad ,
		_w255_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name160 (
		\e1_pad ,
		\m0_pad ,
		\y1_pad ,
		\z1_pad ,
		_w256_
	);
	LUT4 #(
		.INIT('h04af)
	) name161 (
		_w109_,
		_w111_,
		_w255_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\i0_pad ,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		\i0_pad ,
		\y0_pad ,
		_w259_
	);
	LUT4 #(
		.INIT('h8000)
	) name164 (
		\g0_pad ,
		\m1_pad ,
		u_pad,
		\v2_pad ,
		_w260_
	);
	LUT4 #(
		.INIT('hfb08)
	) name165 (
		\a2_pad ,
		\e1_pad ,
		\m0_pad ,
		\z1_pad ,
		_w261_
	);
	LUT4 #(
		.INIT('h04af)
	) name166 (
		_w109_,
		_w111_,
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\i0_pad ,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		\i0_pad ,
		\z0_pad ,
		_w264_
	);
	LUT4 #(
		.INIT('h8000)
	) name169 (
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		v_pad,
		_w265_
	);
	LUT4 #(
		.INIT('haaca)
	) name170 (
		\a2_pad ,
		\b2_pad ,
		\e1_pad ,
		\m0_pad ,
		_w266_
	);
	LUT4 #(
		.INIT('h04af)
	) name171 (
		_w109_,
		_w111_,
		_w265_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\i0_pad ,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\a1_pad ,
		\i0_pad ,
		_w269_
	);
	LUT4 #(
		.INIT('h8000)
	) name174 (
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		w_pad,
		_w270_
	);
	LUT4 #(
		.INIT('haaca)
	) name175 (
		\b2_pad ,
		\c2_pad ,
		\e1_pad ,
		\m0_pad ,
		_w271_
	);
	LUT4 #(
		.INIT('h04af)
	) name176 (
		_w109_,
		_w111_,
		_w270_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\i0_pad ,
		_w272_,
		_w273_
	);
	LUT3 #(
		.INIT('h07)
	) name178 (
		_w123_,
		_w124_,
		_w138_,
		_w274_
	);
	LUT2 #(
		.INIT('hb)
	) name179 (
		_w159_,
		_w274_,
		_w275_
	);
	LUT4 #(
		.INIT('h8000)
	) name180 (
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		x_pad,
		_w276_
	);
	LUT4 #(
		.INIT('haaca)
	) name181 (
		\c2_pad ,
		\d2_pad ,
		\e1_pad ,
		\m0_pad ,
		_w277_
	);
	LUT4 #(
		.INIT('h04af)
	) name182 (
		_w109_,
		_w111_,
		_w276_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\i0_pad ,
		_w278_,
		_w279_
	);
	LUT4 #(
		.INIT('h0400)
	) name184 (
		\g0_pad ,
		\i0_pad ,
		\m1_pad ,
		\v2_pad ,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		_w109_,
		_w280_,
		_w281_
	);
	LUT4 #(
		.INIT('h8000)
	) name186 (
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		y_pad,
		_w282_
	);
	LUT4 #(
		.INIT('haae2)
	) name187 (
		\d2_pad ,
		\e1_pad ,
		\e2_pad ,
		\m0_pad ,
		_w283_
	);
	LUT4 #(
		.INIT('h04af)
	) name188 (
		_w109_,
		_w111_,
		_w282_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\i0_pad ,
		_w284_,
		_w285_
	);
	LUT3 #(
		.INIT('h54)
	) name190 (
		\c1_pad ,
		\d1_pad ,
		\e1_pad ,
		_w286_
	);
	LUT4 #(
		.INIT('h1000)
	) name191 (
		\c1_pad ,
		\k2_pad ,
		\l2_pad ,
		\m2_pad ,
		_w287_
	);
	LUT2 #(
		.INIT('he)
	) name192 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT4 #(
		.INIT('h8000)
	) name193 (
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		z_pad,
		_w289_
	);
	LUT4 #(
		.INIT('hcce4)
	) name194 (
		\e1_pad ,
		\e2_pad ,
		\f2_pad ,
		\m0_pad ,
		_w290_
	);
	LUT4 #(
		.INIT('h04af)
	) name195 (
		_w109_,
		_w111_,
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		\i0_pad ,
		_w291_,
		_w292_
	);
	LUT3 #(
		.INIT('h15)
	) name197 (
		\f1_pad ,
		_w102_,
		_w103_,
		_w293_
	);
	LUT4 #(
		.INIT('h0001)
	) name198 (
		\o0_pad ,
		\p2_pad ,
		\q2_pad ,
		\r2_pad ,
		_w294_
	);
	LUT3 #(
		.INIT('h15)
	) name199 (
		\c1_pad ,
		_w103_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		_w293_,
		_w295_,
		_w296_
	);
	LUT4 #(
		.INIT('h8000)
	) name201 (
		\a0_pad ,
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		_w297_
	);
	LUT4 #(
		.INIT('hcce4)
	) name202 (
		\e1_pad ,
		\f2_pad ,
		\g2_pad ,
		\m0_pad ,
		_w298_
	);
	LUT4 #(
		.INIT('h04af)
	) name203 (
		_w109_,
		_w111_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		\i0_pad ,
		_w299_,
		_w300_
	);
	LUT3 #(
		.INIT('h15)
	) name205 (
		\g1_pad ,
		_w102_,
		_w103_,
		_w301_
	);
	LUT4 #(
		.INIT('h0001)
	) name206 (
		\p0_pad ,
		\p2_pad ,
		\q2_pad ,
		\r2_pad ,
		_w302_
	);
	LUT3 #(
		.INIT('h15)
	) name207 (
		\c1_pad ,
		_w103_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w301_,
		_w303_,
		_w304_
	);
	LUT4 #(
		.INIT('h8000)
	) name209 (
		\b0_pad ,
		\g0_pad ,
		\m1_pad ,
		\v2_pad ,
		_w305_
	);
	LUT4 #(
		.INIT('hcce4)
	) name210 (
		\e1_pad ,
		\g2_pad ,
		\h2_pad ,
		\m0_pad ,
		_w306_
	);
	LUT4 #(
		.INIT('h04af)
	) name211 (
		_w109_,
		_w111_,
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		\i0_pad ,
		_w307_,
		_w308_
	);
	assign \a3_pad  = _w39_ ;
	assign \a4_pad  = _w107_ ;
	assign \a5_pad  = _w114_ ;
	assign \b3_pad  = _w43_ ;
	assign \b4_pad  = _w118_ ;
	assign \b5_pad  = _w122_ ;
	assign \c3_pad  = _w127_ ;
	assign \c4_pad  = _w131_ ;
	assign \c5_pad  = _w137_ ;
	assign \d3_pad  = _w141_ ;
	assign \d4_pad  = _w145_ ;
	assign \d5_pad  = _w150_ ;
	assign \e3_pad  = _w151_ ;
	assign \e4_pad  = _w152_ ;
	assign \e5_pad  = _w157_ ;
	assign \f3_pad  = _w161_ ;
	assign \f4_pad  = _w163_ ;
	assign \f5_pad  = _w170_ ;
	assign \g3_pad  = _w172_ ;
	assign \g4_pad  = _w177_ ;
	assign \g5_pad  = _w183_ ;
	assign \h3_pad  = _w184_ ;
	assign \h4_pad  = _w186_ ;
	assign \h5_pad  = _w187_ ;
	assign \i3_pad  = _w188_ ;
	assign \i4_pad  = _w192_ ;
	assign \i5_pad  = _w196_ ;
	assign \j3_pad  = _w197_ ;
	assign \j4_pad  = _w201_ ;
	assign \j5_pad  = _w205_ ;
	assign \k3_pad  = _w206_ ;
	assign \k4_pad  = _w210_ ;
	assign \k5_pad  = _w215_ ;
	assign \l3_pad  = _w216_ ;
	assign \l4_pad  = _w220_ ;
	assign \l5_pad  = _w223_ ;
	assign \m3_pad  = _w224_ ;
	assign \m4_pad  = _w228_ ;
	assign \m5_pad  = _w229_ ;
	assign \n3_pad  = _w230_ ;
	assign \n4_pad  = _w234_ ;
	assign \n5_pad  = _w236_ ;
	assign \o3_pad  = _w237_ ;
	assign \o4_pad  = _w241_ ;
	assign \o5_pad  = _w243_ ;
	assign \p3_pad  = _w244_ ;
	assign \p4_pad  = _w248_ ;
	assign \q3_pad  = _w249_ ;
	assign \q4_pad  = _w253_ ;
	assign \r3_pad  = _w254_ ;
	assign \r4_pad  = _w258_ ;
	assign \s3_pad  = _w259_ ;
	assign \s4_pad  = _w263_ ;
	assign \t3_pad  = _w264_ ;
	assign \t4_pad  = _w268_ ;
	assign \u3_pad  = _w269_ ;
	assign \u4_pad  = _w273_ ;
	assign \v3_pad  = _w275_ ;
	assign \v4_pad  = _w279_ ;
	assign \w2_pad  = _w21_ ;
	assign \w3_pad  = _w281_ ;
	assign \w4_pad  = _w285_ ;
	assign \x2_pad  = _w25_ ;
	assign \x3_pad  = _w288_ ;
	assign \x4_pad  = _w292_ ;
	assign \y2_pad  = _w30_ ;
	assign \y3_pad  = _w296_ ;
	assign \y4_pad  = _w300_ ;
	assign \z2_pad  = _w35_ ;
	assign \z3_pad  = _w304_ ;
	assign \z4_pad  = _w308_ ;
endmodule;