module top( \din_i[0]_pad  , \din_i[1]_pad  , \din_i[2]_pad  , \din_i[3]_pad  , \din_i[4]_pad  , \din_i[5]_pad  , \din_i[6]_pad  , \din_i[7]_pad  , \pclk_r_reg/NET0131  , \pclk_s_reg/NET0131  , pcm_din_i_pad , pcm_dout_o_pad , pcm_sync_i_pad , \pcm_sync_r1_reg/P0001  , \pcm_sync_r2_reg/P0001  , \pcm_sync_r3_reg/P0001  , \psa_reg[0]/P0001  , \psa_reg[1]/P0001  , \psa_reg[2]/P0001  , \psa_reg[3]/P0001  , \psa_reg[4]/P0001  , \psa_reg[5]/P0001  , \psa_reg[6]/P0001  , \psa_reg[7]/P0001  , \psync_reg/P0001  , re_i_pad , rst_pad , \rx_hold_reg_reg[0]/P0001  , \rx_hold_reg_reg[10]/P0001  , \rx_hold_reg_reg[11]/P0001  , \rx_hold_reg_reg[12]/P0001  , \rx_hold_reg_reg[13]/P0001  , \rx_hold_reg_reg[14]/P0001  , \rx_hold_reg_reg[15]/P0001  , \rx_hold_reg_reg[1]/P0001  , \rx_hold_reg_reg[2]/P0001  , \rx_hold_reg_reg[3]/P0001  , \rx_hold_reg_reg[4]/P0001  , \rx_hold_reg_reg[5]/P0001  , \rx_hold_reg_reg[6]/P0001  , \rx_hold_reg_reg[7]/P0001  , \rx_hold_reg_reg[8]/P0001  , \rx_hold_reg_reg[9]/P0001  , \rx_reg_reg[0]/P0001  , \rx_reg_reg[10]/P0001  , \rx_reg_reg[11]/P0001  , \rx_reg_reg[12]/P0001  , \rx_reg_reg[13]/P0001  , \rx_reg_reg[14]/P0001  , \rx_reg_reg[15]/P0001  , \rx_reg_reg[1]/P0001  , \rx_reg_reg[2]/P0001  , \rx_reg_reg[3]/P0001  , \rx_reg_reg[4]/P0001  , \rx_reg_reg[5]/P0001  , \rx_reg_reg[6]/P0001  , \rx_reg_reg[7]/P0001  , \rx_reg_reg[8]/P0001  , \rx_reg_reg[9]/P0001  , \rxd_reg/P0001  , \rxd_t_reg/P0001  , \ssel[0]_pad  , \ssel[1]_pad  , \ssel[2]_pad  , \tx_cnt_reg[0]/NET0131  , \tx_cnt_reg[1]/NET0131  , \tx_cnt_reg[2]/NET0131  , \tx_cnt_reg[3]/P0001  , \tx_go_r1_reg/NET0131  , \tx_go_reg/NET0131  , \tx_hold_byte_h_reg[0]/P0001  , \tx_hold_byte_h_reg[1]/P0001  , \tx_hold_byte_h_reg[2]/P0001  , \tx_hold_byte_h_reg[3]/P0001  , \tx_hold_byte_h_reg[4]/P0001  , \tx_hold_byte_h_reg[5]/P0001  , \tx_hold_byte_h_reg[6]/P0001  , \tx_hold_byte_h_reg[7]/P0001  , \tx_hold_byte_l_reg[0]/P0001  , \tx_hold_byte_l_reg[1]/P0001  , \tx_hold_byte_l_reg[2]/P0001  , \tx_hold_byte_l_reg[3]/P0001  , \tx_hold_byte_l_reg[4]/P0001  , \tx_hold_byte_l_reg[5]/P0001  , \tx_hold_byte_l_reg[6]/P0001  , \tx_hold_byte_l_reg[7]/P0001  , \tx_hold_reg_reg[0]/P0001  , \tx_hold_reg_reg[10]/P0001  , \tx_hold_reg_reg[11]/P0001  , \tx_hold_reg_reg[12]/P0001  , \tx_hold_reg_reg[13]/P0001  , \tx_hold_reg_reg[14]/P0001  , \tx_hold_reg_reg[1]/P0001  , \tx_hold_reg_reg[2]/P0001  , \tx_hold_reg_reg[3]/P0001  , \tx_hold_reg_reg[4]/P0001  , \tx_hold_reg_reg[5]/P0001  , \tx_hold_reg_reg[6]/P0001  , \tx_hold_reg_reg[7]/P0001  , \tx_hold_reg_reg[8]/P0001  , \tx_hold_reg_reg[9]/P0001  , \we_i[0]_pad  , \we_i[1]_pad  , \_al_n0  , \_al_n1  , \dout_o[0]_pad  , \dout_o[1]_pad  , \dout_o[2]_pad  , \dout_o[3]_pad  , \dout_o[4]_pad  , \dout_o[5]_pad  , \dout_o[6]_pad  , \dout_o[7]_pad  , \g1173/_0_  , \g1174/_0_  , \g1175/_0_  , \g1176/_0_  , \g1177/_0_  , \g1178/_0_  , \g1179/_0_  , \g1180/_0_  , \g1181/_0_  , \g1182/_0_  , \g1183/_0_  , \g1184/_0_  , \g1185/_0_  , \g1186/_0_  , \g1187/_0_  , \g1188/_0_  , \g1189/_0_  , \g1265/_0_  , \g1266/_0_  , \g1267/_0_  , \g1268/_0_  , \g1269/_0_  , \g1270/_0_  , \g1271/_0_  , \g1272/_0_  , \g1273/_0_  , \g1274/_0_  , \g1275/_0_  , \g1276/_0_  , \g1277/_0_  , \g1278/_0_  , \g1279/_0_  , \g1280/_0_  , \g1281/_0_  , \g1282/_0_  , \g1284/_0_  , \g1285/_0_  , \g1286/_0_  , \g1287/_0_  , \g1288/_0_  , \g1289/_0_  , \g1290/_0_  , \g1291/_0_  , \g1292/_0_  , \g1293/_0_  , \g1294/_0_  , \g1295/_0_  , \g1296/_0_  , \g1297/_0_  , \g1298/_0_  , \g1299/_0_  , \g1300/_0_  , \g1301/_0_  , \g1441/_0_  , \g1442/_3_  , \g1479_dup/_1_  , \g1504/_0_  , \g1505/_0_  , \g1506/_0_  , \g1508/_0_  , \g1511/_0_  , \g1516/_0_  , \g1518/_0_  , \g1521/_0_  , \g1522/_0_  , \g1523/_0_  , \g1524/_0_  , \g1526/_0_  , \g1527/_0_  , \g1528/_0_  , \g1529/_0_  , \g24/_0_  , \pcm_sync_r1_reg/P0001_reg_syn_3  , \rxd_t_reg/P0001_reg_syn_3  , \tx_hold_byte_l_reg[0]/P0001_reg_syn_3  );
  input \din_i[0]_pad  ;
  input \din_i[1]_pad  ;
  input \din_i[2]_pad  ;
  input \din_i[3]_pad  ;
  input \din_i[4]_pad  ;
  input \din_i[5]_pad  ;
  input \din_i[6]_pad  ;
  input \din_i[7]_pad  ;
  input \pclk_r_reg/NET0131  ;
  input \pclk_s_reg/NET0131  ;
  input pcm_din_i_pad ;
  input pcm_dout_o_pad ;
  input pcm_sync_i_pad ;
  input \pcm_sync_r1_reg/P0001  ;
  input \pcm_sync_r2_reg/P0001  ;
  input \pcm_sync_r3_reg/P0001  ;
  input \psa_reg[0]/P0001  ;
  input \psa_reg[1]/P0001  ;
  input \psa_reg[2]/P0001  ;
  input \psa_reg[3]/P0001  ;
  input \psa_reg[4]/P0001  ;
  input \psa_reg[5]/P0001  ;
  input \psa_reg[6]/P0001  ;
  input \psa_reg[7]/P0001  ;
  input \psync_reg/P0001  ;
  input re_i_pad ;
  input rst_pad ;
  input \rx_hold_reg_reg[0]/P0001  ;
  input \rx_hold_reg_reg[10]/P0001  ;
  input \rx_hold_reg_reg[11]/P0001  ;
  input \rx_hold_reg_reg[12]/P0001  ;
  input \rx_hold_reg_reg[13]/P0001  ;
  input \rx_hold_reg_reg[14]/P0001  ;
  input \rx_hold_reg_reg[15]/P0001  ;
  input \rx_hold_reg_reg[1]/P0001  ;
  input \rx_hold_reg_reg[2]/P0001  ;
  input \rx_hold_reg_reg[3]/P0001  ;
  input \rx_hold_reg_reg[4]/P0001  ;
  input \rx_hold_reg_reg[5]/P0001  ;
  input \rx_hold_reg_reg[6]/P0001  ;
  input \rx_hold_reg_reg[7]/P0001  ;
  input \rx_hold_reg_reg[8]/P0001  ;
  input \rx_hold_reg_reg[9]/P0001  ;
  input \rx_reg_reg[0]/P0001  ;
  input \rx_reg_reg[10]/P0001  ;
  input \rx_reg_reg[11]/P0001  ;
  input \rx_reg_reg[12]/P0001  ;
  input \rx_reg_reg[13]/P0001  ;
  input \rx_reg_reg[14]/P0001  ;
  input \rx_reg_reg[15]/P0001  ;
  input \rx_reg_reg[1]/P0001  ;
  input \rx_reg_reg[2]/P0001  ;
  input \rx_reg_reg[3]/P0001  ;
  input \rx_reg_reg[4]/P0001  ;
  input \rx_reg_reg[5]/P0001  ;
  input \rx_reg_reg[6]/P0001  ;
  input \rx_reg_reg[7]/P0001  ;
  input \rx_reg_reg[8]/P0001  ;
  input \rx_reg_reg[9]/P0001  ;
  input \rxd_reg/P0001  ;
  input \rxd_t_reg/P0001  ;
  input \ssel[0]_pad  ;
  input \ssel[1]_pad  ;
  input \ssel[2]_pad  ;
  input \tx_cnt_reg[0]/NET0131  ;
  input \tx_cnt_reg[1]/NET0131  ;
  input \tx_cnt_reg[2]/NET0131  ;
  input \tx_cnt_reg[3]/P0001  ;
  input \tx_go_r1_reg/NET0131  ;
  input \tx_go_reg/NET0131  ;
  input \tx_hold_byte_h_reg[0]/P0001  ;
  input \tx_hold_byte_h_reg[1]/P0001  ;
  input \tx_hold_byte_h_reg[2]/P0001  ;
  input \tx_hold_byte_h_reg[3]/P0001  ;
  input \tx_hold_byte_h_reg[4]/P0001  ;
  input \tx_hold_byte_h_reg[5]/P0001  ;
  input \tx_hold_byte_h_reg[6]/P0001  ;
  input \tx_hold_byte_h_reg[7]/P0001  ;
  input \tx_hold_byte_l_reg[0]/P0001  ;
  input \tx_hold_byte_l_reg[1]/P0001  ;
  input \tx_hold_byte_l_reg[2]/P0001  ;
  input \tx_hold_byte_l_reg[3]/P0001  ;
  input \tx_hold_byte_l_reg[4]/P0001  ;
  input \tx_hold_byte_l_reg[5]/P0001  ;
  input \tx_hold_byte_l_reg[6]/P0001  ;
  input \tx_hold_byte_l_reg[7]/P0001  ;
  input \tx_hold_reg_reg[0]/P0001  ;
  input \tx_hold_reg_reg[10]/P0001  ;
  input \tx_hold_reg_reg[11]/P0001  ;
  input \tx_hold_reg_reg[12]/P0001  ;
  input \tx_hold_reg_reg[13]/P0001  ;
  input \tx_hold_reg_reg[14]/P0001  ;
  input \tx_hold_reg_reg[1]/P0001  ;
  input \tx_hold_reg_reg[2]/P0001  ;
  input \tx_hold_reg_reg[3]/P0001  ;
  input \tx_hold_reg_reg[4]/P0001  ;
  input \tx_hold_reg_reg[5]/P0001  ;
  input \tx_hold_reg_reg[6]/P0001  ;
  input \tx_hold_reg_reg[7]/P0001  ;
  input \tx_hold_reg_reg[8]/P0001  ;
  input \tx_hold_reg_reg[9]/P0001  ;
  input \we_i[0]_pad  ;
  input \we_i[1]_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \dout_o[0]_pad  ;
  output \dout_o[1]_pad  ;
  output \dout_o[2]_pad  ;
  output \dout_o[3]_pad  ;
  output \dout_o[4]_pad  ;
  output \dout_o[5]_pad  ;
  output \dout_o[6]_pad  ;
  output \dout_o[7]_pad  ;
  output \g1173/_0_  ;
  output \g1174/_0_  ;
  output \g1175/_0_  ;
  output \g1176/_0_  ;
  output \g1177/_0_  ;
  output \g1178/_0_  ;
  output \g1179/_0_  ;
  output \g1180/_0_  ;
  output \g1181/_0_  ;
  output \g1182/_0_  ;
  output \g1183/_0_  ;
  output \g1184/_0_  ;
  output \g1185/_0_  ;
  output \g1186/_0_  ;
  output \g1187/_0_  ;
  output \g1188/_0_  ;
  output \g1189/_0_  ;
  output \g1265/_0_  ;
  output \g1266/_0_  ;
  output \g1267/_0_  ;
  output \g1268/_0_  ;
  output \g1269/_0_  ;
  output \g1270/_0_  ;
  output \g1271/_0_  ;
  output \g1272/_0_  ;
  output \g1273/_0_  ;
  output \g1274/_0_  ;
  output \g1275/_0_  ;
  output \g1276/_0_  ;
  output \g1277/_0_  ;
  output \g1278/_0_  ;
  output \g1279/_0_  ;
  output \g1280/_0_  ;
  output \g1281/_0_  ;
  output \g1282/_0_  ;
  output \g1284/_0_  ;
  output \g1285/_0_  ;
  output \g1286/_0_  ;
  output \g1287/_0_  ;
  output \g1288/_0_  ;
  output \g1289/_0_  ;
  output \g1290/_0_  ;
  output \g1291/_0_  ;
  output \g1292/_0_  ;
  output \g1293/_0_  ;
  output \g1294/_0_  ;
  output \g1295/_0_  ;
  output \g1296/_0_  ;
  output \g1297/_0_  ;
  output \g1298/_0_  ;
  output \g1299/_0_  ;
  output \g1300/_0_  ;
  output \g1301/_0_  ;
  output \g1441/_0_  ;
  output \g1442/_3_  ;
  output \g1479_dup/_1_  ;
  output \g1504/_0_  ;
  output \g1505/_0_  ;
  output \g1506/_0_  ;
  output \g1508/_0_  ;
  output \g1511/_0_  ;
  output \g1516/_0_  ;
  output \g1518/_0_  ;
  output \g1521/_0_  ;
  output \g1522/_0_  ;
  output \g1523/_0_  ;
  output \g1524/_0_  ;
  output \g1526/_0_  ;
  output \g1527/_0_  ;
  output \g1528/_0_  ;
  output \g1529/_0_  ;
  output \g24/_0_  ;
  output \pcm_sync_r1_reg/P0001_reg_syn_3  ;
  output \rxd_t_reg/P0001_reg_syn_3  ;
  output \tx_hold_byte_l_reg[0]/P0001_reg_syn_3  ;
  wire n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 ;
  assign n104 = re_i_pad & \rx_reg_reg[8]/P0001  ;
  assign n105 = ~re_i_pad & \rx_reg_reg[0]/P0001  ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = re_i_pad & \rx_reg_reg[9]/P0001  ;
  assign n108 = ~re_i_pad & \rx_reg_reg[1]/P0001  ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = re_i_pad & \rx_reg_reg[10]/P0001  ;
  assign n111 = ~re_i_pad & \rx_reg_reg[2]/P0001  ;
  assign n112 = ~n110 & ~n111 ;
  assign n113 = re_i_pad & \rx_reg_reg[11]/P0001  ;
  assign n114 = ~re_i_pad & \rx_reg_reg[3]/P0001  ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = re_i_pad & \rx_reg_reg[12]/P0001  ;
  assign n117 = ~re_i_pad & \rx_reg_reg[4]/P0001  ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = re_i_pad & \rx_reg_reg[13]/P0001  ;
  assign n120 = ~re_i_pad & \rx_reg_reg[5]/P0001  ;
  assign n121 = ~n119 & ~n120 ;
  assign n122 = re_i_pad & \rx_reg_reg[14]/P0001  ;
  assign n123 = ~re_i_pad & \rx_reg_reg[6]/P0001  ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = re_i_pad & \rx_reg_reg[15]/P0001  ;
  assign n126 = ~re_i_pad & \rx_reg_reg[7]/P0001  ;
  assign n127 = ~n125 & ~n126 ;
  assign n129 = ~\pclk_r_reg/NET0131  & \pclk_s_reg/NET0131  ;
  assign n130 = \tx_go_reg/NET0131  & n129 ;
  assign n132 = \tx_hold_reg_reg[2]/P0001  & ~n130 ;
  assign n131 = \tx_hold_reg_reg[1]/P0001  & n130 ;
  assign n133 = ~\psync_reg/P0001  & ~n131 ;
  assign n134 = ~n132 & n133 ;
  assign n128 = \psync_reg/P0001  & ~\tx_hold_byte_l_reg[2]/P0001  ;
  assign n135 = rst_pad & ~n128 ;
  assign n136 = ~n134 & n135 ;
  assign n139 = \tx_hold_reg_reg[3]/P0001  & ~n130 ;
  assign n138 = \tx_hold_reg_reg[2]/P0001  & n130 ;
  assign n140 = ~\psync_reg/P0001  & ~n138 ;
  assign n141 = ~n139 & n140 ;
  assign n137 = \psync_reg/P0001  & ~\tx_hold_byte_l_reg[3]/P0001  ;
  assign n142 = rst_pad & ~n137 ;
  assign n143 = ~n141 & n142 ;
  assign n146 = \tx_hold_reg_reg[1]/P0001  & ~n130 ;
  assign n145 = \tx_hold_reg_reg[0]/P0001  & n130 ;
  assign n147 = ~\psync_reg/P0001  & ~n145 ;
  assign n148 = ~n146 & n147 ;
  assign n144 = \psync_reg/P0001  & ~\tx_hold_byte_l_reg[1]/P0001  ;
  assign n149 = rst_pad & ~n144 ;
  assign n150 = ~n148 & n149 ;
  assign n153 = \tx_hold_reg_reg[4]/P0001  & ~n130 ;
  assign n152 = \tx_hold_reg_reg[3]/P0001  & n130 ;
  assign n154 = ~\psync_reg/P0001  & ~n152 ;
  assign n155 = ~n153 & n154 ;
  assign n151 = \psync_reg/P0001  & ~\tx_hold_byte_l_reg[4]/P0001  ;
  assign n156 = rst_pad & ~n151 ;
  assign n157 = ~n155 & n156 ;
  assign n160 = \tx_hold_reg_reg[5]/P0001  & ~n130 ;
  assign n159 = \tx_hold_reg_reg[4]/P0001  & n130 ;
  assign n161 = ~\psync_reg/P0001  & ~n159 ;
  assign n162 = ~n160 & n161 ;
  assign n158 = \psync_reg/P0001  & ~\tx_hold_byte_l_reg[5]/P0001  ;
  assign n163 = rst_pad & ~n158 ;
  assign n164 = ~n162 & n163 ;
  assign n167 = \tx_hold_reg_reg[6]/P0001  & ~n130 ;
  assign n166 = \tx_hold_reg_reg[5]/P0001  & n130 ;
  assign n168 = ~\psync_reg/P0001  & ~n166 ;
  assign n169 = ~n167 & n168 ;
  assign n165 = \psync_reg/P0001  & ~\tx_hold_byte_l_reg[6]/P0001  ;
  assign n170 = rst_pad & ~n165 ;
  assign n171 = ~n169 & n170 ;
  assign n174 = \tx_hold_reg_reg[7]/P0001  & ~n130 ;
  assign n173 = \tx_hold_reg_reg[6]/P0001  & n130 ;
  assign n175 = ~\psync_reg/P0001  & ~n173 ;
  assign n176 = ~n174 & n175 ;
  assign n172 = \psync_reg/P0001  & ~\tx_hold_byte_l_reg[7]/P0001  ;
  assign n177 = rst_pad & ~n172 ;
  assign n178 = ~n176 & n177 ;
  assign n181 = \tx_hold_reg_reg[8]/P0001  & ~n130 ;
  assign n180 = \tx_hold_reg_reg[7]/P0001  & n130 ;
  assign n182 = ~\psync_reg/P0001  & ~n180 ;
  assign n183 = ~n181 & n182 ;
  assign n179 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[0]/P0001  ;
  assign n184 = rst_pad & ~n179 ;
  assign n185 = ~n183 & n184 ;
  assign n188 = \tx_hold_reg_reg[9]/P0001  & ~n130 ;
  assign n187 = \tx_hold_reg_reg[8]/P0001  & n130 ;
  assign n189 = ~\psync_reg/P0001  & ~n187 ;
  assign n190 = ~n188 & n189 ;
  assign n186 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[1]/P0001  ;
  assign n191 = rst_pad & ~n186 ;
  assign n192 = ~n190 & n191 ;
  assign n195 = \tx_hold_reg_reg[10]/P0001  & ~n130 ;
  assign n194 = \tx_hold_reg_reg[9]/P0001  & n130 ;
  assign n196 = ~\psync_reg/P0001  & ~n194 ;
  assign n197 = ~n195 & n196 ;
  assign n193 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[2]/P0001  ;
  assign n198 = rst_pad & ~n193 ;
  assign n199 = ~n197 & n198 ;
  assign n202 = \tx_hold_reg_reg[11]/P0001  & ~n130 ;
  assign n201 = \tx_hold_reg_reg[10]/P0001  & n130 ;
  assign n203 = ~\psync_reg/P0001  & ~n201 ;
  assign n204 = ~n202 & n203 ;
  assign n200 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[3]/P0001  ;
  assign n205 = rst_pad & ~n200 ;
  assign n206 = ~n204 & n205 ;
  assign n209 = \tx_hold_reg_reg[12]/P0001  & ~n130 ;
  assign n208 = \tx_hold_reg_reg[11]/P0001  & n130 ;
  assign n210 = ~\psync_reg/P0001  & ~n208 ;
  assign n211 = ~n209 & n210 ;
  assign n207 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[4]/P0001  ;
  assign n212 = rst_pad & ~n207 ;
  assign n213 = ~n211 & n212 ;
  assign n216 = \tx_hold_reg_reg[13]/P0001  & ~n130 ;
  assign n215 = \tx_hold_reg_reg[12]/P0001  & n130 ;
  assign n217 = ~\psync_reg/P0001  & ~n215 ;
  assign n218 = ~n216 & n217 ;
  assign n214 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[5]/P0001  ;
  assign n219 = rst_pad & ~n214 ;
  assign n220 = ~n218 & n219 ;
  assign n223 = \tx_hold_reg_reg[14]/P0001  & ~n130 ;
  assign n222 = \tx_hold_reg_reg[13]/P0001  & n130 ;
  assign n224 = ~\psync_reg/P0001  & ~n222 ;
  assign n225 = ~n223 & n224 ;
  assign n221 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[6]/P0001  ;
  assign n226 = rst_pad & ~n221 ;
  assign n227 = ~n225 & n226 ;
  assign n230 = pcm_dout_o_pad & ~n130 ;
  assign n229 = \tx_hold_reg_reg[14]/P0001  & n130 ;
  assign n231 = ~\psync_reg/P0001  & ~n229 ;
  assign n232 = ~n230 & n231 ;
  assign n228 = \psync_reg/P0001  & ~\tx_hold_byte_h_reg[7]/P0001  ;
  assign n233 = rst_pad & ~n228 ;
  assign n234 = ~n232 & n233 ;
  assign n235 = \psync_reg/P0001  & \tx_hold_byte_l_reg[0]/P0001  ;
  assign n236 = ~\psync_reg/P0001  & \tx_hold_reg_reg[0]/P0001  ;
  assign n237 = ~n130 & n236 ;
  assign n238 = ~n235 & ~n237 ;
  assign n239 = rst_pad & ~n238 ;
  assign n240 = \tx_cnt_reg[0]/NET0131  & \tx_cnt_reg[1]/NET0131  ;
  assign n241 = \tx_cnt_reg[2]/NET0131  & n240 ;
  assign n242 = \tx_cnt_reg[3]/P0001  & n129 ;
  assign n243 = n241 & n242 ;
  assign n244 = \tx_go_reg/NET0131  & ~n243 ;
  assign n245 = ~\psync_reg/P0001  & ~n244 ;
  assign n246 = rst_pad & ~n245 ;
  assign n247 = \tx_cnt_reg[0]/NET0131  & n130 ;
  assign n248 = \tx_cnt_reg[1]/NET0131  & n247 ;
  assign n249 = ~\tx_cnt_reg[2]/NET0131  & ~n248 ;
  assign n250 = n130 & n241 ;
  assign n251 = rst_pad & ~n250 ;
  assign n252 = ~n249 & n251 ;
  assign n253 = \tx_go_r1_reg/NET0131  & ~\tx_go_reg/NET0131  ;
  assign n254 = n129 & n253 ;
  assign n256 = ~\rx_hold_reg_reg[14]/P0001  & n254 ;
  assign n255 = ~\rx_reg_reg[14]/P0001  & ~n254 ;
  assign n257 = rst_pad & ~n255 ;
  assign n258 = ~n256 & n257 ;
  assign n260 = ~\rx_hold_reg_reg[3]/P0001  & n254 ;
  assign n259 = ~\rx_reg_reg[3]/P0001  & ~n254 ;
  assign n261 = rst_pad & ~n259 ;
  assign n262 = ~n260 & n261 ;
  assign n264 = ~\rx_hold_reg_reg[13]/P0001  & n254 ;
  assign n263 = ~\rx_reg_reg[13]/P0001  & ~n254 ;
  assign n265 = rst_pad & ~n263 ;
  assign n266 = ~n264 & n265 ;
  assign n268 = ~\rx_hold_reg_reg[15]/P0001  & n254 ;
  assign n267 = ~\rx_reg_reg[15]/P0001  & ~n254 ;
  assign n269 = rst_pad & ~n267 ;
  assign n270 = ~n268 & n269 ;
  assign n272 = ~\rx_hold_reg_reg[1]/P0001  & n254 ;
  assign n271 = ~\rx_reg_reg[1]/P0001  & ~n254 ;
  assign n273 = rst_pad & ~n271 ;
  assign n274 = ~n272 & n273 ;
  assign n276 = ~\rx_hold_reg_reg[2]/P0001  & n254 ;
  assign n275 = ~\rx_reg_reg[2]/P0001  & ~n254 ;
  assign n277 = rst_pad & ~n275 ;
  assign n278 = ~n276 & n277 ;
  assign n280 = ~\rx_hold_reg_reg[5]/P0001  & n254 ;
  assign n279 = ~\rx_reg_reg[5]/P0001  & ~n254 ;
  assign n281 = rst_pad & ~n279 ;
  assign n282 = ~n280 & n281 ;
  assign n284 = ~\rx_hold_reg_reg[6]/P0001  & n254 ;
  assign n283 = ~\rx_reg_reg[6]/P0001  & ~n254 ;
  assign n285 = rst_pad & ~n283 ;
  assign n286 = ~n284 & n285 ;
  assign n288 = ~\rx_hold_reg_reg[7]/P0001  & n254 ;
  assign n287 = ~\rx_reg_reg[7]/P0001  & ~n254 ;
  assign n289 = rst_pad & ~n287 ;
  assign n290 = ~n288 & n289 ;
  assign n292 = ~\rx_hold_reg_reg[8]/P0001  & n254 ;
  assign n291 = ~\rx_reg_reg[8]/P0001  & ~n254 ;
  assign n293 = rst_pad & ~n291 ;
  assign n294 = ~n292 & n293 ;
  assign n296 = ~\rx_hold_reg_reg[9]/P0001  & n254 ;
  assign n295 = ~\rx_reg_reg[9]/P0001  & ~n254 ;
  assign n297 = rst_pad & ~n295 ;
  assign n298 = ~n296 & n297 ;
  assign n300 = ~\rx_hold_reg_reg[0]/P0001  & n254 ;
  assign n299 = ~\rx_reg_reg[0]/P0001  & ~n254 ;
  assign n301 = rst_pad & ~n299 ;
  assign n302 = ~n300 & n301 ;
  assign n304 = ~\rx_hold_reg_reg[4]/P0001  & n254 ;
  assign n303 = ~\rx_reg_reg[4]/P0001  & ~n254 ;
  assign n305 = rst_pad & ~n303 ;
  assign n306 = ~n304 & n305 ;
  assign n308 = ~\rx_hold_reg_reg[10]/P0001  & n254 ;
  assign n307 = ~\rx_reg_reg[10]/P0001  & ~n254 ;
  assign n309 = rst_pad & ~n307 ;
  assign n310 = ~n308 & n309 ;
  assign n312 = ~\rx_hold_reg_reg[11]/P0001  & n254 ;
  assign n311 = ~\rx_reg_reg[11]/P0001  & ~n254 ;
  assign n313 = rst_pad & ~n311 ;
  assign n314 = ~n312 & n313 ;
  assign n316 = ~\rx_hold_reg_reg[12]/P0001  & n254 ;
  assign n315 = ~\rx_reg_reg[12]/P0001  & ~n254 ;
  assign n317 = rst_pad & ~n315 ;
  assign n318 = ~n316 & n317 ;
  assign n319 = \pcm_sync_r2_reg/P0001  & ~\pcm_sync_r3_reg/P0001  ;
  assign n320 = ~\tx_cnt_reg[0]/NET0131  & ~n130 ;
  assign n321 = rst_pad & ~n247 ;
  assign n322 = ~n320 & n321 ;
  assign n323 = ~\tx_go_r1_reg/NET0131  & ~\tx_go_reg/NET0131  ;
  assign n324 = \pclk_r_reg/NET0131  & ~\pclk_s_reg/NET0131  ;
  assign n325 = ~n323 & n324 ;
  assign n327 = ~\rxd_reg/P0001  & n325 ;
  assign n326 = ~\rx_hold_reg_reg[0]/P0001  & ~n325 ;
  assign n328 = rst_pad & ~n326 ;
  assign n329 = ~n327 & n328 ;
  assign n331 = ~\rx_hold_reg_reg[9]/P0001  & n325 ;
  assign n330 = ~\rx_hold_reg_reg[10]/P0001  & ~n325 ;
  assign n332 = rst_pad & ~n330 ;
  assign n333 = ~n331 & n332 ;
  assign n335 = ~\rx_hold_reg_reg[10]/P0001  & n325 ;
  assign n334 = ~\rx_hold_reg_reg[11]/P0001  & ~n325 ;
  assign n336 = rst_pad & ~n334 ;
  assign n337 = ~n335 & n336 ;
  assign n339 = ~\rx_hold_reg_reg[11]/P0001  & n325 ;
  assign n338 = ~\rx_hold_reg_reg[12]/P0001  & ~n325 ;
  assign n340 = rst_pad & ~n338 ;
  assign n341 = ~n339 & n340 ;
  assign n343 = ~\rx_hold_reg_reg[12]/P0001  & n325 ;
  assign n342 = ~\rx_hold_reg_reg[13]/P0001  & ~n325 ;
  assign n344 = rst_pad & ~n342 ;
  assign n345 = ~n343 & n344 ;
  assign n346 = ~\tx_cnt_reg[1]/NET0131  & ~n247 ;
  assign n347 = rst_pad & ~n248 ;
  assign n348 = ~n346 & n347 ;
  assign n350 = ~\rx_hold_reg_reg[13]/P0001  & n325 ;
  assign n349 = ~\rx_hold_reg_reg[14]/P0001  & ~n325 ;
  assign n351 = rst_pad & ~n349 ;
  assign n352 = ~n350 & n351 ;
  assign n354 = ~\rx_hold_reg_reg[14]/P0001  & n325 ;
  assign n353 = ~\rx_hold_reg_reg[15]/P0001  & ~n325 ;
  assign n355 = rst_pad & ~n353 ;
  assign n356 = ~n354 & n355 ;
  assign n358 = ~\rx_hold_reg_reg[0]/P0001  & n325 ;
  assign n357 = ~\rx_hold_reg_reg[1]/P0001  & ~n325 ;
  assign n359 = rst_pad & ~n357 ;
  assign n360 = ~n358 & n359 ;
  assign n362 = ~\rx_hold_reg_reg[1]/P0001  & n325 ;
  assign n361 = ~\rx_hold_reg_reg[2]/P0001  & ~n325 ;
  assign n363 = rst_pad & ~n361 ;
  assign n364 = ~n362 & n363 ;
  assign n366 = ~\rx_hold_reg_reg[2]/P0001  & n325 ;
  assign n365 = ~\rx_hold_reg_reg[3]/P0001  & ~n325 ;
  assign n367 = rst_pad & ~n365 ;
  assign n368 = ~n366 & n367 ;
  assign n370 = ~\rx_hold_reg_reg[3]/P0001  & n325 ;
  assign n369 = ~\rx_hold_reg_reg[4]/P0001  & ~n325 ;
  assign n371 = rst_pad & ~n369 ;
  assign n372 = ~n370 & n371 ;
  assign n374 = ~\rx_hold_reg_reg[4]/P0001  & n325 ;
  assign n373 = ~\rx_hold_reg_reg[5]/P0001  & ~n325 ;
  assign n375 = rst_pad & ~n373 ;
  assign n376 = ~n374 & n375 ;
  assign n378 = ~\rx_hold_reg_reg[5]/P0001  & n325 ;
  assign n377 = ~\rx_hold_reg_reg[6]/P0001  & ~n325 ;
  assign n379 = rst_pad & ~n377 ;
  assign n380 = ~n378 & n379 ;
  assign n382 = ~\rx_hold_reg_reg[6]/P0001  & n325 ;
  assign n381 = ~\rx_hold_reg_reg[7]/P0001  & ~n325 ;
  assign n383 = rst_pad & ~n381 ;
  assign n384 = ~n382 & n383 ;
  assign n386 = ~\rx_hold_reg_reg[8]/P0001  & n325 ;
  assign n385 = ~\rx_hold_reg_reg[9]/P0001  & ~n325 ;
  assign n387 = rst_pad & ~n385 ;
  assign n388 = ~n386 & n387 ;
  assign n390 = ~\rx_hold_reg_reg[7]/P0001  & n325 ;
  assign n389 = ~\rx_hold_reg_reg[8]/P0001  & ~n325 ;
  assign n391 = rst_pad & ~n389 ;
  assign n392 = ~n390 & n391 ;
  assign n393 = \tx_go_r1_reg/NET0131  & ~n129 ;
  assign n394 = ~n130 & ~n393 ;
  assign n396 = ~\psa_reg[4]/P0001  & ~\ssel[0]_pad  ;
  assign n395 = ~\psa_reg[5]/P0001  & \ssel[0]_pad  ;
  assign n397 = ~\ssel[1]_pad  & ~n395 ;
  assign n398 = ~n396 & n397 ;
  assign n400 = ~\psa_reg[6]/P0001  & ~\ssel[0]_pad  ;
  assign n399 = ~\psa_reg[7]/P0001  & \ssel[0]_pad  ;
  assign n401 = \ssel[1]_pad  & ~n399 ;
  assign n402 = ~n400 & n401 ;
  assign n403 = ~n398 & ~n402 ;
  assign n404 = \ssel[2]_pad  & ~n403 ;
  assign n406 = ~\psa_reg[0]/P0001  & ~\ssel[0]_pad  ;
  assign n405 = ~\psa_reg[1]/P0001  & \ssel[0]_pad  ;
  assign n407 = ~\ssel[1]_pad  & ~n405 ;
  assign n408 = ~n406 & n407 ;
  assign n410 = ~\psa_reg[2]/P0001  & ~\ssel[0]_pad  ;
  assign n409 = ~\psa_reg[3]/P0001  & \ssel[0]_pad  ;
  assign n411 = \ssel[1]_pad  & ~n409 ;
  assign n412 = ~n410 & n411 ;
  assign n413 = ~n408 & ~n412 ;
  assign n414 = ~\ssel[2]_pad  & ~n413 ;
  assign n415 = ~n404 & ~n414 ;
  assign n416 = \tx_hold_byte_l_reg[7]/P0001  & ~\we_i[0]_pad  ;
  assign n417 = \din_i[7]_pad  & \we_i[0]_pad  ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = \tx_hold_byte_l_reg[3]/P0001  & ~\we_i[0]_pad  ;
  assign n420 = \din_i[3]_pad  & \we_i[0]_pad  ;
  assign n421 = ~n419 & ~n420 ;
  assign n422 = \tx_hold_byte_h_reg[2]/P0001  & ~\we_i[1]_pad  ;
  assign n423 = \din_i[2]_pad  & \we_i[1]_pad  ;
  assign n424 = ~n422 & ~n423 ;
  assign n425 = \tx_hold_byte_h_reg[5]/P0001  & ~\we_i[1]_pad  ;
  assign n426 = \din_i[5]_pad  & \we_i[1]_pad  ;
  assign n427 = ~n425 & ~n426 ;
  assign n428 = \tx_hold_byte_h_reg[1]/P0001  & ~\we_i[1]_pad  ;
  assign n429 = \din_i[1]_pad  & \we_i[1]_pad  ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = \tx_hold_byte_l_reg[1]/P0001  & ~\we_i[0]_pad  ;
  assign n432 = \din_i[1]_pad  & \we_i[0]_pad  ;
  assign n433 = ~n431 & ~n432 ;
  assign n434 = \tx_hold_byte_h_reg[0]/P0001  & ~\we_i[1]_pad  ;
  assign n435 = \din_i[0]_pad  & \we_i[1]_pad  ;
  assign n436 = ~n434 & ~n435 ;
  assign n437 = \tx_hold_byte_h_reg[3]/P0001  & ~\we_i[1]_pad  ;
  assign n438 = \din_i[3]_pad  & \we_i[1]_pad  ;
  assign n439 = ~n437 & ~n438 ;
  assign n440 = \tx_hold_byte_h_reg[4]/P0001  & ~\we_i[1]_pad  ;
  assign n441 = \din_i[4]_pad  & \we_i[1]_pad  ;
  assign n442 = ~n440 & ~n441 ;
  assign n443 = \tx_hold_byte_h_reg[7]/P0001  & ~\we_i[1]_pad  ;
  assign n444 = \din_i[7]_pad  & \we_i[1]_pad  ;
  assign n445 = ~n443 & ~n444 ;
  assign n446 = \tx_hold_byte_h_reg[6]/P0001  & ~\we_i[1]_pad  ;
  assign n447 = \din_i[6]_pad  & \we_i[1]_pad  ;
  assign n448 = ~n446 & ~n447 ;
  assign n449 = \tx_hold_byte_l_reg[2]/P0001  & ~\we_i[0]_pad  ;
  assign n450 = \din_i[2]_pad  & \we_i[0]_pad  ;
  assign n451 = ~n449 & ~n450 ;
  assign n452 = \tx_hold_byte_l_reg[4]/P0001  & ~\we_i[0]_pad  ;
  assign n453 = \din_i[4]_pad  & \we_i[0]_pad  ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = \tx_hold_byte_l_reg[6]/P0001  & ~\we_i[0]_pad  ;
  assign n456 = \din_i[6]_pad  & \we_i[0]_pad  ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = \tx_hold_byte_l_reg[5]/P0001  & ~\we_i[0]_pad  ;
  assign n459 = \din_i[5]_pad  & \we_i[0]_pad  ;
  assign n460 = ~n458 & ~n459 ;
  assign n462 = \tx_cnt_reg[3]/P0001  & n250 ;
  assign n461 = ~\tx_cnt_reg[3]/P0001  & ~n250 ;
  assign n463 = rst_pad & ~n461 ;
  assign n464 = ~n462 & n463 ;
  assign n465 = \pcm_sync_r1_reg/P0001  & ~n324 ;
  assign n466 = pcm_sync_i_pad & n324 ;
  assign n467 = ~n465 & ~n466 ;
  assign n468 = \rxd_t_reg/P0001  & ~n324 ;
  assign n469 = pcm_din_i_pad & n324 ;
  assign n470 = ~n468 & ~n469 ;
  assign n471 = \din_i[0]_pad  & \we_i[0]_pad  ;
  assign n472 = \tx_hold_byte_l_reg[0]/P0001  & ~\we_i[0]_pad  ;
  assign n473 = ~n471 & ~n472 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \dout_o[0]_pad  = ~n106 ;
  assign \dout_o[1]_pad  = ~n109 ;
  assign \dout_o[2]_pad  = ~n112 ;
  assign \dout_o[3]_pad  = ~n115 ;
  assign \dout_o[4]_pad  = ~n118 ;
  assign \dout_o[5]_pad  = ~n121 ;
  assign \dout_o[6]_pad  = ~n124 ;
  assign \dout_o[7]_pad  = ~n127 ;
  assign \g1173/_0_  = n136 ;
  assign \g1174/_0_  = n143 ;
  assign \g1175/_0_  = n150 ;
  assign \g1176/_0_  = n157 ;
  assign \g1177/_0_  = n164 ;
  assign \g1178/_0_  = n171 ;
  assign \g1179/_0_  = n178 ;
  assign \g1180/_0_  = n185 ;
  assign \g1181/_0_  = n192 ;
  assign \g1182/_0_  = n199 ;
  assign \g1183/_0_  = n206 ;
  assign \g1184/_0_  = n213 ;
  assign \g1185/_0_  = n220 ;
  assign \g1186/_0_  = n227 ;
  assign \g1187/_0_  = n234 ;
  assign \g1188/_0_  = n239 ;
  assign \g1189/_0_  = n246 ;
  assign \g1265/_0_  = n252 ;
  assign \g1266/_0_  = n258 ;
  assign \g1267/_0_  = n262 ;
  assign \g1268/_0_  = n266 ;
  assign \g1269/_0_  = n270 ;
  assign \g1270/_0_  = n274 ;
  assign \g1271/_0_  = n278 ;
  assign \g1272/_0_  = n282 ;
  assign \g1273/_0_  = n286 ;
  assign \g1274/_0_  = n290 ;
  assign \g1275/_0_  = n294 ;
  assign \g1276/_0_  = n298 ;
  assign \g1277/_0_  = n302 ;
  assign \g1278/_0_  = n306 ;
  assign \g1279/_0_  = n310 ;
  assign \g1280/_0_  = n314 ;
  assign \g1281/_0_  = n318 ;
  assign \g1282/_0_  = n319 ;
  assign \g1284/_0_  = n322 ;
  assign \g1285/_0_  = n329 ;
  assign \g1286/_0_  = n333 ;
  assign \g1287/_0_  = n337 ;
  assign \g1288/_0_  = n341 ;
  assign \g1289/_0_  = n345 ;
  assign \g1290/_0_  = n348 ;
  assign \g1291/_0_  = n352 ;
  assign \g1292/_0_  = n356 ;
  assign \g1293/_0_  = n360 ;
  assign \g1294/_0_  = n364 ;
  assign \g1295/_0_  = n368 ;
  assign \g1296/_0_  = n372 ;
  assign \g1297/_0_  = n376 ;
  assign \g1298/_0_  = n380 ;
  assign \g1299/_0_  = n384 ;
  assign \g1300/_0_  = n388 ;
  assign \g1301/_0_  = n392 ;
  assign \g1441/_0_  = ~n394 ;
  assign \g1442/_3_  = ~n415 ;
  assign \g1479_dup/_1_  = n129 ;
  assign \g1504/_0_  = ~n418 ;
  assign \g1505/_0_  = ~n421 ;
  assign \g1506/_0_  = ~n424 ;
  assign \g1508/_0_  = ~n427 ;
  assign \g1511/_0_  = ~n430 ;
  assign \g1516/_0_  = ~n433 ;
  assign \g1518/_0_  = ~n436 ;
  assign \g1521/_0_  = ~n439 ;
  assign \g1522/_0_  = ~n442 ;
  assign \g1523/_0_  = ~n445 ;
  assign \g1524/_0_  = ~n448 ;
  assign \g1526/_0_  = ~n451 ;
  assign \g1527/_0_  = ~n454 ;
  assign \g1528/_0_  = ~n457 ;
  assign \g1529/_0_  = ~n460 ;
  assign \g24/_0_  = n464 ;
  assign \pcm_sync_r1_reg/P0001_reg_syn_3  = ~n467 ;
  assign \rxd_t_reg/P0001_reg_syn_3  = ~n470 ;
  assign \tx_hold_byte_l_reg[0]/P0001_reg_syn_3  = ~n473 ;
endmodule
