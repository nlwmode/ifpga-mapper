module top (\106GAT(15)_pad , \113GAT(16)_pad , \120GAT(17)_pad , \127GAT(18)_pad , \134GAT(19)_pad , \141GAT(20)_pad , \148GAT(21)_pad , \155GAT(22)_pad , \15GAT(2)_pad , \162GAT(23)_pad , \169GAT(24)_pad , \176GAT(25)_pad , \183GAT(26)_pad , \190GAT(27)_pad , \197GAT(28)_pad , \1GAT(0)_pad , \204GAT(29)_pad , \211GAT(30)_pad , \218GAT(31)_pad , \225GAT(32)_pad , \226GAT(33)_pad , \227GAT(34)_pad , \228GAT(35)_pad , \229GAT(36)_pad , \22GAT(3)_pad , \230GAT(37)_pad , \231GAT(38)_pad , \232GAT(39)_pad , \233GAT(40)_pad , \29GAT(4)_pad , \36GAT(5)_pad , \43GAT(6)_pad , \50GAT(7)_pad , \57GAT(8)_pad , \64GAT(9)_pad , \71GAT(10)_pad , \78GAT(11)_pad , \85GAT(12)_pad , \8GAT(1)_pad , \92GAT(13)_pad , \99GAT(14)_pad , \1324GAT(583)_pad , \1325GAT(579)_pad , \1326GAT(575)_pad , \1327GAT(571)_pad , \1328GAT(584)_pad , \1329GAT(580)_pad , \1330GAT(576)_pad , \1331GAT(572)_pad , \1332GAT(585)_pad , \1333GAT(581)_pad , \1334GAT(577)_pad , \1335GAT(573)_pad , \1336GAT(586)_pad , \1337GAT(582)_pad , \1338GAT(578)_pad , \1339GAT(574)_pad , \1340GAT(567)_pad , \1341GAT(563)_pad , \1342GAT(559)_pad , \1343GAT(555)_pad , \1344GAT(568)_pad , \1345GAT(564)_pad , \1346GAT(560)_pad , \1347GAT(556)_pad , \1348GAT(569)_pad , \1349GAT(565)_pad , \1350GAT(561)_pad , \1351GAT(557)_pad , \1352GAT(570)_pad , \1353GAT(566)_pad , \1354GAT(562)_pad , \1355GAT(558)_pad );
	input \106GAT(15)_pad  ;
	input \113GAT(16)_pad  ;
	input \120GAT(17)_pad  ;
	input \127GAT(18)_pad  ;
	input \134GAT(19)_pad  ;
	input \141GAT(20)_pad  ;
	input \148GAT(21)_pad  ;
	input \155GAT(22)_pad  ;
	input \15GAT(2)_pad  ;
	input \162GAT(23)_pad  ;
	input \169GAT(24)_pad  ;
	input \176GAT(25)_pad  ;
	input \183GAT(26)_pad  ;
	input \190GAT(27)_pad  ;
	input \197GAT(28)_pad  ;
	input \1GAT(0)_pad  ;
	input \204GAT(29)_pad  ;
	input \211GAT(30)_pad  ;
	input \218GAT(31)_pad  ;
	input \225GAT(32)_pad  ;
	input \226GAT(33)_pad  ;
	input \227GAT(34)_pad  ;
	input \228GAT(35)_pad  ;
	input \229GAT(36)_pad  ;
	input \22GAT(3)_pad  ;
	input \230GAT(37)_pad  ;
	input \231GAT(38)_pad  ;
	input \232GAT(39)_pad  ;
	input \233GAT(40)_pad  ;
	input \29GAT(4)_pad  ;
	input \36GAT(5)_pad  ;
	input \43GAT(6)_pad  ;
	input \50GAT(7)_pad  ;
	input \57GAT(8)_pad  ;
	input \64GAT(9)_pad  ;
	input \71GAT(10)_pad  ;
	input \78GAT(11)_pad  ;
	input \85GAT(12)_pad  ;
	input \8GAT(1)_pad  ;
	input \92GAT(13)_pad  ;
	input \99GAT(14)_pad  ;
	output \1324GAT(583)_pad  ;
	output \1325GAT(579)_pad  ;
	output \1326GAT(575)_pad  ;
	output \1327GAT(571)_pad  ;
	output \1328GAT(584)_pad  ;
	output \1329GAT(580)_pad  ;
	output \1330GAT(576)_pad  ;
	output \1331GAT(572)_pad  ;
	output \1332GAT(585)_pad  ;
	output \1333GAT(581)_pad  ;
	output \1334GAT(577)_pad  ;
	output \1335GAT(573)_pad  ;
	output \1336GAT(586)_pad  ;
	output \1337GAT(582)_pad  ;
	output \1338GAT(578)_pad  ;
	output \1339GAT(574)_pad  ;
	output \1340GAT(567)_pad  ;
	output \1341GAT(563)_pad  ;
	output \1342GAT(559)_pad  ;
	output \1343GAT(555)_pad  ;
	output \1344GAT(568)_pad  ;
	output \1345GAT(564)_pad  ;
	output \1346GAT(560)_pad  ;
	output \1347GAT(556)_pad  ;
	output \1348GAT(569)_pad  ;
	output \1349GAT(565)_pad  ;
	output \1350GAT(561)_pad  ;
	output \1351GAT(557)_pad  ;
	output \1352GAT(570)_pad  ;
	output \1353GAT(566)_pad  ;
	output \1354GAT(562)_pad  ;
	output \1355GAT(558)_pad  ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\225GAT(32)_pad ,
		\233GAT(40)_pad ,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\57GAT(8)_pad ,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\57GAT(8)_pad ,
		_w42_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w43_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\120GAT(17)_pad ,
		\127GAT(18)_pad ,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\120GAT(17)_pad ,
		\127GAT(18)_pad ,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\113GAT(16)_pad ,
		\134GAT(19)_pad ,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\113GAT(16)_pad ,
		\134GAT(19)_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w48_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w48_,
		_w51_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w45_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w45_,
		_w54_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\1GAT(0)_pad ,
		\29GAT(4)_pad ,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\1GAT(0)_pad ,
		\29GAT(4)_pad ,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w57_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w57_,
		_w60_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\148GAT(21)_pad ,
		\155GAT(22)_pad ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\148GAT(21)_pad ,
		\155GAT(22)_pad ,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w64_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\141GAT(20)_pad ,
		\162GAT(23)_pad ,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		\141GAT(20)_pad ,
		\162GAT(23)_pad ,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w66_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w66_,
		_w69_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\85GAT(12)_pad ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\85GAT(12)_pad ,
		_w72_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w63_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w63_,
		_w75_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\36GAT(5)_pad ,
		\43GAT(6)_pad ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\36GAT(5)_pad ,
		\43GAT(6)_pad ,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\29GAT(4)_pad ,
		\50GAT(7)_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\29GAT(4)_pad ,
		\50GAT(7)_pad ,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w81_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w81_,
		_w84_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w85_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\134GAT(19)_pad ,
		\162GAT(23)_pad ,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\134GAT(19)_pad ,
		\162GAT(23)_pad ,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w88_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		\190GAT(27)_pad ,
		\218GAT(31)_pad ,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\190GAT(27)_pad ,
		\218GAT(31)_pad ,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w91_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w90_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w90_,
		_w93_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\232GAT(39)_pad ,
		\233GAT(40)_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\106GAT(15)_pad ,
		\99GAT(14)_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\106GAT(15)_pad ,
		\99GAT(14)_pad ,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w98_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\85GAT(12)_pad ,
		\92GAT(13)_pad ,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		\85GAT(12)_pad ,
		\92GAT(13)_pad ,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w100_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w100_,
		_w103_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w104_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w97_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w97_,
		_w106_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w107_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		_w96_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w96_,
		_w109_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w87_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w87_,
		_w112_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w113_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\127GAT(18)_pad ,
		\155GAT(22)_pad ,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\127GAT(18)_pad ,
		\155GAT(22)_pad ,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\183GAT(26)_pad ,
		\211GAT(30)_pad ,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\183GAT(26)_pad ,
		\211GAT(30)_pad ,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		_w118_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w118_,
		_w121_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\1GAT(0)_pad ,
		\22GAT(3)_pad ,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\1GAT(0)_pad ,
		\22GAT(3)_pad ,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\15GAT(2)_pad ,
		\8GAT(1)_pad ,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		\15GAT(2)_pad ,
		\8GAT(1)_pad ,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w127_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w127_,
		_w130_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w131_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		\231GAT(38)_pad ,
		\233GAT(40)_pad ,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\64GAT(9)_pad ,
		\71GAT(10)_pad ,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\64GAT(9)_pad ,
		\71GAT(10)_pad ,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w135_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\57GAT(8)_pad ,
		\78GAT(11)_pad ,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		\57GAT(8)_pad ,
		\78GAT(11)_pad ,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w137_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w137_,
		_w140_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w141_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w134_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w134_,
		_w143_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w144_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		_w133_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		_w133_,
		_w146_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w147_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w124_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w124_,
		_w149_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w150_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		\197GAT(28)_pad ,
		\218GAT(31)_pad ,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		\197GAT(28)_pad ,
		\218GAT(31)_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\204GAT(29)_pad ,
		\211GAT(30)_pad ,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		\204GAT(29)_pad ,
		\211GAT(30)_pad ,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w155_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w155_,
		_w158_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		\106GAT(15)_pad ,
		\78GAT(11)_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		\106GAT(15)_pad ,
		\78GAT(11)_pad ,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		\22GAT(3)_pad ,
		\50GAT(7)_pad ,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		\22GAT(3)_pad ,
		\50GAT(7)_pad ,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w165_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w164_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w164_,
		_w167_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\228GAT(35)_pad ,
		\233GAT(40)_pad ,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w72_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w72_,
		_w171_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w172_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		_w170_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w170_,
		_w174_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w175_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w161_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w161_,
		_w177_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\226GAT(33)_pad ,
		\233GAT(40)_pad ,
		_w181_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\64GAT(9)_pad ,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		\64GAT(9)_pad ,
		_w181_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		\176GAT(25)_pad ,
		\183GAT(26)_pad ,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\176GAT(25)_pad ,
		\183GAT(26)_pad ,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\169GAT(24)_pad ,
		\190GAT(27)_pad ,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		\169GAT(24)_pad ,
		\190GAT(27)_pad ,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w187_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w187_,
		_w190_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w184_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w184_,
		_w193_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\36GAT(5)_pad ,
		\8GAT(1)_pad ,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\36GAT(5)_pad ,
		\8GAT(1)_pad ,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w197_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w196_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		_w196_,
		_w199_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		\92GAT(13)_pad ,
		_w161_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		\92GAT(13)_pad ,
		_w161_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w202_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w202_,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w78_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		_w54_,
		_w193_,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		_w54_,
		_w193_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\227GAT(34)_pad ,
		\233GAT(40)_pad ,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\15GAT(2)_pad ,
		\43GAT(6)_pad ,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\15GAT(2)_pad ,
		\43GAT(6)_pad ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w213_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w213_,
		_w216_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		\71GAT(10)_pad ,
		\99GAT(14)_pad ,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		\71GAT(10)_pad ,
		\99GAT(14)_pad ,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w220_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		_w219_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w219_,
		_w222_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w212_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w212_,
		_w225_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w209_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		_w78_,
		_w208_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w228_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w78_,
		_w208_,
		_w232_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w228_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w229_,
		_w231_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w233_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		_w180_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w180_,
		_w228_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w209_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w236_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w115_,
		_w152_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w239_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\230GAT(37)_pad ,
		\233GAT(40)_pad ,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w106_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		_w106_,
		_w242_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w243_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		\120GAT(17)_pad ,
		\148GAT(21)_pad ,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\120GAT(17)_pad ,
		\148GAT(21)_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w246_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w143_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w143_,
		_w248_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w249_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		\176GAT(25)_pad ,
		\204GAT(29)_pad ,
		_w252_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		\176GAT(25)_pad ,
		\204GAT(29)_pad ,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w252_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		_w251_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w251_,
		_w254_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w255_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w245_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w245_,
		_w257_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w258_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		\113GAT(16)_pad ,
		\141GAT(20)_pad ,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\113GAT(16)_pad ,
		\141GAT(20)_pad ,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w261_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w87_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name223 (
		_w87_,
		_w263_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\229GAT(36)_pad ,
		\233GAT(40)_pad ,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w133_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w133_,
		_w267_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w268_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\169GAT(24)_pad ,
		\197GAT(28)_pad ,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		\169GAT(24)_pad ,
		\197GAT(28)_pad ,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		_w270_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w270_,
		_w273_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w274_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w266_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w266_,
		_w276_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		_w260_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w241_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		_w78_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		\1GAT(0)_pad ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		\1GAT(0)_pad ,
		_w282_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w283_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w208_,
		_w281_,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\8GAT(1)_pad ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		\8GAT(1)_pad ,
		_w286_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w228_,
		_w281_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\15GAT(2)_pad ,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\15GAT(2)_pad ,
		_w290_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w291_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w180_,
		_w281_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		\22GAT(3)_pad ,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		\22GAT(3)_pad ,
		_w294_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w115_,
		_w239_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w152_,
		_w280_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w78_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		\29GAT(4)_pad ,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name261 (
		\29GAT(4)_pad ,
		_w301_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w208_,
		_w300_,
		_w305_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\36GAT(5)_pad ,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		\36GAT(5)_pad ,
		_w305_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w228_,
		_w300_,
		_w309_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		\43GAT(6)_pad ,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		\43GAT(6)_pad ,
		_w309_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w310_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name271 (
		_w180_,
		_w300_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		\50GAT(7)_pad ,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		\50GAT(7)_pad ,
		_w313_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w260_,
		_w279_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w241_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		_w78_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		\57GAT(8)_pad ,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		\57GAT(8)_pad ,
		_w319_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w208_,
		_w318_,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		\64GAT(9)_pad ,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		\64GAT(9)_pad ,
		_w323_,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w228_,
		_w318_,
		_w327_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		\71GAT(10)_pad ,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		\71GAT(10)_pad ,
		_w327_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w328_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w180_,
		_w318_,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\78GAT(11)_pad ,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		\78GAT(11)_pad ,
		_w331_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w332_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		_w152_,
		_w317_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		_w298_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		_w78_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\85GAT(12)_pad ,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		\85GAT(12)_pad ,
		_w337_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w338_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w208_,
		_w336_,
		_w341_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\92GAT(13)_pad ,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		\92GAT(13)_pad ,
		_w341_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w228_,
		_w336_,
		_w345_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		\99GAT(14)_pad ,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		\99GAT(14)_pad ,
		_w345_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w180_,
		_w336_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		\106GAT(15)_pad ,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		\106GAT(15)_pad ,
		_w349_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w350_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h2)
	) name311 (
		_w260_,
		_w279_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name312 (
		_w152_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w299_,
		_w335_,
		_w355_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w115_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w115_,
		_w152_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w353_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w357_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w180_,
		_w228_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w360_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w232_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w279_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		\113GAT(16)_pad ,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		\113GAT(16)_pad ,
		_w364_,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w365_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w260_,
		_w363_,
		_w368_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		\120GAT(17)_pad ,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		\120GAT(17)_pad ,
		_w368_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		_w152_,
		_w363_,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		\127GAT(18)_pad ,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h4)
	) name332 (
		\127GAT(18)_pad ,
		_w372_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w373_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w115_,
		_w363_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		\134GAT(19)_pad ,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		\134GAT(19)_pad ,
		_w376_,
		_w378_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w377_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w180_,
		_w360_,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w233_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w279_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\141GAT(20)_pad ,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\141GAT(20)_pad ,
		_w382_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w260_,
		_w381_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		\148GAT(21)_pad ,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		\148GAT(21)_pad ,
		_w386_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w387_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		_w152_,
		_w381_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		\155GAT(22)_pad ,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		\155GAT(22)_pad ,
		_w390_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		_w115_,
		_w381_,
		_w394_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\162GAT(23)_pad ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\162GAT(23)_pad ,
		_w394_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w395_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w230_,
		_w362_,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w279_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\169GAT(24)_pad ,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		\169GAT(24)_pad ,
		_w399_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w400_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w260_,
		_w398_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		\176GAT(25)_pad ,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\176GAT(25)_pad ,
		_w403_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w404_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w152_,
		_w398_,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		\183GAT(26)_pad ,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		\183GAT(26)_pad ,
		_w407_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w408_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		_w115_,
		_w398_,
		_w411_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\190GAT(27)_pad ,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		\190GAT(27)_pad ,
		_w411_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w412_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w231_,
		_w380_,
		_w415_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		_w279_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\197GAT(28)_pad ,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		\197GAT(28)_pad ,
		_w416_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w417_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w260_,
		_w415_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name379 (
		\204GAT(29)_pad ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		\204GAT(29)_pad ,
		_w420_,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w421_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name382 (
		_w152_,
		_w415_,
		_w424_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\211GAT(30)_pad ,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		\211GAT(30)_pad ,
		_w424_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w115_,
		_w415_,
		_w428_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		\218GAT(31)_pad ,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		\218GAT(31)_pad ,
		_w428_,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w429_,
		_w430_,
		_w431_
	);
	assign \1324GAT(583)_pad  = _w285_ ;
	assign \1325GAT(579)_pad  = _w289_ ;
	assign \1326GAT(575)_pad  = _w293_ ;
	assign \1327GAT(571)_pad  = _w297_ ;
	assign \1328GAT(584)_pad  = _w304_ ;
	assign \1329GAT(580)_pad  = _w308_ ;
	assign \1330GAT(576)_pad  = _w312_ ;
	assign \1331GAT(572)_pad  = _w316_ ;
	assign \1332GAT(585)_pad  = _w322_ ;
	assign \1333GAT(581)_pad  = _w326_ ;
	assign \1334GAT(577)_pad  = _w330_ ;
	assign \1335GAT(573)_pad  = _w334_ ;
	assign \1336GAT(586)_pad  = _w340_ ;
	assign \1337GAT(582)_pad  = _w344_ ;
	assign \1338GAT(578)_pad  = _w348_ ;
	assign \1339GAT(574)_pad  = _w352_ ;
	assign \1340GAT(567)_pad  = _w367_ ;
	assign \1341GAT(563)_pad  = _w371_ ;
	assign \1342GAT(559)_pad  = _w375_ ;
	assign \1343GAT(555)_pad  = _w379_ ;
	assign \1344GAT(568)_pad  = _w385_ ;
	assign \1345GAT(564)_pad  = _w389_ ;
	assign \1346GAT(560)_pad  = _w393_ ;
	assign \1347GAT(556)_pad  = _w397_ ;
	assign \1348GAT(569)_pad  = _w402_ ;
	assign \1349GAT(565)_pad  = _w406_ ;
	assign \1350GAT(561)_pad  = _w410_ ;
	assign \1351GAT(557)_pad  = _w414_ ;
	assign \1352GAT(570)_pad  = _w419_ ;
	assign \1353GAT(566)_pad  = _w423_ ;
	assign \1354GAT(562)_pad  = _w427_ ;
	assign \1355GAT(558)_pad  = _w431_ ;
endmodule;