module top( cont_eql_pad , eql_pad , \state_reg[0]/NET0131  , \state_reg[1]/NET0131  , \state_reg[2]/NET0131  , \_al_n0  , \_al_n1  , \g211/_0_  , \g212/_0_  , \g213/_0_  , \g218/_0_  , \g219/_0_  , \g220/_0_  , \g223/_0_  , \g227/_0_  );
  input cont_eql_pad ;
  input eql_pad ;
  input \state_reg[0]/NET0131  ;
  input \state_reg[1]/NET0131  ;
  input \state_reg[2]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g211/_0_  ;
  output \g212/_0_  ;
  output \g213/_0_  ;
  output \g218/_0_  ;
  output \g219/_0_  ;
  output \g220/_0_  ;
  output \g223/_0_  ;
  output \g227/_0_  ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 ;
  assign n6 = eql_pad & \state_reg[1]/NET0131  ;
  assign n7 = ~\state_reg[0]/NET0131  & ~\state_reg[2]/NET0131  ;
  assign n8 = n6 & n7 ;
  assign n9 = \state_reg[0]/NET0131  & \state_reg[1]/NET0131  ;
  assign n10 = \state_reg[2]/NET0131  & n9 ;
  assign n11 = ~n8 & ~n10 ;
  assign n12 = eql_pad & \state_reg[0]/NET0131  ;
  assign n13 = ~\state_reg[1]/NET0131  & n12 ;
  assign n14 = eql_pad & ~\state_reg[1]/NET0131  ;
  assign n15 = \state_reg[2]/NET0131  & n14 ;
  assign n16 = ~n13 & ~n15 ;
  assign n17 = n11 & n16 ;
  assign n18 = \state_reg[0]/NET0131  & ~\state_reg[2]/NET0131  ;
  assign n19 = ~eql_pad & ~\state_reg[1]/NET0131  ;
  assign n20 = n18 & n19 ;
  assign n21 = ~n10 & ~n20 ;
  assign n22 = ~\state_reg[0]/NET0131  & \state_reg[2]/NET0131  ;
  assign n23 = n19 & n22 ;
  assign n24 = \state_reg[2]/NET0131  & n6 ;
  assign n25 = ~n23 & ~n24 ;
  assign n26 = n21 & n25 ;
  assign n27 = ~\state_reg[0]/NET0131  & \state_reg[1]/NET0131  ;
  assign n28 = ~eql_pad & ~\state_reg[2]/NET0131  ;
  assign n29 = n27 & n28 ;
  assign n30 = ~cont_eql_pad & ~n10 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = ~\state_reg[0]/NET0131  & ~\state_reg[1]/NET0131  ;
  assign n33 = ~eql_pad & ~n32 ;
  assign n34 = \state_reg[2]/NET0131  & ~n9 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = \state_reg[0]/NET0131  & ~\state_reg[1]/NET0131  ;
  assign n37 = ~\state_reg[2]/NET0131  & n36 ;
  assign n38 = eql_pad & ~\state_reg[2]/NET0131  ;
  assign n39 = n27 & n38 ;
  assign n40 = ~n37 & ~n39 ;
  assign n41 = ~n35 & n40 ;
  assign n42 = \state_reg[2]/NET0131  & n32 ;
  assign n43 = ~n13 & ~n42 ;
  assign n44 = eql_pad & ~\state_reg[0]/NET0131  ;
  assign n45 = \state_reg[1]/NET0131  & n44 ;
  assign n46 = ~n10 & ~n45 ;
  assign n47 = n43 & n46 ;
  assign n48 = ~eql_pad & \state_reg[2]/NET0131  ;
  assign n49 = n32 & n48 ;
  assign n50 = eql_pad & \state_reg[2]/NET0131  ;
  assign n51 = n27 & n50 ;
  assign n52 = ~n49 & ~n51 ;
  assign n53 = ~eql_pad & \state_reg[0]/NET0131  ;
  assign n54 = ~\state_reg[2]/NET0131  & ~n32 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = n52 & ~n55 ;
  assign n57 = ~n15 & ~n20 ;
  assign n58 = \state_reg[2]/NET0131  & n44 ;
  assign n59 = ~n42 & ~n58 ;
  assign n60 = n57 & n59 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g211/_0_  = n17 ;
  assign \g212/_0_  = n26 ;
  assign \g213/_0_  = ~n31 ;
  assign \g218/_0_  = ~n41 ;
  assign \g219/_0_  = n47 ;
  assign \g220/_0_  = ~n56 ;
  assign \g223/_0_  = ~n60 ;
  assign \g227/_0_  = ~n52 ;
endmodule
