module top (\in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] , \result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] , \result[32] , \result[33] , \result[34] , \result[35] , \result[36] , \result[37] , \result[38] , \result[39] , \result[40] , \result[41] , \result[42] , \result[43] , \result[44] , \result[45] , \result[46] , \result[47] , \result[48] , \result[49] , \result[50] , \result[51] , \result[52] , \result[53] , \result[54] , \result[55] , \result[56] , \result[57] , \result[58] , \result[59] , \result[60] , \result[61] , \result[62] , \result[63] , \result[64] , \result[65] , \result[66] , \result[67] , \result[68] , \result[69] , \result[70] , \result[71] , \result[72] , \result[73] , \result[74] , \result[75] , \result[76] , \result[77] , \result[78] , \result[79] , \result[80] , \result[81] , \result[82] , \result[83] , \result[84] , \result[85] , \result[86] , \result[87] , \result[88] , \result[89] , \result[90] , \result[91] , \result[92] , \result[93] , \result[94] , \result[95] , \result[96] , \result[97] , \result[98] , \result[99] , \result[100] , \result[101] , \result[102] , \result[103] , \result[104] , \result[105] , \result[106] , \result[107] , \result[108] , \result[109] , \result[110] , \result[111] , \result[112] , \result[113] , \result[114] , \result[115] , \result[116] , \result[117] , \result[118] , \result[119] , \result[120] , \result[121] , \result[122] , \result[123] , \result[124] , \result[125] , \result[126] , \result[127] , \address[0] , \address[1] );
	input \in0[0]  ;
	input \in0[1]  ;
	input \in0[2]  ;
	input \in0[3]  ;
	input \in0[4]  ;
	input \in0[5]  ;
	input \in0[6]  ;
	input \in0[7]  ;
	input \in0[8]  ;
	input \in0[9]  ;
	input \in0[10]  ;
	input \in0[11]  ;
	input \in0[12]  ;
	input \in0[13]  ;
	input \in0[14]  ;
	input \in0[15]  ;
	input \in0[16]  ;
	input \in0[17]  ;
	input \in0[18]  ;
	input \in0[19]  ;
	input \in0[20]  ;
	input \in0[21]  ;
	input \in0[22]  ;
	input \in0[23]  ;
	input \in0[24]  ;
	input \in0[25]  ;
	input \in0[26]  ;
	input \in0[27]  ;
	input \in0[28]  ;
	input \in0[29]  ;
	input \in0[30]  ;
	input \in0[31]  ;
	input \in0[32]  ;
	input \in0[33]  ;
	input \in0[34]  ;
	input \in0[35]  ;
	input \in0[36]  ;
	input \in0[37]  ;
	input \in0[38]  ;
	input \in0[39]  ;
	input \in0[40]  ;
	input \in0[41]  ;
	input \in0[42]  ;
	input \in0[43]  ;
	input \in0[44]  ;
	input \in0[45]  ;
	input \in0[46]  ;
	input \in0[47]  ;
	input \in0[48]  ;
	input \in0[49]  ;
	input \in0[50]  ;
	input \in0[51]  ;
	input \in0[52]  ;
	input \in0[53]  ;
	input \in0[54]  ;
	input \in0[55]  ;
	input \in0[56]  ;
	input \in0[57]  ;
	input \in0[58]  ;
	input \in0[59]  ;
	input \in0[60]  ;
	input \in0[61]  ;
	input \in0[62]  ;
	input \in0[63]  ;
	input \in0[64]  ;
	input \in0[65]  ;
	input \in0[66]  ;
	input \in0[67]  ;
	input \in0[68]  ;
	input \in0[69]  ;
	input \in0[70]  ;
	input \in0[71]  ;
	input \in0[72]  ;
	input \in0[73]  ;
	input \in0[74]  ;
	input \in0[75]  ;
	input \in0[76]  ;
	input \in0[77]  ;
	input \in0[78]  ;
	input \in0[79]  ;
	input \in0[80]  ;
	input \in0[81]  ;
	input \in0[82]  ;
	input \in0[83]  ;
	input \in0[84]  ;
	input \in0[85]  ;
	input \in0[86]  ;
	input \in0[87]  ;
	input \in0[88]  ;
	input \in0[89]  ;
	input \in0[90]  ;
	input \in0[91]  ;
	input \in0[92]  ;
	input \in0[93]  ;
	input \in0[94]  ;
	input \in0[95]  ;
	input \in0[96]  ;
	input \in0[97]  ;
	input \in0[98]  ;
	input \in0[99]  ;
	input \in0[100]  ;
	input \in0[101]  ;
	input \in0[102]  ;
	input \in0[103]  ;
	input \in0[104]  ;
	input \in0[105]  ;
	input \in0[106]  ;
	input \in0[107]  ;
	input \in0[108]  ;
	input \in0[109]  ;
	input \in0[110]  ;
	input \in0[111]  ;
	input \in0[112]  ;
	input \in0[113]  ;
	input \in0[114]  ;
	input \in0[115]  ;
	input \in0[116]  ;
	input \in0[117]  ;
	input \in0[118]  ;
	input \in0[119]  ;
	input \in0[120]  ;
	input \in0[121]  ;
	input \in0[122]  ;
	input \in0[123]  ;
	input \in0[124]  ;
	input \in0[125]  ;
	input \in0[126]  ;
	input \in0[127]  ;
	input \in1[0]  ;
	input \in1[1]  ;
	input \in1[2]  ;
	input \in1[3]  ;
	input \in1[4]  ;
	input \in1[5]  ;
	input \in1[6]  ;
	input \in1[7]  ;
	input \in1[8]  ;
	input \in1[9]  ;
	input \in1[10]  ;
	input \in1[11]  ;
	input \in1[12]  ;
	input \in1[13]  ;
	input \in1[14]  ;
	input \in1[15]  ;
	input \in1[16]  ;
	input \in1[17]  ;
	input \in1[18]  ;
	input \in1[19]  ;
	input \in1[20]  ;
	input \in1[21]  ;
	input \in1[22]  ;
	input \in1[23]  ;
	input \in1[24]  ;
	input \in1[25]  ;
	input \in1[26]  ;
	input \in1[27]  ;
	input \in1[28]  ;
	input \in1[29]  ;
	input \in1[30]  ;
	input \in1[31]  ;
	input \in1[32]  ;
	input \in1[33]  ;
	input \in1[34]  ;
	input \in1[35]  ;
	input \in1[36]  ;
	input \in1[37]  ;
	input \in1[38]  ;
	input \in1[39]  ;
	input \in1[40]  ;
	input \in1[41]  ;
	input \in1[42]  ;
	input \in1[43]  ;
	input \in1[44]  ;
	input \in1[45]  ;
	input \in1[46]  ;
	input \in1[47]  ;
	input \in1[48]  ;
	input \in1[49]  ;
	input \in1[50]  ;
	input \in1[51]  ;
	input \in1[52]  ;
	input \in1[53]  ;
	input \in1[54]  ;
	input \in1[55]  ;
	input \in1[56]  ;
	input \in1[57]  ;
	input \in1[58]  ;
	input \in1[59]  ;
	input \in1[60]  ;
	input \in1[61]  ;
	input \in1[62]  ;
	input \in1[63]  ;
	input \in1[64]  ;
	input \in1[65]  ;
	input \in1[66]  ;
	input \in1[67]  ;
	input \in1[68]  ;
	input \in1[69]  ;
	input \in1[70]  ;
	input \in1[71]  ;
	input \in1[72]  ;
	input \in1[73]  ;
	input \in1[74]  ;
	input \in1[75]  ;
	input \in1[76]  ;
	input \in1[77]  ;
	input \in1[78]  ;
	input \in1[79]  ;
	input \in1[80]  ;
	input \in1[81]  ;
	input \in1[82]  ;
	input \in1[83]  ;
	input \in1[84]  ;
	input \in1[85]  ;
	input \in1[86]  ;
	input \in1[87]  ;
	input \in1[88]  ;
	input \in1[89]  ;
	input \in1[90]  ;
	input \in1[91]  ;
	input \in1[92]  ;
	input \in1[93]  ;
	input \in1[94]  ;
	input \in1[95]  ;
	input \in1[96]  ;
	input \in1[97]  ;
	input \in1[98]  ;
	input \in1[99]  ;
	input \in1[100]  ;
	input \in1[101]  ;
	input \in1[102]  ;
	input \in1[103]  ;
	input \in1[104]  ;
	input \in1[105]  ;
	input \in1[106]  ;
	input \in1[107]  ;
	input \in1[108]  ;
	input \in1[109]  ;
	input \in1[110]  ;
	input \in1[111]  ;
	input \in1[112]  ;
	input \in1[113]  ;
	input \in1[114]  ;
	input \in1[115]  ;
	input \in1[116]  ;
	input \in1[117]  ;
	input \in1[118]  ;
	input \in1[119]  ;
	input \in1[120]  ;
	input \in1[121]  ;
	input \in1[122]  ;
	input \in1[123]  ;
	input \in1[124]  ;
	input \in1[125]  ;
	input \in1[126]  ;
	input \in1[127]  ;
	input \in2[0]  ;
	input \in2[1]  ;
	input \in2[2]  ;
	input \in2[3]  ;
	input \in2[4]  ;
	input \in2[5]  ;
	input \in2[6]  ;
	input \in2[7]  ;
	input \in2[8]  ;
	input \in2[9]  ;
	input \in2[10]  ;
	input \in2[11]  ;
	input \in2[12]  ;
	input \in2[13]  ;
	input \in2[14]  ;
	input \in2[15]  ;
	input \in2[16]  ;
	input \in2[17]  ;
	input \in2[18]  ;
	input \in2[19]  ;
	input \in2[20]  ;
	input \in2[21]  ;
	input \in2[22]  ;
	input \in2[23]  ;
	input \in2[24]  ;
	input \in2[25]  ;
	input \in2[26]  ;
	input \in2[27]  ;
	input \in2[28]  ;
	input \in2[29]  ;
	input \in2[30]  ;
	input \in2[31]  ;
	input \in2[32]  ;
	input \in2[33]  ;
	input \in2[34]  ;
	input \in2[35]  ;
	input \in2[36]  ;
	input \in2[37]  ;
	input \in2[38]  ;
	input \in2[39]  ;
	input \in2[40]  ;
	input \in2[41]  ;
	input \in2[42]  ;
	input \in2[43]  ;
	input \in2[44]  ;
	input \in2[45]  ;
	input \in2[46]  ;
	input \in2[47]  ;
	input \in2[48]  ;
	input \in2[49]  ;
	input \in2[50]  ;
	input \in2[51]  ;
	input \in2[52]  ;
	input \in2[53]  ;
	input \in2[54]  ;
	input \in2[55]  ;
	input \in2[56]  ;
	input \in2[57]  ;
	input \in2[58]  ;
	input \in2[59]  ;
	input \in2[60]  ;
	input \in2[61]  ;
	input \in2[62]  ;
	input \in2[63]  ;
	input \in2[64]  ;
	input \in2[65]  ;
	input \in2[66]  ;
	input \in2[67]  ;
	input \in2[68]  ;
	input \in2[69]  ;
	input \in2[70]  ;
	input \in2[71]  ;
	input \in2[72]  ;
	input \in2[73]  ;
	input \in2[74]  ;
	input \in2[75]  ;
	input \in2[76]  ;
	input \in2[77]  ;
	input \in2[78]  ;
	input \in2[79]  ;
	input \in2[80]  ;
	input \in2[81]  ;
	input \in2[82]  ;
	input \in2[83]  ;
	input \in2[84]  ;
	input \in2[85]  ;
	input \in2[86]  ;
	input \in2[87]  ;
	input \in2[88]  ;
	input \in2[89]  ;
	input \in2[90]  ;
	input \in2[91]  ;
	input \in2[92]  ;
	input \in2[93]  ;
	input \in2[94]  ;
	input \in2[95]  ;
	input \in2[96]  ;
	input \in2[97]  ;
	input \in2[98]  ;
	input \in2[99]  ;
	input \in2[100]  ;
	input \in2[101]  ;
	input \in2[102]  ;
	input \in2[103]  ;
	input \in2[104]  ;
	input \in2[105]  ;
	input \in2[106]  ;
	input \in2[107]  ;
	input \in2[108]  ;
	input \in2[109]  ;
	input \in2[110]  ;
	input \in2[111]  ;
	input \in2[112]  ;
	input \in2[113]  ;
	input \in2[114]  ;
	input \in2[115]  ;
	input \in2[116]  ;
	input \in2[117]  ;
	input \in2[118]  ;
	input \in2[119]  ;
	input \in2[120]  ;
	input \in2[121]  ;
	input \in2[122]  ;
	input \in2[123]  ;
	input \in2[124]  ;
	input \in2[125]  ;
	input \in2[126]  ;
	input \in2[127]  ;
	input \in3[0]  ;
	input \in3[1]  ;
	input \in3[2]  ;
	input \in3[3]  ;
	input \in3[4]  ;
	input \in3[5]  ;
	input \in3[6]  ;
	input \in3[7]  ;
	input \in3[8]  ;
	input \in3[9]  ;
	input \in3[10]  ;
	input \in3[11]  ;
	input \in3[12]  ;
	input \in3[13]  ;
	input \in3[14]  ;
	input \in3[15]  ;
	input \in3[16]  ;
	input \in3[17]  ;
	input \in3[18]  ;
	input \in3[19]  ;
	input \in3[20]  ;
	input \in3[21]  ;
	input \in3[22]  ;
	input \in3[23]  ;
	input \in3[24]  ;
	input \in3[25]  ;
	input \in3[26]  ;
	input \in3[27]  ;
	input \in3[28]  ;
	input \in3[29]  ;
	input \in3[30]  ;
	input \in3[31]  ;
	input \in3[32]  ;
	input \in3[33]  ;
	input \in3[34]  ;
	input \in3[35]  ;
	input \in3[36]  ;
	input \in3[37]  ;
	input \in3[38]  ;
	input \in3[39]  ;
	input \in3[40]  ;
	input \in3[41]  ;
	input \in3[42]  ;
	input \in3[43]  ;
	input \in3[44]  ;
	input \in3[45]  ;
	input \in3[46]  ;
	input \in3[47]  ;
	input \in3[48]  ;
	input \in3[49]  ;
	input \in3[50]  ;
	input \in3[51]  ;
	input \in3[52]  ;
	input \in3[53]  ;
	input \in3[54]  ;
	input \in3[55]  ;
	input \in3[56]  ;
	input \in3[57]  ;
	input \in3[58]  ;
	input \in3[59]  ;
	input \in3[60]  ;
	input \in3[61]  ;
	input \in3[62]  ;
	input \in3[63]  ;
	input \in3[64]  ;
	input \in3[65]  ;
	input \in3[66]  ;
	input \in3[67]  ;
	input \in3[68]  ;
	input \in3[69]  ;
	input \in3[70]  ;
	input \in3[71]  ;
	input \in3[72]  ;
	input \in3[73]  ;
	input \in3[74]  ;
	input \in3[75]  ;
	input \in3[76]  ;
	input \in3[77]  ;
	input \in3[78]  ;
	input \in3[79]  ;
	input \in3[80]  ;
	input \in3[81]  ;
	input \in3[82]  ;
	input \in3[83]  ;
	input \in3[84]  ;
	input \in3[85]  ;
	input \in3[86]  ;
	input \in3[87]  ;
	input \in3[88]  ;
	input \in3[89]  ;
	input \in3[90]  ;
	input \in3[91]  ;
	input \in3[92]  ;
	input \in3[93]  ;
	input \in3[94]  ;
	input \in3[95]  ;
	input \in3[96]  ;
	input \in3[97]  ;
	input \in3[98]  ;
	input \in3[99]  ;
	input \in3[100]  ;
	input \in3[101]  ;
	input \in3[102]  ;
	input \in3[103]  ;
	input \in3[104]  ;
	input \in3[105]  ;
	input \in3[106]  ;
	input \in3[107]  ;
	input \in3[108]  ;
	input \in3[109]  ;
	input \in3[110]  ;
	input \in3[111]  ;
	input \in3[112]  ;
	input \in3[113]  ;
	input \in3[114]  ;
	input \in3[115]  ;
	input \in3[116]  ;
	input \in3[117]  ;
	input \in3[118]  ;
	input \in3[119]  ;
	input \in3[120]  ;
	input \in3[121]  ;
	input \in3[122]  ;
	input \in3[123]  ;
	input \in3[124]  ;
	input \in3[125]  ;
	input \in3[126]  ;
	input \in3[127]  ;
	output \result[0]  ;
	output \result[1]  ;
	output \result[2]  ;
	output \result[3]  ;
	output \result[4]  ;
	output \result[5]  ;
	output \result[6]  ;
	output \result[7]  ;
	output \result[8]  ;
	output \result[9]  ;
	output \result[10]  ;
	output \result[11]  ;
	output \result[12]  ;
	output \result[13]  ;
	output \result[14]  ;
	output \result[15]  ;
	output \result[16]  ;
	output \result[17]  ;
	output \result[18]  ;
	output \result[19]  ;
	output \result[20]  ;
	output \result[21]  ;
	output \result[22]  ;
	output \result[23]  ;
	output \result[24]  ;
	output \result[25]  ;
	output \result[26]  ;
	output \result[27]  ;
	output \result[28]  ;
	output \result[29]  ;
	output \result[30]  ;
	output \result[31]  ;
	output \result[32]  ;
	output \result[33]  ;
	output \result[34]  ;
	output \result[35]  ;
	output \result[36]  ;
	output \result[37]  ;
	output \result[38]  ;
	output \result[39]  ;
	output \result[40]  ;
	output \result[41]  ;
	output \result[42]  ;
	output \result[43]  ;
	output \result[44]  ;
	output \result[45]  ;
	output \result[46]  ;
	output \result[47]  ;
	output \result[48]  ;
	output \result[49]  ;
	output \result[50]  ;
	output \result[51]  ;
	output \result[52]  ;
	output \result[53]  ;
	output \result[54]  ;
	output \result[55]  ;
	output \result[56]  ;
	output \result[57]  ;
	output \result[58]  ;
	output \result[59]  ;
	output \result[60]  ;
	output \result[61]  ;
	output \result[62]  ;
	output \result[63]  ;
	output \result[64]  ;
	output \result[65]  ;
	output \result[66]  ;
	output \result[67]  ;
	output \result[68]  ;
	output \result[69]  ;
	output \result[70]  ;
	output \result[71]  ;
	output \result[72]  ;
	output \result[73]  ;
	output \result[74]  ;
	output \result[75]  ;
	output \result[76]  ;
	output \result[77]  ;
	output \result[78]  ;
	output \result[79]  ;
	output \result[80]  ;
	output \result[81]  ;
	output \result[82]  ;
	output \result[83]  ;
	output \result[84]  ;
	output \result[85]  ;
	output \result[86]  ;
	output \result[87]  ;
	output \result[88]  ;
	output \result[89]  ;
	output \result[90]  ;
	output \result[91]  ;
	output \result[92]  ;
	output \result[93]  ;
	output \result[94]  ;
	output \result[95]  ;
	output \result[96]  ;
	output \result[97]  ;
	output \result[98]  ;
	output \result[99]  ;
	output \result[100]  ;
	output \result[101]  ;
	output \result[102]  ;
	output \result[103]  ;
	output \result[104]  ;
	output \result[105]  ;
	output \result[106]  ;
	output \result[107]  ;
	output \result[108]  ;
	output \result[109]  ;
	output \result[110]  ;
	output \result[111]  ;
	output \result[112]  ;
	output \result[113]  ;
	output \result[114]  ;
	output \result[115]  ;
	output \result[116]  ;
	output \result[117]  ;
	output \result[118]  ;
	output \result[119]  ;
	output \result[120]  ;
	output \result[121]  ;
	output \result[122]  ;
	output \result[123]  ;
	output \result[124]  ;
	output \result[125]  ;
	output \result[126]  ;
	output \result[127]  ;
	output \address[0]  ;
	output \address[1]  ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\in2[127] ,
		\in3[127] ,
		_w513_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\in2[126] ,
		\in3[126] ,
		_w514_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\in2[125] ,
		\in3[125] ,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\in2[124] ,
		\in3[124] ,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\in2[125] ,
		\in3[125] ,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w517_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		_w516_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\in2[126] ,
		\in3[126] ,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w520_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w513_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\in2[127] ,
		\in3[127] ,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\in2[123] ,
		\in3[123] ,
		_w525_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\in2[123] ,
		\in3[123] ,
		_w526_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\in2[122] ,
		\in3[122] ,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w526_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\in2[121] ,
		\in3[121] ,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\in2[122] ,
		\in3[122] ,
		_w530_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\in2[121] ,
		\in3[121] ,
		_w531_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\in2[120] ,
		\in3[120] ,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w531_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w529_,
		_w530_,
		_w534_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w533_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		_w528_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\in2[119] ,
		\in3[119] ,
		_w537_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\in2[119] ,
		\in3[119] ,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		\in2[118] ,
		\in3[118] ,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\in2[118] ,
		\in3[118] ,
		_w541_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\in2[117] ,
		\in3[117] ,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		\in2[117] ,
		\in3[117] ,
		_w543_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\in2[116] ,
		\in3[116] ,
		_w544_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w543_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w541_,
		_w542_,
		_w546_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w545_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w540_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\in2[115] ,
		\in3[115] ,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\in2[115] ,
		\in3[115] ,
		_w550_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\in2[114] ,
		\in3[114] ,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w550_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\in2[113] ,
		\in3[113] ,
		_w553_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\in2[114] ,
		\in3[114] ,
		_w554_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\in2[113] ,
		\in3[113] ,
		_w555_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\in2[112] ,
		\in3[112] ,
		_w556_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w555_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w553_,
		_w554_,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		_w552_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\in2[111] ,
		\in3[111] ,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		\in2[111] ,
		\in3[111] ,
		_w562_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\in2[110] ,
		\in3[110] ,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w562_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\in2[110] ,
		\in3[110] ,
		_w565_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\in2[109] ,
		\in3[109] ,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\in2[109] ,
		\in3[109] ,
		_w567_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\in2[108] ,
		\in3[108] ,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w567_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w565_,
		_w566_,
		_w570_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w564_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\in2[107] ,
		\in3[107] ,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\in2[107] ,
		\in3[107] ,
		_w574_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\in2[106] ,
		\in3[106] ,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w574_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\in2[105] ,
		\in3[105] ,
		_w577_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\in2[106] ,
		\in3[106] ,
		_w578_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\in2[105] ,
		\in3[105] ,
		_w579_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\in2[104] ,
		\in3[104] ,
		_w580_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w579_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w577_,
		_w578_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w581_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		_w576_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\in2[103] ,
		\in3[103] ,
		_w585_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\in2[103] ,
		\in3[103] ,
		_w586_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\in2[102] ,
		\in3[102] ,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\in2[102] ,
		\in3[102] ,
		_w589_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\in2[101] ,
		\in3[101] ,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\in2[101] ,
		\in3[101] ,
		_w591_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\in2[100] ,
		\in3[100] ,
		_w592_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w589_,
		_w590_,
		_w594_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		_w588_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\in2[99] ,
		\in3[99] ,
		_w597_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\in2[99] ,
		\in3[99] ,
		_w598_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\in2[98] ,
		\in3[98] ,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\in2[97] ,
		\in3[97] ,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\in2[98] ,
		\in3[98] ,
		_w602_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\in2[97] ,
		\in3[97] ,
		_w603_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\in2[96] ,
		\in3[96] ,
		_w604_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w603_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w601_,
		_w602_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w605_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w600_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\in2[95] ,
		\in3[95] ,
		_w609_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		\in2[95] ,
		\in3[95] ,
		_w610_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		\in2[94] ,
		\in3[94] ,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w610_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\in2[94] ,
		\in3[94] ,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\in2[93] ,
		\in3[93] ,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\in2[93] ,
		\in3[93] ,
		_w615_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\in2[92] ,
		\in3[92] ,
		_w616_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w615_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w613_,
		_w614_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		_w617_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		_w612_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\in2[91] ,
		\in3[91] ,
		_w621_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		\in2[91] ,
		\in3[91] ,
		_w622_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\in2[90] ,
		\in3[90] ,
		_w623_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w622_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\in2[89] ,
		\in3[89] ,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		\in2[90] ,
		\in3[90] ,
		_w626_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		\in2[89] ,
		\in3[89] ,
		_w627_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\in2[88] ,
		\in3[88] ,
		_w628_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w627_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w625_,
		_w626_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w629_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		_w624_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\in2[87] ,
		\in3[87] ,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		\in2[87] ,
		\in3[87] ,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		\in2[86] ,
		\in3[86] ,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w634_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\in2[86] ,
		\in3[86] ,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\in2[85] ,
		\in3[85] ,
		_w638_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		\in2[85] ,
		\in3[85] ,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\in2[84] ,
		\in3[84] ,
		_w640_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w637_,
		_w638_,
		_w642_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w641_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w636_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		\in2[83] ,
		\in3[83] ,
		_w645_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		\in2[83] ,
		\in3[83] ,
		_w646_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		\in2[82] ,
		\in3[82] ,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w646_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\in2[81] ,
		\in3[81] ,
		_w649_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		\in2[82] ,
		\in3[82] ,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		\in2[81] ,
		\in3[81] ,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\in2[80] ,
		\in3[80] ,
		_w652_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w651_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w649_,
		_w650_,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w653_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		_w648_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\in2[79] ,
		\in3[79] ,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		\in2[79] ,
		\in3[79] ,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		\in2[78] ,
		\in3[78] ,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w658_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\in2[78] ,
		\in3[78] ,
		_w661_
	);
	LUT2 #(
		.INIT('h2)
	) name149 (
		\in2[77] ,
		\in3[77] ,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		\in2[77] ,
		\in3[77] ,
		_w663_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\in2[76] ,
		\in3[76] ,
		_w664_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w663_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w661_,
		_w662_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w665_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		_w660_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\in2[75] ,
		\in3[75] ,
		_w669_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		\in2[75] ,
		\in3[75] ,
		_w670_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		\in2[74] ,
		\in3[74] ,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		_w670_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h2)
	) name160 (
		\in2[73] ,
		\in3[73] ,
		_w673_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		\in2[74] ,
		\in3[74] ,
		_w674_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		\in2[73] ,
		\in3[73] ,
		_w675_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		\in2[72] ,
		\in3[72] ,
		_w676_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w675_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w673_,
		_w674_,
		_w678_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		_w677_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w672_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\in2[71] ,
		\in3[71] ,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\in2[71] ,
		\in3[71] ,
		_w682_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		\in2[70] ,
		\in3[70] ,
		_w683_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\in2[70] ,
		\in3[70] ,
		_w685_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\in2[69] ,
		\in3[69] ,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		\in2[69] ,
		\in3[69] ,
		_w687_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		\in2[68] ,
		\in3[68] ,
		_w688_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w687_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w685_,
		_w686_,
		_w690_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h2)
	) name179 (
		_w684_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h2)
	) name180 (
		\in2[67] ,
		\in3[67] ,
		_w693_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		\in2[67] ,
		\in3[67] ,
		_w694_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		\in2[66] ,
		\in3[66] ,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		\in2[65] ,
		\in3[65] ,
		_w697_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\in2[66] ,
		\in3[66] ,
		_w698_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		\in2[65] ,
		\in3[65] ,
		_w699_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		\in2[64] ,
		\in3[64] ,
		_w700_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w699_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w697_,
		_w698_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w701_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		_w696_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		\in2[63] ,
		\in3[63] ,
		_w705_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		\in2[63] ,
		\in3[63] ,
		_w706_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		\in2[62] ,
		\in3[62] ,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		\in2[61] ,
		\in3[61] ,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\in3[60] ,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\in2[60] ,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		\in2[59] ,
		\in3[59] ,
		_w712_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		\in2[59] ,
		\in3[59] ,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		\in2[58] ,
		\in3[58] ,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w713_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\in2[57] ,
		\in3[57] ,
		_w716_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		\in2[58] ,
		\in3[58] ,
		_w717_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		\in2[57] ,
		\in3[57] ,
		_w718_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		\in2[56] ,
		\in3[56] ,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w718_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w716_,
		_w717_,
		_w721_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		_w720_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w715_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w712_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		\in2[60] ,
		_w709_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w710_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w724_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		\in2[62] ,
		\in3[62] ,
		_w728_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\in2[61] ,
		\in3[61] ,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w728_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w711_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		_w727_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h2)
	) name220 (
		_w708_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\in2[55] ,
		\in3[55] ,
		_w734_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		\in2[55] ,
		\in3[55] ,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		\in2[54] ,
		\in3[54] ,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w735_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		\in2[53] ,
		\in3[53] ,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		\in3[52] ,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		\in2[52] ,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		\in2[51] ,
		\in3[51] ,
		_w741_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		\in2[51] ,
		\in3[51] ,
		_w742_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		\in2[50] ,
		\in3[50] ,
		_w743_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		\in2[49] ,
		\in3[49] ,
		_w745_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		\in2[50] ,
		\in3[50] ,
		_w746_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\in2[49] ,
		\in3[49] ,
		_w747_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		\in2[48] ,
		\in3[48] ,
		_w748_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w747_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w745_,
		_w746_,
		_w750_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w749_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		_w744_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w741_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		\in2[52] ,
		_w738_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w739_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w753_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h2)
	) name244 (
		\in2[53] ,
		\in3[53] ,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\in2[54] ,
		\in3[54] ,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w757_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w740_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		_w756_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		_w737_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\in2[47] ,
		\in3[47] ,
		_w763_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		\in2[47] ,
		\in3[47] ,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		\in2[46] ,
		\in3[46] ,
		_w765_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w764_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		\in2[45] ,
		\in3[45] ,
		_w767_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		\in3[44] ,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\in2[44] ,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		\in2[43] ,
		\in3[43] ,
		_w770_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		\in2[43] ,
		\in3[43] ,
		_w771_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		\in2[42] ,
		\in3[42] ,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w771_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		\in2[41] ,
		\in3[41] ,
		_w774_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		\in2[42] ,
		\in3[42] ,
		_w775_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		\in2[41] ,
		\in3[41] ,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\in2[40] ,
		\in3[40] ,
		_w777_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w776_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w774_,
		_w775_,
		_w779_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w778_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		_w773_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w770_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		\in2[44] ,
		_w767_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w768_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w782_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\in2[46] ,
		\in3[46] ,
		_w786_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		\in2[45] ,
		\in3[45] ,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w786_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		_w769_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		_w785_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		_w766_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\in2[1] ,
		\in3[1] ,
		_w792_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\in2[0] ,
		\in3[0] ,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w792_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		\in2[1] ,
		\in3[1] ,
		_w795_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		\in2[2] ,
		\in3[2] ,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h4)
	) name285 (
		_w794_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		\in2[2] ,
		\in3[2] ,
		_w799_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\in2[3] ,
		\in3[3] ,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w799_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w798_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		\in2[3] ,
		\in3[3] ,
		_w803_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		\in2[4] ,
		\in3[4] ,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w803_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		_w802_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		\in2[4] ,
		\in3[4] ,
		_w807_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		\in2[5] ,
		\in3[5] ,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w807_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w806_,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		\in2[5] ,
		\in3[5] ,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		\in2[6] ,
		\in3[6] ,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w811_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w810_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		\in2[6] ,
		\in3[6] ,
		_w815_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		\in2[7] ,
		\in3[7] ,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w815_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w814_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		\in2[7] ,
		\in3[7] ,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		\in2[8] ,
		\in3[8] ,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w819_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w818_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\in2[8] ,
		\in3[8] ,
		_w823_
	);
	LUT2 #(
		.INIT('h2)
	) name311 (
		\in2[9] ,
		\in3[9] ,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w823_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		_w822_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		\in2[9] ,
		\in3[9] ,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		\in2[10] ,
		\in3[10] ,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w827_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w826_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		\in2[10] ,
		\in3[10] ,
		_w831_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		\in2[11] ,
		\in3[11] ,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w831_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h4)
	) name321 (
		_w830_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		\in2[11] ,
		\in3[11] ,
		_w835_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		\in2[12] ,
		\in3[12] ,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w835_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h4)
	) name325 (
		_w834_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		\in2[12] ,
		\in3[12] ,
		_w839_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		\in2[13] ,
		\in3[13] ,
		_w840_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w839_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w838_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		\in2[13] ,
		\in3[13] ,
		_w843_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		\in2[14] ,
		\in3[14] ,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w843_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w842_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		\in2[14] ,
		\in3[14] ,
		_w847_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		\in2[15] ,
		\in3[15] ,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w846_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		\in2[15] ,
		\in3[15] ,
		_w851_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		\in2[16] ,
		\in3[16] ,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w851_,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w850_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h2)
	) name342 (
		\in2[16] ,
		\in3[16] ,
		_w855_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\in2[17] ,
		\in3[17] ,
		_w856_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w855_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		_w854_,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		\in2[17] ,
		\in3[17] ,
		_w859_
	);
	LUT2 #(
		.INIT('h4)
	) name347 (
		\in2[18] ,
		\in3[18] ,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w859_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w858_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		\in2[18] ,
		\in3[18] ,
		_w863_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\in2[19] ,
		\in3[19] ,
		_w864_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w863_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w862_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\in2[19] ,
		\in3[19] ,
		_w867_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		\in2[20] ,
		\in3[20] ,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w867_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h4)
	) name357 (
		_w866_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\in2[20] ,
		\in3[20] ,
		_w871_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\in2[21] ,
		\in3[21] ,
		_w872_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w871_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w870_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h4)
	) name362 (
		\in2[21] ,
		\in3[21] ,
		_w875_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\in2[22] ,
		\in3[22] ,
		_w876_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w875_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w874_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		\in2[22] ,
		\in3[22] ,
		_w879_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\in2[23] ,
		\in3[23] ,
		_w880_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w879_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		_w878_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		\in2[23] ,
		\in3[23] ,
		_w883_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		\in2[24] ,
		\in3[24] ,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w883_,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		_w882_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		\in2[24] ,
		\in3[24] ,
		_w887_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\in2[25] ,
		\in3[25] ,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w887_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w886_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		\in2[25] ,
		\in3[25] ,
		_w891_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		\in2[26] ,
		\in3[26] ,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w891_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w890_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\in2[26] ,
		\in3[26] ,
		_w895_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\in2[27] ,
		\in3[27] ,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		_w894_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		\in2[27] ,
		\in3[27] ,
		_w899_
	);
	LUT2 #(
		.INIT('h4)
	) name387 (
		\in2[28] ,
		\in3[28] ,
		_w900_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w899_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		_w898_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		\in2[28] ,
		\in3[28] ,
		_w903_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		\in2[29] ,
		\in3[29] ,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w903_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h4)
	) name393 (
		_w902_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		\in2[29] ,
		\in3[29] ,
		_w907_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		\in2[30] ,
		\in3[30] ,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w907_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w906_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h2)
	) name398 (
		\in2[30] ,
		\in3[30] ,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		\in2[31] ,
		\in3[31] ,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w911_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		_w910_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		\in2[32] ,
		\in3[32] ,
		_w915_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		\in2[35] ,
		\in3[35] ,
		_w916_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		\in2[34] ,
		\in3[34] ,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w916_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name406 (
		\in2[39] ,
		\in3[39] ,
		_w919_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		\in2[38] ,
		\in3[38] ,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w919_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		\in2[33] ,
		\in3[33] ,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name410 (
		\in2[31] ,
		\in3[31] ,
		_w923_
	);
	LUT2 #(
		.INIT('h4)
	) name411 (
		\in2[37] ,
		\in3[37] ,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		\in3[36] ,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\in2[36] ,
		_w924_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w925_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w915_,
		_w922_,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w923_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		_w918_,
		_w921_,
		_w930_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		_w929_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		_w927_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w914_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		\in2[39] ,
		\in3[39] ,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\in2[36] ,
		_w925_,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		\in2[35] ,
		\in3[35] ,
		_w936_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		\in2[33] ,
		\in3[33] ,
		_w937_
	);
	LUT2 #(
		.INIT('h2)
	) name425 (
		\in2[34] ,
		\in3[34] ,
		_w938_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		\in2[32] ,
		\in3[32] ,
		_w939_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w922_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w937_,
		_w938_,
		_w941_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		_w940_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		_w918_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w936_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w927_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		\in2[38] ,
		\in3[38] ,
		_w946_
	);
	LUT2 #(
		.INIT('h2)
	) name434 (
		\in2[37] ,
		\in3[37] ,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w946_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		_w935_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w945_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		_w921_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w934_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w933_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h4)
	) name441 (
		\in2[40] ,
		\in3[40] ,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w776_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w766_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w773_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w784_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w953_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w763_,
		_w791_,
		_w960_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		\in2[48] ,
		\in3[48] ,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w747_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w737_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		_w744_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		_w755_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		_w961_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		_w734_,
		_w762_,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		_w967_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		\in2[56] ,
		\in3[56] ,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w718_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w708_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h8)
	) name460 (
		_w715_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		_w726_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w969_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w705_,
		_w733_,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		_w975_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h4)
	) name465 (
		\in2[64] ,
		\in3[64] ,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w699_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w696_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		_w977_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w693_,
		_w704_,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		_w981_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		\in2[68] ,
		\in3[68] ,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w687_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w684_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		_w983_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w681_,
		_w692_,
		_w988_
	);
	LUT2 #(
		.INIT('h4)
	) name476 (
		_w987_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		\in2[72] ,
		\in3[72] ,
		_w990_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w675_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w672_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h4)
	) name480 (
		_w989_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w669_,
		_w680_,
		_w994_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		_w993_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		\in2[76] ,
		\in3[76] ,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w663_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		_w660_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		_w995_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w657_,
		_w668_,
		_w1000_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		\in2[80] ,
		\in3[80] ,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w651_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		_w648_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h4)
	) name492 (
		_w1001_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w645_,
		_w656_,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		_w1005_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		\in2[84] ,
		\in3[84] ,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w639_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w636_,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		_w1007_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		_w633_,
		_w644_,
		_w1012_
	);
	LUT2 #(
		.INIT('h4)
	) name500 (
		_w1011_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		\in2[88] ,
		\in3[88] ,
		_w1014_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w627_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		_w624_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h4)
	) name504 (
		_w1013_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w621_,
		_w632_,
		_w1018_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		\in2[92] ,
		\in3[92] ,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w615_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		_w612_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		_w1019_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w609_,
		_w620_,
		_w1024_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		\in2[96] ,
		\in3[96] ,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w603_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		_w600_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w1025_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w597_,
		_w608_,
		_w1030_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		_w1029_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		\in2[100] ,
		\in3[100] ,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w591_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		_w588_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		_w1031_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w585_,
		_w596_,
		_w1036_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w1035_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		\in2[104] ,
		\in3[104] ,
		_w1038_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w579_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		_w576_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		_w1037_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w573_,
		_w584_,
		_w1042_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w1041_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		\in2[108] ,
		\in3[108] ,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w567_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		_w564_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		_w1043_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w561_,
		_w572_,
		_w1048_
	);
	LUT2 #(
		.INIT('h4)
	) name536 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		\in2[112] ,
		\in3[112] ,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w555_,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		_w552_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w1049_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w549_,
		_w560_,
		_w1054_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w1053_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		\in2[116] ,
		\in3[116] ,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w543_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		_w540_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w1055_,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w537_,
		_w548_,
		_w1060_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w1059_,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h4)
	) name549 (
		\in2[120] ,
		\in3[120] ,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w531_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		_w528_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w1061_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w525_,
		_w536_,
		_w1066_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w1065_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		\in2[124] ,
		\in3[124] ,
		_w1068_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w513_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		_w516_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		_w1067_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		_w523_,
		_w524_,
		_w1072_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		\in2[0] ,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h8)
	) name562 (
		\in3[0] ,
		_w1073_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w1074_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h2)
	) name564 (
		\in0[127] ,
		\in1[127] ,
		_w1077_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		\in0[126] ,
		\in1[126] ,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		\in0[125] ,
		\in1[125] ,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h2)
	) name568 (
		\in0[124] ,
		\in1[124] ,
		_w1081_
	);
	LUT2 #(
		.INIT('h2)
	) name569 (
		\in0[125] ,
		\in1[125] ,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w1081_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w1080_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		\in0[126] ,
		\in1[126] ,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w1084_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w1077_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		\in0[127] ,
		\in1[127] ,
		_w1088_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		\in0[123] ,
		\in1[123] ,
		_w1089_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\in0[123] ,
		\in1[123] ,
		_w1090_
	);
	LUT2 #(
		.INIT('h4)
	) name578 (
		\in0[122] ,
		\in1[122] ,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		\in0[121] ,
		\in1[121] ,
		_w1093_
	);
	LUT2 #(
		.INIT('h2)
	) name581 (
		\in0[122] ,
		\in1[122] ,
		_w1094_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		\in0[121] ,
		\in1[121] ,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		\in0[120] ,
		\in1[120] ,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w1093_,
		_w1094_,
		_w1098_
	);
	LUT2 #(
		.INIT('h4)
	) name586 (
		_w1097_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		_w1092_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		\in0[119] ,
		\in1[119] ,
		_w1101_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		\in0[119] ,
		\in1[119] ,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		\in0[118] ,
		\in1[118] ,
		_w1103_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		\in0[118] ,
		\in1[118] ,
		_w1105_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		\in0[117] ,
		\in1[117] ,
		_w1106_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		\in0[117] ,
		\in1[117] ,
		_w1107_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		\in0[116] ,
		\in1[116] ,
		_w1108_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w1105_,
		_w1106_,
		_w1110_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		_w1104_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		\in0[115] ,
		\in1[115] ,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		\in0[115] ,
		\in1[115] ,
		_w1114_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		\in0[114] ,
		\in1[114] ,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w1114_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		\in0[113] ,
		\in1[113] ,
		_w1117_
	);
	LUT2 #(
		.INIT('h2)
	) name605 (
		\in0[114] ,
		\in1[114] ,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		\in0[113] ,
		\in1[113] ,
		_w1119_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		\in0[112] ,
		\in1[112] ,
		_w1120_
	);
	LUT2 #(
		.INIT('h4)
	) name608 (
		_w1119_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w1117_,
		_w1118_,
		_w1122_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h2)
	) name611 (
		_w1116_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h2)
	) name612 (
		\in0[111] ,
		\in1[111] ,
		_w1125_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		\in0[111] ,
		\in1[111] ,
		_w1126_
	);
	LUT2 #(
		.INIT('h4)
	) name614 (
		\in0[110] ,
		\in1[110] ,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w1126_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		\in0[110] ,
		\in1[110] ,
		_w1129_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		\in0[109] ,
		\in1[109] ,
		_w1130_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		\in0[109] ,
		\in1[109] ,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name619 (
		\in0[108] ,
		\in1[108] ,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w1129_,
		_w1130_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		_w1133_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		_w1128_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h2)
	) name624 (
		\in0[107] ,
		\in1[107] ,
		_w1137_
	);
	LUT2 #(
		.INIT('h4)
	) name625 (
		\in0[107] ,
		\in1[107] ,
		_w1138_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		\in0[106] ,
		\in1[106] ,
		_w1139_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		_w1138_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		\in0[105] ,
		\in1[105] ,
		_w1141_
	);
	LUT2 #(
		.INIT('h2)
	) name629 (
		\in0[106] ,
		\in1[106] ,
		_w1142_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		\in0[105] ,
		\in1[105] ,
		_w1143_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		\in0[104] ,
		\in1[104] ,
		_w1144_
	);
	LUT2 #(
		.INIT('h4)
	) name632 (
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w1141_,
		_w1142_,
		_w1146_
	);
	LUT2 #(
		.INIT('h4)
	) name634 (
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h2)
	) name635 (
		_w1140_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h2)
	) name636 (
		\in0[103] ,
		\in1[103] ,
		_w1149_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		\in0[103] ,
		\in1[103] ,
		_w1150_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		\in0[102] ,
		\in1[102] ,
		_w1151_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w1150_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		\in0[102] ,
		\in1[102] ,
		_w1153_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		\in0[101] ,
		\in1[101] ,
		_w1154_
	);
	LUT2 #(
		.INIT('h4)
	) name642 (
		\in0[101] ,
		\in1[101] ,
		_w1155_
	);
	LUT2 #(
		.INIT('h2)
	) name643 (
		\in0[100] ,
		\in1[100] ,
		_w1156_
	);
	LUT2 #(
		.INIT('h4)
	) name644 (
		_w1155_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w1153_,
		_w1154_,
		_w1158_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w1157_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h2)
	) name647 (
		_w1152_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		\in0[99] ,
		\in1[99] ,
		_w1161_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		\in0[99] ,
		\in1[99] ,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name650 (
		\in0[98] ,
		\in1[98] ,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w1162_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		\in0[97] ,
		\in1[97] ,
		_w1165_
	);
	LUT2 #(
		.INIT('h2)
	) name653 (
		\in0[98] ,
		\in1[98] ,
		_w1166_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		\in0[97] ,
		\in1[97] ,
		_w1167_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		\in0[96] ,
		\in1[96] ,
		_w1168_
	);
	LUT2 #(
		.INIT('h4)
	) name656 (
		_w1167_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w1165_,
		_w1166_,
		_w1170_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w1169_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		_w1164_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h2)
	) name660 (
		\in0[95] ,
		\in1[95] ,
		_w1173_
	);
	LUT2 #(
		.INIT('h4)
	) name661 (
		\in0[95] ,
		\in1[95] ,
		_w1174_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		\in0[94] ,
		\in1[94] ,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w1174_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		\in0[94] ,
		\in1[94] ,
		_w1177_
	);
	LUT2 #(
		.INIT('h2)
	) name665 (
		\in0[93] ,
		\in1[93] ,
		_w1178_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		\in0[93] ,
		\in1[93] ,
		_w1179_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		\in0[92] ,
		\in1[92] ,
		_w1180_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		_w1179_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		_w1177_,
		_w1178_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name670 (
		_w1181_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		_w1176_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		\in0[91] ,
		\in1[91] ,
		_w1185_
	);
	LUT2 #(
		.INIT('h4)
	) name673 (
		\in0[91] ,
		\in1[91] ,
		_w1186_
	);
	LUT2 #(
		.INIT('h4)
	) name674 (
		\in0[90] ,
		\in1[90] ,
		_w1187_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w1186_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		\in0[89] ,
		\in1[89] ,
		_w1189_
	);
	LUT2 #(
		.INIT('h2)
	) name677 (
		\in0[90] ,
		\in1[90] ,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name678 (
		\in0[89] ,
		\in1[89] ,
		_w1191_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		\in0[88] ,
		\in1[88] ,
		_w1192_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w1189_,
		_w1190_,
		_w1194_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		_w1193_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		_w1188_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		\in0[87] ,
		\in1[87] ,
		_w1197_
	);
	LUT2 #(
		.INIT('h4)
	) name685 (
		\in0[87] ,
		\in1[87] ,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		\in0[86] ,
		\in1[86] ,
		_w1199_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w1198_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h2)
	) name688 (
		\in0[86] ,
		\in1[86] ,
		_w1201_
	);
	LUT2 #(
		.INIT('h2)
	) name689 (
		\in0[85] ,
		\in1[85] ,
		_w1202_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		\in0[85] ,
		\in1[85] ,
		_w1203_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		\in0[84] ,
		\in1[84] ,
		_w1204_
	);
	LUT2 #(
		.INIT('h4)
	) name692 (
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w1201_,
		_w1202_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		_w1200_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		\in0[83] ,
		\in1[83] ,
		_w1209_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		\in0[83] ,
		\in1[83] ,
		_w1210_
	);
	LUT2 #(
		.INIT('h4)
	) name698 (
		\in0[82] ,
		\in1[82] ,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w1210_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		\in0[81] ,
		\in1[81] ,
		_w1213_
	);
	LUT2 #(
		.INIT('h2)
	) name701 (
		\in0[82] ,
		\in1[82] ,
		_w1214_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		\in0[81] ,
		\in1[81] ,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name703 (
		\in0[80] ,
		\in1[80] ,
		_w1216_
	);
	LUT2 #(
		.INIT('h4)
	) name704 (
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		_w1213_,
		_w1214_,
		_w1218_
	);
	LUT2 #(
		.INIT('h4)
	) name706 (
		_w1217_,
		_w1218_,
		_w1219_
	);
	LUT2 #(
		.INIT('h2)
	) name707 (
		_w1212_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h2)
	) name708 (
		\in0[79] ,
		\in1[79] ,
		_w1221_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		\in0[79] ,
		\in1[79] ,
		_w1222_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		\in0[78] ,
		\in1[78] ,
		_w1223_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w1222_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		\in0[78] ,
		\in1[78] ,
		_w1225_
	);
	LUT2 #(
		.INIT('h2)
	) name713 (
		\in0[77] ,
		\in1[77] ,
		_w1226_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		\in0[77] ,
		\in1[77] ,
		_w1227_
	);
	LUT2 #(
		.INIT('h2)
	) name715 (
		\in0[76] ,
		\in1[76] ,
		_w1228_
	);
	LUT2 #(
		.INIT('h4)
	) name716 (
		_w1227_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w1225_,
		_w1226_,
		_w1230_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		_w1224_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h2)
	) name720 (
		\in0[75] ,
		\in1[75] ,
		_w1233_
	);
	LUT2 #(
		.INIT('h4)
	) name721 (
		\in0[75] ,
		\in1[75] ,
		_w1234_
	);
	LUT2 #(
		.INIT('h4)
	) name722 (
		\in0[74] ,
		\in1[74] ,
		_w1235_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w1234_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h2)
	) name724 (
		\in0[73] ,
		\in1[73] ,
		_w1237_
	);
	LUT2 #(
		.INIT('h2)
	) name725 (
		\in0[74] ,
		\in1[74] ,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		\in0[73] ,
		\in1[73] ,
		_w1239_
	);
	LUT2 #(
		.INIT('h2)
	) name727 (
		\in0[72] ,
		\in1[72] ,
		_w1240_
	);
	LUT2 #(
		.INIT('h4)
	) name728 (
		_w1239_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		_w1237_,
		_w1238_,
		_w1242_
	);
	LUT2 #(
		.INIT('h4)
	) name730 (
		_w1241_,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		_w1236_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h2)
	) name732 (
		\in0[71] ,
		\in1[71] ,
		_w1245_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		\in0[71] ,
		\in1[71] ,
		_w1246_
	);
	LUT2 #(
		.INIT('h4)
	) name734 (
		\in0[70] ,
		\in1[70] ,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w1246_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h2)
	) name736 (
		\in0[70] ,
		\in1[70] ,
		_w1249_
	);
	LUT2 #(
		.INIT('h2)
	) name737 (
		\in0[69] ,
		\in1[69] ,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		\in0[69] ,
		\in1[69] ,
		_w1251_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		\in0[68] ,
		\in1[68] ,
		_w1252_
	);
	LUT2 #(
		.INIT('h4)
	) name740 (
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w1249_,
		_w1250_,
		_w1254_
	);
	LUT2 #(
		.INIT('h4)
	) name742 (
		_w1253_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h2)
	) name743 (
		_w1248_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		\in0[67] ,
		\in1[67] ,
		_w1257_
	);
	LUT2 #(
		.INIT('h4)
	) name745 (
		\in0[67] ,
		\in1[67] ,
		_w1258_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		\in0[66] ,
		\in1[66] ,
		_w1259_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h2)
	) name748 (
		\in0[65] ,
		\in1[65] ,
		_w1261_
	);
	LUT2 #(
		.INIT('h2)
	) name749 (
		\in0[66] ,
		\in1[66] ,
		_w1262_
	);
	LUT2 #(
		.INIT('h4)
	) name750 (
		\in0[65] ,
		\in1[65] ,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		\in0[64] ,
		\in1[64] ,
		_w1264_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w1261_,
		_w1262_,
		_w1266_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		_w1265_,
		_w1266_,
		_w1267_
	);
	LUT2 #(
		.INIT('h2)
	) name755 (
		_w1260_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h2)
	) name756 (
		\in0[63] ,
		\in1[63] ,
		_w1269_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		\in0[63] ,
		\in1[63] ,
		_w1270_
	);
	LUT2 #(
		.INIT('h4)
	) name758 (
		\in0[62] ,
		\in1[62] ,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w1270_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h4)
	) name760 (
		\in0[61] ,
		\in1[61] ,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		\in1[60] ,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name762 (
		\in0[60] ,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h2)
	) name763 (
		\in0[59] ,
		\in1[59] ,
		_w1276_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		\in0[59] ,
		\in1[59] ,
		_w1277_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		\in0[58] ,
		\in1[58] ,
		_w1278_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		_w1277_,
		_w1278_,
		_w1279_
	);
	LUT2 #(
		.INIT('h2)
	) name767 (
		\in0[57] ,
		\in1[57] ,
		_w1280_
	);
	LUT2 #(
		.INIT('h2)
	) name768 (
		\in0[58] ,
		\in1[58] ,
		_w1281_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		\in0[57] ,
		\in1[57] ,
		_w1282_
	);
	LUT2 #(
		.INIT('h2)
	) name770 (
		\in0[56] ,
		\in1[56] ,
		_w1283_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w1282_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w1280_,
		_w1281_,
		_w1285_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT2 #(
		.INIT('h2)
	) name774 (
		_w1279_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w1276_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h2)
	) name776 (
		\in0[60] ,
		_w1273_,
		_w1289_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w1274_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		_w1288_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		\in0[62] ,
		\in1[62] ,
		_w1292_
	);
	LUT2 #(
		.INIT('h2)
	) name780 (
		\in0[61] ,
		\in1[61] ,
		_w1293_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w1292_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w1275_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		_w1291_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h2)
	) name784 (
		_w1272_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h2)
	) name785 (
		\in0[55] ,
		\in1[55] ,
		_w1298_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		\in0[55] ,
		\in1[55] ,
		_w1299_
	);
	LUT2 #(
		.INIT('h4)
	) name787 (
		\in0[54] ,
		\in1[54] ,
		_w1300_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		_w1299_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h4)
	) name789 (
		\in0[53] ,
		\in1[53] ,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		\in1[52] ,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		\in0[52] ,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		\in0[51] ,
		\in1[51] ,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name793 (
		\in0[51] ,
		\in1[51] ,
		_w1306_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		\in0[50] ,
		\in1[50] ,
		_w1307_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w1306_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\in0[49] ,
		\in1[49] ,
		_w1309_
	);
	LUT2 #(
		.INIT('h2)
	) name797 (
		\in0[50] ,
		\in1[50] ,
		_w1310_
	);
	LUT2 #(
		.INIT('h4)
	) name798 (
		\in0[49] ,
		\in1[49] ,
		_w1311_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		\in0[48] ,
		\in1[48] ,
		_w1312_
	);
	LUT2 #(
		.INIT('h4)
	) name800 (
		_w1311_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w1309_,
		_w1310_,
		_w1314_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		_w1313_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		_w1308_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w1305_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h2)
	) name805 (
		\in0[52] ,
		_w1302_,
		_w1318_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		_w1303_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w1317_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h2)
	) name808 (
		\in0[53] ,
		\in1[53] ,
		_w1321_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\in0[54] ,
		\in1[54] ,
		_w1322_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w1321_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h4)
	) name811 (
		_w1304_,
		_w1323_,
		_w1324_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		_w1320_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h2)
	) name813 (
		_w1301_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h2)
	) name814 (
		\in0[47] ,
		\in1[47] ,
		_w1327_
	);
	LUT2 #(
		.INIT('h4)
	) name815 (
		\in0[47] ,
		\in1[47] ,
		_w1328_
	);
	LUT2 #(
		.INIT('h4)
	) name816 (
		\in0[46] ,
		\in1[46] ,
		_w1329_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w1328_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		\in0[45] ,
		\in1[45] ,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		\in1[44] ,
		_w1331_,
		_w1332_
	);
	LUT2 #(
		.INIT('h8)
	) name820 (
		\in0[44] ,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h2)
	) name821 (
		\in0[43] ,
		\in1[43] ,
		_w1334_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		\in0[43] ,
		\in1[43] ,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name823 (
		\in0[42] ,
		\in1[42] ,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h2)
	) name825 (
		\in0[41] ,
		\in1[41] ,
		_w1338_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		\in0[42] ,
		\in1[42] ,
		_w1339_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		\in0[41] ,
		\in1[41] ,
		_w1340_
	);
	LUT2 #(
		.INIT('h2)
	) name828 (
		\in0[40] ,
		\in1[40] ,
		_w1341_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		_w1340_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w1338_,
		_w1339_,
		_w1343_
	);
	LUT2 #(
		.INIT('h4)
	) name831 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		_w1337_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w1334_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		\in0[44] ,
		_w1331_,
		_w1347_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w1332_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w1346_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		\in0[46] ,
		\in1[46] ,
		_w1350_
	);
	LUT2 #(
		.INIT('h2)
	) name838 (
		\in0[45] ,
		\in1[45] ,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w1350_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w1333_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		_w1349_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		_w1330_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h2)
	) name843 (
		\in0[1] ,
		\in1[1] ,
		_w1356_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		\in0[0] ,
		\in1[0] ,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		\in0[1] ,
		\in1[1] ,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name847 (
		\in0[2] ,
		\in1[2] ,
		_w1360_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w1358_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		\in0[2] ,
		\in1[2] ,
		_w1363_
	);
	LUT2 #(
		.INIT('h2)
	) name851 (
		\in0[3] ,
		\in1[3] ,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w1363_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h4)
	) name853 (
		_w1362_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		\in0[3] ,
		\in1[3] ,
		_w1367_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		\in0[4] ,
		\in1[4] ,
		_w1368_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w1367_,
		_w1368_,
		_w1369_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w1366_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		\in0[4] ,
		\in1[4] ,
		_w1371_
	);
	LUT2 #(
		.INIT('h2)
	) name859 (
		\in0[5] ,
		\in1[5] ,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h4)
	) name861 (
		_w1370_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h4)
	) name862 (
		\in0[5] ,
		\in1[5] ,
		_w1375_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		\in0[6] ,
		\in1[6] ,
		_w1376_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w1375_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h4)
	) name865 (
		_w1374_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h2)
	) name866 (
		\in0[6] ,
		\in1[6] ,
		_w1379_
	);
	LUT2 #(
		.INIT('h2)
	) name867 (
		\in0[7] ,
		\in1[7] ,
		_w1380_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1379_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w1378_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		\in0[7] ,
		\in1[7] ,
		_w1383_
	);
	LUT2 #(
		.INIT('h4)
	) name871 (
		\in0[8] ,
		\in1[8] ,
		_w1384_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h4)
	) name873 (
		_w1382_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		\in0[8] ,
		\in1[8] ,
		_w1387_
	);
	LUT2 #(
		.INIT('h2)
	) name875 (
		\in0[9] ,
		\in1[9] ,
		_w1388_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w1387_,
		_w1388_,
		_w1389_
	);
	LUT2 #(
		.INIT('h4)
	) name877 (
		_w1386_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		\in0[9] ,
		\in1[9] ,
		_w1391_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		\in0[10] ,
		\in1[10] ,
		_w1392_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		_w1391_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h4)
	) name881 (
		_w1390_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		\in0[10] ,
		\in1[10] ,
		_w1395_
	);
	LUT2 #(
		.INIT('h2)
	) name883 (
		\in0[11] ,
		\in1[11] ,
		_w1396_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1395_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		_w1394_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		\in0[11] ,
		\in1[11] ,
		_w1399_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		\in0[12] ,
		\in1[12] ,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		_w1399_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		_w1398_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name890 (
		\in0[12] ,
		\in1[12] ,
		_w1403_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		\in0[13] ,
		\in1[13] ,
		_w1404_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1403_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		_w1402_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		\in0[13] ,
		\in1[13] ,
		_w1407_
	);
	LUT2 #(
		.INIT('h4)
	) name895 (
		\in0[14] ,
		\in1[14] ,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w1406_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		\in0[14] ,
		\in1[14] ,
		_w1411_
	);
	LUT2 #(
		.INIT('h2)
	) name899 (
		\in0[15] ,
		\in1[15] ,
		_w1412_
	);
	LUT2 #(
		.INIT('h1)
	) name900 (
		_w1411_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h4)
	) name901 (
		_w1410_,
		_w1413_,
		_w1414_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		\in0[15] ,
		\in1[15] ,
		_w1415_
	);
	LUT2 #(
		.INIT('h4)
	) name903 (
		\in0[16] ,
		\in1[16] ,
		_w1416_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		_w1415_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h4)
	) name905 (
		_w1414_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h2)
	) name906 (
		\in0[16] ,
		\in1[16] ,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name907 (
		\in0[17] ,
		\in1[17] ,
		_w1420_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w1419_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h4)
	) name909 (
		_w1418_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		\in0[17] ,
		\in1[17] ,
		_w1423_
	);
	LUT2 #(
		.INIT('h4)
	) name911 (
		\in0[18] ,
		\in1[18] ,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name913 (
		_w1422_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h2)
	) name914 (
		\in0[18] ,
		\in1[18] ,
		_w1427_
	);
	LUT2 #(
		.INIT('h2)
	) name915 (
		\in0[19] ,
		\in1[19] ,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w1427_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		_w1426_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name918 (
		\in0[19] ,
		\in1[19] ,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name919 (
		\in0[20] ,
		\in1[20] ,
		_w1432_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		_w1430_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h2)
	) name922 (
		\in0[20] ,
		\in1[20] ,
		_w1435_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		\in0[21] ,
		\in1[21] ,
		_w1436_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1435_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h4)
	) name925 (
		_w1434_,
		_w1437_,
		_w1438_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		\in0[21] ,
		\in1[21] ,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name927 (
		\in0[22] ,
		\in1[22] ,
		_w1440_
	);
	LUT2 #(
		.INIT('h1)
	) name928 (
		_w1439_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		_w1438_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h2)
	) name930 (
		\in0[22] ,
		\in1[22] ,
		_w1443_
	);
	LUT2 #(
		.INIT('h2)
	) name931 (
		\in0[23] ,
		\in1[23] ,
		_w1444_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h4)
	) name933 (
		_w1442_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		\in0[23] ,
		\in1[23] ,
		_w1447_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		\in0[24] ,
		\in1[24] ,
		_w1448_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1447_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h4)
	) name937 (
		_w1446_,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		\in0[24] ,
		\in1[24] ,
		_w1451_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\in0[25] ,
		\in1[25] ,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w1451_,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w1450_,
		_w1453_,
		_w1454_
	);
	LUT2 #(
		.INIT('h4)
	) name942 (
		\in0[25] ,
		\in1[25] ,
		_w1455_
	);
	LUT2 #(
		.INIT('h4)
	) name943 (
		\in0[26] ,
		\in1[26] ,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w1455_,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h4)
	) name945 (
		_w1454_,
		_w1457_,
		_w1458_
	);
	LUT2 #(
		.INIT('h2)
	) name946 (
		\in0[26] ,
		\in1[26] ,
		_w1459_
	);
	LUT2 #(
		.INIT('h2)
	) name947 (
		\in0[27] ,
		\in1[27] ,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w1459_,
		_w1460_,
		_w1461_
	);
	LUT2 #(
		.INIT('h4)
	) name949 (
		_w1458_,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		\in0[27] ,
		\in1[27] ,
		_w1463_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		\in0[28] ,
		\in1[28] ,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w1463_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h4)
	) name953 (
		_w1462_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		\in0[28] ,
		\in1[28] ,
		_w1467_
	);
	LUT2 #(
		.INIT('h2)
	) name955 (
		\in0[29] ,
		\in1[29] ,
		_w1468_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w1467_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h4)
	) name957 (
		_w1466_,
		_w1469_,
		_w1470_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		\in0[29] ,
		\in1[29] ,
		_w1471_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		\in0[30] ,
		\in1[30] ,
		_w1472_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT2 #(
		.INIT('h4)
	) name961 (
		_w1470_,
		_w1473_,
		_w1474_
	);
	LUT2 #(
		.INIT('h2)
	) name962 (
		\in0[30] ,
		\in1[30] ,
		_w1475_
	);
	LUT2 #(
		.INIT('h2)
	) name963 (
		\in0[31] ,
		\in1[31] ,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		_w1475_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w1474_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h4)
	) name966 (
		\in0[32] ,
		\in1[32] ,
		_w1479_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		\in0[35] ,
		\in1[35] ,
		_w1480_
	);
	LUT2 #(
		.INIT('h4)
	) name968 (
		\in0[34] ,
		\in1[34] ,
		_w1481_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		_w1480_,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h4)
	) name970 (
		\in0[39] ,
		\in1[39] ,
		_w1483_
	);
	LUT2 #(
		.INIT('h4)
	) name971 (
		\in0[38] ,
		\in1[38] ,
		_w1484_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		_w1483_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h4)
	) name973 (
		\in0[33] ,
		\in1[33] ,
		_w1486_
	);
	LUT2 #(
		.INIT('h4)
	) name974 (
		\in0[31] ,
		\in1[31] ,
		_w1487_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		\in0[37] ,
		\in1[37] ,
		_w1488_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		\in1[36] ,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h2)
	) name977 (
		\in0[36] ,
		_w1488_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		_w1489_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1479_,
		_w1486_,
		_w1492_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		_w1487_,
		_w1492_,
		_w1493_
	);
	LUT2 #(
		.INIT('h8)
	) name981 (
		_w1482_,
		_w1485_,
		_w1494_
	);
	LUT2 #(
		.INIT('h8)
	) name982 (
		_w1493_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h4)
	) name983 (
		_w1491_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h4)
	) name984 (
		_w1478_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h2)
	) name985 (
		\in0[39] ,
		\in1[39] ,
		_w1498_
	);
	LUT2 #(
		.INIT('h8)
	) name986 (
		\in0[36] ,
		_w1489_,
		_w1499_
	);
	LUT2 #(
		.INIT('h2)
	) name987 (
		\in0[35] ,
		\in1[35] ,
		_w1500_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		\in0[33] ,
		\in1[33] ,
		_w1501_
	);
	LUT2 #(
		.INIT('h2)
	) name989 (
		\in0[34] ,
		\in1[34] ,
		_w1502_
	);
	LUT2 #(
		.INIT('h2)
	) name990 (
		\in0[32] ,
		\in1[32] ,
		_w1503_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		_w1486_,
		_w1503_,
		_w1504_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		_w1501_,
		_w1502_,
		_w1505_
	);
	LUT2 #(
		.INIT('h4)
	) name993 (
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h2)
	) name994 (
		_w1482_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w1500_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		_w1491_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h2)
	) name997 (
		\in0[38] ,
		\in1[38] ,
		_w1510_
	);
	LUT2 #(
		.INIT('h2)
	) name998 (
		\in0[37] ,
		\in1[37] ,
		_w1511_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h4)
	) name1000 (
		_w1499_,
		_w1512_,
		_w1513_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w1509_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h2)
	) name1002 (
		_w1485_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1498_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		_w1497_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		\in0[40] ,
		\in1[40] ,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w1340_,
		_w1518_,
		_w1519_
	);
	LUT2 #(
		.INIT('h8)
	) name1007 (
		_w1330_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		_w1337_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h4)
	) name1009 (
		_w1348_,
		_w1521_,
		_w1522_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w1517_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w1327_,
		_w1355_,
		_w1524_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		_w1523_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		\in0[48] ,
		\in1[48] ,
		_w1526_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		_w1311_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		_w1301_,
		_w1527_,
		_w1528_
	);
	LUT2 #(
		.INIT('h8)
	) name1016 (
		_w1308_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h4)
	) name1017 (
		_w1319_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		_w1525_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		_w1298_,
		_w1326_,
		_w1532_
	);
	LUT2 #(
		.INIT('h4)
	) name1020 (
		_w1531_,
		_w1532_,
		_w1533_
	);
	LUT2 #(
		.INIT('h4)
	) name1021 (
		\in0[56] ,
		\in1[56] ,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		_w1282_,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name1023 (
		_w1272_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name1024 (
		_w1279_,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h4)
	) name1025 (
		_w1290_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		_w1533_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w1269_,
		_w1297_,
		_w1540_
	);
	LUT2 #(
		.INIT('h4)
	) name1028 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		\in0[64] ,
		\in1[64] ,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w1263_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h8)
	) name1031 (
		_w1260_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		_w1541_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		_w1257_,
		_w1268_,
		_w1546_
	);
	LUT2 #(
		.INIT('h4)
	) name1034 (
		_w1545_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		\in0[68] ,
		\in1[68] ,
		_w1548_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w1251_,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		_w1248_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h4)
	) name1038 (
		_w1547_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name1039 (
		_w1245_,
		_w1256_,
		_w1552_
	);
	LUT2 #(
		.INIT('h4)
	) name1040 (
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h4)
	) name1041 (
		\in0[72] ,
		\in1[72] ,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w1239_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		_w1236_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h4)
	) name1044 (
		_w1553_,
		_w1556_,
		_w1557_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w1233_,
		_w1244_,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name1046 (
		_w1557_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		\in0[76] ,
		\in1[76] ,
		_w1560_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		_w1227_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		_w1224_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h4)
	) name1050 (
		_w1559_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		_w1221_,
		_w1232_,
		_w1564_
	);
	LUT2 #(
		.INIT('h4)
	) name1052 (
		_w1563_,
		_w1564_,
		_w1565_
	);
	LUT2 #(
		.INIT('h4)
	) name1053 (
		\in0[80] ,
		\in1[80] ,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		_w1215_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		_w1212_,
		_w1567_,
		_w1568_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		_w1565_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w1209_,
		_w1220_,
		_w1570_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		\in0[84] ,
		\in1[84] ,
		_w1572_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w1203_,
		_w1572_,
		_w1573_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		_w1200_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		_w1571_,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h1)
	) name1063 (
		_w1197_,
		_w1208_,
		_w1576_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w1575_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		\in0[88] ,
		\in1[88] ,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		_w1191_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		_w1188_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h4)
	) name1068 (
		_w1577_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h1)
	) name1069 (
		_w1185_,
		_w1196_,
		_w1582_
	);
	LUT2 #(
		.INIT('h4)
	) name1070 (
		_w1581_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h4)
	) name1071 (
		\in0[92] ,
		\in1[92] ,
		_w1584_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w1179_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		_w1176_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		_w1583_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h1)
	) name1075 (
		_w1173_,
		_w1184_,
		_w1588_
	);
	LUT2 #(
		.INIT('h4)
	) name1076 (
		_w1587_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h4)
	) name1077 (
		\in0[96] ,
		\in1[96] ,
		_w1590_
	);
	LUT2 #(
		.INIT('h1)
	) name1078 (
		_w1167_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('h8)
	) name1079 (
		_w1164_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		_w1589_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w1161_,
		_w1172_,
		_w1594_
	);
	LUT2 #(
		.INIT('h4)
	) name1082 (
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h4)
	) name1083 (
		\in0[100] ,
		\in1[100] ,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w1155_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h8)
	) name1085 (
		_w1152_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		_w1595_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w1149_,
		_w1160_,
		_w1600_
	);
	LUT2 #(
		.INIT('h4)
	) name1088 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		\in0[104] ,
		\in1[104] ,
		_w1602_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		_w1143_,
		_w1602_,
		_w1603_
	);
	LUT2 #(
		.INIT('h8)
	) name1091 (
		_w1140_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h4)
	) name1092 (
		_w1601_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		_w1137_,
		_w1148_,
		_w1606_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w1605_,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h4)
	) name1095 (
		\in0[108] ,
		\in1[108] ,
		_w1608_
	);
	LUT2 #(
		.INIT('h1)
	) name1096 (
		_w1131_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h8)
	) name1097 (
		_w1128_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		_w1607_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w1125_,
		_w1136_,
		_w1612_
	);
	LUT2 #(
		.INIT('h4)
	) name1100 (
		_w1611_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name1101 (
		\in0[112] ,
		\in1[112] ,
		_w1614_
	);
	LUT2 #(
		.INIT('h1)
	) name1102 (
		_w1119_,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		_w1116_,
		_w1615_,
		_w1616_
	);
	LUT2 #(
		.INIT('h4)
	) name1104 (
		_w1613_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		_w1113_,
		_w1124_,
		_w1618_
	);
	LUT2 #(
		.INIT('h4)
	) name1106 (
		_w1617_,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h4)
	) name1107 (
		\in0[116] ,
		\in1[116] ,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w1107_,
		_w1620_,
		_w1621_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w1104_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		_w1619_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w1101_,
		_w1112_,
		_w1624_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		_w1623_,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		\in0[120] ,
		\in1[120] ,
		_w1626_
	);
	LUT2 #(
		.INIT('h1)
	) name1114 (
		_w1095_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		_w1092_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w1625_,
		_w1628_,
		_w1629_
	);
	LUT2 #(
		.INIT('h1)
	) name1117 (
		_w1089_,
		_w1100_,
		_w1630_
	);
	LUT2 #(
		.INIT('h4)
	) name1118 (
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h4)
	) name1119 (
		\in0[124] ,
		\in1[124] ,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1120 (
		_w1077_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h8)
	) name1121 (
		_w1080_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h4)
	) name1122 (
		_w1631_,
		_w1634_,
		_w1635_
	);
	LUT2 #(
		.INIT('h1)
	) name1123 (
		_w1087_,
		_w1088_,
		_w1636_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		_w1635_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h2)
	) name1125 (
		\in0[123] ,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		\in1[123] ,
		_w1637_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h2)
	) name1128 (
		\in2[123] ,
		_w1073_,
		_w1641_
	);
	LUT2 #(
		.INIT('h8)
	) name1129 (
		\in3[123] ,
		_w1073_,
		_w1642_
	);
	LUT2 #(
		.INIT('h1)
	) name1130 (
		_w1641_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h4)
	) name1131 (
		_w1640_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h2)
	) name1132 (
		_w1640_,
		_w1643_,
		_w1645_
	);
	LUT2 #(
		.INIT('h2)
	) name1133 (
		\in2[122] ,
		_w1073_,
		_w1646_
	);
	LUT2 #(
		.INIT('h8)
	) name1134 (
		\in3[122] ,
		_w1073_,
		_w1647_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w1646_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h2)
	) name1136 (
		\in0[122] ,
		_w1637_,
		_w1649_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		\in1[122] ,
		_w1637_,
		_w1650_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		_w1649_,
		_w1650_,
		_w1651_
	);
	LUT2 #(
		.INIT('h4)
	) name1139 (
		_w1648_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w1645_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h2)
	) name1141 (
		\in0[121] ,
		_w1637_,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		\in1[121] ,
		_w1637_,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w1654_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h2)
	) name1144 (
		\in2[121] ,
		_w1073_,
		_w1657_
	);
	LUT2 #(
		.INIT('h8)
	) name1145 (
		\in3[121] ,
		_w1073_,
		_w1658_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		_w1656_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		_w1648_,
		_w1651_,
		_w1661_
	);
	LUT2 #(
		.INIT('h2)
	) name1149 (
		\in2[120] ,
		_w1073_,
		_w1662_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\in3[120] ,
		_w1073_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h2)
	) name1152 (
		_w1656_,
		_w1659_,
		_w1665_
	);
	LUT2 #(
		.INIT('h2)
	) name1153 (
		\in0[120] ,
		_w1637_,
		_w1666_
	);
	LUT2 #(
		.INIT('h8)
	) name1154 (
		\in1[120] ,
		_w1637_,
		_w1667_
	);
	LUT2 #(
		.INIT('h1)
	) name1155 (
		_w1666_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		_w1664_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		_w1665_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name1158 (
		_w1660_,
		_w1661_,
		_w1671_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w1670_,
		_w1671_,
		_w1672_
	);
	LUT2 #(
		.INIT('h2)
	) name1160 (
		_w1653_,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\in0[119] ,
		_w1637_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name1162 (
		\in1[119] ,
		_w1637_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w1674_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		\in2[119] ,
		_w1073_,
		_w1677_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		\in3[119] ,
		_w1073_,
		_w1678_
	);
	LUT2 #(
		.INIT('h1)
	) name1166 (
		_w1677_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		_w1676_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h2)
	) name1168 (
		_w1676_,
		_w1679_,
		_w1681_
	);
	LUT2 #(
		.INIT('h2)
	) name1169 (
		\in2[118] ,
		_w1073_,
		_w1682_
	);
	LUT2 #(
		.INIT('h8)
	) name1170 (
		\in3[118] ,
		_w1073_,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name1171 (
		_w1682_,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h2)
	) name1172 (
		\in0[118] ,
		_w1637_,
		_w1685_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		\in1[118] ,
		_w1637_,
		_w1686_
	);
	LUT2 #(
		.INIT('h1)
	) name1174 (
		_w1685_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1175 (
		_w1684_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h1)
	) name1176 (
		_w1681_,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h2)
	) name1177 (
		_w1684_,
		_w1687_,
		_w1690_
	);
	LUT2 #(
		.INIT('h2)
	) name1178 (
		\in0[117] ,
		_w1637_,
		_w1691_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		\in1[117] ,
		_w1637_,
		_w1692_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w1691_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h2)
	) name1181 (
		\in2[117] ,
		_w1073_,
		_w1694_
	);
	LUT2 #(
		.INIT('h8)
	) name1182 (
		\in3[117] ,
		_w1073_,
		_w1695_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w1694_,
		_w1695_,
		_w1696_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		_w1693_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h2)
	) name1185 (
		\in2[116] ,
		_w1073_,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name1186 (
		\in3[116] ,
		_w1073_,
		_w1699_
	);
	LUT2 #(
		.INIT('h1)
	) name1187 (
		_w1698_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h2)
	) name1188 (
		_w1693_,
		_w1696_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		\in0[116] ,
		_w1637_,
		_w1702_
	);
	LUT2 #(
		.INIT('h8)
	) name1190 (
		\in1[116] ,
		_w1637_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		_w1700_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h4)
	) name1193 (
		_w1701_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w1690_,
		_w1697_,
		_w1707_
	);
	LUT2 #(
		.INIT('h4)
	) name1195 (
		_w1706_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h2)
	) name1196 (
		_w1689_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h2)
	) name1197 (
		\in0[115] ,
		_w1637_,
		_w1710_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		\in1[115] ,
		_w1637_,
		_w1711_
	);
	LUT2 #(
		.INIT('h1)
	) name1199 (
		_w1710_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h2)
	) name1200 (
		\in2[115] ,
		_w1073_,
		_w1713_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		\in3[115] ,
		_w1073_,
		_w1714_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w1713_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w1712_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h2)
	) name1204 (
		_w1712_,
		_w1715_,
		_w1717_
	);
	LUT2 #(
		.INIT('h2)
	) name1205 (
		\in2[114] ,
		_w1073_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name1206 (
		\in3[114] ,
		_w1073_,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h2)
	) name1208 (
		\in0[114] ,
		_w1637_,
		_w1721_
	);
	LUT2 #(
		.INIT('h8)
	) name1209 (
		\in1[114] ,
		_w1637_,
		_w1722_
	);
	LUT2 #(
		.INIT('h1)
	) name1210 (
		_w1721_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h4)
	) name1211 (
		_w1720_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1717_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		\in0[113] ,
		_w1637_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		\in1[113] ,
		_w1637_,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name1215 (
		_w1726_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h2)
	) name1216 (
		\in2[113] ,
		_w1073_,
		_w1729_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		\in3[113] ,
		_w1073_,
		_w1730_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1729_,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h4)
	) name1219 (
		_w1728_,
		_w1731_,
		_w1732_
	);
	LUT2 #(
		.INIT('h2)
	) name1220 (
		_w1720_,
		_w1723_,
		_w1733_
	);
	LUT2 #(
		.INIT('h2)
	) name1221 (
		\in2[112] ,
		_w1073_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name1222 (
		\in3[112] ,
		_w1073_,
		_w1735_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w1734_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h2)
	) name1224 (
		_w1728_,
		_w1731_,
		_w1737_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		\in0[112] ,
		_w1637_,
		_w1738_
	);
	LUT2 #(
		.INIT('h8)
	) name1226 (
		\in1[112] ,
		_w1637_,
		_w1739_
	);
	LUT2 #(
		.INIT('h1)
	) name1227 (
		_w1738_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h2)
	) name1228 (
		_w1736_,
		_w1740_,
		_w1741_
	);
	LUT2 #(
		.INIT('h4)
	) name1229 (
		_w1737_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w1732_,
		_w1733_,
		_w1743_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		_w1742_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name1232 (
		_w1725_,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name1233 (
		\in0[111] ,
		_w1637_,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		\in1[111] ,
		_w1637_,
		_w1747_
	);
	LUT2 #(
		.INIT('h1)
	) name1235 (
		_w1746_,
		_w1747_,
		_w1748_
	);
	LUT2 #(
		.INIT('h2)
	) name1236 (
		\in2[111] ,
		_w1073_,
		_w1749_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		\in3[111] ,
		_w1073_,
		_w1750_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		_w1749_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w1748_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h2)
	) name1240 (
		_w1748_,
		_w1751_,
		_w1753_
	);
	LUT2 #(
		.INIT('h2)
	) name1241 (
		\in2[110] ,
		_w1073_,
		_w1754_
	);
	LUT2 #(
		.INIT('h8)
	) name1242 (
		\in3[110] ,
		_w1073_,
		_w1755_
	);
	LUT2 #(
		.INIT('h1)
	) name1243 (
		_w1754_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h2)
	) name1244 (
		\in0[110] ,
		_w1637_,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		\in1[110] ,
		_w1637_,
		_w1758_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w1757_,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		_w1756_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1753_,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h2)
	) name1249 (
		_w1756_,
		_w1759_,
		_w1762_
	);
	LUT2 #(
		.INIT('h2)
	) name1250 (
		\in0[109] ,
		_w1637_,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		\in1[109] ,
		_w1637_,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		\in2[109] ,
		_w1073_,
		_w1766_
	);
	LUT2 #(
		.INIT('h8)
	) name1254 (
		\in3[109] ,
		_w1073_,
		_w1767_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w1766_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h4)
	) name1256 (
		_w1765_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		\in2[108] ,
		_w1073_,
		_w1770_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		\in3[108] ,
		_w1073_,
		_w1771_
	);
	LUT2 #(
		.INIT('h1)
	) name1259 (
		_w1770_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h2)
	) name1260 (
		_w1765_,
		_w1768_,
		_w1773_
	);
	LUT2 #(
		.INIT('h2)
	) name1261 (
		\in0[108] ,
		_w1637_,
		_w1774_
	);
	LUT2 #(
		.INIT('h8)
	) name1262 (
		\in1[108] ,
		_w1637_,
		_w1775_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w1774_,
		_w1775_,
		_w1776_
	);
	LUT2 #(
		.INIT('h2)
	) name1264 (
		_w1772_,
		_w1776_,
		_w1777_
	);
	LUT2 #(
		.INIT('h4)
	) name1265 (
		_w1773_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w1762_,
		_w1769_,
		_w1779_
	);
	LUT2 #(
		.INIT('h4)
	) name1267 (
		_w1778_,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('h2)
	) name1268 (
		_w1761_,
		_w1780_,
		_w1781_
	);
	LUT2 #(
		.INIT('h2)
	) name1269 (
		\in0[107] ,
		_w1637_,
		_w1782_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		\in1[107] ,
		_w1637_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w1782_,
		_w1783_,
		_w1784_
	);
	LUT2 #(
		.INIT('h2)
	) name1272 (
		\in2[107] ,
		_w1073_,
		_w1785_
	);
	LUT2 #(
		.INIT('h8)
	) name1273 (
		\in3[107] ,
		_w1073_,
		_w1786_
	);
	LUT2 #(
		.INIT('h1)
	) name1274 (
		_w1785_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('h4)
	) name1275 (
		_w1784_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h2)
	) name1276 (
		_w1784_,
		_w1787_,
		_w1789_
	);
	LUT2 #(
		.INIT('h2)
	) name1277 (
		\in2[106] ,
		_w1073_,
		_w1790_
	);
	LUT2 #(
		.INIT('h8)
	) name1278 (
		\in3[106] ,
		_w1073_,
		_w1791_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w1790_,
		_w1791_,
		_w1792_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		\in0[106] ,
		_w1637_,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name1281 (
		\in1[106] ,
		_w1637_,
		_w1794_
	);
	LUT2 #(
		.INIT('h1)
	) name1282 (
		_w1793_,
		_w1794_,
		_w1795_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w1792_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w1789_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h2)
	) name1285 (
		\in0[105] ,
		_w1637_,
		_w1798_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		\in1[105] ,
		_w1637_,
		_w1799_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w1798_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		\in2[105] ,
		_w1073_,
		_w1801_
	);
	LUT2 #(
		.INIT('h8)
	) name1289 (
		\in3[105] ,
		_w1073_,
		_w1802_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w1801_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		_w1800_,
		_w1803_,
		_w1804_
	);
	LUT2 #(
		.INIT('h2)
	) name1292 (
		_w1792_,
		_w1795_,
		_w1805_
	);
	LUT2 #(
		.INIT('h2)
	) name1293 (
		\in2[104] ,
		_w1073_,
		_w1806_
	);
	LUT2 #(
		.INIT('h8)
	) name1294 (
		\in3[104] ,
		_w1073_,
		_w1807_
	);
	LUT2 #(
		.INIT('h1)
	) name1295 (
		_w1806_,
		_w1807_,
		_w1808_
	);
	LUT2 #(
		.INIT('h2)
	) name1296 (
		_w1800_,
		_w1803_,
		_w1809_
	);
	LUT2 #(
		.INIT('h2)
	) name1297 (
		\in0[104] ,
		_w1637_,
		_w1810_
	);
	LUT2 #(
		.INIT('h8)
	) name1298 (
		\in1[104] ,
		_w1637_,
		_w1811_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		_w1810_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h2)
	) name1300 (
		_w1808_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		_w1809_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w1804_,
		_w1805_,
		_w1815_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		_w1814_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		_w1797_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h2)
	) name1305 (
		\in0[103] ,
		_w1637_,
		_w1818_
	);
	LUT2 #(
		.INIT('h8)
	) name1306 (
		\in1[103] ,
		_w1637_,
		_w1819_
	);
	LUT2 #(
		.INIT('h1)
	) name1307 (
		_w1818_,
		_w1819_,
		_w1820_
	);
	LUT2 #(
		.INIT('h2)
	) name1308 (
		\in2[103] ,
		_w1073_,
		_w1821_
	);
	LUT2 #(
		.INIT('h8)
	) name1309 (
		\in3[103] ,
		_w1073_,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name1310 (
		_w1821_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h4)
	) name1311 (
		_w1820_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h2)
	) name1312 (
		_w1820_,
		_w1823_,
		_w1825_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		\in2[102] ,
		_w1073_,
		_w1826_
	);
	LUT2 #(
		.INIT('h8)
	) name1314 (
		\in3[102] ,
		_w1073_,
		_w1827_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h2)
	) name1316 (
		\in0[102] ,
		_w1637_,
		_w1829_
	);
	LUT2 #(
		.INIT('h8)
	) name1317 (
		\in1[102] ,
		_w1637_,
		_w1830_
	);
	LUT2 #(
		.INIT('h1)
	) name1318 (
		_w1829_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h4)
	) name1319 (
		_w1828_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w1825_,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h2)
	) name1321 (
		_w1828_,
		_w1831_,
		_w1834_
	);
	LUT2 #(
		.INIT('h2)
	) name1322 (
		\in0[101] ,
		_w1637_,
		_w1835_
	);
	LUT2 #(
		.INIT('h8)
	) name1323 (
		\in1[101] ,
		_w1637_,
		_w1836_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w1835_,
		_w1836_,
		_w1837_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		\in2[101] ,
		_w1073_,
		_w1838_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		\in3[101] ,
		_w1073_,
		_w1839_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w1838_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h4)
	) name1328 (
		_w1837_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h2)
	) name1329 (
		\in2[100] ,
		_w1073_,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name1330 (
		\in3[100] ,
		_w1073_,
		_w1843_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w1842_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h2)
	) name1332 (
		_w1837_,
		_w1840_,
		_w1845_
	);
	LUT2 #(
		.INIT('h2)
	) name1333 (
		\in0[100] ,
		_w1637_,
		_w1846_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		\in1[100] ,
		_w1637_,
		_w1847_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w1846_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name1336 (
		_w1844_,
		_w1848_,
		_w1849_
	);
	LUT2 #(
		.INIT('h4)
	) name1337 (
		_w1845_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		_w1834_,
		_w1841_,
		_w1851_
	);
	LUT2 #(
		.INIT('h4)
	) name1339 (
		_w1850_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h2)
	) name1340 (
		_w1833_,
		_w1852_,
		_w1853_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		\in0[99] ,
		_w1637_,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name1342 (
		\in1[99] ,
		_w1637_,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w1854_,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h2)
	) name1344 (
		\in2[99] ,
		_w1073_,
		_w1857_
	);
	LUT2 #(
		.INIT('h8)
	) name1345 (
		\in3[99] ,
		_w1073_,
		_w1858_
	);
	LUT2 #(
		.INIT('h1)
	) name1346 (
		_w1857_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h4)
	) name1347 (
		_w1856_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h2)
	) name1348 (
		_w1856_,
		_w1859_,
		_w1861_
	);
	LUT2 #(
		.INIT('h2)
	) name1349 (
		\in2[98] ,
		_w1073_,
		_w1862_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		\in3[98] ,
		_w1073_,
		_w1863_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		_w1862_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h2)
	) name1352 (
		\in0[98] ,
		_w1637_,
		_w1865_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		\in1[98] ,
		_w1637_,
		_w1866_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		_w1865_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h4)
	) name1355 (
		_w1864_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		_w1861_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h2)
	) name1357 (
		\in0[97] ,
		_w1637_,
		_w1870_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		\in1[97] ,
		_w1637_,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		_w1870_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h2)
	) name1360 (
		\in2[97] ,
		_w1073_,
		_w1873_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		\in3[97] ,
		_w1073_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name1362 (
		_w1873_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h4)
	) name1363 (
		_w1872_,
		_w1875_,
		_w1876_
	);
	LUT2 #(
		.INIT('h2)
	) name1364 (
		_w1864_,
		_w1867_,
		_w1877_
	);
	LUT2 #(
		.INIT('h2)
	) name1365 (
		\in2[96] ,
		_w1073_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		\in3[96] ,
		_w1073_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w1878_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h2)
	) name1368 (
		_w1872_,
		_w1875_,
		_w1881_
	);
	LUT2 #(
		.INIT('h2)
	) name1369 (
		\in0[96] ,
		_w1637_,
		_w1882_
	);
	LUT2 #(
		.INIT('h8)
	) name1370 (
		\in1[96] ,
		_w1637_,
		_w1883_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w1882_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h2)
	) name1372 (
		_w1880_,
		_w1884_,
		_w1885_
	);
	LUT2 #(
		.INIT('h4)
	) name1373 (
		_w1881_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		_w1876_,
		_w1877_,
		_w1887_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		_w1886_,
		_w1887_,
		_w1888_
	);
	LUT2 #(
		.INIT('h2)
	) name1376 (
		_w1869_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h2)
	) name1377 (
		\in0[95] ,
		_w1637_,
		_w1890_
	);
	LUT2 #(
		.INIT('h8)
	) name1378 (
		\in1[95] ,
		_w1637_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w1890_,
		_w1891_,
		_w1892_
	);
	LUT2 #(
		.INIT('h2)
	) name1380 (
		\in2[95] ,
		_w1073_,
		_w1893_
	);
	LUT2 #(
		.INIT('h8)
	) name1381 (
		\in3[95] ,
		_w1073_,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w1893_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h4)
	) name1383 (
		_w1892_,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('h2)
	) name1384 (
		_w1892_,
		_w1895_,
		_w1897_
	);
	LUT2 #(
		.INIT('h2)
	) name1385 (
		\in2[94] ,
		_w1073_,
		_w1898_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		\in3[94] ,
		_w1073_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h2)
	) name1388 (
		\in0[94] ,
		_w1637_,
		_w1901_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		\in1[94] ,
		_w1637_,
		_w1902_
	);
	LUT2 #(
		.INIT('h1)
	) name1390 (
		_w1901_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h4)
	) name1391 (
		_w1900_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h1)
	) name1392 (
		_w1897_,
		_w1904_,
		_w1905_
	);
	LUT2 #(
		.INIT('h2)
	) name1393 (
		_w1900_,
		_w1903_,
		_w1906_
	);
	LUT2 #(
		.INIT('h2)
	) name1394 (
		\in0[93] ,
		_w1637_,
		_w1907_
	);
	LUT2 #(
		.INIT('h8)
	) name1395 (
		\in1[93] ,
		_w1637_,
		_w1908_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		_w1907_,
		_w1908_,
		_w1909_
	);
	LUT2 #(
		.INIT('h2)
	) name1397 (
		\in2[93] ,
		_w1073_,
		_w1910_
	);
	LUT2 #(
		.INIT('h8)
	) name1398 (
		\in3[93] ,
		_w1073_,
		_w1911_
	);
	LUT2 #(
		.INIT('h1)
	) name1399 (
		_w1910_,
		_w1911_,
		_w1912_
	);
	LUT2 #(
		.INIT('h4)
	) name1400 (
		_w1909_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h2)
	) name1401 (
		\in2[92] ,
		_w1073_,
		_w1914_
	);
	LUT2 #(
		.INIT('h8)
	) name1402 (
		\in3[92] ,
		_w1073_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name1403 (
		_w1914_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h2)
	) name1404 (
		_w1909_,
		_w1912_,
		_w1917_
	);
	LUT2 #(
		.INIT('h2)
	) name1405 (
		\in0[92] ,
		_w1637_,
		_w1918_
	);
	LUT2 #(
		.INIT('h8)
	) name1406 (
		\in1[92] ,
		_w1637_,
		_w1919_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		_w1918_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h2)
	) name1408 (
		_w1916_,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h4)
	) name1409 (
		_w1917_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		_w1906_,
		_w1913_,
		_w1923_
	);
	LUT2 #(
		.INIT('h4)
	) name1411 (
		_w1922_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h2)
	) name1412 (
		_w1905_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h2)
	) name1413 (
		\in0[91] ,
		_w1637_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name1414 (
		\in1[91] ,
		_w1637_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w1926_,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('h2)
	) name1416 (
		\in2[91] ,
		_w1073_,
		_w1929_
	);
	LUT2 #(
		.INIT('h8)
	) name1417 (
		\in3[91] ,
		_w1073_,
		_w1930_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		_w1929_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('h4)
	) name1419 (
		_w1928_,
		_w1931_,
		_w1932_
	);
	LUT2 #(
		.INIT('h2)
	) name1420 (
		_w1928_,
		_w1931_,
		_w1933_
	);
	LUT2 #(
		.INIT('h2)
	) name1421 (
		\in2[90] ,
		_w1073_,
		_w1934_
	);
	LUT2 #(
		.INIT('h8)
	) name1422 (
		\in3[90] ,
		_w1073_,
		_w1935_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h2)
	) name1424 (
		\in0[90] ,
		_w1637_,
		_w1937_
	);
	LUT2 #(
		.INIT('h8)
	) name1425 (
		\in1[90] ,
		_w1637_,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		_w1937_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h4)
	) name1427 (
		_w1936_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		_w1933_,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		\in0[89] ,
		_w1637_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name1430 (
		\in1[89] ,
		_w1637_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name1431 (
		_w1942_,
		_w1943_,
		_w1944_
	);
	LUT2 #(
		.INIT('h2)
	) name1432 (
		\in2[89] ,
		_w1073_,
		_w1945_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		\in3[89] ,
		_w1073_,
		_w1946_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w1945_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h4)
	) name1435 (
		_w1944_,
		_w1947_,
		_w1948_
	);
	LUT2 #(
		.INIT('h2)
	) name1436 (
		_w1936_,
		_w1939_,
		_w1949_
	);
	LUT2 #(
		.INIT('h2)
	) name1437 (
		\in2[88] ,
		_w1073_,
		_w1950_
	);
	LUT2 #(
		.INIT('h8)
	) name1438 (
		\in3[88] ,
		_w1073_,
		_w1951_
	);
	LUT2 #(
		.INIT('h1)
	) name1439 (
		_w1950_,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h2)
	) name1440 (
		_w1944_,
		_w1947_,
		_w1953_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		\in0[88] ,
		_w1637_,
		_w1954_
	);
	LUT2 #(
		.INIT('h8)
	) name1442 (
		\in1[88] ,
		_w1637_,
		_w1955_
	);
	LUT2 #(
		.INIT('h1)
	) name1443 (
		_w1954_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h2)
	) name1444 (
		_w1952_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h4)
	) name1445 (
		_w1953_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h1)
	) name1446 (
		_w1948_,
		_w1949_,
		_w1959_
	);
	LUT2 #(
		.INIT('h4)
	) name1447 (
		_w1958_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h2)
	) name1448 (
		_w1941_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		\in0[87] ,
		_w1637_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name1450 (
		\in1[87] ,
		_w1637_,
		_w1963_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w1962_,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h2)
	) name1452 (
		\in2[87] ,
		_w1073_,
		_w1965_
	);
	LUT2 #(
		.INIT('h8)
	) name1453 (
		\in3[87] ,
		_w1073_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		_w1964_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		_w1964_,
		_w1967_,
		_w1969_
	);
	LUT2 #(
		.INIT('h2)
	) name1457 (
		\in2[86] ,
		_w1073_,
		_w1970_
	);
	LUT2 #(
		.INIT('h8)
	) name1458 (
		\in3[86] ,
		_w1073_,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		_w1970_,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h2)
	) name1460 (
		\in0[86] ,
		_w1637_,
		_w1973_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		\in1[86] ,
		_w1637_,
		_w1974_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h4)
	) name1463 (
		_w1972_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h1)
	) name1464 (
		_w1969_,
		_w1976_,
		_w1977_
	);
	LUT2 #(
		.INIT('h2)
	) name1465 (
		_w1972_,
		_w1975_,
		_w1978_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		\in0[85] ,
		_w1637_,
		_w1979_
	);
	LUT2 #(
		.INIT('h8)
	) name1467 (
		\in1[85] ,
		_w1637_,
		_w1980_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		_w1979_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h2)
	) name1469 (
		\in2[85] ,
		_w1073_,
		_w1982_
	);
	LUT2 #(
		.INIT('h8)
	) name1470 (
		\in3[85] ,
		_w1073_,
		_w1983_
	);
	LUT2 #(
		.INIT('h1)
	) name1471 (
		_w1982_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h4)
	) name1472 (
		_w1981_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h2)
	) name1473 (
		\in2[84] ,
		_w1073_,
		_w1986_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		\in3[84] ,
		_w1073_,
		_w1987_
	);
	LUT2 #(
		.INIT('h1)
	) name1475 (
		_w1986_,
		_w1987_,
		_w1988_
	);
	LUT2 #(
		.INIT('h2)
	) name1476 (
		_w1981_,
		_w1984_,
		_w1989_
	);
	LUT2 #(
		.INIT('h2)
	) name1477 (
		\in0[84] ,
		_w1637_,
		_w1990_
	);
	LUT2 #(
		.INIT('h8)
	) name1478 (
		\in1[84] ,
		_w1637_,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name1479 (
		_w1990_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h2)
	) name1480 (
		_w1988_,
		_w1992_,
		_w1993_
	);
	LUT2 #(
		.INIT('h4)
	) name1481 (
		_w1989_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1482 (
		_w1978_,
		_w1985_,
		_w1995_
	);
	LUT2 #(
		.INIT('h4)
	) name1483 (
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h2)
	) name1484 (
		_w1977_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h2)
	) name1485 (
		\in0[83] ,
		_w1637_,
		_w1998_
	);
	LUT2 #(
		.INIT('h8)
	) name1486 (
		\in1[83] ,
		_w1637_,
		_w1999_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		_w1998_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h2)
	) name1488 (
		\in2[83] ,
		_w1073_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name1489 (
		\in3[83] ,
		_w1073_,
		_w2002_
	);
	LUT2 #(
		.INIT('h1)
	) name1490 (
		_w2001_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('h4)
	) name1491 (
		_w2000_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h2)
	) name1492 (
		_w2000_,
		_w2003_,
		_w2005_
	);
	LUT2 #(
		.INIT('h2)
	) name1493 (
		\in2[82] ,
		_w1073_,
		_w2006_
	);
	LUT2 #(
		.INIT('h8)
	) name1494 (
		\in3[82] ,
		_w1073_,
		_w2007_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h2)
	) name1496 (
		\in0[82] ,
		_w1637_,
		_w2009_
	);
	LUT2 #(
		.INIT('h8)
	) name1497 (
		\in1[82] ,
		_w1637_,
		_w2010_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		_w2009_,
		_w2010_,
		_w2011_
	);
	LUT2 #(
		.INIT('h4)
	) name1499 (
		_w2008_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		_w2005_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h2)
	) name1501 (
		\in0[81] ,
		_w1637_,
		_w2014_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		\in1[81] ,
		_w1637_,
		_w2015_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w2014_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name1504 (
		\in2[81] ,
		_w1073_,
		_w2017_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		\in3[81] ,
		_w1073_,
		_w2018_
	);
	LUT2 #(
		.INIT('h1)
	) name1506 (
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h4)
	) name1507 (
		_w2016_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h2)
	) name1508 (
		_w2008_,
		_w2011_,
		_w2021_
	);
	LUT2 #(
		.INIT('h2)
	) name1509 (
		\in2[80] ,
		_w1073_,
		_w2022_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		\in3[80] ,
		_w1073_,
		_w2023_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		_w2022_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h2)
	) name1512 (
		_w2016_,
		_w2019_,
		_w2025_
	);
	LUT2 #(
		.INIT('h2)
	) name1513 (
		\in0[80] ,
		_w1637_,
		_w2026_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		\in1[80] ,
		_w1637_,
		_w2027_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		_w2026_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h2)
	) name1516 (
		_w2024_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h4)
	) name1517 (
		_w2025_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h1)
	) name1518 (
		_w2020_,
		_w2021_,
		_w2031_
	);
	LUT2 #(
		.INIT('h4)
	) name1519 (
		_w2030_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h2)
	) name1520 (
		_w2013_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h2)
	) name1521 (
		\in0[79] ,
		_w1637_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name1522 (
		\in1[79] ,
		_w1637_,
		_w2035_
	);
	LUT2 #(
		.INIT('h1)
	) name1523 (
		_w2034_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('h2)
	) name1524 (
		\in2[79] ,
		_w1073_,
		_w2037_
	);
	LUT2 #(
		.INIT('h8)
	) name1525 (
		\in3[79] ,
		_w1073_,
		_w2038_
	);
	LUT2 #(
		.INIT('h1)
	) name1526 (
		_w2037_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h4)
	) name1527 (
		_w2036_,
		_w2039_,
		_w2040_
	);
	LUT2 #(
		.INIT('h2)
	) name1528 (
		_w2036_,
		_w2039_,
		_w2041_
	);
	LUT2 #(
		.INIT('h2)
	) name1529 (
		\in2[78] ,
		_w1073_,
		_w2042_
	);
	LUT2 #(
		.INIT('h8)
	) name1530 (
		\in3[78] ,
		_w1073_,
		_w2043_
	);
	LUT2 #(
		.INIT('h1)
	) name1531 (
		_w2042_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h2)
	) name1532 (
		\in0[78] ,
		_w1637_,
		_w2045_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		\in1[78] ,
		_w1637_,
		_w2046_
	);
	LUT2 #(
		.INIT('h1)
	) name1534 (
		_w2045_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h4)
	) name1535 (
		_w2044_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h1)
	) name1536 (
		_w2041_,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h2)
	) name1537 (
		_w2044_,
		_w2047_,
		_w2050_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		\in0[77] ,
		_w1637_,
		_w2051_
	);
	LUT2 #(
		.INIT('h8)
	) name1539 (
		\in1[77] ,
		_w1637_,
		_w2052_
	);
	LUT2 #(
		.INIT('h1)
	) name1540 (
		_w2051_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h2)
	) name1541 (
		\in2[77] ,
		_w1073_,
		_w2054_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		\in3[77] ,
		_w1073_,
		_w2055_
	);
	LUT2 #(
		.INIT('h1)
	) name1543 (
		_w2054_,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h4)
	) name1544 (
		_w2053_,
		_w2056_,
		_w2057_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		\in2[76] ,
		_w1073_,
		_w2058_
	);
	LUT2 #(
		.INIT('h8)
	) name1546 (
		\in3[76] ,
		_w1073_,
		_w2059_
	);
	LUT2 #(
		.INIT('h1)
	) name1547 (
		_w2058_,
		_w2059_,
		_w2060_
	);
	LUT2 #(
		.INIT('h2)
	) name1548 (
		_w2053_,
		_w2056_,
		_w2061_
	);
	LUT2 #(
		.INIT('h2)
	) name1549 (
		\in0[76] ,
		_w1637_,
		_w2062_
	);
	LUT2 #(
		.INIT('h8)
	) name1550 (
		\in1[76] ,
		_w1637_,
		_w2063_
	);
	LUT2 #(
		.INIT('h1)
	) name1551 (
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h2)
	) name1552 (
		_w2060_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h4)
	) name1553 (
		_w2061_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w2050_,
		_w2057_,
		_w2067_
	);
	LUT2 #(
		.INIT('h4)
	) name1555 (
		_w2066_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h2)
	) name1556 (
		_w2049_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h2)
	) name1557 (
		\in0[75] ,
		_w1637_,
		_w2070_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		\in1[75] ,
		_w1637_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name1559 (
		_w2070_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name1560 (
		\in2[75] ,
		_w1073_,
		_w2073_
	);
	LUT2 #(
		.INIT('h8)
	) name1561 (
		\in3[75] ,
		_w1073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name1562 (
		_w2073_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h4)
	) name1563 (
		_w2072_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h2)
	) name1564 (
		_w2072_,
		_w2075_,
		_w2077_
	);
	LUT2 #(
		.INIT('h2)
	) name1565 (
		\in2[74] ,
		_w1073_,
		_w2078_
	);
	LUT2 #(
		.INIT('h8)
	) name1566 (
		\in3[74] ,
		_w1073_,
		_w2079_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		_w2078_,
		_w2079_,
		_w2080_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		\in0[74] ,
		_w1637_,
		_w2081_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		\in1[74] ,
		_w1637_,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w2081_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h4)
	) name1571 (
		_w2080_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w2077_,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h2)
	) name1573 (
		\in0[73] ,
		_w1637_,
		_w2086_
	);
	LUT2 #(
		.INIT('h8)
	) name1574 (
		\in1[73] ,
		_w1637_,
		_w2087_
	);
	LUT2 #(
		.INIT('h1)
	) name1575 (
		_w2086_,
		_w2087_,
		_w2088_
	);
	LUT2 #(
		.INIT('h2)
	) name1576 (
		\in2[73] ,
		_w1073_,
		_w2089_
	);
	LUT2 #(
		.INIT('h8)
	) name1577 (
		\in3[73] ,
		_w1073_,
		_w2090_
	);
	LUT2 #(
		.INIT('h1)
	) name1578 (
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h4)
	) name1579 (
		_w2088_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		_w2080_,
		_w2083_,
		_w2093_
	);
	LUT2 #(
		.INIT('h2)
	) name1581 (
		\in2[72] ,
		_w1073_,
		_w2094_
	);
	LUT2 #(
		.INIT('h8)
	) name1582 (
		\in3[72] ,
		_w1073_,
		_w2095_
	);
	LUT2 #(
		.INIT('h1)
	) name1583 (
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h2)
	) name1584 (
		_w2088_,
		_w2091_,
		_w2097_
	);
	LUT2 #(
		.INIT('h2)
	) name1585 (
		\in0[72] ,
		_w1637_,
		_w2098_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		\in1[72] ,
		_w1637_,
		_w2099_
	);
	LUT2 #(
		.INIT('h1)
	) name1587 (
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h2)
	) name1588 (
		_w2096_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h4)
	) name1589 (
		_w2097_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w2092_,
		_w2093_,
		_w2103_
	);
	LUT2 #(
		.INIT('h4)
	) name1591 (
		_w2102_,
		_w2103_,
		_w2104_
	);
	LUT2 #(
		.INIT('h2)
	) name1592 (
		_w2085_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h2)
	) name1593 (
		\in0[71] ,
		_w1637_,
		_w2106_
	);
	LUT2 #(
		.INIT('h8)
	) name1594 (
		\in1[71] ,
		_w1637_,
		_w2107_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h2)
	) name1596 (
		\in2[71] ,
		_w1073_,
		_w2109_
	);
	LUT2 #(
		.INIT('h8)
	) name1597 (
		\in3[71] ,
		_w1073_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h4)
	) name1599 (
		_w2108_,
		_w2111_,
		_w2112_
	);
	LUT2 #(
		.INIT('h2)
	) name1600 (
		_w2108_,
		_w2111_,
		_w2113_
	);
	LUT2 #(
		.INIT('h2)
	) name1601 (
		\in2[70] ,
		_w1073_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name1602 (
		\in3[70] ,
		_w1073_,
		_w2115_
	);
	LUT2 #(
		.INIT('h1)
	) name1603 (
		_w2114_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h2)
	) name1604 (
		\in0[70] ,
		_w1637_,
		_w2117_
	);
	LUT2 #(
		.INIT('h8)
	) name1605 (
		\in1[70] ,
		_w1637_,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name1606 (
		_w2117_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('h4)
	) name1607 (
		_w2116_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w2113_,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h2)
	) name1609 (
		_w2116_,
		_w2119_,
		_w2122_
	);
	LUT2 #(
		.INIT('h2)
	) name1610 (
		\in0[69] ,
		_w1637_,
		_w2123_
	);
	LUT2 #(
		.INIT('h8)
	) name1611 (
		\in1[69] ,
		_w1637_,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name1612 (
		_w2123_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('h2)
	) name1613 (
		\in2[69] ,
		_w1073_,
		_w2126_
	);
	LUT2 #(
		.INIT('h8)
	) name1614 (
		\in3[69] ,
		_w1073_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name1615 (
		_w2126_,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		_w2125_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		\in2[68] ,
		_w1073_,
		_w2130_
	);
	LUT2 #(
		.INIT('h8)
	) name1618 (
		\in3[68] ,
		_w1073_,
		_w2131_
	);
	LUT2 #(
		.INIT('h1)
	) name1619 (
		_w2130_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h2)
	) name1620 (
		_w2125_,
		_w2128_,
		_w2133_
	);
	LUT2 #(
		.INIT('h2)
	) name1621 (
		\in0[68] ,
		_w1637_,
		_w2134_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		\in1[68] ,
		_w1637_,
		_w2135_
	);
	LUT2 #(
		.INIT('h1)
	) name1623 (
		_w2134_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h2)
	) name1624 (
		_w2132_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h4)
	) name1625 (
		_w2133_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		_w2122_,
		_w2129_,
		_w2139_
	);
	LUT2 #(
		.INIT('h4)
	) name1627 (
		_w2138_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h2)
	) name1628 (
		_w2121_,
		_w2140_,
		_w2141_
	);
	LUT2 #(
		.INIT('h2)
	) name1629 (
		\in0[67] ,
		_w1637_,
		_w2142_
	);
	LUT2 #(
		.INIT('h8)
	) name1630 (
		\in1[67] ,
		_w1637_,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w2142_,
		_w2143_,
		_w2144_
	);
	LUT2 #(
		.INIT('h2)
	) name1632 (
		\in2[67] ,
		_w1073_,
		_w2145_
	);
	LUT2 #(
		.INIT('h8)
	) name1633 (
		\in3[67] ,
		_w1073_,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name1634 (
		_w2145_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('h4)
	) name1635 (
		_w2144_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h2)
	) name1636 (
		_w2144_,
		_w2147_,
		_w2149_
	);
	LUT2 #(
		.INIT('h2)
	) name1637 (
		\in2[66] ,
		_w1073_,
		_w2150_
	);
	LUT2 #(
		.INIT('h8)
	) name1638 (
		\in3[66] ,
		_w1073_,
		_w2151_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w2150_,
		_w2151_,
		_w2152_
	);
	LUT2 #(
		.INIT('h2)
	) name1640 (
		\in0[66] ,
		_w1637_,
		_w2153_
	);
	LUT2 #(
		.INIT('h8)
	) name1641 (
		\in1[66] ,
		_w1637_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w2153_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h4)
	) name1643 (
		_w2152_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w2149_,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h2)
	) name1645 (
		\in0[65] ,
		_w1637_,
		_w2158_
	);
	LUT2 #(
		.INIT('h8)
	) name1646 (
		\in1[65] ,
		_w1637_,
		_w2159_
	);
	LUT2 #(
		.INIT('h1)
	) name1647 (
		_w2158_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h2)
	) name1648 (
		\in2[65] ,
		_w1073_,
		_w2161_
	);
	LUT2 #(
		.INIT('h8)
	) name1649 (
		\in3[65] ,
		_w1073_,
		_w2162_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		_w2161_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h4)
	) name1651 (
		_w2160_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h2)
	) name1652 (
		_w2152_,
		_w2155_,
		_w2165_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		\in2[64] ,
		_w1073_,
		_w2166_
	);
	LUT2 #(
		.INIT('h8)
	) name1654 (
		\in3[64] ,
		_w1073_,
		_w2167_
	);
	LUT2 #(
		.INIT('h1)
	) name1655 (
		_w2166_,
		_w2167_,
		_w2168_
	);
	LUT2 #(
		.INIT('h2)
	) name1656 (
		_w2160_,
		_w2163_,
		_w2169_
	);
	LUT2 #(
		.INIT('h2)
	) name1657 (
		\in0[64] ,
		_w1637_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name1658 (
		\in1[64] ,
		_w1637_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name1659 (
		_w2170_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		_w2168_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name1661 (
		_w2169_,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		_w2164_,
		_w2165_,
		_w2175_
	);
	LUT2 #(
		.INIT('h4)
	) name1663 (
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name1664 (
		_w2157_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h2)
	) name1665 (
		\in0[27] ,
		_w1637_,
		_w2178_
	);
	LUT2 #(
		.INIT('h8)
	) name1666 (
		\in1[27] ,
		_w1637_,
		_w2179_
	);
	LUT2 #(
		.INIT('h1)
	) name1667 (
		_w2178_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('h2)
	) name1668 (
		\in2[27] ,
		_w1073_,
		_w2181_
	);
	LUT2 #(
		.INIT('h8)
	) name1669 (
		\in3[27] ,
		_w1073_,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		_w2181_,
		_w2182_,
		_w2183_
	);
	LUT2 #(
		.INIT('h4)
	) name1671 (
		_w2180_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h2)
	) name1672 (
		\in0[12] ,
		_w1637_,
		_w2185_
	);
	LUT2 #(
		.INIT('h8)
	) name1673 (
		\in1[12] ,
		_w1637_,
		_w2186_
	);
	LUT2 #(
		.INIT('h1)
	) name1674 (
		_w2185_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h2)
	) name1675 (
		\in2[12] ,
		_w1073_,
		_w2188_
	);
	LUT2 #(
		.INIT('h8)
	) name1676 (
		\in3[12] ,
		_w1073_,
		_w2189_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w2188_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h4)
	) name1678 (
		_w2187_,
		_w2190_,
		_w2191_
	);
	LUT2 #(
		.INIT('h2)
	) name1679 (
		\in2[6] ,
		_w1073_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name1680 (
		\in3[6] ,
		_w1073_,
		_w2193_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w2192_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h2)
	) name1682 (
		\in0[6] ,
		_w1637_,
		_w2195_
	);
	LUT2 #(
		.INIT('h8)
	) name1683 (
		\in1[6] ,
		_w1637_,
		_w2196_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w2195_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h4)
	) name1685 (
		_w2194_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h2)
	) name1686 (
		\in2[1] ,
		_w1073_,
		_w2199_
	);
	LUT2 #(
		.INIT('h8)
	) name1687 (
		\in3[1] ,
		_w1073_,
		_w2200_
	);
	LUT2 #(
		.INIT('h1)
	) name1688 (
		_w2199_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h2)
	) name1689 (
		\in0[1] ,
		_w1637_,
		_w2202_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		\in1[1] ,
		_w1637_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w2202_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h4)
	) name1692 (
		_w2201_,
		_w2204_,
		_w2205_
	);
	LUT2 #(
		.INIT('h2)
	) name1693 (
		\in0[0] ,
		_w1637_,
		_w2206_
	);
	LUT2 #(
		.INIT('h8)
	) name1694 (
		\in1[0] ,
		_w1637_,
		_w2207_
	);
	LUT2 #(
		.INIT('h1)
	) name1695 (
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h2)
	) name1696 (
		_w1076_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h4)
	) name1697 (
		_w2205_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h2)
	) name1698 (
		\in0[2] ,
		_w1637_,
		_w2211_
	);
	LUT2 #(
		.INIT('h8)
	) name1699 (
		\in1[2] ,
		_w1637_,
		_w2212_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w2211_,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h2)
	) name1701 (
		\in2[2] ,
		_w1073_,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name1702 (
		\in3[2] ,
		_w1073_,
		_w2215_
	);
	LUT2 #(
		.INIT('h1)
	) name1703 (
		_w2214_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h4)
	) name1704 (
		_w2213_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w2201_,
		_w2204_,
		_w2218_
	);
	LUT2 #(
		.INIT('h1)
	) name1706 (
		_w2217_,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h4)
	) name1707 (
		_w2210_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h2)
	) name1708 (
		\in0[3] ,
		_w1637_,
		_w2221_
	);
	LUT2 #(
		.INIT('h8)
	) name1709 (
		\in1[3] ,
		_w1637_,
		_w2222_
	);
	LUT2 #(
		.INIT('h1)
	) name1710 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h2)
	) name1711 (
		\in2[3] ,
		_w1073_,
		_w2224_
	);
	LUT2 #(
		.INIT('h8)
	) name1712 (
		\in3[3] ,
		_w1073_,
		_w2225_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h2)
	) name1714 (
		_w2223_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h2)
	) name1715 (
		_w2213_,
		_w2216_,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w2227_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w2220_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h4)
	) name1718 (
		_w2223_,
		_w2226_,
		_w2231_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		\in0[4] ,
		_w1637_,
		_w2232_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\in1[4] ,
		_w1637_,
		_w2233_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		_w2232_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h2)
	) name1722 (
		\in2[4] ,
		_w1073_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name1723 (
		\in3[4] ,
		_w1073_,
		_w2236_
	);
	LUT2 #(
		.INIT('h1)
	) name1724 (
		_w2235_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h4)
	) name1725 (
		_w2234_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w2231_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h4)
	) name1727 (
		_w2230_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		_w2234_,
		_w2237_,
		_w2241_
	);
	LUT2 #(
		.INIT('h2)
	) name1729 (
		\in2[5] ,
		_w1073_,
		_w2242_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		\in3[5] ,
		_w1073_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name1731 (
		_w2242_,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h2)
	) name1732 (
		\in0[5] ,
		_w1637_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name1733 (
		\in1[5] ,
		_w1637_,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h4)
	) name1735 (
		_w2244_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w2241_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h4)
	) name1737 (
		_w2240_,
		_w2249_,
		_w2250_
	);
	LUT2 #(
		.INIT('h2)
	) name1738 (
		_w2244_,
		_w2247_,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name1739 (
		_w2250_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w2198_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h2)
	) name1741 (
		_w2194_,
		_w2197_,
		_w2254_
	);
	LUT2 #(
		.INIT('h2)
	) name1742 (
		\in0[7] ,
		_w1637_,
		_w2255_
	);
	LUT2 #(
		.INIT('h8)
	) name1743 (
		\in1[7] ,
		_w1637_,
		_w2256_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w2255_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h2)
	) name1745 (
		\in2[7] ,
		_w1073_,
		_w2258_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		\in3[7] ,
		_w1073_,
		_w2259_
	);
	LUT2 #(
		.INIT('h1)
	) name1747 (
		_w2258_,
		_w2259_,
		_w2260_
	);
	LUT2 #(
		.INIT('h4)
	) name1748 (
		_w2257_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w2254_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h4)
	) name1750 (
		_w2253_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h2)
	) name1751 (
		_w2257_,
		_w2260_,
		_w2264_
	);
	LUT2 #(
		.INIT('h2)
	) name1752 (
		\in0[8] ,
		_w1637_,
		_w2265_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		\in1[8] ,
		_w1637_,
		_w2266_
	);
	LUT2 #(
		.INIT('h1)
	) name1754 (
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h2)
	) name1755 (
		\in2[8] ,
		_w1073_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		\in3[8] ,
		_w1073_,
		_w2269_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w2268_,
		_w2269_,
		_w2270_
	);
	LUT2 #(
		.INIT('h2)
	) name1758 (
		_w2267_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w2264_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h4)
	) name1760 (
		_w2263_,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h4)
	) name1761 (
		_w2267_,
		_w2270_,
		_w2274_
	);
	LUT2 #(
		.INIT('h2)
	) name1762 (
		\in0[9] ,
		_w1637_,
		_w2275_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		\in1[9] ,
		_w1637_,
		_w2276_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('h2)
	) name1765 (
		\in2[9] ,
		_w1073_,
		_w2278_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		\in3[9] ,
		_w1073_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name1767 (
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT2 #(
		.INIT('h4)
	) name1768 (
		_w2277_,
		_w2280_,
		_w2281_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w2274_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h4)
	) name1770 (
		_w2273_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		\in0[10] ,
		_w1637_,
		_w2284_
	);
	LUT2 #(
		.INIT('h8)
	) name1772 (
		\in1[10] ,
		_w1637_,
		_w2285_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w2284_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h2)
	) name1774 (
		\in2[10] ,
		_w1073_,
		_w2287_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		\in3[10] ,
		_w1073_,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name1776 (
		_w2287_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h2)
	) name1777 (
		_w2286_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h2)
	) name1778 (
		_w2277_,
		_w2280_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1779 (
		_w2290_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h4)
	) name1780 (
		_w2283_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h4)
	) name1781 (
		_w2286_,
		_w2289_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name1782 (
		\in0[11] ,
		_w1637_,
		_w2295_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		\in1[11] ,
		_w1637_,
		_w2296_
	);
	LUT2 #(
		.INIT('h1)
	) name1784 (
		_w2295_,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h2)
	) name1785 (
		\in2[11] ,
		_w1073_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		\in3[11] ,
		_w1073_,
		_w2299_
	);
	LUT2 #(
		.INIT('h1)
	) name1787 (
		_w2298_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('h4)
	) name1788 (
		_w2297_,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1789 (
		_w2294_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h4)
	) name1790 (
		_w2293_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h2)
	) name1791 (
		_w2297_,
		_w2300_,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w2303_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w2191_,
		_w2305_,
		_w2306_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		_w2187_,
		_w2190_,
		_w2307_
	);
	LUT2 #(
		.INIT('h2)
	) name1795 (
		\in0[13] ,
		_w1637_,
		_w2308_
	);
	LUT2 #(
		.INIT('h8)
	) name1796 (
		\in1[13] ,
		_w1637_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		\in2[13] ,
		_w1073_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name1799 (
		\in3[13] ,
		_w1073_,
		_w2312_
	);
	LUT2 #(
		.INIT('h1)
	) name1800 (
		_w2311_,
		_w2312_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name1801 (
		_w2310_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		_w2307_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h4)
	) name1803 (
		_w2306_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h4)
	) name1804 (
		_w2310_,
		_w2313_,
		_w2317_
	);
	LUT2 #(
		.INIT('h2)
	) name1805 (
		\in0[14] ,
		_w1637_,
		_w2318_
	);
	LUT2 #(
		.INIT('h8)
	) name1806 (
		\in1[14] ,
		_w1637_,
		_w2319_
	);
	LUT2 #(
		.INIT('h1)
	) name1807 (
		_w2318_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name1808 (
		\in2[14] ,
		_w1073_,
		_w2321_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		\in3[14] ,
		_w1073_,
		_w2322_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w2321_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w2320_,
		_w2323_,
		_w2324_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w2317_,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h4)
	) name1813 (
		_w2316_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h2)
	) name1814 (
		_w2320_,
		_w2323_,
		_w2327_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		\in0[15] ,
		_w1637_,
		_w2328_
	);
	LUT2 #(
		.INIT('h8)
	) name1816 (
		\in1[15] ,
		_w1637_,
		_w2329_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w2328_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h2)
	) name1818 (
		\in2[15] ,
		_w1073_,
		_w2331_
	);
	LUT2 #(
		.INIT('h8)
	) name1819 (
		\in3[15] ,
		_w1073_,
		_w2332_
	);
	LUT2 #(
		.INIT('h1)
	) name1820 (
		_w2331_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h2)
	) name1821 (
		_w2330_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name1822 (
		_w2327_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h4)
	) name1823 (
		_w2326_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h4)
	) name1824 (
		_w2330_,
		_w2333_,
		_w2337_
	);
	LUT2 #(
		.INIT('h2)
	) name1825 (
		\in0[16] ,
		_w1637_,
		_w2338_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		\in1[16] ,
		_w1637_,
		_w2339_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w2338_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h2)
	) name1828 (
		\in2[16] ,
		_w1073_,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name1829 (
		\in3[16] ,
		_w1073_,
		_w2342_
	);
	LUT2 #(
		.INIT('h1)
	) name1830 (
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT2 #(
		.INIT('h4)
	) name1831 (
		_w2340_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h1)
	) name1832 (
		_w2337_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		_w2336_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h2)
	) name1834 (
		_w2340_,
		_w2343_,
		_w2347_
	);
	LUT2 #(
		.INIT('h2)
	) name1835 (
		\in0[17] ,
		_w1637_,
		_w2348_
	);
	LUT2 #(
		.INIT('h8)
	) name1836 (
		\in1[17] ,
		_w1637_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name1837 (
		_w2348_,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('h2)
	) name1838 (
		\in2[17] ,
		_w1073_,
		_w2351_
	);
	LUT2 #(
		.INIT('h8)
	) name1839 (
		\in3[17] ,
		_w1073_,
		_w2352_
	);
	LUT2 #(
		.INIT('h1)
	) name1840 (
		_w2351_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w2350_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h1)
	) name1842 (
		_w2347_,
		_w2354_,
		_w2355_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w2346_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h4)
	) name1844 (
		_w2350_,
		_w2353_,
		_w2357_
	);
	LUT2 #(
		.INIT('h2)
	) name1845 (
		\in0[18] ,
		_w1637_,
		_w2358_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		\in1[18] ,
		_w1637_,
		_w2359_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w2358_,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h2)
	) name1848 (
		\in2[18] ,
		_w1073_,
		_w2361_
	);
	LUT2 #(
		.INIT('h8)
	) name1849 (
		\in3[18] ,
		_w1073_,
		_w2362_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w2361_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h4)
	) name1851 (
		_w2360_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w2357_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name1853 (
		_w2356_,
		_w2365_,
		_w2366_
	);
	LUT2 #(
		.INIT('h2)
	) name1854 (
		_w2360_,
		_w2363_,
		_w2367_
	);
	LUT2 #(
		.INIT('h2)
	) name1855 (
		\in2[19] ,
		_w1073_,
		_w2368_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		\in3[19] ,
		_w1073_,
		_w2369_
	);
	LUT2 #(
		.INIT('h1)
	) name1857 (
		_w2368_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h2)
	) name1858 (
		\in0[19] ,
		_w1637_,
		_w2371_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		\in1[19] ,
		_w1637_,
		_w2372_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w2371_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		_w2370_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w2367_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h4)
	) name1863 (
		_w2366_,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('h2)
	) name1864 (
		\in0[20] ,
		_w1637_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name1865 (
		\in1[20] ,
		_w1637_,
		_w2378_
	);
	LUT2 #(
		.INIT('h1)
	) name1866 (
		_w2377_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h2)
	) name1867 (
		\in2[20] ,
		_w1073_,
		_w2380_
	);
	LUT2 #(
		.INIT('h8)
	) name1868 (
		\in3[20] ,
		_w1073_,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w2380_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h4)
	) name1870 (
		_w2379_,
		_w2382_,
		_w2383_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		_w2370_,
		_w2373_,
		_w2384_
	);
	LUT2 #(
		.INIT('h1)
	) name1872 (
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h4)
	) name1873 (
		_w2376_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h2)
	) name1874 (
		\in0[21] ,
		_w1637_,
		_w2387_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		\in1[21] ,
		_w1637_,
		_w2388_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		_w2387_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name1877 (
		\in2[21] ,
		_w1073_,
		_w2390_
	);
	LUT2 #(
		.INIT('h8)
	) name1878 (
		\in3[21] ,
		_w1073_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name1879 (
		_w2390_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h2)
	) name1880 (
		_w2389_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		_w2379_,
		_w2382_,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		_w2393_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h4)
	) name1883 (
		_w2386_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h4)
	) name1884 (
		_w2389_,
		_w2392_,
		_w2397_
	);
	LUT2 #(
		.INIT('h2)
	) name1885 (
		\in0[22] ,
		_w1637_,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name1886 (
		\in1[22] ,
		_w1637_,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name1887 (
		_w2398_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name1888 (
		\in2[22] ,
		_w1073_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name1889 (
		\in3[22] ,
		_w1073_,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2401_,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h4)
	) name1891 (
		_w2400_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h1)
	) name1892 (
		_w2397_,
		_w2404_,
		_w2405_
	);
	LUT2 #(
		.INIT('h4)
	) name1893 (
		_w2396_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h2)
	) name1894 (
		_w2400_,
		_w2403_,
		_w2407_
	);
	LUT2 #(
		.INIT('h2)
	) name1895 (
		\in0[23] ,
		_w1637_,
		_w2408_
	);
	LUT2 #(
		.INIT('h8)
	) name1896 (
		\in1[23] ,
		_w1637_,
		_w2409_
	);
	LUT2 #(
		.INIT('h1)
	) name1897 (
		_w2408_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h2)
	) name1898 (
		\in2[23] ,
		_w1073_,
		_w2411_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		\in3[23] ,
		_w1073_,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name1900 (
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		_w2410_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name1902 (
		_w2407_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name1903 (
		_w2406_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h4)
	) name1904 (
		_w2410_,
		_w2413_,
		_w2417_
	);
	LUT2 #(
		.INIT('h2)
	) name1905 (
		\in0[24] ,
		_w1637_,
		_w2418_
	);
	LUT2 #(
		.INIT('h8)
	) name1906 (
		\in1[24] ,
		_w1637_,
		_w2419_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		_w2418_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h2)
	) name1908 (
		\in2[24] ,
		_w1073_,
		_w2421_
	);
	LUT2 #(
		.INIT('h8)
	) name1909 (
		\in3[24] ,
		_w1073_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name1910 (
		_w2421_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h4)
	) name1911 (
		_w2420_,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h1)
	) name1912 (
		_w2417_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h4)
	) name1913 (
		_w2416_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h2)
	) name1914 (
		_w2420_,
		_w2423_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name1915 (
		\in0[25] ,
		_w1637_,
		_w2428_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		\in1[25] ,
		_w1637_,
		_w2429_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h2)
	) name1918 (
		\in2[25] ,
		_w1073_,
		_w2431_
	);
	LUT2 #(
		.INIT('h8)
	) name1919 (
		\in3[25] ,
		_w1073_,
		_w2432_
	);
	LUT2 #(
		.INIT('h1)
	) name1920 (
		_w2431_,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		_w2430_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h1)
	) name1922 (
		_w2427_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h4)
	) name1923 (
		_w2426_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		_w2430_,
		_w2433_,
		_w2437_
	);
	LUT2 #(
		.INIT('h2)
	) name1925 (
		\in0[26] ,
		_w1637_,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name1926 (
		\in1[26] ,
		_w1637_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name1927 (
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name1928 (
		\in2[26] ,
		_w1073_,
		_w2441_
	);
	LUT2 #(
		.INIT('h8)
	) name1929 (
		\in3[26] ,
		_w1073_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name1930 (
		_w2441_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name1931 (
		_w2440_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name1932 (
		_w2437_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h4)
	) name1933 (
		_w2436_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h2)
	) name1934 (
		_w2440_,
		_w2443_,
		_w2447_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w2446_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h1)
	) name1936 (
		_w2184_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h2)
	) name1937 (
		_w2180_,
		_w2183_,
		_w2450_
	);
	LUT2 #(
		.INIT('h2)
	) name1938 (
		\in0[28] ,
		_w1637_,
		_w2451_
	);
	LUT2 #(
		.INIT('h8)
	) name1939 (
		\in1[28] ,
		_w1637_,
		_w2452_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w2451_,
		_w2452_,
		_w2453_
	);
	LUT2 #(
		.INIT('h2)
	) name1941 (
		\in2[28] ,
		_w1073_,
		_w2454_
	);
	LUT2 #(
		.INIT('h8)
	) name1942 (
		\in3[28] ,
		_w1073_,
		_w2455_
	);
	LUT2 #(
		.INIT('h1)
	) name1943 (
		_w2454_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		_w2453_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h1)
	) name1945 (
		_w2450_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h4)
	) name1946 (
		_w2449_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h4)
	) name1947 (
		_w2453_,
		_w2456_,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name1948 (
		\in0[29] ,
		_w1637_,
		_w2461_
	);
	LUT2 #(
		.INIT('h8)
	) name1949 (
		\in1[29] ,
		_w1637_,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w2461_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		\in2[29] ,
		_w1073_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name1952 (
		\in3[29] ,
		_w1073_,
		_w2465_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w2464_,
		_w2465_,
		_w2466_
	);
	LUT2 #(
		.INIT('h4)
	) name1954 (
		_w2463_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name1955 (
		_w2460_,
		_w2467_,
		_w2468_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		_w2459_,
		_w2468_,
		_w2469_
	);
	LUT2 #(
		.INIT('h2)
	) name1957 (
		_w2463_,
		_w2466_,
		_w2470_
	);
	LUT2 #(
		.INIT('h2)
	) name1958 (
		\in0[30] ,
		_w1637_,
		_w2471_
	);
	LUT2 #(
		.INIT('h8)
	) name1959 (
		\in1[30] ,
		_w1637_,
		_w2472_
	);
	LUT2 #(
		.INIT('h1)
	) name1960 (
		_w2471_,
		_w2472_,
		_w2473_
	);
	LUT2 #(
		.INIT('h2)
	) name1961 (
		\in2[30] ,
		_w1073_,
		_w2474_
	);
	LUT2 #(
		.INIT('h8)
	) name1962 (
		\in3[30] ,
		_w1073_,
		_w2475_
	);
	LUT2 #(
		.INIT('h1)
	) name1963 (
		_w2474_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h2)
	) name1964 (
		_w2473_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		_w2470_,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w2469_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h4)
	) name1967 (
		_w2473_,
		_w2476_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		\in0[31] ,
		_w1637_,
		_w2481_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		\in1[31] ,
		_w1637_,
		_w2482_
	);
	LUT2 #(
		.INIT('h1)
	) name1970 (
		_w2481_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h2)
	) name1971 (
		\in2[31] ,
		_w1073_,
		_w2484_
	);
	LUT2 #(
		.INIT('h8)
	) name1972 (
		\in3[31] ,
		_w1073_,
		_w2485_
	);
	LUT2 #(
		.INIT('h1)
	) name1973 (
		_w2484_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h4)
	) name1974 (
		_w2483_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h1)
	) name1975 (
		_w2480_,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h4)
	) name1976 (
		_w2479_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h2)
	) name1977 (
		_w2483_,
		_w2486_,
		_w2490_
	);
	LUT2 #(
		.INIT('h2)
	) name1978 (
		\in0[35] ,
		_w1637_,
		_w2491_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		\in1[35] ,
		_w1637_,
		_w2492_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		_w2491_,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h2)
	) name1981 (
		\in2[35] ,
		_w1073_,
		_w2494_
	);
	LUT2 #(
		.INIT('h8)
	) name1982 (
		\in3[35] ,
		_w1073_,
		_w2495_
	);
	LUT2 #(
		.INIT('h1)
	) name1983 (
		_w2494_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h2)
	) name1984 (
		_w2493_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('h2)
	) name1985 (
		\in2[34] ,
		_w1073_,
		_w2498_
	);
	LUT2 #(
		.INIT('h8)
	) name1986 (
		\in3[34] ,
		_w1073_,
		_w2499_
	);
	LUT2 #(
		.INIT('h1)
	) name1987 (
		_w2498_,
		_w2499_,
		_w2500_
	);
	LUT2 #(
		.INIT('h2)
	) name1988 (
		\in0[34] ,
		_w1637_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name1989 (
		\in1[34] ,
		_w1637_,
		_w2502_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w2501_,
		_w2502_,
		_w2503_
	);
	LUT2 #(
		.INIT('h4)
	) name1991 (
		_w2500_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h2)
	) name1992 (
		\in0[33] ,
		_w1637_,
		_w2505_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		\in1[33] ,
		_w1637_,
		_w2506_
	);
	LUT2 #(
		.INIT('h1)
	) name1994 (
		_w2505_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('h2)
	) name1995 (
		\in2[33] ,
		_w1073_,
		_w2508_
	);
	LUT2 #(
		.INIT('h8)
	) name1996 (
		\in3[33] ,
		_w1073_,
		_w2509_
	);
	LUT2 #(
		.INIT('h1)
	) name1997 (
		_w2508_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		_w2507_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		_w2497_,
		_w2504_,
		_w2512_
	);
	LUT2 #(
		.INIT('h4)
	) name2000 (
		_w2511_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h2)
	) name2001 (
		\in0[37] ,
		_w1637_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name2002 (
		\in1[37] ,
		_w1637_,
		_w2515_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		_w2514_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		\in2[37] ,
		_w1073_,
		_w2517_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		\in3[37] ,
		_w1073_,
		_w2518_
	);
	LUT2 #(
		.INIT('h1)
	) name2006 (
		_w2517_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h2)
	) name2007 (
		_w2516_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		\in2[38] ,
		_w1073_,
		_w2521_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		\in3[38] ,
		_w1073_,
		_w2522_
	);
	LUT2 #(
		.INIT('h1)
	) name2010 (
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h2)
	) name2011 (
		\in0[38] ,
		_w1637_,
		_w2524_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		\in1[38] ,
		_w1637_,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name2013 (
		_w2524_,
		_w2525_,
		_w2526_
	);
	LUT2 #(
		.INIT('h4)
	) name2014 (
		_w2523_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h2)
	) name2015 (
		\in0[39] ,
		_w1637_,
		_w2528_
	);
	LUT2 #(
		.INIT('h8)
	) name2016 (
		\in1[39] ,
		_w1637_,
		_w2529_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w2528_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h2)
	) name2018 (
		\in2[39] ,
		_w1073_,
		_w2531_
	);
	LUT2 #(
		.INIT('h8)
	) name2019 (
		\in3[39] ,
		_w1073_,
		_w2532_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w2531_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h2)
	) name2021 (
		_w2530_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name2022 (
		_w2520_,
		_w2527_,
		_w2535_
	);
	LUT2 #(
		.INIT('h4)
	) name2023 (
		_w2534_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('h2)
	) name2024 (
		\in0[36] ,
		_w1637_,
		_w2537_
	);
	LUT2 #(
		.INIT('h8)
	) name2025 (
		\in1[36] ,
		_w1637_,
		_w2538_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		_w2537_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h2)
	) name2027 (
		\in2[36] ,
		_w1073_,
		_w2540_
	);
	LUT2 #(
		.INIT('h8)
	) name2028 (
		\in3[36] ,
		_w1073_,
		_w2541_
	);
	LUT2 #(
		.INIT('h1)
	) name2029 (
		_w2540_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name2030 (
		_w2539_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h2)
	) name2031 (
		\in2[32] ,
		_w1073_,
		_w2544_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		\in3[32] ,
		_w1073_,
		_w2545_
	);
	LUT2 #(
		.INIT('h1)
	) name2033 (
		_w2544_,
		_w2545_,
		_w2546_
	);
	LUT2 #(
		.INIT('h2)
	) name2034 (
		\in0[32] ,
		_w1637_,
		_w2547_
	);
	LUT2 #(
		.INIT('h8)
	) name2035 (
		\in1[32] ,
		_w1637_,
		_w2548_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		_w2547_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h4)
	) name2037 (
		_w2546_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h1)
	) name2038 (
		_w2490_,
		_w2543_,
		_w2551_
	);
	LUT2 #(
		.INIT('h4)
	) name2039 (
		_w2550_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h8)
	) name2040 (
		_w2513_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h8)
	) name2041 (
		_w2536_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w2489_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h2)
	) name2043 (
		_w2523_,
		_w2526_,
		_w2556_
	);
	LUT2 #(
		.INIT('h4)
	) name2044 (
		_w2534_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		_w2530_,
		_w2533_,
		_w2558_
	);
	LUT2 #(
		.INIT('h4)
	) name2046 (
		_w2539_,
		_w2542_,
		_w2559_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w2516_,
		_w2519_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		_w2500_,
		_w2503_,
		_w2561_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		_w2497_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		_w2493_,
		_w2496_,
		_w2563_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		_w2546_,
		_w2549_,
		_w2564_
	);
	LUT2 #(
		.INIT('h4)
	) name2052 (
		_w2507_,
		_w2510_,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w2564_,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h2)
	) name2054 (
		_w2513_,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name2055 (
		_w2562_,
		_w2563_,
		_w2568_
	);
	LUT2 #(
		.INIT('h4)
	) name2056 (
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		_w2543_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name2058 (
		_w2559_,
		_w2560_,
		_w2571_
	);
	LUT2 #(
		.INIT('h4)
	) name2059 (
		_w2570_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h2)
	) name2060 (
		_w2536_,
		_w2572_,
		_w2573_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		_w2557_,
		_w2558_,
		_w2574_
	);
	LUT2 #(
		.INIT('h4)
	) name2062 (
		_w2573_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h4)
	) name2063 (
		_w2555_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		\in0[43] ,
		_w1637_,
		_w2577_
	);
	LUT2 #(
		.INIT('h8)
	) name2065 (
		\in1[43] ,
		_w1637_,
		_w2578_
	);
	LUT2 #(
		.INIT('h1)
	) name2066 (
		_w2577_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\in2[43] ,
		_w1073_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name2068 (
		\in3[43] ,
		_w1073_,
		_w2581_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		_w2580_,
		_w2581_,
		_w2582_
	);
	LUT2 #(
		.INIT('h2)
	) name2070 (
		_w2579_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h2)
	) name2071 (
		\in0[42] ,
		_w1637_,
		_w2584_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		\in1[42] ,
		_w1637_,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name2073 (
		_w2584_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h2)
	) name2074 (
		\in2[42] ,
		_w1073_,
		_w2587_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		\in3[42] ,
		_w1073_,
		_w2588_
	);
	LUT2 #(
		.INIT('h1)
	) name2076 (
		_w2587_,
		_w2588_,
		_w2589_
	);
	LUT2 #(
		.INIT('h2)
	) name2077 (
		_w2586_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h1)
	) name2078 (
		_w2583_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h2)
	) name2079 (
		\in0[40] ,
		_w1637_,
		_w2592_
	);
	LUT2 #(
		.INIT('h8)
	) name2080 (
		\in1[40] ,
		_w1637_,
		_w2593_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w2592_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h2)
	) name2082 (
		\in2[40] ,
		_w1073_,
		_w2595_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		\in3[40] ,
		_w1073_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w2595_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h2)
	) name2085 (
		_w2594_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h2)
	) name2086 (
		\in0[44] ,
		_w1637_,
		_w2599_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		\in1[44] ,
		_w1637_,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('h2)
	) name2089 (
		\in2[44] ,
		_w1073_,
		_w2602_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		\in3[44] ,
		_w1073_,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name2091 (
		_w2602_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h2)
	) name2092 (
		_w2601_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h2)
	) name2093 (
		\in0[41] ,
		_w1637_,
		_w2606_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		\in1[41] ,
		_w1637_,
		_w2607_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		_w2606_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h2)
	) name2096 (
		\in2[41] ,
		_w1073_,
		_w2609_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		\in3[41] ,
		_w1073_,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name2098 (
		_w2609_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h2)
	) name2099 (
		_w2608_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		\in0[45] ,
		_w1637_,
		_w2613_
	);
	LUT2 #(
		.INIT('h8)
	) name2101 (
		\in1[45] ,
		_w1637_,
		_w2614_
	);
	LUT2 #(
		.INIT('h1)
	) name2102 (
		_w2613_,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h2)
	) name2103 (
		\in2[45] ,
		_w1073_,
		_w2616_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		\in3[45] ,
		_w1073_,
		_w2617_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w2616_,
		_w2617_,
		_w2618_
	);
	LUT2 #(
		.INIT('h2)
	) name2106 (
		_w2615_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h2)
	) name2107 (
		\in2[46] ,
		_w1073_,
		_w2620_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		\in3[46] ,
		_w1073_,
		_w2621_
	);
	LUT2 #(
		.INIT('h1)
	) name2109 (
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h2)
	) name2110 (
		\in0[46] ,
		_w1637_,
		_w2623_
	);
	LUT2 #(
		.INIT('h8)
	) name2111 (
		\in1[46] ,
		_w1637_,
		_w2624_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w2623_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h4)
	) name2113 (
		_w2622_,
		_w2625_,
		_w2626_
	);
	LUT2 #(
		.INIT('h2)
	) name2114 (
		\in0[47] ,
		_w1637_,
		_w2627_
	);
	LUT2 #(
		.INIT('h8)
	) name2115 (
		\in1[47] ,
		_w1637_,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h2)
	) name2117 (
		\in2[47] ,
		_w1073_,
		_w2630_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		\in3[47] ,
		_w1073_,
		_w2631_
	);
	LUT2 #(
		.INIT('h1)
	) name2119 (
		_w2630_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h2)
	) name2120 (
		_w2629_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name2121 (
		_w2619_,
		_w2626_,
		_w2634_
	);
	LUT2 #(
		.INIT('h4)
	) name2122 (
		_w2633_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h1)
	) name2123 (
		_w2598_,
		_w2605_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name2124 (
		_w2612_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('h8)
	) name2125 (
		_w2591_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		_w2635_,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h4)
	) name2127 (
		_w2576_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h2)
	) name2128 (
		_w2622_,
		_w2625_,
		_w2641_
	);
	LUT2 #(
		.INIT('h4)
	) name2129 (
		_w2633_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h4)
	) name2130 (
		_w2629_,
		_w2632_,
		_w2643_
	);
	LUT2 #(
		.INIT('h4)
	) name2131 (
		_w2601_,
		_w2604_,
		_w2644_
	);
	LUT2 #(
		.INIT('h4)
	) name2132 (
		_w2615_,
		_w2618_,
		_w2645_
	);
	LUT2 #(
		.INIT('h4)
	) name2133 (
		_w2579_,
		_w2582_,
		_w2646_
	);
	LUT2 #(
		.INIT('h4)
	) name2134 (
		_w2586_,
		_w2589_,
		_w2647_
	);
	LUT2 #(
		.INIT('h4)
	) name2135 (
		_w2608_,
		_w2611_,
		_w2648_
	);
	LUT2 #(
		.INIT('h4)
	) name2136 (
		_w2594_,
		_w2597_,
		_w2649_
	);
	LUT2 #(
		.INIT('h4)
	) name2137 (
		_w2612_,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		_w2647_,
		_w2648_,
		_w2651_
	);
	LUT2 #(
		.INIT('h4)
	) name2139 (
		_w2650_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		_w2591_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h1)
	) name2141 (
		_w2646_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		_w2605_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w2644_,
		_w2645_,
		_w2656_
	);
	LUT2 #(
		.INIT('h4)
	) name2144 (
		_w2655_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h2)
	) name2145 (
		_w2635_,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h1)
	) name2146 (
		_w2642_,
		_w2643_,
		_w2659_
	);
	LUT2 #(
		.INIT('h4)
	) name2147 (
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT2 #(
		.INIT('h4)
	) name2148 (
		_w2640_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h2)
	) name2149 (
		\in0[51] ,
		_w1637_,
		_w2662_
	);
	LUT2 #(
		.INIT('h8)
	) name2150 (
		\in1[51] ,
		_w1637_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		_w2662_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		\in2[51] ,
		_w1073_,
		_w2665_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		\in3[51] ,
		_w1073_,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w2665_,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h2)
	) name2155 (
		_w2664_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h2)
	) name2156 (
		\in2[50] ,
		_w1073_,
		_w2669_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		\in3[50] ,
		_w1073_,
		_w2670_
	);
	LUT2 #(
		.INIT('h1)
	) name2158 (
		_w2669_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h2)
	) name2159 (
		\in0[50] ,
		_w1637_,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		\in1[50] ,
		_w1637_,
		_w2673_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w2672_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h4)
	) name2162 (
		_w2671_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name2163 (
		\in0[49] ,
		_w1637_,
		_w2676_
	);
	LUT2 #(
		.INIT('h8)
	) name2164 (
		\in1[49] ,
		_w1637_,
		_w2677_
	);
	LUT2 #(
		.INIT('h1)
	) name2165 (
		_w2676_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h2)
	) name2166 (
		\in2[49] ,
		_w1073_,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		\in3[49] ,
		_w1073_,
		_w2680_
	);
	LUT2 #(
		.INIT('h1)
	) name2168 (
		_w2679_,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h2)
	) name2169 (
		_w2678_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w2668_,
		_w2675_,
		_w2683_
	);
	LUT2 #(
		.INIT('h4)
	) name2171 (
		_w2682_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h2)
	) name2172 (
		\in2[48] ,
		_w1073_,
		_w2685_
	);
	LUT2 #(
		.INIT('h8)
	) name2173 (
		\in3[48] ,
		_w1073_,
		_w2686_
	);
	LUT2 #(
		.INIT('h1)
	) name2174 (
		_w2685_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h2)
	) name2175 (
		\in0[48] ,
		_w1637_,
		_w2688_
	);
	LUT2 #(
		.INIT('h8)
	) name2176 (
		\in1[48] ,
		_w1637_,
		_w2689_
	);
	LUT2 #(
		.INIT('h1)
	) name2177 (
		_w2688_,
		_w2689_,
		_w2690_
	);
	LUT2 #(
		.INIT('h4)
	) name2178 (
		_w2687_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h2)
	) name2179 (
		\in0[55] ,
		_w1637_,
		_w2692_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		\in1[55] ,
		_w1637_,
		_w2693_
	);
	LUT2 #(
		.INIT('h1)
	) name2181 (
		_w2692_,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		\in2[55] ,
		_w1073_,
		_w2695_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		\in3[55] ,
		_w1073_,
		_w2696_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		_w2695_,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h2)
	) name2185 (
		_w2694_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h2)
	) name2186 (
		\in2[54] ,
		_w1073_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		\in3[54] ,
		_w1073_,
		_w2700_
	);
	LUT2 #(
		.INIT('h1)
	) name2188 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h2)
	) name2189 (
		\in0[54] ,
		_w1637_,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name2190 (
		\in1[54] ,
		_w1637_,
		_w2703_
	);
	LUT2 #(
		.INIT('h1)
	) name2191 (
		_w2702_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h4)
	) name2192 (
		_w2701_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name2193 (
		_w2698_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h2)
	) name2194 (
		\in0[53] ,
		_w1637_,
		_w2707_
	);
	LUT2 #(
		.INIT('h8)
	) name2195 (
		\in1[53] ,
		_w1637_,
		_w2708_
	);
	LUT2 #(
		.INIT('h1)
	) name2196 (
		_w2707_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h2)
	) name2197 (
		\in2[53] ,
		_w1073_,
		_w2710_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		\in3[53] ,
		_w1073_,
		_w2711_
	);
	LUT2 #(
		.INIT('h1)
	) name2199 (
		_w2710_,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h2)
	) name2200 (
		_w2709_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h2)
	) name2201 (
		\in2[52] ,
		_w1073_,
		_w2714_
	);
	LUT2 #(
		.INIT('h8)
	) name2202 (
		\in3[52] ,
		_w1073_,
		_w2715_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w2714_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h2)
	) name2204 (
		\in0[52] ,
		_w1637_,
		_w2717_
	);
	LUT2 #(
		.INIT('h8)
	) name2205 (
		\in1[52] ,
		_w1637_,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w2717_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h4)
	) name2207 (
		_w2716_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		_w2713_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		_w2706_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h2)
	) name2210 (
		_w2684_,
		_w2691_,
		_w2723_
	);
	LUT2 #(
		.INIT('h8)
	) name2211 (
		_w2722_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h4)
	) name2212 (
		_w2661_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h4)
	) name2213 (
		_w2694_,
		_w2697_,
		_w2726_
	);
	LUT2 #(
		.INIT('h4)
	) name2214 (
		_w2664_,
		_w2667_,
		_w2727_
	);
	LUT2 #(
		.INIT('h2)
	) name2215 (
		_w2687_,
		_w2690_,
		_w2728_
	);
	LUT2 #(
		.INIT('h4)
	) name2216 (
		_w2678_,
		_w2681_,
		_w2729_
	);
	LUT2 #(
		.INIT('h1)
	) name2217 (
		_w2728_,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h2)
	) name2218 (
		_w2684_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name2219 (
		_w2671_,
		_w2674_,
		_w2732_
	);
	LUT2 #(
		.INIT('h4)
	) name2220 (
		_w2668_,
		_w2732_,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name2221 (
		_w2727_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h4)
	) name2222 (
		_w2731_,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		_w2722_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h4)
	) name2224 (
		_w2709_,
		_w2712_,
		_w2737_
	);
	LUT2 #(
		.INIT('h2)
	) name2225 (
		_w2701_,
		_w2704_,
		_w2738_
	);
	LUT2 #(
		.INIT('h2)
	) name2226 (
		_w2716_,
		_w2719_,
		_w2739_
	);
	LUT2 #(
		.INIT('h4)
	) name2227 (
		_w2713_,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		_w2737_,
		_w2738_,
		_w2741_
	);
	LUT2 #(
		.INIT('h4)
	) name2229 (
		_w2740_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h2)
	) name2230 (
		_w2706_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		_w2726_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h4)
	) name2232 (
		_w2736_,
		_w2744_,
		_w2745_
	);
	LUT2 #(
		.INIT('h4)
	) name2233 (
		_w2725_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h2)
	) name2234 (
		\in0[59] ,
		_w1637_,
		_w2747_
	);
	LUT2 #(
		.INIT('h8)
	) name2235 (
		\in1[59] ,
		_w1637_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name2236 (
		_w2747_,
		_w2748_,
		_w2749_
	);
	LUT2 #(
		.INIT('h2)
	) name2237 (
		\in2[59] ,
		_w1073_,
		_w2750_
	);
	LUT2 #(
		.INIT('h8)
	) name2238 (
		\in3[59] ,
		_w1073_,
		_w2751_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w2750_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h2)
	) name2240 (
		_w2749_,
		_w2752_,
		_w2753_
	);
	LUT2 #(
		.INIT('h2)
	) name2241 (
		\in0[58] ,
		_w1637_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		\in1[58] ,
		_w1637_,
		_w2755_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		_w2754_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h2)
	) name2244 (
		\in2[58] ,
		_w1073_,
		_w2757_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		\in3[58] ,
		_w1073_,
		_w2758_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		_w2757_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h2)
	) name2247 (
		_w2756_,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h1)
	) name2248 (
		_w2753_,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h2)
	) name2249 (
		\in0[56] ,
		_w1637_,
		_w2762_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		\in1[56] ,
		_w1637_,
		_w2763_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		_w2762_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		\in2[56] ,
		_w1073_,
		_w2765_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		\in3[56] ,
		_w1073_,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name2254 (
		_w2765_,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name2255 (
		_w2764_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h2)
	) name2256 (
		\in0[60] ,
		_w1637_,
		_w2769_
	);
	LUT2 #(
		.INIT('h8)
	) name2257 (
		\in1[60] ,
		_w1637_,
		_w2770_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		_w2769_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name2259 (
		\in2[60] ,
		_w1073_,
		_w2772_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		\in3[60] ,
		_w1073_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		_w2772_,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h2)
	) name2262 (
		_w2771_,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h2)
	) name2263 (
		\in0[57] ,
		_w1637_,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		\in1[57] ,
		_w1637_,
		_w2777_
	);
	LUT2 #(
		.INIT('h1)
	) name2265 (
		_w2776_,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h2)
	) name2266 (
		\in2[57] ,
		_w1073_,
		_w2779_
	);
	LUT2 #(
		.INIT('h8)
	) name2267 (
		\in3[57] ,
		_w1073_,
		_w2780_
	);
	LUT2 #(
		.INIT('h1)
	) name2268 (
		_w2779_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h2)
	) name2269 (
		_w2778_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h2)
	) name2270 (
		\in0[61] ,
		_w1637_,
		_w2783_
	);
	LUT2 #(
		.INIT('h8)
	) name2271 (
		\in1[61] ,
		_w1637_,
		_w2784_
	);
	LUT2 #(
		.INIT('h1)
	) name2272 (
		_w2783_,
		_w2784_,
		_w2785_
	);
	LUT2 #(
		.INIT('h2)
	) name2273 (
		\in2[61] ,
		_w1073_,
		_w2786_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		\in3[61] ,
		_w1073_,
		_w2787_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w2786_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h2)
	) name2276 (
		_w2785_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h2)
	) name2277 (
		\in2[62] ,
		_w1073_,
		_w2790_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		\in3[62] ,
		_w1073_,
		_w2791_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		_w2790_,
		_w2791_,
		_w2792_
	);
	LUT2 #(
		.INIT('h2)
	) name2280 (
		\in0[62] ,
		_w1637_,
		_w2793_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		\in1[62] ,
		_w1637_,
		_w2794_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w2793_,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h4)
	) name2283 (
		_w2792_,
		_w2795_,
		_w2796_
	);
	LUT2 #(
		.INIT('h2)
	) name2284 (
		\in0[63] ,
		_w1637_,
		_w2797_
	);
	LUT2 #(
		.INIT('h8)
	) name2285 (
		\in1[63] ,
		_w1637_,
		_w2798_
	);
	LUT2 #(
		.INIT('h1)
	) name2286 (
		_w2797_,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h2)
	) name2287 (
		\in2[63] ,
		_w1073_,
		_w2800_
	);
	LUT2 #(
		.INIT('h8)
	) name2288 (
		\in3[63] ,
		_w1073_,
		_w2801_
	);
	LUT2 #(
		.INIT('h1)
	) name2289 (
		_w2800_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h2)
	) name2290 (
		_w2799_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w2789_,
		_w2796_,
		_w2804_
	);
	LUT2 #(
		.INIT('h4)
	) name2292 (
		_w2803_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		_w2768_,
		_w2775_,
		_w2806_
	);
	LUT2 #(
		.INIT('h4)
	) name2294 (
		_w2782_,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		_w2761_,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		_w2805_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h4)
	) name2297 (
		_w2746_,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h2)
	) name2298 (
		_w2792_,
		_w2795_,
		_w2811_
	);
	LUT2 #(
		.INIT('h4)
	) name2299 (
		_w2803_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h4)
	) name2300 (
		_w2799_,
		_w2802_,
		_w2813_
	);
	LUT2 #(
		.INIT('h4)
	) name2301 (
		_w2771_,
		_w2774_,
		_w2814_
	);
	LUT2 #(
		.INIT('h4)
	) name2302 (
		_w2785_,
		_w2788_,
		_w2815_
	);
	LUT2 #(
		.INIT('h4)
	) name2303 (
		_w2749_,
		_w2752_,
		_w2816_
	);
	LUT2 #(
		.INIT('h4)
	) name2304 (
		_w2756_,
		_w2759_,
		_w2817_
	);
	LUT2 #(
		.INIT('h4)
	) name2305 (
		_w2778_,
		_w2781_,
		_w2818_
	);
	LUT2 #(
		.INIT('h4)
	) name2306 (
		_w2764_,
		_w2767_,
		_w2819_
	);
	LUT2 #(
		.INIT('h4)
	) name2307 (
		_w2782_,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		_w2817_,
		_w2818_,
		_w2821_
	);
	LUT2 #(
		.INIT('h4)
	) name2309 (
		_w2820_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h2)
	) name2310 (
		_w2761_,
		_w2822_,
		_w2823_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		_w2816_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h1)
	) name2312 (
		_w2775_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		_w2814_,
		_w2815_,
		_w2826_
	);
	LUT2 #(
		.INIT('h4)
	) name2314 (
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name2315 (
		_w2805_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h1)
	) name2316 (
		_w2812_,
		_w2813_,
		_w2829_
	);
	LUT2 #(
		.INIT('h4)
	) name2317 (
		_w2828_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h4)
	) name2318 (
		_w2810_,
		_w2830_,
		_w2831_
	);
	LUT2 #(
		.INIT('h4)
	) name2319 (
		_w2168_,
		_w2172_,
		_w2832_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		_w2169_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w2157_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h4)
	) name2322 (
		_w2831_,
		_w2834_,
		_w2835_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		_w2148_,
		_w2177_,
		_w2836_
	);
	LUT2 #(
		.INIT('h4)
	) name2324 (
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h4)
	) name2325 (
		_w2132_,
		_w2136_,
		_w2838_
	);
	LUT2 #(
		.INIT('h1)
	) name2326 (
		_w2133_,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('h8)
	) name2327 (
		_w2121_,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h4)
	) name2328 (
		_w2837_,
		_w2840_,
		_w2841_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w2112_,
		_w2141_,
		_w2842_
	);
	LUT2 #(
		.INIT('h4)
	) name2330 (
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h4)
	) name2331 (
		_w2096_,
		_w2100_,
		_w2844_
	);
	LUT2 #(
		.INIT('h1)
	) name2332 (
		_w2097_,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h8)
	) name2333 (
		_w2085_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h4)
	) name2334 (
		_w2843_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h1)
	) name2335 (
		_w2076_,
		_w2105_,
		_w2848_
	);
	LUT2 #(
		.INIT('h4)
	) name2336 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h4)
	) name2337 (
		_w2060_,
		_w2064_,
		_w2850_
	);
	LUT2 #(
		.INIT('h1)
	) name2338 (
		_w2061_,
		_w2850_,
		_w2851_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		_w2049_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h4)
	) name2340 (
		_w2849_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w2040_,
		_w2069_,
		_w2854_
	);
	LUT2 #(
		.INIT('h4)
	) name2342 (
		_w2853_,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h4)
	) name2343 (
		_w2024_,
		_w2028_,
		_w2856_
	);
	LUT2 #(
		.INIT('h1)
	) name2344 (
		_w2025_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		_w2013_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h4)
	) name2346 (
		_w2855_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h1)
	) name2347 (
		_w2004_,
		_w2033_,
		_w2860_
	);
	LUT2 #(
		.INIT('h4)
	) name2348 (
		_w2859_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h4)
	) name2349 (
		_w1988_,
		_w1992_,
		_w2862_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		_w1989_,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		_w1977_,
		_w2863_,
		_w2864_
	);
	LUT2 #(
		.INIT('h4)
	) name2352 (
		_w2861_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w1968_,
		_w1997_,
		_w2866_
	);
	LUT2 #(
		.INIT('h4)
	) name2354 (
		_w2865_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h4)
	) name2355 (
		_w1952_,
		_w1956_,
		_w2868_
	);
	LUT2 #(
		.INIT('h1)
	) name2356 (
		_w1953_,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h8)
	) name2357 (
		_w1941_,
		_w2869_,
		_w2870_
	);
	LUT2 #(
		.INIT('h4)
	) name2358 (
		_w2867_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		_w1932_,
		_w1961_,
		_w2872_
	);
	LUT2 #(
		.INIT('h4)
	) name2360 (
		_w2871_,
		_w2872_,
		_w2873_
	);
	LUT2 #(
		.INIT('h4)
	) name2361 (
		_w1916_,
		_w1920_,
		_w2874_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w1917_,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name2363 (
		_w1905_,
		_w2875_,
		_w2876_
	);
	LUT2 #(
		.INIT('h4)
	) name2364 (
		_w2873_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w1896_,
		_w1925_,
		_w2878_
	);
	LUT2 #(
		.INIT('h4)
	) name2366 (
		_w2877_,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h4)
	) name2367 (
		_w1880_,
		_w1884_,
		_w2880_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		_w1881_,
		_w2880_,
		_w2881_
	);
	LUT2 #(
		.INIT('h8)
	) name2369 (
		_w1869_,
		_w2881_,
		_w2882_
	);
	LUT2 #(
		.INIT('h4)
	) name2370 (
		_w2879_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w1860_,
		_w1889_,
		_w2884_
	);
	LUT2 #(
		.INIT('h4)
	) name2372 (
		_w2883_,
		_w2884_,
		_w2885_
	);
	LUT2 #(
		.INIT('h4)
	) name2373 (
		_w1844_,
		_w1848_,
		_w2886_
	);
	LUT2 #(
		.INIT('h1)
	) name2374 (
		_w1845_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		_w1833_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('h4)
	) name2376 (
		_w2885_,
		_w2888_,
		_w2889_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w1824_,
		_w1853_,
		_w2890_
	);
	LUT2 #(
		.INIT('h4)
	) name2378 (
		_w2889_,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h4)
	) name2379 (
		_w1808_,
		_w1812_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name2380 (
		_w1809_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h8)
	) name2381 (
		_w1797_,
		_w2893_,
		_w2894_
	);
	LUT2 #(
		.INIT('h4)
	) name2382 (
		_w2891_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w1788_,
		_w1817_,
		_w2896_
	);
	LUT2 #(
		.INIT('h4)
	) name2384 (
		_w2895_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h4)
	) name2385 (
		_w1772_,
		_w1776_,
		_w2898_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		_w1773_,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h8)
	) name2387 (
		_w1761_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h4)
	) name2388 (
		_w2897_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		_w1752_,
		_w1781_,
		_w2902_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		_w2901_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h4)
	) name2391 (
		_w1736_,
		_w1740_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name2392 (
		_w1737_,
		_w2904_,
		_w2905_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		_w1725_,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h4)
	) name2394 (
		_w2903_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h1)
	) name2395 (
		_w1716_,
		_w1745_,
		_w2908_
	);
	LUT2 #(
		.INIT('h4)
	) name2396 (
		_w2907_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h4)
	) name2397 (
		_w1700_,
		_w1704_,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name2398 (
		_w1701_,
		_w2910_,
		_w2911_
	);
	LUT2 #(
		.INIT('h8)
	) name2399 (
		_w1689_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h4)
	) name2400 (
		_w2909_,
		_w2912_,
		_w2913_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w1680_,
		_w1709_,
		_w2914_
	);
	LUT2 #(
		.INIT('h4)
	) name2402 (
		_w2913_,
		_w2914_,
		_w2915_
	);
	LUT2 #(
		.INIT('h4)
	) name2403 (
		_w1664_,
		_w1668_,
		_w2916_
	);
	LUT2 #(
		.INIT('h1)
	) name2404 (
		_w1665_,
		_w2916_,
		_w2917_
	);
	LUT2 #(
		.INIT('h8)
	) name2405 (
		_w1653_,
		_w2917_,
		_w2918_
	);
	LUT2 #(
		.INIT('h4)
	) name2406 (
		_w2915_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name2407 (
		_w1644_,
		_w1673_,
		_w2920_
	);
	LUT2 #(
		.INIT('h4)
	) name2408 (
		_w2919_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name2409 (
		\in2[127] ,
		\in3[127] ,
		_w2922_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		\in0[127] ,
		\in1[127] ,
		_w2923_
	);
	LUT2 #(
		.INIT('h4)
	) name2411 (
		_w2922_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h2)
	) name2412 (
		\in0[126] ,
		_w1637_,
		_w2925_
	);
	LUT2 #(
		.INIT('h8)
	) name2413 (
		\in1[126] ,
		_w1637_,
		_w2926_
	);
	LUT2 #(
		.INIT('h1)
	) name2414 (
		_w2925_,
		_w2926_,
		_w2927_
	);
	LUT2 #(
		.INIT('h2)
	) name2415 (
		\in2[126] ,
		_w1073_,
		_w2928_
	);
	LUT2 #(
		.INIT('h8)
	) name2416 (
		\in3[126] ,
		_w1073_,
		_w2929_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		_w2928_,
		_w2929_,
		_w2930_
	);
	LUT2 #(
		.INIT('h2)
	) name2418 (
		_w2927_,
		_w2930_,
		_w2931_
	);
	LUT2 #(
		.INIT('h2)
	) name2419 (
		\in0[125] ,
		_w1637_,
		_w2932_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		\in1[125] ,
		_w1637_,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name2421 (
		_w2932_,
		_w2933_,
		_w2934_
	);
	LUT2 #(
		.INIT('h2)
	) name2422 (
		\in2[125] ,
		_w1073_,
		_w2935_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		\in3[125] ,
		_w1073_,
		_w2936_
	);
	LUT2 #(
		.INIT('h1)
	) name2424 (
		_w2935_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('h2)
	) name2425 (
		_w2934_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name2426 (
		_w2931_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h2)
	) name2427 (
		\in0[124] ,
		_w1637_,
		_w2940_
	);
	LUT2 #(
		.INIT('h8)
	) name2428 (
		\in1[124] ,
		_w1637_,
		_w2941_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w2940_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h2)
	) name2430 (
		\in2[124] ,
		_w1073_,
		_w2943_
	);
	LUT2 #(
		.INIT('h8)
	) name2431 (
		\in3[124] ,
		_w1073_,
		_w2944_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		_w2943_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h2)
	) name2433 (
		_w2942_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w2924_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h8)
	) name2435 (
		_w2939_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h4)
	) name2436 (
		_w2921_,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h2)
	) name2437 (
		_w2922_,
		_w2923_,
		_w2950_
	);
	LUT2 #(
		.INIT('h4)
	) name2438 (
		_w2942_,
		_w2945_,
		_w2951_
	);
	LUT2 #(
		.INIT('h4)
	) name2439 (
		_w2934_,
		_w2937_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		_w2951_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h2)
	) name2441 (
		_w2939_,
		_w2953_,
		_w2954_
	);
	LUT2 #(
		.INIT('h4)
	) name2442 (
		_w2927_,
		_w2930_,
		_w2955_
	);
	LUT2 #(
		.INIT('h1)
	) name2443 (
		_w2950_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h4)
	) name2444 (
		_w2954_,
		_w2956_,
		_w2957_
	);
	LUT2 #(
		.INIT('h1)
	) name2445 (
		_w2924_,
		_w2957_,
		_w2958_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		_w2949_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h4)
	) name2447 (
		_w1076_,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name2448 (
		_w2208_,
		_w2959_,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name2449 (
		_w2960_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h4)
	) name2450 (
		_w2201_,
		_w2959_,
		_w2963_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		_w2204_,
		_w2959_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		_w2963_,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h4)
	) name2453 (
		_w2216_,
		_w2959_,
		_w2966_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		_w2213_,
		_w2959_,
		_w2967_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w2966_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h4)
	) name2456 (
		_w2226_,
		_w2959_,
		_w2969_
	);
	LUT2 #(
		.INIT('h1)
	) name2457 (
		_w2223_,
		_w2959_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name2458 (
		_w2969_,
		_w2970_,
		_w2971_
	);
	LUT2 #(
		.INIT('h2)
	) name2459 (
		_w2234_,
		_w2959_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		_w2237_,
		_w2959_,
		_w2973_
	);
	LUT2 #(
		.INIT('h1)
	) name2461 (
		_w2972_,
		_w2973_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name2462 (
		_w2247_,
		_w2959_,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name2463 (
		_w2244_,
		_w2959_,
		_w2976_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w2975_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h2)
	) name2465 (
		_w2197_,
		_w2959_,
		_w2978_
	);
	LUT2 #(
		.INIT('h8)
	) name2466 (
		_w2194_,
		_w2959_,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name2467 (
		_w2978_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h4)
	) name2468 (
		_w2260_,
		_w2959_,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name2469 (
		_w2257_,
		_w2959_,
		_w2982_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		_w2981_,
		_w2982_,
		_w2983_
	);
	LUT2 #(
		.INIT('h4)
	) name2471 (
		_w2270_,
		_w2959_,
		_w2984_
	);
	LUT2 #(
		.INIT('h1)
	) name2472 (
		_w2267_,
		_w2959_,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w2984_,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('h4)
	) name2474 (
		_w2280_,
		_w2959_,
		_w2987_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		_w2277_,
		_w2959_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name2476 (
		_w2987_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h4)
	) name2477 (
		_w2289_,
		_w2959_,
		_w2990_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		_w2286_,
		_w2959_,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name2479 (
		_w2990_,
		_w2991_,
		_w2992_
	);
	LUT2 #(
		.INIT('h4)
	) name2480 (
		_w2300_,
		_w2959_,
		_w2993_
	);
	LUT2 #(
		.INIT('h1)
	) name2481 (
		_w2297_,
		_w2959_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		_w2993_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h4)
	) name2483 (
		_w2190_,
		_w2959_,
		_w2996_
	);
	LUT2 #(
		.INIT('h1)
	) name2484 (
		_w2187_,
		_w2959_,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w2996_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h4)
	) name2486 (
		_w2313_,
		_w2959_,
		_w2999_
	);
	LUT2 #(
		.INIT('h1)
	) name2487 (
		_w2310_,
		_w2959_,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name2488 (
		_w2999_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h4)
	) name2489 (
		_w2323_,
		_w2959_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name2490 (
		_w2320_,
		_w2959_,
		_w3003_
	);
	LUT2 #(
		.INIT('h1)
	) name2491 (
		_w3002_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h4)
	) name2492 (
		_w2333_,
		_w2959_,
		_w3005_
	);
	LUT2 #(
		.INIT('h1)
	) name2493 (
		_w2330_,
		_w2959_,
		_w3006_
	);
	LUT2 #(
		.INIT('h1)
	) name2494 (
		_w3005_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h4)
	) name2495 (
		_w2343_,
		_w2959_,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name2496 (
		_w2340_,
		_w2959_,
		_w3009_
	);
	LUT2 #(
		.INIT('h1)
	) name2497 (
		_w3008_,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h4)
	) name2498 (
		_w2353_,
		_w2959_,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name2499 (
		_w2350_,
		_w2959_,
		_w3012_
	);
	LUT2 #(
		.INIT('h1)
	) name2500 (
		_w3011_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h4)
	) name2501 (
		_w2363_,
		_w2959_,
		_w3014_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w2360_,
		_w2959_,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2503 (
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h4)
	) name2504 (
		_w2370_,
		_w2959_,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		_w2373_,
		_w2959_,
		_w3018_
	);
	LUT2 #(
		.INIT('h1)
	) name2506 (
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h4)
	) name2507 (
		_w2382_,
		_w2959_,
		_w3020_
	);
	LUT2 #(
		.INIT('h1)
	) name2508 (
		_w2379_,
		_w2959_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name2509 (
		_w3020_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h4)
	) name2510 (
		_w2392_,
		_w2959_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name2511 (
		_w2389_,
		_w2959_,
		_w3024_
	);
	LUT2 #(
		.INIT('h1)
	) name2512 (
		_w3023_,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h4)
	) name2513 (
		_w2403_,
		_w2959_,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name2514 (
		_w2400_,
		_w2959_,
		_w3027_
	);
	LUT2 #(
		.INIT('h1)
	) name2515 (
		_w3026_,
		_w3027_,
		_w3028_
	);
	LUT2 #(
		.INIT('h4)
	) name2516 (
		_w2413_,
		_w2959_,
		_w3029_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w2410_,
		_w2959_,
		_w3030_
	);
	LUT2 #(
		.INIT('h1)
	) name2518 (
		_w3029_,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h4)
	) name2519 (
		_w2423_,
		_w2959_,
		_w3032_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w2420_,
		_w2959_,
		_w3033_
	);
	LUT2 #(
		.INIT('h1)
	) name2521 (
		_w3032_,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h4)
	) name2522 (
		_w2433_,
		_w2959_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2523 (
		_w2430_,
		_w2959_,
		_w3036_
	);
	LUT2 #(
		.INIT('h1)
	) name2524 (
		_w3035_,
		_w3036_,
		_w3037_
	);
	LUT2 #(
		.INIT('h4)
	) name2525 (
		_w2443_,
		_w2959_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name2526 (
		_w2440_,
		_w2959_,
		_w3039_
	);
	LUT2 #(
		.INIT('h1)
	) name2527 (
		_w3038_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h4)
	) name2528 (
		_w2183_,
		_w2959_,
		_w3041_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		_w2180_,
		_w2959_,
		_w3042_
	);
	LUT2 #(
		.INIT('h1)
	) name2530 (
		_w3041_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h4)
	) name2531 (
		_w2456_,
		_w2959_,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		_w2453_,
		_w2959_,
		_w3045_
	);
	LUT2 #(
		.INIT('h1)
	) name2533 (
		_w3044_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h4)
	) name2534 (
		_w2466_,
		_w2959_,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name2535 (
		_w2463_,
		_w2959_,
		_w3048_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w3047_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h4)
	) name2537 (
		_w2476_,
		_w2959_,
		_w3050_
	);
	LUT2 #(
		.INIT('h1)
	) name2538 (
		_w2473_,
		_w2959_,
		_w3051_
	);
	LUT2 #(
		.INIT('h1)
	) name2539 (
		_w3050_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h4)
	) name2540 (
		_w2486_,
		_w2959_,
		_w3053_
	);
	LUT2 #(
		.INIT('h1)
	) name2541 (
		_w2483_,
		_w2959_,
		_w3054_
	);
	LUT2 #(
		.INIT('h1)
	) name2542 (
		_w3053_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h4)
	) name2543 (
		_w2546_,
		_w2959_,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name2544 (
		_w2549_,
		_w2959_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name2545 (
		_w3056_,
		_w3057_,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		_w2510_,
		_w2959_,
		_w3059_
	);
	LUT2 #(
		.INIT('h1)
	) name2547 (
		_w2507_,
		_w2959_,
		_w3060_
	);
	LUT2 #(
		.INIT('h1)
	) name2548 (
		_w3059_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h4)
	) name2549 (
		_w2500_,
		_w2959_,
		_w3062_
	);
	LUT2 #(
		.INIT('h1)
	) name2550 (
		_w2503_,
		_w2959_,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name2551 (
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h4)
	) name2552 (
		_w2496_,
		_w2959_,
		_w3065_
	);
	LUT2 #(
		.INIT('h1)
	) name2553 (
		_w2493_,
		_w2959_,
		_w3066_
	);
	LUT2 #(
		.INIT('h1)
	) name2554 (
		_w3065_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h4)
	) name2555 (
		_w2542_,
		_w2959_,
		_w3068_
	);
	LUT2 #(
		.INIT('h1)
	) name2556 (
		_w2539_,
		_w2959_,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w3068_,
		_w3069_,
		_w3070_
	);
	LUT2 #(
		.INIT('h4)
	) name2558 (
		_w2519_,
		_w2959_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name2559 (
		_w2516_,
		_w2959_,
		_w3072_
	);
	LUT2 #(
		.INIT('h1)
	) name2560 (
		_w3071_,
		_w3072_,
		_w3073_
	);
	LUT2 #(
		.INIT('h4)
	) name2561 (
		_w2523_,
		_w2959_,
		_w3074_
	);
	LUT2 #(
		.INIT('h1)
	) name2562 (
		_w2526_,
		_w2959_,
		_w3075_
	);
	LUT2 #(
		.INIT('h1)
	) name2563 (
		_w3074_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('h4)
	) name2564 (
		_w2533_,
		_w2959_,
		_w3077_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w2530_,
		_w2959_,
		_w3078_
	);
	LUT2 #(
		.INIT('h1)
	) name2566 (
		_w3077_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h4)
	) name2567 (
		_w2597_,
		_w2959_,
		_w3080_
	);
	LUT2 #(
		.INIT('h1)
	) name2568 (
		_w2594_,
		_w2959_,
		_w3081_
	);
	LUT2 #(
		.INIT('h1)
	) name2569 (
		_w3080_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h4)
	) name2570 (
		_w2611_,
		_w2959_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2571 (
		_w2608_,
		_w2959_,
		_w3084_
	);
	LUT2 #(
		.INIT('h1)
	) name2572 (
		_w3083_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h4)
	) name2573 (
		_w2589_,
		_w2959_,
		_w3086_
	);
	LUT2 #(
		.INIT('h1)
	) name2574 (
		_w2586_,
		_w2959_,
		_w3087_
	);
	LUT2 #(
		.INIT('h1)
	) name2575 (
		_w3086_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h4)
	) name2576 (
		_w2582_,
		_w2959_,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w2579_,
		_w2959_,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name2578 (
		_w3089_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h4)
	) name2579 (
		_w2604_,
		_w2959_,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name2580 (
		_w2601_,
		_w2959_,
		_w3093_
	);
	LUT2 #(
		.INIT('h1)
	) name2581 (
		_w3092_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h4)
	) name2582 (
		_w2618_,
		_w2959_,
		_w3095_
	);
	LUT2 #(
		.INIT('h1)
	) name2583 (
		_w2615_,
		_w2959_,
		_w3096_
	);
	LUT2 #(
		.INIT('h1)
	) name2584 (
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h4)
	) name2585 (
		_w2622_,
		_w2959_,
		_w3098_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w2625_,
		_w2959_,
		_w3099_
	);
	LUT2 #(
		.INIT('h1)
	) name2587 (
		_w3098_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h4)
	) name2588 (
		_w2632_,
		_w2959_,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name2589 (
		_w2629_,
		_w2959_,
		_w3102_
	);
	LUT2 #(
		.INIT('h1)
	) name2590 (
		_w3101_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h4)
	) name2591 (
		_w2687_,
		_w2959_,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w2690_,
		_w2959_,
		_w3105_
	);
	LUT2 #(
		.INIT('h1)
	) name2593 (
		_w3104_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h4)
	) name2594 (
		_w2681_,
		_w2959_,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name2595 (
		_w2678_,
		_w2959_,
		_w3108_
	);
	LUT2 #(
		.INIT('h1)
	) name2596 (
		_w3107_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h4)
	) name2597 (
		_w2671_,
		_w2959_,
		_w3110_
	);
	LUT2 #(
		.INIT('h1)
	) name2598 (
		_w2674_,
		_w2959_,
		_w3111_
	);
	LUT2 #(
		.INIT('h1)
	) name2599 (
		_w3110_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h4)
	) name2600 (
		_w2667_,
		_w2959_,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name2601 (
		_w2664_,
		_w2959_,
		_w3114_
	);
	LUT2 #(
		.INIT('h1)
	) name2602 (
		_w3113_,
		_w3114_,
		_w3115_
	);
	LUT2 #(
		.INIT('h4)
	) name2603 (
		_w2716_,
		_w2959_,
		_w3116_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w2719_,
		_w2959_,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name2605 (
		_w3116_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h4)
	) name2606 (
		_w2712_,
		_w2959_,
		_w3119_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		_w2709_,
		_w2959_,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h4)
	) name2609 (
		_w2701_,
		_w2959_,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name2610 (
		_w2704_,
		_w2959_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name2611 (
		_w3122_,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h4)
	) name2612 (
		_w2697_,
		_w2959_,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name2613 (
		_w2694_,
		_w2959_,
		_w3126_
	);
	LUT2 #(
		.INIT('h1)
	) name2614 (
		_w3125_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h4)
	) name2615 (
		_w2767_,
		_w2959_,
		_w3128_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w2764_,
		_w2959_,
		_w3129_
	);
	LUT2 #(
		.INIT('h1)
	) name2617 (
		_w3128_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h4)
	) name2618 (
		_w2781_,
		_w2959_,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name2619 (
		_w2778_,
		_w2959_,
		_w3132_
	);
	LUT2 #(
		.INIT('h1)
	) name2620 (
		_w3131_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h4)
	) name2621 (
		_w2759_,
		_w2959_,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name2622 (
		_w2756_,
		_w2959_,
		_w3135_
	);
	LUT2 #(
		.INIT('h1)
	) name2623 (
		_w3134_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h4)
	) name2624 (
		_w2752_,
		_w2959_,
		_w3137_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		_w2749_,
		_w2959_,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w3137_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h4)
	) name2627 (
		_w2774_,
		_w2959_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w2771_,
		_w2959_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name2629 (
		_w3140_,
		_w3141_,
		_w3142_
	);
	LUT2 #(
		.INIT('h4)
	) name2630 (
		_w2788_,
		_w2959_,
		_w3143_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w2785_,
		_w2959_,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		_w3143_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('h4)
	) name2633 (
		_w2792_,
		_w2959_,
		_w3146_
	);
	LUT2 #(
		.INIT('h1)
	) name2634 (
		_w2795_,
		_w2959_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name2635 (
		_w3146_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h4)
	) name2636 (
		_w2802_,
		_w2959_,
		_w3149_
	);
	LUT2 #(
		.INIT('h1)
	) name2637 (
		_w2799_,
		_w2959_,
		_w3150_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w3149_,
		_w3150_,
		_w3151_
	);
	LUT2 #(
		.INIT('h4)
	) name2639 (
		_w2168_,
		_w2959_,
		_w3152_
	);
	LUT2 #(
		.INIT('h1)
	) name2640 (
		_w2172_,
		_w2959_,
		_w3153_
	);
	LUT2 #(
		.INIT('h1)
	) name2641 (
		_w3152_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h4)
	) name2642 (
		_w2163_,
		_w2959_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name2643 (
		_w2160_,
		_w2959_,
		_w3156_
	);
	LUT2 #(
		.INIT('h1)
	) name2644 (
		_w3155_,
		_w3156_,
		_w3157_
	);
	LUT2 #(
		.INIT('h4)
	) name2645 (
		_w2152_,
		_w2959_,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name2646 (
		_w2155_,
		_w2959_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name2647 (
		_w3158_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		_w2147_,
		_w2959_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w2144_,
		_w2959_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		_w3161_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h4)
	) name2651 (
		_w2132_,
		_w2959_,
		_w3164_
	);
	LUT2 #(
		.INIT('h1)
	) name2652 (
		_w2136_,
		_w2959_,
		_w3165_
	);
	LUT2 #(
		.INIT('h1)
	) name2653 (
		_w3164_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h4)
	) name2654 (
		_w2128_,
		_w2959_,
		_w3167_
	);
	LUT2 #(
		.INIT('h1)
	) name2655 (
		_w2125_,
		_w2959_,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name2656 (
		_w3167_,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h4)
	) name2657 (
		_w2116_,
		_w2959_,
		_w3170_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w2119_,
		_w2959_,
		_w3171_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w3170_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h4)
	) name2660 (
		_w2111_,
		_w2959_,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name2661 (
		_w2108_,
		_w2959_,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name2662 (
		_w3173_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h4)
	) name2663 (
		_w2096_,
		_w2959_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w2100_,
		_w2959_,
		_w3177_
	);
	LUT2 #(
		.INIT('h1)
	) name2665 (
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w2091_,
		_w2959_,
		_w3179_
	);
	LUT2 #(
		.INIT('h1)
	) name2667 (
		_w2088_,
		_w2959_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name2668 (
		_w3179_,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h4)
	) name2669 (
		_w2080_,
		_w2959_,
		_w3182_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w2083_,
		_w2959_,
		_w3183_
	);
	LUT2 #(
		.INIT('h1)
	) name2671 (
		_w3182_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h4)
	) name2672 (
		_w2075_,
		_w2959_,
		_w3185_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		_w2072_,
		_w2959_,
		_w3186_
	);
	LUT2 #(
		.INIT('h1)
	) name2674 (
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('h4)
	) name2675 (
		_w2060_,
		_w2959_,
		_w3188_
	);
	LUT2 #(
		.INIT('h1)
	) name2676 (
		_w2064_,
		_w2959_,
		_w3189_
	);
	LUT2 #(
		.INIT('h1)
	) name2677 (
		_w3188_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h4)
	) name2678 (
		_w2056_,
		_w2959_,
		_w3191_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w2053_,
		_w2959_,
		_w3192_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w3191_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h4)
	) name2681 (
		_w2044_,
		_w2959_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name2682 (
		_w2047_,
		_w2959_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name2683 (
		_w3194_,
		_w3195_,
		_w3196_
	);
	LUT2 #(
		.INIT('h4)
	) name2684 (
		_w2039_,
		_w2959_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w2036_,
		_w2959_,
		_w3198_
	);
	LUT2 #(
		.INIT('h1)
	) name2686 (
		_w3197_,
		_w3198_,
		_w3199_
	);
	LUT2 #(
		.INIT('h4)
	) name2687 (
		_w2024_,
		_w2959_,
		_w3200_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w2028_,
		_w2959_,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name2689 (
		_w3200_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h4)
	) name2690 (
		_w2019_,
		_w2959_,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name2691 (
		_w2016_,
		_w2959_,
		_w3204_
	);
	LUT2 #(
		.INIT('h1)
	) name2692 (
		_w3203_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h4)
	) name2693 (
		_w2008_,
		_w2959_,
		_w3206_
	);
	LUT2 #(
		.INIT('h1)
	) name2694 (
		_w2011_,
		_w2959_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2695 (
		_w3206_,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h4)
	) name2696 (
		_w2003_,
		_w2959_,
		_w3209_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w2000_,
		_w2959_,
		_w3210_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		_w3209_,
		_w3210_,
		_w3211_
	);
	LUT2 #(
		.INIT('h4)
	) name2699 (
		_w1988_,
		_w2959_,
		_w3212_
	);
	LUT2 #(
		.INIT('h1)
	) name2700 (
		_w1992_,
		_w2959_,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name2701 (
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT2 #(
		.INIT('h4)
	) name2702 (
		_w1984_,
		_w2959_,
		_w3215_
	);
	LUT2 #(
		.INIT('h1)
	) name2703 (
		_w1981_,
		_w2959_,
		_w3216_
	);
	LUT2 #(
		.INIT('h1)
	) name2704 (
		_w3215_,
		_w3216_,
		_w3217_
	);
	LUT2 #(
		.INIT('h4)
	) name2705 (
		_w1972_,
		_w2959_,
		_w3218_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w1975_,
		_w2959_,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w3218_,
		_w3219_,
		_w3220_
	);
	LUT2 #(
		.INIT('h4)
	) name2708 (
		_w1967_,
		_w2959_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w1964_,
		_w2959_,
		_w3222_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w3221_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h4)
	) name2711 (
		_w1952_,
		_w2959_,
		_w3224_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		_w1956_,
		_w2959_,
		_w3225_
	);
	LUT2 #(
		.INIT('h1)
	) name2713 (
		_w3224_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		_w1947_,
		_w2959_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w1944_,
		_w2959_,
		_w3228_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		_w3227_,
		_w3228_,
		_w3229_
	);
	LUT2 #(
		.INIT('h4)
	) name2717 (
		_w1936_,
		_w2959_,
		_w3230_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w1939_,
		_w2959_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name2719 (
		_w3230_,
		_w3231_,
		_w3232_
	);
	LUT2 #(
		.INIT('h4)
	) name2720 (
		_w1931_,
		_w2959_,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name2721 (
		_w1928_,
		_w2959_,
		_w3234_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w3233_,
		_w3234_,
		_w3235_
	);
	LUT2 #(
		.INIT('h4)
	) name2723 (
		_w1916_,
		_w2959_,
		_w3236_
	);
	LUT2 #(
		.INIT('h1)
	) name2724 (
		_w1920_,
		_w2959_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		_w3236_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h4)
	) name2726 (
		_w1912_,
		_w2959_,
		_w3239_
	);
	LUT2 #(
		.INIT('h1)
	) name2727 (
		_w1909_,
		_w2959_,
		_w3240_
	);
	LUT2 #(
		.INIT('h1)
	) name2728 (
		_w3239_,
		_w3240_,
		_w3241_
	);
	LUT2 #(
		.INIT('h4)
	) name2729 (
		_w1900_,
		_w2959_,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name2730 (
		_w1903_,
		_w2959_,
		_w3243_
	);
	LUT2 #(
		.INIT('h1)
	) name2731 (
		_w3242_,
		_w3243_,
		_w3244_
	);
	LUT2 #(
		.INIT('h4)
	) name2732 (
		_w1895_,
		_w2959_,
		_w3245_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w1892_,
		_w2959_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name2734 (
		_w3245_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		_w1880_,
		_w2959_,
		_w3248_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w1884_,
		_w2959_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name2737 (
		_w3248_,
		_w3249_,
		_w3250_
	);
	LUT2 #(
		.INIT('h4)
	) name2738 (
		_w1875_,
		_w2959_,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		_w1872_,
		_w2959_,
		_w3252_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		_w3251_,
		_w3252_,
		_w3253_
	);
	LUT2 #(
		.INIT('h4)
	) name2741 (
		_w1864_,
		_w2959_,
		_w3254_
	);
	LUT2 #(
		.INIT('h1)
	) name2742 (
		_w1867_,
		_w2959_,
		_w3255_
	);
	LUT2 #(
		.INIT('h1)
	) name2743 (
		_w3254_,
		_w3255_,
		_w3256_
	);
	LUT2 #(
		.INIT('h4)
	) name2744 (
		_w1859_,
		_w2959_,
		_w3257_
	);
	LUT2 #(
		.INIT('h1)
	) name2745 (
		_w1856_,
		_w2959_,
		_w3258_
	);
	LUT2 #(
		.INIT('h1)
	) name2746 (
		_w3257_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('h4)
	) name2747 (
		_w1844_,
		_w2959_,
		_w3260_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w1848_,
		_w2959_,
		_w3261_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w3260_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h4)
	) name2750 (
		_w1840_,
		_w2959_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w1837_,
		_w2959_,
		_w3264_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w3263_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h4)
	) name2753 (
		_w1828_,
		_w2959_,
		_w3266_
	);
	LUT2 #(
		.INIT('h1)
	) name2754 (
		_w1831_,
		_w2959_,
		_w3267_
	);
	LUT2 #(
		.INIT('h1)
	) name2755 (
		_w3266_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h4)
	) name2756 (
		_w1823_,
		_w2959_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w1820_,
		_w2959_,
		_w3270_
	);
	LUT2 #(
		.INIT('h1)
	) name2758 (
		_w3269_,
		_w3270_,
		_w3271_
	);
	LUT2 #(
		.INIT('h4)
	) name2759 (
		_w1808_,
		_w2959_,
		_w3272_
	);
	LUT2 #(
		.INIT('h1)
	) name2760 (
		_w1812_,
		_w2959_,
		_w3273_
	);
	LUT2 #(
		.INIT('h1)
	) name2761 (
		_w3272_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h4)
	) name2762 (
		_w1803_,
		_w2959_,
		_w3275_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w1800_,
		_w2959_,
		_w3276_
	);
	LUT2 #(
		.INIT('h1)
	) name2764 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h4)
	) name2765 (
		_w1792_,
		_w2959_,
		_w3278_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		_w1795_,
		_w2959_,
		_w3279_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		_w3278_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h4)
	) name2768 (
		_w1787_,
		_w2959_,
		_w3281_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		_w1784_,
		_w2959_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name2770 (
		_w3281_,
		_w3282_,
		_w3283_
	);
	LUT2 #(
		.INIT('h4)
	) name2771 (
		_w1772_,
		_w2959_,
		_w3284_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w1776_,
		_w2959_,
		_w3285_
	);
	LUT2 #(
		.INIT('h1)
	) name2773 (
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h4)
	) name2774 (
		_w1768_,
		_w2959_,
		_w3287_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		_w1765_,
		_w2959_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name2776 (
		_w3287_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('h4)
	) name2777 (
		_w1756_,
		_w2959_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		_w1759_,
		_w2959_,
		_w3291_
	);
	LUT2 #(
		.INIT('h1)
	) name2779 (
		_w3290_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h4)
	) name2780 (
		_w1751_,
		_w2959_,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		_w1748_,
		_w2959_,
		_w3294_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		_w3293_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h4)
	) name2783 (
		_w1736_,
		_w2959_,
		_w3296_
	);
	LUT2 #(
		.INIT('h1)
	) name2784 (
		_w1740_,
		_w2959_,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w3296_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h4)
	) name2786 (
		_w1731_,
		_w2959_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name2787 (
		_w1728_,
		_w2959_,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w3299_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h4)
	) name2789 (
		_w1720_,
		_w2959_,
		_w3302_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		_w1723_,
		_w2959_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h4)
	) name2792 (
		_w1715_,
		_w2959_,
		_w3305_
	);
	LUT2 #(
		.INIT('h1)
	) name2793 (
		_w1712_,
		_w2959_,
		_w3306_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		_w3305_,
		_w3306_,
		_w3307_
	);
	LUT2 #(
		.INIT('h4)
	) name2795 (
		_w1700_,
		_w2959_,
		_w3308_
	);
	LUT2 #(
		.INIT('h1)
	) name2796 (
		_w1704_,
		_w2959_,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w3308_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h4)
	) name2798 (
		_w1696_,
		_w2959_,
		_w3311_
	);
	LUT2 #(
		.INIT('h1)
	) name2799 (
		_w1693_,
		_w2959_,
		_w3312_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w3311_,
		_w3312_,
		_w3313_
	);
	LUT2 #(
		.INIT('h4)
	) name2801 (
		_w1684_,
		_w2959_,
		_w3314_
	);
	LUT2 #(
		.INIT('h1)
	) name2802 (
		_w1687_,
		_w2959_,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name2803 (
		_w3314_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h4)
	) name2804 (
		_w1679_,
		_w2959_,
		_w3317_
	);
	LUT2 #(
		.INIT('h1)
	) name2805 (
		_w1676_,
		_w2959_,
		_w3318_
	);
	LUT2 #(
		.INIT('h1)
	) name2806 (
		_w3317_,
		_w3318_,
		_w3319_
	);
	LUT2 #(
		.INIT('h4)
	) name2807 (
		_w1664_,
		_w2959_,
		_w3320_
	);
	LUT2 #(
		.INIT('h1)
	) name2808 (
		_w1668_,
		_w2959_,
		_w3321_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w3320_,
		_w3321_,
		_w3322_
	);
	LUT2 #(
		.INIT('h4)
	) name2810 (
		_w1659_,
		_w2959_,
		_w3323_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w1656_,
		_w2959_,
		_w3324_
	);
	LUT2 #(
		.INIT('h1)
	) name2812 (
		_w3323_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h4)
	) name2813 (
		_w1648_,
		_w2959_,
		_w3326_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		_w1651_,
		_w2959_,
		_w3327_
	);
	LUT2 #(
		.INIT('h1)
	) name2815 (
		_w3326_,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h4)
	) name2816 (
		_w1643_,
		_w2959_,
		_w3329_
	);
	LUT2 #(
		.INIT('h1)
	) name2817 (
		_w1640_,
		_w2959_,
		_w3330_
	);
	LUT2 #(
		.INIT('h1)
	) name2818 (
		_w3329_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h4)
	) name2819 (
		_w2945_,
		_w2959_,
		_w3332_
	);
	LUT2 #(
		.INIT('h1)
	) name2820 (
		_w2942_,
		_w2959_,
		_w3333_
	);
	LUT2 #(
		.INIT('h1)
	) name2821 (
		_w3332_,
		_w3333_,
		_w3334_
	);
	LUT2 #(
		.INIT('h4)
	) name2822 (
		_w2937_,
		_w2959_,
		_w3335_
	);
	LUT2 #(
		.INIT('h1)
	) name2823 (
		_w2934_,
		_w2959_,
		_w3336_
	);
	LUT2 #(
		.INIT('h1)
	) name2824 (
		_w3335_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('h4)
	) name2825 (
		_w2930_,
		_w2959_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w2927_,
		_w2959_,
		_w3339_
	);
	LUT2 #(
		.INIT('h1)
	) name2827 (
		_w3338_,
		_w3339_,
		_w3340_
	);
	LUT2 #(
		.INIT('h8)
	) name2828 (
		_w2922_,
		_w2923_,
		_w3341_
	);
	LUT2 #(
		.INIT('h2)
	) name2829 (
		_w1637_,
		_w2959_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name2830 (
		_w1073_,
		_w2959_,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		_w3342_,
		_w3343_,
		_w3344_
	);
	assign \result[0]  = _w2962_ ;
	assign \result[1]  = _w2965_ ;
	assign \result[2]  = _w2968_ ;
	assign \result[3]  = _w2971_ ;
	assign \result[4]  = _w2974_ ;
	assign \result[5]  = _w2977_ ;
	assign \result[6]  = _w2980_ ;
	assign \result[7]  = _w2983_ ;
	assign \result[8]  = _w2986_ ;
	assign \result[9]  = _w2989_ ;
	assign \result[10]  = _w2992_ ;
	assign \result[11]  = _w2995_ ;
	assign \result[12]  = _w2998_ ;
	assign \result[13]  = _w3001_ ;
	assign \result[14]  = _w3004_ ;
	assign \result[15]  = _w3007_ ;
	assign \result[16]  = _w3010_ ;
	assign \result[17]  = _w3013_ ;
	assign \result[18]  = _w3016_ ;
	assign \result[19]  = _w3019_ ;
	assign \result[20]  = _w3022_ ;
	assign \result[21]  = _w3025_ ;
	assign \result[22]  = _w3028_ ;
	assign \result[23]  = _w3031_ ;
	assign \result[24]  = _w3034_ ;
	assign \result[25]  = _w3037_ ;
	assign \result[26]  = _w3040_ ;
	assign \result[27]  = _w3043_ ;
	assign \result[28]  = _w3046_ ;
	assign \result[29]  = _w3049_ ;
	assign \result[30]  = _w3052_ ;
	assign \result[31]  = _w3055_ ;
	assign \result[32]  = _w3058_ ;
	assign \result[33]  = _w3061_ ;
	assign \result[34]  = _w3064_ ;
	assign \result[35]  = _w3067_ ;
	assign \result[36]  = _w3070_ ;
	assign \result[37]  = _w3073_ ;
	assign \result[38]  = _w3076_ ;
	assign \result[39]  = _w3079_ ;
	assign \result[40]  = _w3082_ ;
	assign \result[41]  = _w3085_ ;
	assign \result[42]  = _w3088_ ;
	assign \result[43]  = _w3091_ ;
	assign \result[44]  = _w3094_ ;
	assign \result[45]  = _w3097_ ;
	assign \result[46]  = _w3100_ ;
	assign \result[47]  = _w3103_ ;
	assign \result[48]  = _w3106_ ;
	assign \result[49]  = _w3109_ ;
	assign \result[50]  = _w3112_ ;
	assign \result[51]  = _w3115_ ;
	assign \result[52]  = _w3118_ ;
	assign \result[53]  = _w3121_ ;
	assign \result[54]  = _w3124_ ;
	assign \result[55]  = _w3127_ ;
	assign \result[56]  = _w3130_ ;
	assign \result[57]  = _w3133_ ;
	assign \result[58]  = _w3136_ ;
	assign \result[59]  = _w3139_ ;
	assign \result[60]  = _w3142_ ;
	assign \result[61]  = _w3145_ ;
	assign \result[62]  = _w3148_ ;
	assign \result[63]  = _w3151_ ;
	assign \result[64]  = _w3154_ ;
	assign \result[65]  = _w3157_ ;
	assign \result[66]  = _w3160_ ;
	assign \result[67]  = _w3163_ ;
	assign \result[68]  = _w3166_ ;
	assign \result[69]  = _w3169_ ;
	assign \result[70]  = _w3172_ ;
	assign \result[71]  = _w3175_ ;
	assign \result[72]  = _w3178_ ;
	assign \result[73]  = _w3181_ ;
	assign \result[74]  = _w3184_ ;
	assign \result[75]  = _w3187_ ;
	assign \result[76]  = _w3190_ ;
	assign \result[77]  = _w3193_ ;
	assign \result[78]  = _w3196_ ;
	assign \result[79]  = _w3199_ ;
	assign \result[80]  = _w3202_ ;
	assign \result[81]  = _w3205_ ;
	assign \result[82]  = _w3208_ ;
	assign \result[83]  = _w3211_ ;
	assign \result[84]  = _w3214_ ;
	assign \result[85]  = _w3217_ ;
	assign \result[86]  = _w3220_ ;
	assign \result[87]  = _w3223_ ;
	assign \result[88]  = _w3226_ ;
	assign \result[89]  = _w3229_ ;
	assign \result[90]  = _w3232_ ;
	assign \result[91]  = _w3235_ ;
	assign \result[92]  = _w3238_ ;
	assign \result[93]  = _w3241_ ;
	assign \result[94]  = _w3244_ ;
	assign \result[95]  = _w3247_ ;
	assign \result[96]  = _w3250_ ;
	assign \result[97]  = _w3253_ ;
	assign \result[98]  = _w3256_ ;
	assign \result[99]  = _w3259_ ;
	assign \result[100]  = _w3262_ ;
	assign \result[101]  = _w3265_ ;
	assign \result[102]  = _w3268_ ;
	assign \result[103]  = _w3271_ ;
	assign \result[104]  = _w3274_ ;
	assign \result[105]  = _w3277_ ;
	assign \result[106]  = _w3280_ ;
	assign \result[107]  = _w3283_ ;
	assign \result[108]  = _w3286_ ;
	assign \result[109]  = _w3289_ ;
	assign \result[110]  = _w3292_ ;
	assign \result[111]  = _w3295_ ;
	assign \result[112]  = _w3298_ ;
	assign \result[113]  = _w3301_ ;
	assign \result[114]  = _w3304_ ;
	assign \result[115]  = _w3307_ ;
	assign \result[116]  = _w3310_ ;
	assign \result[117]  = _w3313_ ;
	assign \result[118]  = _w3316_ ;
	assign \result[119]  = _w3319_ ;
	assign \result[120]  = _w3322_ ;
	assign \result[121]  = _w3325_ ;
	assign \result[122]  = _w3328_ ;
	assign \result[123]  = _w3331_ ;
	assign \result[124]  = _w3334_ ;
	assign \result[125]  = _w3337_ ;
	assign \result[126]  = _w3340_ ;
	assign \result[127]  = _w3341_ ;
	assign \address[0]  = _w3344_ ;
	assign \address[1]  = _w2959_ ;
endmodule;