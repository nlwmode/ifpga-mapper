module top( \106GAT(15)_pad  , \113GAT(16)_pad  , \120GAT(17)_pad  , \127GAT(18)_pad  , \134GAT(19)_pad  , \141GAT(20)_pad  , \148GAT(21)_pad  , \155GAT(22)_pad  , \15GAT(2)_pad  , \162GAT(23)_pad  , \169GAT(24)_pad  , \176GAT(25)_pad  , \183GAT(26)_pad  , \190GAT(27)_pad  , \197GAT(28)_pad  , \1GAT(0)_pad  , \204GAT(29)_pad  , \211GAT(30)_pad  , \218GAT(31)_pad  , \225GAT(32)_pad  , \226GAT(33)_pad  , \227GAT(34)_pad  , \228GAT(35)_pad  , \229GAT(36)_pad  , \22GAT(3)_pad  , \230GAT(37)_pad  , \231GAT(38)_pad  , \232GAT(39)_pad  , \233GAT(40)_pad  , \29GAT(4)_pad  , \36GAT(5)_pad  , \43GAT(6)_pad  , \50GAT(7)_pad  , \57GAT(8)_pad  , \64GAT(9)_pad  , \71GAT(10)_pad  , \78GAT(11)_pad  , \85GAT(12)_pad  , \8GAT(1)_pad  , \92GAT(13)_pad  , \99GAT(14)_pad  , \1324GAT(583)_pad  , \1325GAT(579)_pad  , \1326GAT(575)_pad  , \1327GAT(571)_pad  , \1328GAT(584)_pad  , \1329GAT(580)_pad  , \1330GAT(576)_pad  , \1331GAT(572)_pad  , \1332GAT(585)_pad  , \1333GAT(581)_pad  , \1334GAT(577)_pad  , \1335GAT(573)_pad  , \1336GAT(586)_pad  , \1337GAT(582)_pad  , \1338GAT(578)_pad  , \1339GAT(574)_pad  , \1340GAT(567)_pad  , \1341GAT(563)_pad  , \1342GAT(559)_pad  , \1343GAT(555)_pad  , \1344GAT(568)_pad  , \1345GAT(564)_pad  , \1346GAT(560)_pad  , \1347GAT(556)_pad  , \1348GAT(569)_pad  , \1349GAT(565)_pad  , \1350GAT(561)_pad  , \1351GAT(557)_pad  , \1352GAT(570)_pad  , \1353GAT(566)_pad  , \1354GAT(562)_pad  , \1355GAT(558)_pad  );
  input \106GAT(15)_pad  ;
  input \113GAT(16)_pad  ;
  input \120GAT(17)_pad  ;
  input \127GAT(18)_pad  ;
  input \134GAT(19)_pad  ;
  input \141GAT(20)_pad  ;
  input \148GAT(21)_pad  ;
  input \155GAT(22)_pad  ;
  input \15GAT(2)_pad  ;
  input \162GAT(23)_pad  ;
  input \169GAT(24)_pad  ;
  input \176GAT(25)_pad  ;
  input \183GAT(26)_pad  ;
  input \190GAT(27)_pad  ;
  input \197GAT(28)_pad  ;
  input \1GAT(0)_pad  ;
  input \204GAT(29)_pad  ;
  input \211GAT(30)_pad  ;
  input \218GAT(31)_pad  ;
  input \225GAT(32)_pad  ;
  input \226GAT(33)_pad  ;
  input \227GAT(34)_pad  ;
  input \228GAT(35)_pad  ;
  input \229GAT(36)_pad  ;
  input \22GAT(3)_pad  ;
  input \230GAT(37)_pad  ;
  input \231GAT(38)_pad  ;
  input \232GAT(39)_pad  ;
  input \233GAT(40)_pad  ;
  input \29GAT(4)_pad  ;
  input \36GAT(5)_pad  ;
  input \43GAT(6)_pad  ;
  input \50GAT(7)_pad  ;
  input \57GAT(8)_pad  ;
  input \64GAT(9)_pad  ;
  input \71GAT(10)_pad  ;
  input \78GAT(11)_pad  ;
  input \85GAT(12)_pad  ;
  input \8GAT(1)_pad  ;
  input \92GAT(13)_pad  ;
  input \99GAT(14)_pad  ;
  output \1324GAT(583)_pad  ;
  output \1325GAT(579)_pad  ;
  output \1326GAT(575)_pad  ;
  output \1327GAT(571)_pad  ;
  output \1328GAT(584)_pad  ;
  output \1329GAT(580)_pad  ;
  output \1330GAT(576)_pad  ;
  output \1331GAT(572)_pad  ;
  output \1332GAT(585)_pad  ;
  output \1333GAT(581)_pad  ;
  output \1334GAT(577)_pad  ;
  output \1335GAT(573)_pad  ;
  output \1336GAT(586)_pad  ;
  output \1337GAT(582)_pad  ;
  output \1338GAT(578)_pad  ;
  output \1339GAT(574)_pad  ;
  output \1340GAT(567)_pad  ;
  output \1341GAT(563)_pad  ;
  output \1342GAT(559)_pad  ;
  output \1343GAT(555)_pad  ;
  output \1344GAT(568)_pad  ;
  output \1345GAT(564)_pad  ;
  output \1346GAT(560)_pad  ;
  output \1347GAT(556)_pad  ;
  output \1348GAT(569)_pad  ;
  output \1349GAT(565)_pad  ;
  output \1350GAT(561)_pad  ;
  output \1351GAT(557)_pad  ;
  output \1352GAT(570)_pad  ;
  output \1353GAT(566)_pad  ;
  output \1354GAT(562)_pad  ;
  output \1355GAT(558)_pad  ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 ;
  assign n42 = ~\176GAT(25)_pad  & ~\183GAT(26)_pad  ;
  assign n43 = \176GAT(25)_pad  & \183GAT(26)_pad  ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = \169GAT(24)_pad  & ~\190GAT(27)_pad  ;
  assign n46 = ~\169GAT(24)_pad  & \190GAT(27)_pad  ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = n44 & n47 ;
  assign n49 = ~n44 & ~n47 ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = \226GAT(33)_pad  & \233GAT(40)_pad  ;
  assign n52 = \64GAT(9)_pad  & ~n51 ;
  assign n53 = ~\64GAT(9)_pad  & n51 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = \36GAT(5)_pad  & ~\8GAT(1)_pad  ;
  assign n56 = ~\36GAT(5)_pad  & \8GAT(1)_pad  ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = n54 & n57 ;
  assign n59 = ~n50 & n58 ;
  assign n60 = ~n54 & n57 ;
  assign n61 = n50 & n60 ;
  assign n62 = ~n59 & ~n61 ;
  assign n63 = ~n54 & ~n57 ;
  assign n64 = ~n50 & n63 ;
  assign n65 = n54 & ~n57 ;
  assign n66 = n50 & n65 ;
  assign n67 = ~n64 & ~n66 ;
  assign n68 = n62 & n67 ;
  assign n69 = \197GAT(28)_pad  & ~\218GAT(31)_pad  ;
  assign n70 = ~\197GAT(28)_pad  & \218GAT(31)_pad  ;
  assign n71 = ~n69 & ~n70 ;
  assign n72 = \204GAT(29)_pad  & ~\211GAT(30)_pad  ;
  assign n73 = ~\204GAT(29)_pad  & \211GAT(30)_pad  ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = n71 & n74 ;
  assign n76 = ~n71 & ~n74 ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = \92GAT(13)_pad  & ~n77 ;
  assign n79 = ~\92GAT(13)_pad  & n77 ;
  assign n80 = ~n78 & ~n79 ;
  assign n81 = n68 & n80 ;
  assign n82 = ~n68 & ~n80 ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = ~\120GAT(17)_pad  & ~\127GAT(18)_pad  ;
  assign n85 = \120GAT(17)_pad  & \127GAT(18)_pad  ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = \113GAT(16)_pad  & ~\134GAT(19)_pad  ;
  assign n88 = ~\113GAT(16)_pad  & \134GAT(19)_pad  ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = n86 & n89 ;
  assign n91 = ~n86 & ~n89 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = ~n50 & n92 ;
  assign n94 = n50 & ~n92 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = \227GAT(34)_pad  & \233GAT(40)_pad  ;
  assign n97 = \15GAT(2)_pad  & ~\43GAT(6)_pad  ;
  assign n98 = ~\15GAT(2)_pad  & \43GAT(6)_pad  ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = n96 & n99 ;
  assign n101 = ~n96 & ~n99 ;
  assign n102 = ~n100 & ~n101 ;
  assign n103 = \71GAT(10)_pad  & ~\99GAT(14)_pad  ;
  assign n104 = ~\71GAT(10)_pad  & \99GAT(14)_pad  ;
  assign n105 = ~n103 & ~n104 ;
  assign n106 = n102 & ~n105 ;
  assign n107 = ~n102 & n105 ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = n95 & n108 ;
  assign n110 = ~n95 & ~n108 ;
  assign n111 = ~n109 & ~n110 ;
  assign n112 = ~n83 & n111 ;
  assign n113 = \225GAT(32)_pad  & \233GAT(40)_pad  ;
  assign n114 = \57GAT(8)_pad  & ~n113 ;
  assign n115 = ~\57GAT(8)_pad  & n113 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = \1GAT(0)_pad  & ~\29GAT(4)_pad  ;
  assign n118 = ~\1GAT(0)_pad  & \29GAT(4)_pad  ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = n116 & n119 ;
  assign n121 = ~n92 & n120 ;
  assign n122 = ~n116 & n119 ;
  assign n123 = n92 & n122 ;
  assign n124 = ~n121 & ~n123 ;
  assign n125 = ~n116 & ~n119 ;
  assign n126 = ~n92 & n125 ;
  assign n127 = n116 & ~n119 ;
  assign n128 = n92 & n127 ;
  assign n129 = ~n126 & ~n128 ;
  assign n130 = n124 & n129 ;
  assign n131 = ~\148GAT(21)_pad  & ~\155GAT(22)_pad  ;
  assign n132 = \148GAT(21)_pad  & \155GAT(22)_pad  ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = \141GAT(20)_pad  & ~\162GAT(23)_pad  ;
  assign n135 = ~\141GAT(20)_pad  & \162GAT(23)_pad  ;
  assign n136 = ~n134 & ~n135 ;
  assign n137 = n133 & n136 ;
  assign n138 = ~n133 & ~n136 ;
  assign n139 = ~n137 & ~n138 ;
  assign n140 = \85GAT(12)_pad  & ~n139 ;
  assign n141 = ~\85GAT(12)_pad  & n139 ;
  assign n142 = ~n140 & ~n141 ;
  assign n143 = n130 & n142 ;
  assign n144 = ~n130 & ~n142 ;
  assign n145 = ~n143 & ~n144 ;
  assign n146 = \228GAT(35)_pad  & \233GAT(40)_pad  ;
  assign n147 = n139 & n146 ;
  assign n148 = ~n139 & ~n146 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = ~\106GAT(15)_pad  & ~\78GAT(11)_pad  ;
  assign n151 = \106GAT(15)_pad  & \78GAT(11)_pad  ;
  assign n152 = ~n150 & ~n151 ;
  assign n153 = \22GAT(3)_pad  & ~\50GAT(7)_pad  ;
  assign n154 = ~\22GAT(3)_pad  & \50GAT(7)_pad  ;
  assign n155 = ~n153 & ~n154 ;
  assign n156 = n152 & n155 ;
  assign n157 = ~n152 & ~n155 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = n77 & ~n158 ;
  assign n160 = ~n149 & n159 ;
  assign n161 = n77 & n158 ;
  assign n162 = n149 & n161 ;
  assign n163 = ~n160 & ~n162 ;
  assign n164 = ~n77 & n158 ;
  assign n165 = ~n149 & n164 ;
  assign n166 = ~n77 & ~n158 ;
  assign n167 = n149 & n166 ;
  assign n168 = ~n165 & ~n167 ;
  assign n169 = n163 & n168 ;
  assign n170 = n145 & n169 ;
  assign n171 = n112 & n170 ;
  assign n172 = ~n83 & ~n111 ;
  assign n173 = ~n145 & n169 ;
  assign n174 = n172 & n173 ;
  assign n175 = n83 & ~n111 ;
  assign n176 = n170 & n175 ;
  assign n177 = ~n174 & ~n176 ;
  assign n178 = ~n171 & n177 ;
  assign n179 = ~n83 & n145 ;
  assign n180 = ~n111 & ~n169 ;
  assign n181 = n179 & n180 ;
  assign n182 = n178 & ~n181 ;
  assign n183 = ~\106GAT(15)_pad  & ~\99GAT(14)_pad  ;
  assign n184 = \106GAT(15)_pad  & \99GAT(14)_pad  ;
  assign n185 = ~n183 & ~n184 ;
  assign n186 = \85GAT(12)_pad  & ~\92GAT(13)_pad  ;
  assign n187 = ~\85GAT(12)_pad  & \92GAT(13)_pad  ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = n185 & n188 ;
  assign n190 = ~n185 & ~n188 ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = \230GAT(37)_pad  & \233GAT(40)_pad  ;
  assign n193 = ~n191 & n192 ;
  assign n194 = n191 & ~n192 ;
  assign n195 = ~n193 & ~n194 ;
  assign n196 = ~\64GAT(9)_pad  & ~\71GAT(10)_pad  ;
  assign n197 = \64GAT(9)_pad  & \71GAT(10)_pad  ;
  assign n198 = ~n196 & ~n197 ;
  assign n199 = \57GAT(8)_pad  & ~\78GAT(11)_pad  ;
  assign n200 = ~\57GAT(8)_pad  & \78GAT(11)_pad  ;
  assign n201 = ~n199 & ~n200 ;
  assign n202 = n198 & n201 ;
  assign n203 = ~n198 & ~n201 ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = ~\120GAT(17)_pad  & ~\148GAT(21)_pad  ;
  assign n206 = \120GAT(17)_pad  & \148GAT(21)_pad  ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = \176GAT(25)_pad  & ~\204GAT(29)_pad  ;
  assign n209 = ~\176GAT(25)_pad  & \204GAT(29)_pad  ;
  assign n210 = ~n208 & ~n209 ;
  assign n211 = ~n207 & ~n210 ;
  assign n212 = n204 & n211 ;
  assign n213 = n207 & ~n210 ;
  assign n214 = ~n204 & n213 ;
  assign n215 = ~n212 & ~n214 ;
  assign n216 = ~n207 & n210 ;
  assign n217 = ~n204 & n216 ;
  assign n218 = n207 & n210 ;
  assign n219 = n204 & n218 ;
  assign n220 = ~n217 & ~n219 ;
  assign n221 = n215 & n220 ;
  assign n222 = n195 & n221 ;
  assign n223 = ~n195 & ~n221 ;
  assign n224 = ~n222 & ~n223 ;
  assign n225 = ~\36GAT(5)_pad  & ~\43GAT(6)_pad  ;
  assign n226 = \36GAT(5)_pad  & \43GAT(6)_pad  ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = \29GAT(4)_pad  & ~\50GAT(7)_pad  ;
  assign n229 = ~\29GAT(4)_pad  & \50GAT(7)_pad  ;
  assign n230 = ~n228 & ~n229 ;
  assign n231 = n227 & n230 ;
  assign n232 = ~n227 & ~n230 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = \113GAT(16)_pad  & ~\141GAT(20)_pad  ;
  assign n235 = ~\113GAT(16)_pad  & \141GAT(20)_pad  ;
  assign n236 = ~n234 & ~n235 ;
  assign n237 = ~n233 & n236 ;
  assign n238 = n233 & ~n236 ;
  assign n239 = ~n237 & ~n238 ;
  assign n240 = ~\1GAT(0)_pad  & ~\22GAT(3)_pad  ;
  assign n241 = \1GAT(0)_pad  & \22GAT(3)_pad  ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = \15GAT(2)_pad  & ~\8GAT(1)_pad  ;
  assign n244 = ~\15GAT(2)_pad  & \8GAT(1)_pad  ;
  assign n245 = ~n243 & ~n244 ;
  assign n246 = n242 & n245 ;
  assign n247 = ~n242 & ~n245 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = \229GAT(36)_pad  & \233GAT(40)_pad  ;
  assign n250 = \169GAT(24)_pad  & ~\197GAT(28)_pad  ;
  assign n251 = ~\169GAT(24)_pad  & \197GAT(28)_pad  ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = ~n249 & ~n252 ;
  assign n254 = n248 & n253 ;
  assign n255 = n249 & ~n252 ;
  assign n256 = ~n248 & n255 ;
  assign n257 = ~n254 & ~n256 ;
  assign n258 = ~n249 & n252 ;
  assign n259 = ~n248 & n258 ;
  assign n260 = n249 & n252 ;
  assign n261 = n248 & n260 ;
  assign n262 = ~n259 & ~n261 ;
  assign n263 = n257 & n262 ;
  assign n264 = n239 & n263 ;
  assign n265 = ~n239 & ~n263 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n224 & n266 ;
  assign n268 = \232GAT(39)_pad  & \233GAT(40)_pad  ;
  assign n269 = n191 & n268 ;
  assign n270 = ~n191 & ~n268 ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = ~\134GAT(19)_pad  & ~\162GAT(23)_pad  ;
  assign n273 = \134GAT(19)_pad  & \162GAT(23)_pad  ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = \190GAT(27)_pad  & ~\218GAT(31)_pad  ;
  assign n276 = ~\190GAT(27)_pad  & \218GAT(31)_pad  ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = n274 & n277 ;
  assign n279 = ~n274 & ~n277 ;
  assign n280 = ~n278 & ~n279 ;
  assign n281 = n233 & ~n280 ;
  assign n282 = ~n271 & n281 ;
  assign n283 = n233 & n280 ;
  assign n284 = n271 & n283 ;
  assign n285 = ~n282 & ~n284 ;
  assign n286 = ~n233 & n280 ;
  assign n287 = ~n271 & n286 ;
  assign n288 = ~n233 & ~n280 ;
  assign n289 = n271 & n288 ;
  assign n290 = ~n287 & ~n289 ;
  assign n291 = n285 & n290 ;
  assign n292 = \231GAT(38)_pad  & \233GAT(40)_pad  ;
  assign n293 = n204 & n292 ;
  assign n294 = ~n204 & ~n292 ;
  assign n295 = ~n293 & ~n294 ;
  assign n296 = ~\127GAT(18)_pad  & ~\155GAT(22)_pad  ;
  assign n297 = \127GAT(18)_pad  & \155GAT(22)_pad  ;
  assign n298 = ~n296 & ~n297 ;
  assign n299 = \183GAT(26)_pad  & ~\211GAT(30)_pad  ;
  assign n300 = ~\183GAT(26)_pad  & \211GAT(30)_pad  ;
  assign n301 = ~n299 & ~n300 ;
  assign n302 = n298 & ~n301 ;
  assign n303 = ~n298 & n301 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = ~n248 & n304 ;
  assign n306 = ~n295 & n305 ;
  assign n307 = n248 & n304 ;
  assign n308 = n295 & n307 ;
  assign n309 = ~n306 & ~n308 ;
  assign n310 = n248 & ~n304 ;
  assign n311 = ~n295 & n310 ;
  assign n312 = ~n248 & ~n304 ;
  assign n313 = n295 & n312 ;
  assign n314 = ~n311 & ~n313 ;
  assign n315 = n309 & n314 ;
  assign n316 = ~n291 & ~n315 ;
  assign n317 = ~n145 & n316 ;
  assign n318 = n267 & n317 ;
  assign n319 = ~n182 & n318 ;
  assign n320 = \1GAT(0)_pad  & ~n319 ;
  assign n321 = ~\1GAT(0)_pad  & n319 ;
  assign n322 = ~n320 & ~n321 ;
  assign n323 = n83 & n316 ;
  assign n324 = n267 & n323 ;
  assign n325 = ~n182 & n324 ;
  assign n326 = \8GAT(1)_pad  & ~n325 ;
  assign n327 = ~\8GAT(1)_pad  & n325 ;
  assign n328 = ~n326 & ~n327 ;
  assign n329 = n111 & n316 ;
  assign n330 = n267 & n329 ;
  assign n331 = ~n182 & n330 ;
  assign n332 = \15GAT(2)_pad  & ~n331 ;
  assign n333 = ~\15GAT(2)_pad  & n331 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = ~n169 & n316 ;
  assign n336 = n267 & n335 ;
  assign n337 = ~n182 & n336 ;
  assign n338 = \22GAT(3)_pad  & ~n337 ;
  assign n339 = ~\22GAT(3)_pad  & n337 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = n267 & n315 ;
  assign n342 = ~n145 & n291 ;
  assign n343 = n341 & n342 ;
  assign n344 = ~n182 & n343 ;
  assign n345 = \29GAT(4)_pad  & ~n344 ;
  assign n346 = ~\29GAT(4)_pad  & n344 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = n83 & n291 ;
  assign n349 = n341 & n348 ;
  assign n350 = ~n182 & n349 ;
  assign n351 = \36GAT(5)_pad  & ~n350 ;
  assign n352 = ~\36GAT(5)_pad  & n350 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = n111 & n291 ;
  assign n355 = n341 & n354 ;
  assign n356 = ~n182 & n355 ;
  assign n357 = \43GAT(6)_pad  & ~n356 ;
  assign n358 = ~\43GAT(6)_pad  & n356 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = ~n169 & n291 ;
  assign n361 = n341 & n360 ;
  assign n362 = ~n182 & n361 ;
  assign n363 = \50GAT(7)_pad  & ~n362 ;
  assign n364 = ~\50GAT(7)_pad  & n362 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = ~n224 & ~n266 ;
  assign n367 = n317 & n366 ;
  assign n368 = ~n182 & n367 ;
  assign n369 = \57GAT(8)_pad  & ~n368 ;
  assign n370 = ~\57GAT(8)_pad  & n368 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = n323 & n366 ;
  assign n373 = ~n182 & n372 ;
  assign n374 = \64GAT(9)_pad  & ~n373 ;
  assign n375 = ~\64GAT(9)_pad  & n373 ;
  assign n376 = ~n374 & ~n375 ;
  assign n377 = n329 & n366 ;
  assign n378 = ~n182 & n377 ;
  assign n379 = \71GAT(10)_pad  & ~n378 ;
  assign n380 = ~\71GAT(10)_pad  & n378 ;
  assign n381 = ~n379 & ~n380 ;
  assign n382 = n335 & n366 ;
  assign n383 = ~n182 & n382 ;
  assign n384 = \78GAT(11)_pad  & ~n383 ;
  assign n385 = ~\78GAT(11)_pad  & n383 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = n315 & n366 ;
  assign n388 = n342 & n387 ;
  assign n389 = ~n182 & n388 ;
  assign n390 = \85GAT(12)_pad  & ~n389 ;
  assign n391 = ~\85GAT(12)_pad  & n389 ;
  assign n392 = ~n390 & ~n391 ;
  assign n393 = n348 & n387 ;
  assign n394 = ~n182 & n393 ;
  assign n395 = \92GAT(13)_pad  & ~n394 ;
  assign n396 = ~\92GAT(13)_pad  & n394 ;
  assign n397 = ~n395 & ~n396 ;
  assign n398 = n354 & n387 ;
  assign n399 = ~n182 & n398 ;
  assign n400 = \99GAT(14)_pad  & ~n399 ;
  assign n401 = ~\99GAT(14)_pad  & n399 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = n360 & n387 ;
  assign n404 = ~n182 & n403 ;
  assign n405 = \106GAT(15)_pad  & ~n404 ;
  assign n406 = ~\106GAT(15)_pad  & n404 ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = n224 & ~n291 ;
  assign n409 = n266 & n315 ;
  assign n410 = n408 & n409 ;
  assign n411 = ~n266 & n315 ;
  assign n412 = ~n224 & ~n291 ;
  assign n413 = n411 & n412 ;
  assign n414 = ~n266 & ~n315 ;
  assign n415 = n408 & n414 ;
  assign n416 = ~n413 & ~n415 ;
  assign n417 = ~n410 & n416 ;
  assign n418 = n224 & ~n266 ;
  assign n419 = n291 & n315 ;
  assign n420 = n418 & n419 ;
  assign n421 = n417 & ~n420 ;
  assign n422 = n111 & n169 ;
  assign n423 = ~n83 & ~n145 ;
  assign n424 = n266 & n423 ;
  assign n425 = n422 & n424 ;
  assign n426 = ~n421 & n425 ;
  assign n427 = \113GAT(16)_pad  & ~n426 ;
  assign n428 = ~\113GAT(16)_pad  & n426 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = ~n224 & n423 ;
  assign n431 = n422 & n430 ;
  assign n432 = ~n421 & n431 ;
  assign n433 = \120GAT(17)_pad  & ~n432 ;
  assign n434 = ~\120GAT(17)_pad  & n432 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = ~n315 & n423 ;
  assign n437 = n422 & n436 ;
  assign n438 = ~n421 & n437 ;
  assign n439 = \127GAT(18)_pad  & ~n438 ;
  assign n440 = ~\127GAT(18)_pad  & n438 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = n291 & n423 ;
  assign n443 = n422 & n442 ;
  assign n444 = ~n421 & n443 ;
  assign n445 = \134GAT(19)_pad  & ~n444 ;
  assign n446 = ~\134GAT(19)_pad  & n444 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = ~n111 & n423 ;
  assign n449 = ~n169 & n266 ;
  assign n450 = n448 & n449 ;
  assign n451 = ~n421 & n450 ;
  assign n452 = \141GAT(20)_pad  & ~n451 ;
  assign n453 = ~\141GAT(20)_pad  & n451 ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = ~n169 & ~n224 ;
  assign n456 = n448 & n455 ;
  assign n457 = ~n421 & n456 ;
  assign n458 = \148GAT(21)_pad  & ~n457 ;
  assign n459 = ~\148GAT(21)_pad  & n457 ;
  assign n460 = ~n458 & ~n459 ;
  assign n461 = ~n169 & ~n315 ;
  assign n462 = n448 & n461 ;
  assign n463 = ~n421 & n462 ;
  assign n464 = \155GAT(22)_pad  & ~n463 ;
  assign n465 = ~\155GAT(22)_pad  & n463 ;
  assign n466 = ~n464 & ~n465 ;
  assign n467 = n360 & n448 ;
  assign n468 = ~n421 & n467 ;
  assign n469 = \162GAT(23)_pad  & ~n468 ;
  assign n470 = ~\162GAT(23)_pad  & n468 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = n83 & n145 ;
  assign n473 = n266 & n472 ;
  assign n474 = n422 & n473 ;
  assign n475 = ~n421 & n474 ;
  assign n476 = \169GAT(24)_pad  & ~n475 ;
  assign n477 = ~\169GAT(24)_pad  & n475 ;
  assign n478 = ~n476 & ~n477 ;
  assign n479 = ~n224 & n472 ;
  assign n480 = n422 & n479 ;
  assign n481 = ~n421 & n480 ;
  assign n482 = \176GAT(25)_pad  & ~n481 ;
  assign n483 = ~\176GAT(25)_pad  & n481 ;
  assign n484 = ~n482 & ~n483 ;
  assign n485 = ~n315 & n472 ;
  assign n486 = n422 & n485 ;
  assign n487 = ~n421 & n486 ;
  assign n488 = \183GAT(26)_pad  & ~n487 ;
  assign n489 = ~\183GAT(26)_pad  & n487 ;
  assign n490 = ~n488 & ~n489 ;
  assign n491 = n291 & n472 ;
  assign n492 = n422 & n491 ;
  assign n493 = ~n421 & n492 ;
  assign n494 = \190GAT(27)_pad  & ~n493 ;
  assign n495 = ~\190GAT(27)_pad  & n493 ;
  assign n496 = ~n494 & ~n495 ;
  assign n497 = ~n111 & n472 ;
  assign n498 = n449 & n497 ;
  assign n499 = ~n421 & n498 ;
  assign n500 = \197GAT(28)_pad  & ~n499 ;
  assign n501 = ~\197GAT(28)_pad  & n499 ;
  assign n502 = ~n500 & ~n501 ;
  assign n503 = n455 & n497 ;
  assign n504 = ~n421 & n503 ;
  assign n505 = \204GAT(29)_pad  & ~n504 ;
  assign n506 = ~\204GAT(29)_pad  & n504 ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = n461 & n497 ;
  assign n509 = ~n421 & n508 ;
  assign n510 = \211GAT(30)_pad  & ~n509 ;
  assign n511 = ~\211GAT(30)_pad  & n509 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = n360 & n497 ;
  assign n514 = ~n421 & n513 ;
  assign n515 = \218GAT(31)_pad  & ~n514 ;
  assign n516 = ~\218GAT(31)_pad  & n514 ;
  assign n517 = ~n515 & ~n516 ;
  assign \1324GAT(583)_pad  = ~n322 ;
  assign \1325GAT(579)_pad  = ~n328 ;
  assign \1326GAT(575)_pad  = ~n334 ;
  assign \1327GAT(571)_pad  = ~n340 ;
  assign \1328GAT(584)_pad  = ~n347 ;
  assign \1329GAT(580)_pad  = ~n353 ;
  assign \1330GAT(576)_pad  = ~n359 ;
  assign \1331GAT(572)_pad  = ~n365 ;
  assign \1332GAT(585)_pad  = ~n371 ;
  assign \1333GAT(581)_pad  = ~n376 ;
  assign \1334GAT(577)_pad  = ~n381 ;
  assign \1335GAT(573)_pad  = ~n386 ;
  assign \1336GAT(586)_pad  = ~n392 ;
  assign \1337GAT(582)_pad  = ~n397 ;
  assign \1338GAT(578)_pad  = ~n402 ;
  assign \1339GAT(574)_pad  = ~n407 ;
  assign \1340GAT(567)_pad  = ~n429 ;
  assign \1341GAT(563)_pad  = ~n435 ;
  assign \1342GAT(559)_pad  = ~n441 ;
  assign \1343GAT(555)_pad  = ~n447 ;
  assign \1344GAT(568)_pad  = ~n454 ;
  assign \1345GAT(564)_pad  = ~n460 ;
  assign \1346GAT(560)_pad  = ~n466 ;
  assign \1347GAT(556)_pad  = ~n471 ;
  assign \1348GAT(569)_pad  = ~n478 ;
  assign \1349GAT(565)_pad  = ~n484 ;
  assign \1350GAT(561)_pad  = ~n490 ;
  assign \1351GAT(557)_pad  = ~n496 ;
  assign \1352GAT(570)_pad  = ~n502 ;
  assign \1353GAT(566)_pad  = ~n507 ;
  assign \1354GAT(562)_pad  = ~n512 ;
  assign \1355GAT(558)_pad  = ~n517 ;
endmodule
