module top (\ccyc_addr_in[0]_pad , \ccyc_addr_in[11]_pad , \ccyc_addr_in[12]_pad , \ccyc_addr_in[13]_pad , \ccyc_addr_in[14]_pad , \ccyc_addr_in[15]_pad , \ccyc_addr_in[16]_pad , \ccyc_addr_in[17]_pad , \ccyc_addr_in[18]_pad , \ccyc_addr_in[19]_pad , \ccyc_addr_in[20]_pad , \ccyc_addr_in[21]_pad , \ccyc_addr_in[22]_pad , \ccyc_addr_in[23]_pad , \ccyc_addr_in[24]_pad , \ccyc_addr_in[25]_pad , \ccyc_addr_in[26]_pad , \ccyc_addr_in[27]_pad , \ccyc_addr_in[28]_pad , \ccyc_addr_in[29]_pad , \ccyc_addr_in[30]_pad , \ccyc_addr_in[31]_pad , \ccyc_addr_out[11]_pad , \ccyc_addr_out[12]_pad , \ccyc_addr_out[13]_pad , \ccyc_addr_out[14]_pad , \ccyc_addr_out[15]_pad , \ccyc_addr_out[16]_pad , \ccyc_addr_out[17]_pad , \ccyc_addr_out[18]_pad , \ccyc_addr_out[19]_pad , \ccyc_addr_out[20]_pad , \ccyc_addr_out[21]_pad , \ccyc_addr_out[22]_pad , \ccyc_addr_out[23]_pad , \ccyc_addr_out[24]_pad , \ccyc_addr_out[25]_pad , \ccyc_addr_out[26]_pad , \ccyc_addr_out[27]_pad , \ccyc_addr_out[28]_pad , \ccyc_addr_out[29]_pad , \ccyc_addr_out[30]_pad , \ccyc_addr_out[31]_pad );
	input \ccyc_addr_in[0]_pad  ;
	input \ccyc_addr_in[11]_pad  ;
	input \ccyc_addr_in[12]_pad  ;
	input \ccyc_addr_in[13]_pad  ;
	input \ccyc_addr_in[14]_pad  ;
	input \ccyc_addr_in[15]_pad  ;
	input \ccyc_addr_in[16]_pad  ;
	input \ccyc_addr_in[17]_pad  ;
	input \ccyc_addr_in[18]_pad  ;
	input \ccyc_addr_in[19]_pad  ;
	input \ccyc_addr_in[20]_pad  ;
	input \ccyc_addr_in[21]_pad  ;
	input \ccyc_addr_in[22]_pad  ;
	input \ccyc_addr_in[23]_pad  ;
	input \ccyc_addr_in[24]_pad  ;
	input \ccyc_addr_in[25]_pad  ;
	input \ccyc_addr_in[26]_pad  ;
	input \ccyc_addr_in[27]_pad  ;
	input \ccyc_addr_in[28]_pad  ;
	input \ccyc_addr_in[29]_pad  ;
	input \ccyc_addr_in[30]_pad  ;
	input \ccyc_addr_in[31]_pad  ;
	output \ccyc_addr_out[11]_pad  ;
	output \ccyc_addr_out[12]_pad  ;
	output \ccyc_addr_out[13]_pad  ;
	output \ccyc_addr_out[14]_pad  ;
	output \ccyc_addr_out[15]_pad  ;
	output \ccyc_addr_out[16]_pad  ;
	output \ccyc_addr_out[17]_pad  ;
	output \ccyc_addr_out[18]_pad  ;
	output \ccyc_addr_out[19]_pad  ;
	output \ccyc_addr_out[20]_pad  ;
	output \ccyc_addr_out[21]_pad  ;
	output \ccyc_addr_out[22]_pad  ;
	output \ccyc_addr_out[23]_pad  ;
	output \ccyc_addr_out[24]_pad  ;
	output \ccyc_addr_out[25]_pad  ;
	output \ccyc_addr_out[26]_pad  ;
	output \ccyc_addr_out[27]_pad  ;
	output \ccyc_addr_out[28]_pad  ;
	output \ccyc_addr_out[29]_pad  ;
	output \ccyc_addr_out[30]_pad  ;
	output \ccyc_addr_out[31]_pad  ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\ccyc_addr_in[13]_pad ,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\ccyc_addr_in[12]_pad ,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\ccyc_addr_in[0]_pad ,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		_w27_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		_w28_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w27_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w26_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\ccyc_addr_in[12]_pad ,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w26_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\ccyc_addr_in[12]_pad ,
		_w24_,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w27_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[13]_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w31_,
		_w34_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[14]_pad ,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w23_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w27_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w41_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w31_,
		_w43_,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[16]_pad ,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w23_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w27_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[17]_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w31_,
		_w50_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[18]_pad ,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		\ccyc_addr_in[13]_pad ,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		\ccyc_addr_in[12]_pad ,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w27_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[19]_pad ,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w31_,
		_w59_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[20]_pad ,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w63_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\ccyc_addr_in[12]_pad ,
		_w58_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w27_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[21]_pad ,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w31_,
		_w66_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[22]_pad ,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[23]_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w42_,
		_w57_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w27_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w73_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w31_,
		_w74_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[24]_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w77_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w49_,
		_w57_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w27_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[25]_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w81_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w31_,
		_w80_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[26]_pad ,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\ccyc_addr_in[13]_pad ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\ccyc_addr_in[12]_pad ,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w27_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[27]_pad ,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w90_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w31_,
		_w89_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[28]_pad ,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\ccyc_addr_in[12]_pad ,
		_w88_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w27_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[29]_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w97_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w31_,
		_w96_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[30]_pad ,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[31]_pad ,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w27_,
		_w42_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w87_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w103_,
		_w105_,
		_w106_
	);
	assign \ccyc_addr_out[11]_pad  = _w30_ ;
	assign \ccyc_addr_out[12]_pad  = _w33_ ;
	assign \ccyc_addr_out[13]_pad  = _w37_ ;
	assign \ccyc_addr_out[14]_pad  = _w40_ ;
	assign \ccyc_addr_out[15]_pad  = _w45_ ;
	assign \ccyc_addr_out[16]_pad  = _w48_ ;
	assign \ccyc_addr_out[17]_pad  = _w53_ ;
	assign \ccyc_addr_out[18]_pad  = _w56_ ;
	assign \ccyc_addr_out[19]_pad  = _w62_ ;
	assign \ccyc_addr_out[20]_pad  = _w65_ ;
	assign \ccyc_addr_out[21]_pad  = _w69_ ;
	assign \ccyc_addr_out[22]_pad  = _w72_ ;
	assign \ccyc_addr_out[23]_pad  = _w76_ ;
	assign \ccyc_addr_out[24]_pad  = _w79_ ;
	assign \ccyc_addr_out[25]_pad  = _w83_ ;
	assign \ccyc_addr_out[26]_pad  = _w86_ ;
	assign \ccyc_addr_out[27]_pad  = _w92_ ;
	assign \ccyc_addr_out[28]_pad  = _w95_ ;
	assign \ccyc_addr_out[29]_pad  = _w99_ ;
	assign \ccyc_addr_out[30]_pad  = _w102_ ;
	assign \ccyc_addr_out[31]_pad  = _w106_ ;
endmodule;