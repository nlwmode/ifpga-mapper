module top( a_pad , \b0_pad  , b_pad , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , f_pad , g_pad , \h0_pad  , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , o_pad , t_pad , v_pad , \a0_pad  , \f0_pad  , \g0_pad  , \i0_pad  , \j0_pad  , \k0_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , w_pad , x_pad , y_pad , z_pad );
  input a_pad ;
  input \b0_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input \h0_pad  ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input o_pad ;
  input t_pad ;
  input v_pad ;
  output \a0_pad  ;
  output \f0_pad  ;
  output \g0_pad  ;
  output \i0_pad  ;
  output \j0_pad  ;
  output \k0_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output w_pad ;
  output x_pad ;
  output y_pad ;
  output z_pad ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 ;
  assign n22 = i_pad & j_pad ;
  assign n23 = i_pad & k_pad ;
  assign n24 = ~\c0_pad  & n23 ;
  assign n26 = ~a_pad & n24 ;
  assign n25 = ~o_pad & ~n24 ;
  assign n27 = m_pad & ~n25 ;
  assign n28 = ~n26 & n27 ;
  assign n31 = b_pad & n24 ;
  assign n29 = \c0_pad  & n23 ;
  assign n30 = ~\h0_pad  & ~n29 ;
  assign n32 = m_pad & ~n30 ;
  assign n33 = ~n31 & n32 ;
  assign n34 = c_pad & n23 ;
  assign n35 = ~\c0_pad  & ~n34 ;
  assign n36 = m_pad & ~n29 ;
  assign n37 = ~n35 & n36 ;
  assign n39 = \e0_pad  & ~\h0_pad  ;
  assign n40 = ~n24 & ~n39 ;
  assign n38 = ~d_pad & n24 ;
  assign n41 = m_pad & ~n38 ;
  assign n42 = ~n40 & n41 ;
  assign n44 = ~e_pad & n24 ;
  assign n43 = ~\d0_pad  & ~n24 ;
  assign n45 = m_pad & ~n43 ;
  assign n46 = ~n44 & n45 ;
  assign n48 = ~f_pad & n24 ;
  assign n47 = ~t_pad & ~n24 ;
  assign n49 = m_pad & ~n47 ;
  assign n50 = ~n48 & n49 ;
  assign n52 = ~g_pad & n24 ;
  assign n51 = ~\b0_pad  & ~n24 ;
  assign n53 = m_pad & ~n51 ;
  assign n54 = ~n52 & n53 ;
  assign n56 = ~h_pad & n24 ;
  assign n55 = ~v_pad & ~n24 ;
  assign n57 = m_pad & ~n55 ;
  assign n58 = ~n56 & n57 ;
  assign n59 = l_pad & v_pad ;
  assign n60 = ~\h0_pad  & n29 ;
  assign n61 = ~\h0_pad  & ~n24 ;
  assign n62 = ~l_pad & m_pad ;
  assign n63 = ~n61 & n62 ;
  assign n64 = m_pad & n60 ;
  assign \a0_pad  = ~t_pad ;
  assign \f0_pad  = n22 ;
  assign \g0_pad  = ~n22 ;
  assign \i0_pad  = n28 ;
  assign \j0_pad  = n33 ;
  assign \k0_pad  = n37 ;
  assign \l0_pad  = n42 ;
  assign \m0_pad  = n46 ;
  assign \n0_pad  = n50 ;
  assign \o0_pad  = n54 ;
  assign \p0_pad  = n58 ;
  assign w_pad = n59 ;
  assign x_pad = n60 ;
  assign y_pad = n63 ;
  assign z_pad = n64 ;
endmodule
