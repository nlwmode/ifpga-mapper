module top (ACCRPY_pad, \BULL0_pad , \BULL1_pad , \BULL2_pad , \BULL3_pad , \BULL4_pad , \BULL5_pad , \BULL6_pad , CAPSD_pad, \CAT0_pad , \CAT1_pad , \CAT2_pad , \CAT3_pad , \CAT4_pad , \CAT5_pad , COMPPAR_pad, \DEL1_pad , END_pad, FBI_pad, \IBT0_pad , \IBT1_pad , \IBT2_pad , ICLR_pad, KBG_N_pad, LSD_pad, MARSSR_pad, MMERR_pad, ORWD_N_pad, OVACC_pad, OWL_N_pad, \PLUTO0_pad , \PLUTO1_pad , \PLUTO2_pad , \PLUTO3_pad , \PLUTO4_pad , \PLUTO5_pad , PY_pad, RATR_pad, SDO_pad, \STAR0_pad , \STAR1_pad , \STAR2_pad , \STAR3_pad , VACC_pad, VERR_N_pad, VLENESR_pad, \VST1_pad , VSUMESR_pad, WATCH_pad, ACCRPY_P_pad, \BULL0_P_pad , \BULL1_P_pad , \BULL2_P_pad , \BULL3_P_pad , \BULL4_P_pad , \BULL5_P_pad , \BULL6_P_pad , COMPPAR_P_pad, \DEL1_P_pad , END_P_pad, KBG_F_pad, LSD_P_pad, MARSSR_P_pad, ORWD_F_pad, OVACC_P_pad, OWL_F_pad, \PLUTO0_P_pad , \PLUTO1_P_pad , \PLUTO2_P_pad , \PLUTO3_P_pad , \PLUTO4_P_pad , \PLUTO5_P_pad , PY_P_pad, RATR_P_pad, \STAR0_P_pad , \STAR1_P_pad , \STAR2_P_pad , \STAR3_P_pad , VERR_F_pad, VLENESR_P_pad, \VST0_P_pad , \VST1_P_pad , VSUMESR_P_pad, WATCH_P_pad, \n1022 );
	input ACCRPY_pad ;
	input \BULL0_pad  ;
	input \BULL1_pad  ;
	input \BULL2_pad  ;
	input \BULL3_pad  ;
	input \BULL4_pad  ;
	input \BULL5_pad  ;
	input \BULL6_pad  ;
	input CAPSD_pad ;
	input \CAT0_pad  ;
	input \CAT1_pad  ;
	input \CAT2_pad  ;
	input \CAT3_pad  ;
	input \CAT4_pad  ;
	input \CAT5_pad  ;
	input COMPPAR_pad ;
	input \DEL1_pad  ;
	input END_pad ;
	input FBI_pad ;
	input \IBT0_pad  ;
	input \IBT1_pad  ;
	input \IBT2_pad  ;
	input ICLR_pad ;
	input KBG_N_pad ;
	input LSD_pad ;
	input MARSSR_pad ;
	input MMERR_pad ;
	input ORWD_N_pad ;
	input OVACC_pad ;
	input OWL_N_pad ;
	input \PLUTO0_pad  ;
	input \PLUTO1_pad  ;
	input \PLUTO2_pad  ;
	input \PLUTO3_pad  ;
	input \PLUTO4_pad  ;
	input \PLUTO5_pad  ;
	input PY_pad ;
	input RATR_pad ;
	input SDO_pad ;
	input \STAR0_pad  ;
	input \STAR1_pad  ;
	input \STAR2_pad  ;
	input \STAR3_pad  ;
	input VACC_pad ;
	input VERR_N_pad ;
	input VLENESR_pad ;
	input \VST1_pad  ;
	input VSUMESR_pad ;
	input WATCH_pad ;
	output ACCRPY_P_pad ;
	output \BULL0_P_pad  ;
	output \BULL1_P_pad  ;
	output \BULL2_P_pad  ;
	output \BULL3_P_pad  ;
	output \BULL4_P_pad  ;
	output \BULL5_P_pad  ;
	output \BULL6_P_pad  ;
	output COMPPAR_P_pad ;
	output \DEL1_P_pad  ;
	output END_P_pad ;
	output KBG_F_pad ;
	output LSD_P_pad ;
	output MARSSR_P_pad ;
	output ORWD_F_pad ;
	output OVACC_P_pad ;
	output OWL_F_pad ;
	output \PLUTO0_P_pad  ;
	output \PLUTO1_P_pad  ;
	output \PLUTO2_P_pad  ;
	output \PLUTO3_P_pad  ;
	output \PLUTO4_P_pad  ;
	output \PLUTO5_P_pad  ;
	output PY_P_pad ;
	output RATR_P_pad ;
	output \STAR0_P_pad  ;
	output \STAR1_P_pad  ;
	output \STAR2_P_pad  ;
	output \STAR3_P_pad  ;
	output VERR_F_pad ;
	output VLENESR_P_pad ;
	output \VST0_P_pad  ;
	output \VST1_P_pad  ;
	output VSUMESR_P_pad ;
	output WATCH_P_pad ;
	output \n1022  ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\CAT4_pad ,
		\IBT0_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\CAT5_pad ,
		\IBT0_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\IBT1_pad ,
		_w50_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\CAT2_pad ,
		\IBT0_pad ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\CAT3_pad ,
		\IBT0_pad ,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\IBT1_pad ,
		_w54_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w53_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\IBT2_pad ,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		\CAT0_pad ,
		\IBT0_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\CAT1_pad ,
		\IBT0_pad ,
		_w61_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\IBT1_pad ,
		\IBT2_pad ,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w60_,
		_w61_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w62_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w59_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		WATCH_pad,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\STAR0_pad ,
		\STAR1_pad ,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\STAR2_pad ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w66_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		FBI_pad,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		ACCRPY_pad,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		OWL_N_pad,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\BULL0_pad ,
		WATCH_pad,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\BULL0_pad ,
		WATCH_pad,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		OWL_N_pad,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\BULL0_pad ,
		\BULL1_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		WATCH_pad,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		OWL_N_pad,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\BULL1_pad ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		OWL_N_pad,
		WATCH_pad,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\BULL0_pad ,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\BULL1_pad ,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w80_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\BULL2_pad ,
		_w78_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\BULL2_pad ,
		_w78_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		OWL_N_pad,
		_w85_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\BULL3_pad ,
		_w85_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\BULL3_pad ,
		_w85_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		OWL_N_pad,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w89_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\BULL4_pad ,
		_w91_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		OWL_N_pad,
		_w90_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		\BULL4_pad ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w93_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\BULL5_pad ,
		_w91_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\BULL4_pad ,
		\BULL5_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\BULL4_pad ,
		\BULL5_pad ,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w98_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w94_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w97_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\BULL2_pad ,
		\BULL3_pad ,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w98_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w79_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\BULL6_pad ,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\BULL6_pad ,
		_w98_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w90_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w106_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		OWL_N_pad,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\DEL1_pad ,
		FBI_pad,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		COMPPAR_pad,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		COMPPAR_pad,
		_w111_,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		OWL_N_pad,
		_w112_,
		_w114_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w113_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		CAPSD_pad,
		ICLR_pad,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		END_pad,
		_w70_,
		_w117_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		OWL_N_pad,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\STAR3_pad ,
		_w68_,
		_w119_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		_w66_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		FBI_pad,
		_w69_,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		KBG_N_pad,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		OWL_N_pad,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		LSD_pad,
		OWL_N_pad,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		FBI_pad,
		_w119_,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		FBI_pad,
		\STAR3_pad ,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w81_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w125_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w68_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w65_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w127_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\BULL1_pad ,
		\BULL2_pad ,
		_w134_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\BULL3_pad ,
		\BULL4_pad ,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\BULL5_pad ,
		\BULL6_pad ,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w135_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w74_,
		_w134_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		MARSSR_pad,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		OWL_N_pad,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		ICLR_pad,
		VACC_pad,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		KBG_N_pad,
		_w139_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		END_pad,
		ICLR_pad,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		OWL_N_pad,
		\PLUTO0_pad ,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		MMERR_pad,
		SDO_pad,
		_w147_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		COMPPAR_pad,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		\VST1_pad ,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		END_pad,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		_w143_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		OWL_N_pad,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w62_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\IBT0_pad ,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w146_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		OWL_N_pad,
		\PLUTO1_pad ,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\IBT0_pad ,
		_w153_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		OWL_N_pad,
		\PLUTO2_pad ,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\IBT2_pad ,
		_w152_,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		\IBT0_pad ,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		\IBT1_pad ,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w159_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		OWL_N_pad,
		\PLUTO3_pad ,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\IBT0_pad ,
		_w160_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		\IBT1_pad ,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w164_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		OWL_N_pad,
		\PLUTO4_pad ,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\IBT1_pad ,
		_w161_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		OWL_N_pad,
		\PLUTO5_pad ,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\IBT1_pad ,
		_w165_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w171_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		FBI_pad,
		PY_pad,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w111_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		ICLR_pad,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		END_pad,
		_w148_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		RATR_pad,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		OWL_N_pad,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		ORWD_N_pad,
		_w66_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		FBI_pad,
		OWL_N_pad,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w180_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\STAR0_pad ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		FBI_pad,
		_w180_,
		_w184_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		OWL_N_pad,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\STAR0_pad ,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w183_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		_w67_,
		_w184_,
		_w188_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		OWL_N_pad,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\STAR1_pad ,
		_w183_,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		\STAR0_pad ,
		\STAR1_pad ,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w185_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w191_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\STAR2_pad ,
		_w189_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w68_,
		_w185_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\STAR2_pad ,
		_w67_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w184_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		\STAR3_pad ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\STAR3_pad ,
		_w199_,
		_w201_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		OWL_N_pad,
		_w200_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		VERR_N_pad,
		_w139_,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w122_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		OWL_N_pad,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name157 (
		KBG_N_pad,
		VLENESR_pad,
		_w207_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		OWL_N_pad,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		FBI_pad,
		ICLR_pad,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\VST1_pad ,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		FBI_pad,
		ICLR_pad,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		SDO_pad,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w210_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\VST1_pad ,
		_w211_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		PY_pad,
		_w209_,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		END_pad,
		\VST1_pad ,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		VSUMESR_pad,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name169 (
		OWL_N_pad,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		OVACC_pad,
		VACC_pad,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		WATCH_pad,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		OWL_N_pad,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		_w69_,
		_w185_,
		_w223_
	);
	assign ACCRPY_P_pad = _w72_ ;
	assign \BULL0_P_pad  = _w76_ ;
	assign \BULL1_P_pad  = _w84_ ;
	assign \BULL2_P_pad  = _w88_ ;
	assign \BULL3_P_pad  = _w92_ ;
	assign \BULL4_P_pad  = _w96_ ;
	assign \BULL5_P_pad  = _w102_ ;
	assign \BULL6_P_pad  = _w110_ ;
	assign COMPPAR_P_pad = _w115_ ;
	assign \DEL1_P_pad  = _w116_ ;
	assign END_P_pad = _w118_ ;
	assign KBG_F_pad = _w124_ ;
	assign LSD_P_pad = _w133_ ;
	assign MARSSR_P_pad = _w141_ ;
	assign ORWD_F_pad = _w66_ ;
	assign OVACC_P_pad = _w142_ ;
	assign OWL_F_pad = _w145_ ;
	assign \PLUTO0_P_pad  = _w155_ ;
	assign \PLUTO1_P_pad  = _w158_ ;
	assign \PLUTO2_P_pad  = _w163_ ;
	assign \PLUTO3_P_pad  = _w167_ ;
	assign \PLUTO4_P_pad  = _w170_ ;
	assign \PLUTO5_P_pad  = _w173_ ;
	assign PY_P_pad = _w176_ ;
	assign RATR_P_pad = _w179_ ;
	assign \STAR0_P_pad  = _w187_ ;
	assign \STAR1_P_pad  = _w194_ ;
	assign \STAR2_P_pad  = _w197_ ;
	assign \STAR3_P_pad  = _w203_ ;
	assign VERR_F_pad = _w206_ ;
	assign VLENESR_P_pad = _w208_ ;
	assign \VST0_P_pad  = _w213_ ;
	assign \VST1_P_pad  = _w216_ ;
	assign VSUMESR_P_pad = _w219_ ;
	assign WATCH_P_pad = _w222_ ;
	assign \n1022  = _w223_ ;
endmodule;