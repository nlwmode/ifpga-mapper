module top( \a[0]  , \a[1]  , \a[2]  , \a[3]  , \a[4]  , \a[5]  , \a[6]  , \a[7]  , \a[8]  , \a[9]  , \a[10]  , \a[11]  , \a[12]  , \a[13]  , \a[14]  , \a[15]  , \a[16]  , \a[17]  , \a[18]  , \a[19]  , \a[20]  , \a[21]  , \a[22]  , \a[23]  , \a[24]  , \a[25]  , \a[26]  , \a[27]  , \a[28]  , \a[29]  , \a[30]  , \a[31]  , \a[32]  , \a[33]  , \a[34]  , \a[35]  , \a[36]  , \a[37]  , \a[38]  , \a[39]  , \a[40]  , \a[41]  , \a[42]  , \a[43]  , \a[44]  , \a[45]  , \a[46]  , \a[47]  , \a[48]  , \a[49]  , \a[50]  , \a[51]  , \a[52]  , \a[53]  , \a[54]  , \a[55]  , \a[56]  , \a[57]  , \a[58]  , \a[59]  , \a[60]  , \a[61]  , \a[62]  , \a[63]  , \b[0]  , \b[1]  , \b[2]  , \b[3]  , \b[4]  , \b[5]  , \b[6]  , \b[7]  , \b[8]  , \b[9]  , \b[10]  , \b[11]  , \b[12]  , \b[13]  , \b[14]  , \b[15]  , \b[16]  , \b[17]  , \b[18]  , \b[19]  , \b[20]  , \b[21]  , \b[22]  , \b[23]  , \b[24]  , \b[25]  , \b[26]  , \b[27]  , \b[28]  , \b[29]  , \b[30]  , \b[31]  , \b[32]  , \b[33]  , \b[34]  , \b[35]  , \b[36]  , \b[37]  , \b[38]  , \b[39]  , \b[40]  , \b[41]  , \b[42]  , \b[43]  , \b[44]  , \b[45]  , \b[46]  , \b[47]  , \b[48]  , \b[49]  , \b[50]  , \b[51]  , \b[52]  , \b[53]  , \b[54]  , \b[55]  , \b[56]  , \b[57]  , \b[58]  , \b[59]  , \b[60]  , \b[61]  , \b[62]  , \b[63]  , \f[0]  , \f[1]  , \f[2]  , \f[3]  , \f[4]  , \f[5]  , \f[6]  , \f[7]  , \f[8]  , \f[9]  , \f[10]  , \f[11]  , \f[12]  , \f[13]  , \f[14]  , \f[15]  , \f[16]  , \f[17]  , \f[18]  , \f[19]  , \f[20]  , \f[21]  , \f[22]  , \f[23]  , \f[24]  , \f[25]  , \f[26]  , \f[27]  , \f[28]  , \f[29]  , \f[30]  , \f[31]  , \f[32]  , \f[33]  , \f[34]  , \f[35]  , \f[36]  , \f[37]  , \f[38]  , \f[39]  , \f[40]  , \f[41]  , \f[42]  , \f[43]  , \f[44]  , \f[45]  , \f[46]  , \f[47]  , \f[48]  , \f[49]  , \f[50]  , \f[51]  , \f[52]  , \f[53]  , \f[54]  , \f[55]  , \f[56]  , \f[57]  , \f[58]  , \f[59]  , \f[60]  , \f[61]  , \f[62]  , \f[63]  , \f[64]  , \f[65]  , \f[66]  , \f[67]  , \f[68]  , \f[69]  , \f[70]  , \f[71]  , \f[72]  , \f[73]  , \f[74]  , \f[75]  , \f[76]  , \f[77]  , \f[78]  , \f[79]  , \f[80]  , \f[81]  , \f[82]  , \f[83]  , \f[84]  , \f[85]  , \f[86]  , \f[87]  , \f[88]  , \f[89]  , \f[90]  , \f[91]  , \f[92]  , \f[93]  , \f[94]  , \f[95]  , \f[96]  , \f[97]  , \f[98]  , \f[99]  , \f[100]  , \f[101]  , \f[102]  , \f[103]  , \f[104]  , \f[105]  , \f[106]  , \f[107]  , \f[108]  , \f[109]  , \f[110]  , \f[111]  , \f[112]  , \f[113]  , \f[114]  , \f[115]  , \f[116]  , \f[117]  , \f[118]  , \f[119]  , \f[120]  , \f[121]  , \f[122]  , \f[123]  , \f[124]  , \f[125]  , \f[126]  , \f[127]  );
  input \a[0]  ;
  input \a[1]  ;
  input \a[2]  ;
  input \a[3]  ;
  input \a[4]  ;
  input \a[5]  ;
  input \a[6]  ;
  input \a[7]  ;
  input \a[8]  ;
  input \a[9]  ;
  input \a[10]  ;
  input \a[11]  ;
  input \a[12]  ;
  input \a[13]  ;
  input \a[14]  ;
  input \a[15]  ;
  input \a[16]  ;
  input \a[17]  ;
  input \a[18]  ;
  input \a[19]  ;
  input \a[20]  ;
  input \a[21]  ;
  input \a[22]  ;
  input \a[23]  ;
  input \a[24]  ;
  input \a[25]  ;
  input \a[26]  ;
  input \a[27]  ;
  input \a[28]  ;
  input \a[29]  ;
  input \a[30]  ;
  input \a[31]  ;
  input \a[32]  ;
  input \a[33]  ;
  input \a[34]  ;
  input \a[35]  ;
  input \a[36]  ;
  input \a[37]  ;
  input \a[38]  ;
  input \a[39]  ;
  input \a[40]  ;
  input \a[41]  ;
  input \a[42]  ;
  input \a[43]  ;
  input \a[44]  ;
  input \a[45]  ;
  input \a[46]  ;
  input \a[47]  ;
  input \a[48]  ;
  input \a[49]  ;
  input \a[50]  ;
  input \a[51]  ;
  input \a[52]  ;
  input \a[53]  ;
  input \a[54]  ;
  input \a[55]  ;
  input \a[56]  ;
  input \a[57]  ;
  input \a[58]  ;
  input \a[59]  ;
  input \a[60]  ;
  input \a[61]  ;
  input \a[62]  ;
  input \a[63]  ;
  input \b[0]  ;
  input \b[1]  ;
  input \b[2]  ;
  input \b[3]  ;
  input \b[4]  ;
  input \b[5]  ;
  input \b[6]  ;
  input \b[7]  ;
  input \b[8]  ;
  input \b[9]  ;
  input \b[10]  ;
  input \b[11]  ;
  input \b[12]  ;
  input \b[13]  ;
  input \b[14]  ;
  input \b[15]  ;
  input \b[16]  ;
  input \b[17]  ;
  input \b[18]  ;
  input \b[19]  ;
  input \b[20]  ;
  input \b[21]  ;
  input \b[22]  ;
  input \b[23]  ;
  input \b[24]  ;
  input \b[25]  ;
  input \b[26]  ;
  input \b[27]  ;
  input \b[28]  ;
  input \b[29]  ;
  input \b[30]  ;
  input \b[31]  ;
  input \b[32]  ;
  input \b[33]  ;
  input \b[34]  ;
  input \b[35]  ;
  input \b[36]  ;
  input \b[37]  ;
  input \b[38]  ;
  input \b[39]  ;
  input \b[40]  ;
  input \b[41]  ;
  input \b[42]  ;
  input \b[43]  ;
  input \b[44]  ;
  input \b[45]  ;
  input \b[46]  ;
  input \b[47]  ;
  input \b[48]  ;
  input \b[49]  ;
  input \b[50]  ;
  input \b[51]  ;
  input \b[52]  ;
  input \b[53]  ;
  input \b[54]  ;
  input \b[55]  ;
  input \b[56]  ;
  input \b[57]  ;
  input \b[58]  ;
  input \b[59]  ;
  input \b[60]  ;
  input \b[61]  ;
  input \b[62]  ;
  input \b[63]  ;
  output \f[0]  ;
  output \f[1]  ;
  output \f[2]  ;
  output \f[3]  ;
  output \f[4]  ;
  output \f[5]  ;
  output \f[6]  ;
  output \f[7]  ;
  output \f[8]  ;
  output \f[9]  ;
  output \f[10]  ;
  output \f[11]  ;
  output \f[12]  ;
  output \f[13]  ;
  output \f[14]  ;
  output \f[15]  ;
  output \f[16]  ;
  output \f[17]  ;
  output \f[18]  ;
  output \f[19]  ;
  output \f[20]  ;
  output \f[21]  ;
  output \f[22]  ;
  output \f[23]  ;
  output \f[24]  ;
  output \f[25]  ;
  output \f[26]  ;
  output \f[27]  ;
  output \f[28]  ;
  output \f[29]  ;
  output \f[30]  ;
  output \f[31]  ;
  output \f[32]  ;
  output \f[33]  ;
  output \f[34]  ;
  output \f[35]  ;
  output \f[36]  ;
  output \f[37]  ;
  output \f[38]  ;
  output \f[39]  ;
  output \f[40]  ;
  output \f[41]  ;
  output \f[42]  ;
  output \f[43]  ;
  output \f[44]  ;
  output \f[45]  ;
  output \f[46]  ;
  output \f[47]  ;
  output \f[48]  ;
  output \f[49]  ;
  output \f[50]  ;
  output \f[51]  ;
  output \f[52]  ;
  output \f[53]  ;
  output \f[54]  ;
  output \f[55]  ;
  output \f[56]  ;
  output \f[57]  ;
  output \f[58]  ;
  output \f[59]  ;
  output \f[60]  ;
  output \f[61]  ;
  output \f[62]  ;
  output \f[63]  ;
  output \f[64]  ;
  output \f[65]  ;
  output \f[66]  ;
  output \f[67]  ;
  output \f[68]  ;
  output \f[69]  ;
  output \f[70]  ;
  output \f[71]  ;
  output \f[72]  ;
  output \f[73]  ;
  output \f[74]  ;
  output \f[75]  ;
  output \f[76]  ;
  output \f[77]  ;
  output \f[78]  ;
  output \f[79]  ;
  output \f[80]  ;
  output \f[81]  ;
  output \f[82]  ;
  output \f[83]  ;
  output \f[84]  ;
  output \f[85]  ;
  output \f[86]  ;
  output \f[87]  ;
  output \f[88]  ;
  output \f[89]  ;
  output \f[90]  ;
  output \f[91]  ;
  output \f[92]  ;
  output \f[93]  ;
  output \f[94]  ;
  output \f[95]  ;
  output \f[96]  ;
  output \f[97]  ;
  output \f[98]  ;
  output \f[99]  ;
  output \f[100]  ;
  output \f[101]  ;
  output \f[102]  ;
  output \f[103]  ;
  output \f[104]  ;
  output \f[105]  ;
  output \f[106]  ;
  output \f[107]  ;
  output \f[108]  ;
  output \f[109]  ;
  output \f[110]  ;
  output \f[111]  ;
  output \f[112]  ;
  output \f[113]  ;
  output \f[114]  ;
  output \f[115]  ;
  output \f[116]  ;
  output \f[117]  ;
  output \f[118]  ;
  output \f[119]  ;
  output \f[120]  ;
  output \f[121]  ;
  output \f[122]  ;
  output \f[123]  ;
  output \f[124]  ;
  output \f[125]  ;
  output \f[126]  ;
  output \f[127]  ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 ;
  assign n129 = \a[0]  & \b[0]  ;
  assign n130 = \a[2]  & n129 ;
  assign n131 = \a[1]  & ~\a[2]  ;
  assign n132 = ~\a[1]  & \a[2]  ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = \a[0]  & ~n133 ;
  assign n135 = ~\b[0]  & \b[1]  ;
  assign n136 = \b[0]  & ~\b[1]  ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = n134 & ~n137 ;
  assign n139 = \a[0]  & \b[1]  ;
  assign n140 = n133 & n139 ;
  assign n141 = ~\a[0]  & \a[1]  ;
  assign n142 = \b[0]  & n141 ;
  assign n143 = ~n140 & ~n142 ;
  assign n144 = ~n138 & n143 ;
  assign n145 = n130 & ~n144 ;
  assign n146 = ~n130 & ~n142 ;
  assign n147 = ~n140 & n146 ;
  assign n148 = ~n138 & n147 ;
  assign n149 = ~n145 & ~n148 ;
  assign n150 = \a[2]  & ~n129 ;
  assign n151 = ~n142 & n150 ;
  assign n152 = ~n140 & n151 ;
  assign n153 = ~n138 & n152 ;
  assign n154 = \a[2]  & ~n153 ;
  assign n155 = ~\b[2]  & ~n135 ;
  assign n156 = \b[2]  & n135 ;
  assign n157 = ~n155 & ~n156 ;
  assign n158 = n134 & n157 ;
  assign n159 = \a[0]  & \b[2]  ;
  assign n160 = n133 & n159 ;
  assign n161 = ~\a[0]  & \b[0]  ;
  assign n162 = n132 & n161 ;
  assign n163 = \b[1]  & n141 ;
  assign n164 = ~n162 & ~n163 ;
  assign n165 = ~n160 & n164 ;
  assign n166 = ~n158 & n165 ;
  assign n167 = ~n154 & n166 ;
  assign n168 = n154 & ~n166 ;
  assign n169 = ~n167 & ~n168 ;
  assign n170 = ~\b[2]  & ~\b[3]  ;
  assign n171 = \b[2]  & \b[3]  ;
  assign n172 = ~n170 & ~n171 ;
  assign n173 = ~\b[0]  & ~\b[2]  ;
  assign n174 = \b[1]  & ~n173 ;
  assign n175 = n172 & n174 ;
  assign n176 = ~n172 & ~n174 ;
  assign n177 = ~n175 & ~n176 ;
  assign n178 = n134 & n177 ;
  assign n179 = \a[0]  & \b[3]  ;
  assign n180 = n133 & n179 ;
  assign n181 = ~\a[0]  & \b[1]  ;
  assign n182 = n132 & n181 ;
  assign n183 = \b[2]  & n141 ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = ~n180 & n184 ;
  assign n186 = \a[2]  & n185 ;
  assign n187 = ~n178 & n186 ;
  assign n188 = ~\a[2]  & ~n185 ;
  assign n189 = \a[0]  & \a[1]  ;
  assign n190 = ~\a[2]  & n189 ;
  assign n191 = n177 & n190 ;
  assign n192 = ~n188 & ~n191 ;
  assign n193 = ~n187 & n192 ;
  assign n194 = \a[2]  & ~\a[3]  ;
  assign n195 = ~\a[2]  & \a[3]  ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = \b[0]  & ~n196 ;
  assign n198 = n153 & n166 ;
  assign n199 = ~n197 & n198 ;
  assign n200 = ~n193 & n199 ;
  assign n201 = n197 & n198 ;
  assign n202 = n193 & n201 ;
  assign n203 = ~n200 & ~n202 ;
  assign n204 = ~n197 & ~n198 ;
  assign n205 = n193 & n204 ;
  assign n206 = n197 & ~n198 ;
  assign n207 = ~n193 & n206 ;
  assign n208 = ~n205 & ~n207 ;
  assign n209 = n203 & n208 ;
  assign n210 = ~n193 & n197 ;
  assign n211 = n203 & ~n210 ;
  assign n212 = ~\b[1]  & ~\b[2]  ;
  assign n213 = ~n170 & ~n212 ;
  assign n214 = ~\b[1]  & ~\b[3]  ;
  assign n215 = ~n173 & ~n214 ;
  assign n216 = n213 & n215 ;
  assign n217 = ~\b[3]  & ~\b[4]  ;
  assign n218 = \b[3]  & \b[4]  ;
  assign n219 = ~n217 & ~n218 ;
  assign n220 = n216 & n219 ;
  assign n221 = ~n216 & ~n219 ;
  assign n222 = ~n220 & ~n221 ;
  assign n223 = n134 & n222 ;
  assign n224 = \a[0]  & \b[4]  ;
  assign n225 = n133 & n224 ;
  assign n226 = ~\a[0]  & \b[2]  ;
  assign n227 = n132 & n226 ;
  assign n228 = \b[3]  & n141 ;
  assign n229 = ~n227 & ~n228 ;
  assign n230 = ~n225 & n229 ;
  assign n231 = ~\a[2]  & n230 ;
  assign n232 = ~n223 & n231 ;
  assign n233 = \a[2]  & ~n230 ;
  assign n234 = \a[2]  & n134 ;
  assign n235 = n222 & n234 ;
  assign n236 = ~n233 & ~n235 ;
  assign n237 = ~n232 & n236 ;
  assign n238 = \a[5]  & \b[0]  ;
  assign n239 = ~n196 & n238 ;
  assign n240 = \a[3]  & \b[0]  ;
  assign n241 = \a[2]  & ~\a[4]  ;
  assign n242 = n240 & n241 ;
  assign n243 = ~\a[3]  & \b[0]  ;
  assign n244 = ~\a[2]  & \a[4]  ;
  assign n245 = n243 & n244 ;
  assign n246 = ~n242 & ~n245 ;
  assign n247 = \a[4]  & ~\a[5]  ;
  assign n248 = ~\a[4]  & \a[5]  ;
  assign n249 = ~n247 & ~n248 ;
  assign n250 = ~n196 & n249 ;
  assign n251 = \b[1]  & n250 ;
  assign n252 = ~n196 & ~n249 ;
  assign n253 = ~n137 & n252 ;
  assign n254 = ~n251 & ~n253 ;
  assign n255 = n246 & n254 ;
  assign n256 = n239 & ~n255 ;
  assign n257 = ~n239 & n246 ;
  assign n258 = n254 & n257 ;
  assign n259 = ~n256 & ~n258 ;
  assign n260 = n237 & n259 ;
  assign n261 = ~n237 & ~n259 ;
  assign n262 = ~n260 & ~n261 ;
  assign n263 = ~n211 & n262 ;
  assign n264 = n211 & ~n262 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = ~n260 & ~n263 ;
  assign n267 = ~n218 & ~n220 ;
  assign n268 = ~\b[4]  & ~\b[5]  ;
  assign n269 = \b[4]  & \b[5]  ;
  assign n270 = ~n268 & ~n269 ;
  assign n271 = ~n267 & n270 ;
  assign n272 = ~n218 & ~n270 ;
  assign n273 = ~n220 & n272 ;
  assign n274 = n134 & ~n273 ;
  assign n275 = ~n271 & n274 ;
  assign n276 = \a[0]  & \b[5]  ;
  assign n277 = n133 & n276 ;
  assign n278 = ~\a[0]  & \b[3]  ;
  assign n279 = n132 & n278 ;
  assign n280 = \b[4]  & n141 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = ~n277 & n281 ;
  assign n283 = ~n275 & n282 ;
  assign n284 = ~\a[2]  & ~n283 ;
  assign n285 = \a[2]  & n282 ;
  assign n286 = ~n275 & n285 ;
  assign n287 = ~n284 & ~n286 ;
  assign n288 = \a[5]  & ~n197 ;
  assign n289 = n246 & n288 ;
  assign n290 = n254 & n289 ;
  assign n291 = \a[5]  & ~n290 ;
  assign n292 = \b[2]  & n250 ;
  assign n293 = ~\a[3]  & \b[1]  ;
  assign n294 = n244 & n293 ;
  assign n295 = \a[3]  & \b[1]  ;
  assign n296 = n241 & n295 ;
  assign n297 = ~n294 & ~n296 ;
  assign n298 = ~n292 & n297 ;
  assign n299 = n157 & n252 ;
  assign n300 = n196 & ~n249 ;
  assign n301 = \a[3]  & ~\a[4]  ;
  assign n302 = ~\a[3]  & \a[4]  ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = \b[0]  & n303 ;
  assign n305 = n300 & n304 ;
  assign n306 = ~n299 & ~n305 ;
  assign n307 = n298 & n306 ;
  assign n308 = ~n291 & ~n307 ;
  assign n309 = n291 & n307 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = ~n287 & ~n310 ;
  assign n312 = n287 & n310 ;
  assign n313 = ~n311 & ~n312 ;
  assign n314 = ~n266 & n313 ;
  assign n315 = n266 & ~n313 ;
  assign n316 = ~n314 & ~n315 ;
  assign n317 = ~n311 & ~n314 ;
  assign n318 = ~n218 & ~n269 ;
  assign n319 = ~n220 & n318 ;
  assign n320 = ~n268 & ~n319 ;
  assign n321 = ~\b[5]  & ~\b[6]  ;
  assign n322 = \b[5]  & \b[6]  ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = ~n320 & ~n323 ;
  assign n325 = ~n268 & n323 ;
  assign n326 = ~n319 & n325 ;
  assign n327 = n134 & ~n326 ;
  assign n328 = ~n324 & n327 ;
  assign n329 = \a[0]  & \b[6]  ;
  assign n330 = n133 & n329 ;
  assign n331 = ~\a[0]  & \b[4]  ;
  assign n332 = n132 & n331 ;
  assign n333 = \b[5]  & n141 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = ~n330 & n334 ;
  assign n336 = ~n328 & n335 ;
  assign n337 = ~\a[2]  & ~n336 ;
  assign n338 = \a[2]  & n335 ;
  assign n339 = ~n328 & n338 ;
  assign n340 = ~n337 & ~n339 ;
  assign n341 = n177 & n252 ;
  assign n342 = \b[3]  & n250 ;
  assign n343 = \a[3]  & \b[2]  ;
  assign n344 = n241 & n343 ;
  assign n345 = ~\a[2]  & \b[2]  ;
  assign n346 = n302 & n345 ;
  assign n347 = ~n344 & ~n346 ;
  assign n348 = ~n342 & n347 ;
  assign n349 = ~n341 & n348 ;
  assign n350 = \b[1]  & n303 ;
  assign n351 = n300 & n350 ;
  assign n352 = ~\a[5]  & ~n351 ;
  assign n353 = n349 & n352 ;
  assign n354 = n349 & ~n351 ;
  assign n355 = \a[5]  & ~n354 ;
  assign n356 = ~n353 & ~n355 ;
  assign n357 = \a[5]  & ~\a[6]  ;
  assign n358 = ~\a[5]  & \a[6]  ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = \b[0]  & ~n359 ;
  assign n361 = n290 & n307 ;
  assign n362 = n360 & n361 ;
  assign n363 = ~n360 & ~n361 ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = n356 & n364 ;
  assign n366 = ~n356 & ~n364 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = ~n340 & n367 ;
  assign n369 = n340 & ~n367 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = ~n317 & n370 ;
  assign n372 = n317 & ~n370 ;
  assign n373 = ~n371 & ~n372 ;
  assign n374 = ~n311 & ~n368 ;
  assign n375 = ~n314 & n374 ;
  assign n376 = ~n369 & ~n375 ;
  assign n377 = ~n322 & ~n326 ;
  assign n378 = ~\b[6]  & ~\b[7]  ;
  assign n379 = \b[6]  & \b[7]  ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n377 & n380 ;
  assign n382 = ~n322 & ~n380 ;
  assign n383 = ~n326 & n382 ;
  assign n384 = n134 & ~n383 ;
  assign n385 = ~n381 & n384 ;
  assign n386 = \a[0]  & \b[7]  ;
  assign n387 = n133 & n386 ;
  assign n388 = ~\a[0]  & \b[5]  ;
  assign n389 = n132 & n388 ;
  assign n390 = \b[6]  & n141 ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = ~n387 & n391 ;
  assign n393 = ~n385 & n392 ;
  assign n394 = ~\a[2]  & ~n393 ;
  assign n395 = \a[2]  & n392 ;
  assign n396 = ~n385 & n395 ;
  assign n397 = ~n394 & ~n396 ;
  assign n398 = ~n362 & ~n365 ;
  assign n399 = n222 & n252 ;
  assign n400 = \b[4]  & n250 ;
  assign n401 = ~\a[2]  & \b[3]  ;
  assign n402 = n302 & n401 ;
  assign n403 = \a[3]  & \b[3]  ;
  assign n404 = n241 & n403 ;
  assign n405 = ~n402 & ~n404 ;
  assign n406 = ~n400 & n405 ;
  assign n407 = \b[2]  & n303 ;
  assign n408 = n300 & n407 ;
  assign n409 = \a[5]  & ~n408 ;
  assign n410 = n406 & n409 ;
  assign n411 = ~n399 & n410 ;
  assign n412 = n406 & ~n408 ;
  assign n413 = ~n399 & n412 ;
  assign n414 = ~\a[5]  & ~n413 ;
  assign n415 = ~n411 & ~n414 ;
  assign n416 = \a[8]  & \b[0]  ;
  assign n417 = ~n359 & n416 ;
  assign n418 = \a[6]  & \b[0]  ;
  assign n419 = \a[5]  & ~\a[7]  ;
  assign n420 = n418 & n419 ;
  assign n421 = ~\a[6]  & \b[0]  ;
  assign n422 = ~\a[5]  & \a[7]  ;
  assign n423 = n421 & n422 ;
  assign n424 = ~n420 & ~n423 ;
  assign n425 = \a[7]  & ~\a[8]  ;
  assign n426 = ~\a[7]  & \a[8]  ;
  assign n427 = ~n425 & ~n426 ;
  assign n428 = ~n359 & n427 ;
  assign n429 = \b[1]  & n428 ;
  assign n430 = ~n359 & ~n427 ;
  assign n431 = ~n137 & n430 ;
  assign n432 = ~n429 & ~n431 ;
  assign n433 = n424 & n432 ;
  assign n434 = n417 & ~n433 ;
  assign n435 = ~n417 & n424 ;
  assign n436 = n432 & n435 ;
  assign n437 = ~n434 & ~n436 ;
  assign n438 = ~n415 & n437 ;
  assign n439 = n415 & ~n437 ;
  assign n440 = ~n438 & ~n439 ;
  assign n441 = ~n398 & n440 ;
  assign n442 = n398 & ~n440 ;
  assign n443 = ~n441 & ~n442 ;
  assign n444 = ~n397 & n443 ;
  assign n445 = n397 & ~n443 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = n376 & n446 ;
  assign n448 = ~n376 & ~n446 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = ~n444 & ~n447 ;
  assign n451 = ~n438 & ~n441 ;
  assign n452 = n252 & ~n273 ;
  assign n453 = ~n271 & n452 ;
  assign n454 = \b[3]  & n303 ;
  assign n455 = n300 & n454 ;
  assign n456 = ~\a[2]  & \b[4]  ;
  assign n457 = n302 & n456 ;
  assign n458 = ~n455 & ~n457 ;
  assign n459 = \b[5]  & n250 ;
  assign n460 = \a[3]  & \b[4]  ;
  assign n461 = n241 & n460 ;
  assign n462 = \a[5]  & ~n461 ;
  assign n463 = ~n459 & n462 ;
  assign n464 = n458 & n463 ;
  assign n465 = ~n453 & n464 ;
  assign n466 = ~n459 & ~n461 ;
  assign n467 = n458 & n466 ;
  assign n468 = ~n453 & n467 ;
  assign n469 = ~\a[5]  & ~n468 ;
  assign n470 = ~n465 & ~n469 ;
  assign n471 = \a[8]  & ~n360 ;
  assign n472 = n424 & n471 ;
  assign n473 = n432 & n472 ;
  assign n474 = \a[8]  & ~n473 ;
  assign n475 = \b[2]  & n428 ;
  assign n476 = ~\a[6]  & \b[1]  ;
  assign n477 = n422 & n476 ;
  assign n478 = \a[6]  & \b[1]  ;
  assign n479 = n419 & n478 ;
  assign n480 = ~n477 & ~n479 ;
  assign n481 = ~n475 & n480 ;
  assign n482 = n157 & n430 ;
  assign n483 = n359 & ~n427 ;
  assign n484 = \a[6]  & ~\a[7]  ;
  assign n485 = ~\a[6]  & \a[7]  ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = \b[0]  & n486 ;
  assign n488 = n483 & n487 ;
  assign n489 = ~n482 & ~n488 ;
  assign n490 = n481 & n489 ;
  assign n491 = ~n474 & ~n490 ;
  assign n492 = n474 & n490 ;
  assign n493 = ~n491 & ~n492 ;
  assign n494 = ~n470 & ~n493 ;
  assign n495 = n470 & n493 ;
  assign n496 = ~n494 & ~n495 ;
  assign n497 = n451 & ~n496 ;
  assign n498 = ~n451 & n496 ;
  assign n499 = ~n497 & ~n498 ;
  assign n500 = ~n322 & ~n379 ;
  assign n501 = ~n326 & n500 ;
  assign n502 = ~n378 & ~n501 ;
  assign n503 = ~\b[7]  & ~\b[8]  ;
  assign n504 = \b[7]  & \b[8]  ;
  assign n505 = ~n503 & ~n504 ;
  assign n506 = ~n502 & ~n505 ;
  assign n507 = ~n378 & n505 ;
  assign n508 = ~n501 & n507 ;
  assign n509 = n134 & ~n508 ;
  assign n510 = ~n506 & n509 ;
  assign n511 = \a[0]  & \b[8]  ;
  assign n512 = n133 & n511 ;
  assign n513 = ~\a[0]  & \b[6]  ;
  assign n514 = n132 & n513 ;
  assign n515 = \b[7]  & n141 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = ~n512 & n516 ;
  assign n518 = ~n510 & n517 ;
  assign n519 = ~\a[2]  & ~n518 ;
  assign n520 = \a[2]  & n517 ;
  assign n521 = ~n510 & n520 ;
  assign n522 = ~n519 & ~n521 ;
  assign n523 = n499 & ~n522 ;
  assign n524 = ~n499 & n522 ;
  assign n525 = ~n523 & ~n524 ;
  assign n526 = ~n450 & n525 ;
  assign n527 = n450 & ~n525 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = ~n523 & ~n526 ;
  assign n530 = ~n438 & ~n494 ;
  assign n531 = ~n441 & n530 ;
  assign n532 = ~n495 & ~n531 ;
  assign n533 = n177 & n430 ;
  assign n534 = \b[3]  & n428 ;
  assign n535 = \a[5]  & \b[2]  ;
  assign n536 = n484 & n535 ;
  assign n537 = ~\a[6]  & \b[2]  ;
  assign n538 = n422 & n537 ;
  assign n539 = ~n536 & ~n538 ;
  assign n540 = ~n534 & n539 ;
  assign n541 = ~n533 & n540 ;
  assign n542 = \b[1]  & n486 ;
  assign n543 = n483 & n542 ;
  assign n544 = ~\a[8]  & ~n543 ;
  assign n545 = n541 & n544 ;
  assign n546 = n541 & ~n543 ;
  assign n547 = \a[8]  & ~n546 ;
  assign n548 = ~n545 & ~n547 ;
  assign n549 = \a[8]  & ~\a[9]  ;
  assign n550 = ~\a[8]  & \a[9]  ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = \b[0]  & ~n551 ;
  assign n553 = n473 & n490 ;
  assign n554 = n552 & n553 ;
  assign n555 = ~n552 & ~n553 ;
  assign n556 = ~n554 & ~n555 ;
  assign n557 = n548 & n556 ;
  assign n558 = ~n548 & ~n556 ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = n252 & ~n326 ;
  assign n561 = ~n324 & n560 ;
  assign n562 = \b[4]  & n303 ;
  assign n563 = n300 & n562 ;
  assign n564 = \b[6]  & n250 ;
  assign n565 = \a[3]  & \b[5]  ;
  assign n566 = n241 & n565 ;
  assign n567 = ~\a[3]  & \b[5]  ;
  assign n568 = n244 & n567 ;
  assign n569 = ~n566 & ~n568 ;
  assign n570 = ~n564 & n569 ;
  assign n571 = ~n563 & n570 ;
  assign n572 = ~n561 & n571 ;
  assign n573 = ~\a[5]  & ~n572 ;
  assign n574 = \a[5]  & n571 ;
  assign n575 = ~n561 & n574 ;
  assign n576 = ~n573 & ~n575 ;
  assign n577 = n559 & ~n576 ;
  assign n578 = ~n559 & n576 ;
  assign n579 = ~n577 & ~n578 ;
  assign n580 = ~n532 & ~n579 ;
  assign n581 = n532 & n579 ;
  assign n582 = ~n580 & ~n581 ;
  assign n583 = ~n504 & ~n508 ;
  assign n584 = ~\b[8]  & ~\b[9]  ;
  assign n585 = \b[8]  & \b[9]  ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~n583 & n586 ;
  assign n588 = ~n504 & ~n586 ;
  assign n589 = ~n508 & n588 ;
  assign n590 = n134 & ~n589 ;
  assign n591 = ~n587 & n590 ;
  assign n592 = \a[0]  & \b[9]  ;
  assign n593 = n133 & n592 ;
  assign n594 = ~\a[0]  & \b[7]  ;
  assign n595 = n132 & n594 ;
  assign n596 = \b[8]  & n141 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = ~n593 & n597 ;
  assign n599 = ~n591 & n598 ;
  assign n600 = ~\a[2]  & ~n599 ;
  assign n601 = \a[2]  & n598 ;
  assign n602 = ~n591 & n601 ;
  assign n603 = ~n600 & ~n602 ;
  assign n604 = n582 & ~n603 ;
  assign n605 = ~n582 & n603 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = ~n529 & n606 ;
  assign n608 = n529 & ~n606 ;
  assign n609 = ~n607 & ~n608 ;
  assign n610 = ~n523 & ~n604 ;
  assign n611 = ~n526 & n610 ;
  assign n612 = ~n605 & ~n611 ;
  assign n613 = ~n577 & ~n581 ;
  assign n614 = ~n554 & ~n557 ;
  assign n615 = n222 & n430 ;
  assign n616 = \b[4]  & n428 ;
  assign n617 = \a[5]  & \b[3]  ;
  assign n618 = n484 & n617 ;
  assign n619 = ~\a[6]  & \b[3]  ;
  assign n620 = n422 & n619 ;
  assign n621 = ~n618 & ~n620 ;
  assign n622 = ~n616 & n621 ;
  assign n623 = \b[2]  & n486 ;
  assign n624 = n483 & n623 ;
  assign n625 = \a[8]  & ~n624 ;
  assign n626 = n622 & n625 ;
  assign n627 = ~n615 & n626 ;
  assign n628 = n622 & ~n624 ;
  assign n629 = ~n615 & n628 ;
  assign n630 = ~\a[8]  & ~n629 ;
  assign n631 = ~n627 & ~n630 ;
  assign n632 = \a[11]  & \b[0]  ;
  assign n633 = ~n551 & n632 ;
  assign n634 = \a[9]  & \b[0]  ;
  assign n635 = \a[8]  & ~\a[10]  ;
  assign n636 = n634 & n635 ;
  assign n637 = ~\a[9]  & \b[0]  ;
  assign n638 = ~\a[8]  & \a[10]  ;
  assign n639 = n637 & n638 ;
  assign n640 = ~n636 & ~n639 ;
  assign n641 = \a[10]  & ~\a[11]  ;
  assign n642 = ~\a[10]  & \a[11]  ;
  assign n643 = ~n641 & ~n642 ;
  assign n644 = ~n551 & n643 ;
  assign n645 = \b[1]  & n644 ;
  assign n646 = ~n551 & ~n643 ;
  assign n647 = ~n137 & n646 ;
  assign n648 = ~n645 & ~n647 ;
  assign n649 = n640 & n648 ;
  assign n650 = n633 & ~n649 ;
  assign n651 = ~n633 & n640 ;
  assign n652 = n648 & n651 ;
  assign n653 = ~n650 & ~n652 ;
  assign n654 = n631 & ~n653 ;
  assign n655 = ~n631 & n653 ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = ~n614 & n656 ;
  assign n658 = n614 & ~n656 ;
  assign n659 = ~n657 & ~n658 ;
  assign n660 = n252 & ~n383 ;
  assign n661 = ~n381 & n660 ;
  assign n662 = \b[5]  & n303 ;
  assign n663 = n300 & n662 ;
  assign n664 = \b[7]  & n250 ;
  assign n665 = \a[3]  & \b[6]  ;
  assign n666 = n241 & n665 ;
  assign n667 = ~\a[3]  & \b[6]  ;
  assign n668 = n244 & n667 ;
  assign n669 = ~n666 & ~n668 ;
  assign n670 = ~n664 & n669 ;
  assign n671 = ~n663 & n670 ;
  assign n672 = ~\a[5]  & n671 ;
  assign n673 = ~n661 & n672 ;
  assign n674 = ~n661 & n671 ;
  assign n675 = \a[5]  & ~n674 ;
  assign n676 = ~n673 & ~n675 ;
  assign n677 = n659 & n676 ;
  assign n678 = ~n659 & ~n676 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = ~n504 & ~n585 ;
  assign n681 = ~n508 & n680 ;
  assign n682 = ~n584 & ~n681 ;
  assign n683 = ~\b[9]  & ~\b[10]  ;
  assign n684 = \b[9]  & \b[10]  ;
  assign n685 = ~n683 & ~n684 ;
  assign n686 = n134 & n685 ;
  assign n687 = ~n682 & n686 ;
  assign n688 = n134 & ~n685 ;
  assign n689 = ~n584 & n688 ;
  assign n690 = ~n681 & n689 ;
  assign n691 = \a[0]  & \b[10]  ;
  assign n692 = n133 & n691 ;
  assign n693 = ~\a[0]  & \b[8]  ;
  assign n694 = n132 & n693 ;
  assign n695 = \b[9]  & n141 ;
  assign n696 = ~n694 & ~n695 ;
  assign n697 = ~n692 & n696 ;
  assign n698 = ~n690 & n697 ;
  assign n699 = ~n687 & n698 ;
  assign n700 = ~\a[2]  & ~n699 ;
  assign n701 = \a[2]  & n697 ;
  assign n702 = ~n690 & n701 ;
  assign n703 = ~n687 & n702 ;
  assign n704 = ~n700 & ~n703 ;
  assign n705 = ~n679 & n704 ;
  assign n706 = n613 & n705 ;
  assign n707 = n679 & n704 ;
  assign n708 = ~n613 & n707 ;
  assign n709 = ~n706 & ~n708 ;
  assign n710 = ~n679 & ~n704 ;
  assign n711 = ~n613 & n710 ;
  assign n712 = n679 & ~n704 ;
  assign n713 = n613 & n712 ;
  assign n714 = ~n711 & ~n713 ;
  assign n715 = n709 & n714 ;
  assign n716 = n612 & n715 ;
  assign n717 = ~n612 & ~n715 ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = n714 & ~n716 ;
  assign n720 = ~n584 & n685 ;
  assign n721 = ~n681 & n720 ;
  assign n722 = ~n684 & ~n721 ;
  assign n723 = ~\b[10]  & ~\b[11]  ;
  assign n724 = \b[10]  & \b[11]  ;
  assign n725 = ~n723 & ~n724 ;
  assign n726 = ~n722 & n725 ;
  assign n727 = ~n684 & ~n725 ;
  assign n728 = ~n721 & n727 ;
  assign n729 = n134 & ~n728 ;
  assign n730 = ~n726 & n729 ;
  assign n731 = \a[0]  & \b[11]  ;
  assign n732 = n133 & n731 ;
  assign n733 = ~\a[0]  & \b[9]  ;
  assign n734 = n132 & n733 ;
  assign n735 = \b[10]  & n141 ;
  assign n736 = ~n734 & ~n735 ;
  assign n737 = ~n732 & n736 ;
  assign n738 = ~n730 & n737 ;
  assign n739 = ~\a[2]  & ~n738 ;
  assign n740 = \a[2]  & n737 ;
  assign n741 = ~n730 & n740 ;
  assign n742 = ~n739 & ~n741 ;
  assign n743 = ~n577 & ~n677 ;
  assign n744 = ~n581 & n743 ;
  assign n745 = ~n678 & ~n744 ;
  assign n746 = n252 & ~n508 ;
  assign n747 = ~n506 & n746 ;
  assign n748 = \b[6]  & n303 ;
  assign n749 = n300 & n748 ;
  assign n750 = \b[8]  & n250 ;
  assign n751 = \a[3]  & \b[7]  ;
  assign n752 = n241 & n751 ;
  assign n753 = ~\a[3]  & \b[7]  ;
  assign n754 = n244 & n753 ;
  assign n755 = ~n752 & ~n754 ;
  assign n756 = ~n750 & n755 ;
  assign n757 = ~n749 & n756 ;
  assign n758 = ~n747 & n757 ;
  assign n759 = ~\a[5]  & ~n758 ;
  assign n760 = \a[5]  & n757 ;
  assign n761 = ~n747 & n760 ;
  assign n762 = ~n759 & ~n761 ;
  assign n763 = ~n655 & ~n657 ;
  assign n764 = ~n273 & n430 ;
  assign n765 = ~n271 & n764 ;
  assign n766 = \b[3]  & n486 ;
  assign n767 = n483 & n766 ;
  assign n768 = \b[5]  & n428 ;
  assign n769 = \a[5]  & \b[4]  ;
  assign n770 = n484 & n769 ;
  assign n771 = ~\a[6]  & \b[4]  ;
  assign n772 = n422 & n771 ;
  assign n773 = ~n770 & ~n772 ;
  assign n774 = ~n768 & n773 ;
  assign n775 = ~n767 & n774 ;
  assign n776 = ~n765 & n775 ;
  assign n777 = ~\a[8]  & ~n776 ;
  assign n778 = \a[8]  & n775 ;
  assign n779 = ~n765 & n778 ;
  assign n780 = ~n777 & ~n779 ;
  assign n781 = \a[11]  & ~n552 ;
  assign n782 = n640 & n781 ;
  assign n783 = n648 & n782 ;
  assign n784 = \a[11]  & ~n783 ;
  assign n785 = \b[2]  & n644 ;
  assign n786 = ~\a[9]  & \b[1]  ;
  assign n787 = n638 & n786 ;
  assign n788 = \a[9]  & \b[1]  ;
  assign n789 = n635 & n788 ;
  assign n790 = ~n787 & ~n789 ;
  assign n791 = ~n785 & n790 ;
  assign n792 = n157 & n646 ;
  assign n793 = n551 & ~n643 ;
  assign n794 = \a[9]  & ~\a[10]  ;
  assign n795 = ~\a[9]  & \a[10]  ;
  assign n796 = ~n794 & ~n795 ;
  assign n797 = \b[0]  & n796 ;
  assign n798 = n793 & n797 ;
  assign n799 = ~n792 & ~n798 ;
  assign n800 = n791 & n799 ;
  assign n801 = ~n784 & ~n800 ;
  assign n802 = n784 & n800 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = ~n780 & ~n803 ;
  assign n805 = n780 & n803 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~n763 & n806 ;
  assign n808 = n763 & ~n806 ;
  assign n809 = ~n807 & ~n808 ;
  assign n810 = ~n762 & n809 ;
  assign n811 = n762 & ~n809 ;
  assign n812 = ~n810 & ~n811 ;
  assign n813 = n745 & n812 ;
  assign n814 = ~n745 & ~n812 ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = ~n742 & n815 ;
  assign n817 = n742 & ~n815 ;
  assign n818 = ~n816 & ~n817 ;
  assign n819 = ~n719 & n818 ;
  assign n820 = n719 & ~n818 ;
  assign n821 = ~n819 & ~n820 ;
  assign n822 = n714 & ~n816 ;
  assign n823 = ~n716 & n822 ;
  assign n824 = ~n817 & ~n823 ;
  assign n825 = ~n810 & ~n813 ;
  assign n826 = ~n655 & ~n804 ;
  assign n827 = ~n657 & n826 ;
  assign n828 = ~n805 & ~n827 ;
  assign n829 = n177 & n646 ;
  assign n830 = \b[3]  & n644 ;
  assign n831 = \a[8]  & \b[2]  ;
  assign n832 = n794 & n831 ;
  assign n833 = ~\a[9]  & \b[2]  ;
  assign n834 = n638 & n833 ;
  assign n835 = ~n832 & ~n834 ;
  assign n836 = ~n830 & n835 ;
  assign n837 = ~n829 & n836 ;
  assign n838 = \b[1]  & n796 ;
  assign n839 = n793 & n838 ;
  assign n840 = ~\a[11]  & ~n839 ;
  assign n841 = n837 & n840 ;
  assign n842 = n837 & ~n839 ;
  assign n843 = \a[11]  & ~n842 ;
  assign n844 = ~n841 & ~n843 ;
  assign n845 = \a[11]  & ~\a[12]  ;
  assign n846 = ~\a[11]  & \a[12]  ;
  assign n847 = ~n845 & ~n846 ;
  assign n848 = \b[0]  & ~n847 ;
  assign n849 = n783 & n800 ;
  assign n850 = n848 & n849 ;
  assign n851 = ~n848 & ~n849 ;
  assign n852 = ~n850 & ~n851 ;
  assign n853 = n844 & n852 ;
  assign n854 = ~n844 & ~n852 ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = ~n323 & ~n359 ;
  assign n857 = ~n427 & n856 ;
  assign n858 = n320 & n857 ;
  assign n859 = n323 & ~n359 ;
  assign n860 = ~n427 & n859 ;
  assign n861 = ~n320 & n860 ;
  assign n862 = ~n858 & ~n861 ;
  assign n863 = \b[4]  & n486 ;
  assign n864 = n483 & n863 ;
  assign n865 = \b[6]  & n428 ;
  assign n866 = \a[5]  & \b[5]  ;
  assign n867 = n484 & n866 ;
  assign n868 = ~\a[6]  & \b[5]  ;
  assign n869 = n422 & n868 ;
  assign n870 = ~n867 & ~n869 ;
  assign n871 = ~n865 & n870 ;
  assign n872 = ~n864 & n871 ;
  assign n873 = n862 & n872 ;
  assign n874 = ~\a[8]  & ~n873 ;
  assign n875 = \a[8]  & n872 ;
  assign n876 = n862 & n875 ;
  assign n877 = ~n874 & ~n876 ;
  assign n878 = n855 & ~n877 ;
  assign n879 = ~n855 & n877 ;
  assign n880 = ~n878 & ~n879 ;
  assign n881 = ~n828 & ~n880 ;
  assign n882 = n828 & n880 ;
  assign n883 = ~n881 & ~n882 ;
  assign n884 = n252 & ~n589 ;
  assign n885 = ~n587 & n884 ;
  assign n886 = \b[7]  & n303 ;
  assign n887 = n300 & n886 ;
  assign n888 = \b[9]  & n250 ;
  assign n889 = \a[3]  & \b[8]  ;
  assign n890 = n241 & n889 ;
  assign n891 = ~\a[3]  & \b[8]  ;
  assign n892 = n244 & n891 ;
  assign n893 = ~n890 & ~n892 ;
  assign n894 = ~n888 & n893 ;
  assign n895 = ~n887 & n894 ;
  assign n896 = ~\a[5]  & n895 ;
  assign n897 = ~n885 & n896 ;
  assign n898 = ~n885 & n895 ;
  assign n899 = \a[5]  & ~n898 ;
  assign n900 = ~n897 & ~n899 ;
  assign n901 = ~n883 & ~n900 ;
  assign n902 = n883 & n900 ;
  assign n903 = ~n901 & ~n902 ;
  assign n904 = ~n684 & ~n724 ;
  assign n905 = ~n721 & n904 ;
  assign n906 = ~n723 & ~n905 ;
  assign n907 = ~\b[11]  & ~\b[12]  ;
  assign n908 = \b[11]  & \b[12]  ;
  assign n909 = ~n907 & ~n908 ;
  assign n910 = ~n906 & ~n909 ;
  assign n911 = ~n723 & n909 ;
  assign n912 = ~n905 & n911 ;
  assign n913 = n134 & ~n912 ;
  assign n914 = ~n910 & n913 ;
  assign n915 = \a[0]  & \b[12]  ;
  assign n916 = n133 & n915 ;
  assign n917 = ~\a[0]  & \b[10]  ;
  assign n918 = n132 & n917 ;
  assign n919 = \b[11]  & n141 ;
  assign n920 = ~n918 & ~n919 ;
  assign n921 = ~n916 & n920 ;
  assign n922 = ~n914 & n921 ;
  assign n923 = ~\a[2]  & ~n922 ;
  assign n924 = \a[2]  & n921 ;
  assign n925 = ~n914 & n924 ;
  assign n926 = ~n923 & ~n925 ;
  assign n927 = ~n903 & ~n926 ;
  assign n928 = ~n825 & n927 ;
  assign n929 = n903 & ~n926 ;
  assign n930 = n825 & n929 ;
  assign n931 = ~n928 & ~n930 ;
  assign n932 = n903 & n926 ;
  assign n933 = ~n825 & n932 ;
  assign n934 = ~n903 & n926 ;
  assign n935 = n825 & n934 ;
  assign n936 = ~n933 & ~n935 ;
  assign n937 = n931 & n936 ;
  assign n938 = n824 & n937 ;
  assign n939 = ~n824 & ~n937 ;
  assign n940 = ~n938 & ~n939 ;
  assign n941 = n931 & ~n938 ;
  assign n942 = ~n810 & ~n902 ;
  assign n943 = ~n813 & n942 ;
  assign n944 = ~n901 & ~n943 ;
  assign n945 = ~n908 & ~n912 ;
  assign n946 = ~\b[12]  & ~\b[13]  ;
  assign n947 = \b[12]  & \b[13]  ;
  assign n948 = ~n946 & ~n947 ;
  assign n949 = ~n945 & n948 ;
  assign n950 = ~n908 & ~n948 ;
  assign n951 = ~n912 & n950 ;
  assign n952 = n134 & ~n951 ;
  assign n953 = ~n949 & n952 ;
  assign n954 = \a[0]  & \b[13]  ;
  assign n955 = n133 & n954 ;
  assign n956 = ~\a[0]  & \b[11]  ;
  assign n957 = n132 & n956 ;
  assign n958 = \b[12]  & n141 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = ~n955 & n959 ;
  assign n961 = ~n953 & n960 ;
  assign n962 = ~\a[2]  & ~n961 ;
  assign n963 = \a[2]  & n960 ;
  assign n964 = ~n953 & n963 ;
  assign n965 = ~n962 & ~n964 ;
  assign n966 = ~n878 & ~n882 ;
  assign n967 = ~n850 & ~n853 ;
  assign n968 = n222 & n646 ;
  assign n969 = \b[4]  & n644 ;
  assign n970 = \a[8]  & \b[3]  ;
  assign n971 = n794 & n970 ;
  assign n972 = ~\a[9]  & \b[3]  ;
  assign n973 = n638 & n972 ;
  assign n974 = ~n971 & ~n973 ;
  assign n975 = ~n969 & n974 ;
  assign n976 = \b[2]  & n796 ;
  assign n977 = n793 & n976 ;
  assign n978 = \a[11]  & ~n977 ;
  assign n979 = n975 & n978 ;
  assign n980 = ~n968 & n979 ;
  assign n981 = n975 & ~n977 ;
  assign n982 = ~n968 & n981 ;
  assign n983 = ~\a[11]  & ~n982 ;
  assign n984 = ~n980 & ~n983 ;
  assign n985 = \a[14]  & \b[0]  ;
  assign n986 = ~n847 & n985 ;
  assign n987 = \a[12]  & \b[0]  ;
  assign n988 = \a[11]  & ~\a[13]  ;
  assign n989 = n987 & n988 ;
  assign n990 = ~\a[12]  & \b[0]  ;
  assign n991 = ~\a[11]  & \a[13]  ;
  assign n992 = n990 & n991 ;
  assign n993 = ~n989 & ~n992 ;
  assign n994 = \a[13]  & ~\a[14]  ;
  assign n995 = ~\a[13]  & \a[14]  ;
  assign n996 = ~n994 & ~n995 ;
  assign n997 = ~n847 & n996 ;
  assign n998 = \b[1]  & n997 ;
  assign n999 = ~n847 & ~n996 ;
  assign n1000 = ~n137 & n999 ;
  assign n1001 = ~n998 & ~n1000 ;
  assign n1002 = n993 & n1001 ;
  assign n1003 = n986 & ~n1002 ;
  assign n1004 = ~n986 & n993 ;
  assign n1005 = n1001 & n1004 ;
  assign n1006 = ~n1003 & ~n1005 ;
  assign n1007 = n984 & ~n1006 ;
  assign n1008 = ~n984 & n1006 ;
  assign n1009 = ~n1007 & ~n1008 ;
  assign n1010 = ~n967 & n1009 ;
  assign n1011 = n967 & ~n1009 ;
  assign n1012 = ~n1010 & ~n1011 ;
  assign n1013 = ~n383 & n430 ;
  assign n1014 = ~n381 & n1013 ;
  assign n1015 = \b[5]  & n486 ;
  assign n1016 = n483 & n1015 ;
  assign n1017 = \b[7]  & n428 ;
  assign n1018 = \a[5]  & \b[6]  ;
  assign n1019 = n484 & n1018 ;
  assign n1020 = ~\a[6]  & \b[6]  ;
  assign n1021 = n422 & n1020 ;
  assign n1022 = ~n1019 & ~n1021 ;
  assign n1023 = ~n1017 & n1022 ;
  assign n1024 = ~n1016 & n1023 ;
  assign n1025 = ~n1014 & n1024 ;
  assign n1026 = ~\a[8]  & ~n1025 ;
  assign n1027 = \a[8]  & n1024 ;
  assign n1028 = ~n1014 & n1027 ;
  assign n1029 = ~n1026 & ~n1028 ;
  assign n1030 = n1012 & ~n1029 ;
  assign n1031 = ~n1012 & n1029 ;
  assign n1032 = ~n1030 & ~n1031 ;
  assign n1033 = ~n682 & ~n685 ;
  assign n1034 = n252 & ~n721 ;
  assign n1035 = ~n1033 & n1034 ;
  assign n1036 = \b[8]  & n303 ;
  assign n1037 = n300 & n1036 ;
  assign n1038 = \b[10]  & n250 ;
  assign n1039 = \a[3]  & \b[9]  ;
  assign n1040 = n241 & n1039 ;
  assign n1041 = ~\a[3]  & \b[9]  ;
  assign n1042 = n244 & n1041 ;
  assign n1043 = ~n1040 & ~n1042 ;
  assign n1044 = ~n1038 & n1043 ;
  assign n1045 = ~n1037 & n1044 ;
  assign n1046 = ~n1035 & n1045 ;
  assign n1047 = ~\a[5]  & ~n1046 ;
  assign n1048 = \a[5]  & n1045 ;
  assign n1049 = ~n1035 & n1048 ;
  assign n1050 = ~n1047 & ~n1049 ;
  assign n1051 = ~n1032 & ~n1050 ;
  assign n1052 = ~n966 & n1051 ;
  assign n1053 = n1032 & ~n1050 ;
  assign n1054 = n966 & n1053 ;
  assign n1055 = ~n1052 & ~n1054 ;
  assign n1056 = ~n1032 & n1050 ;
  assign n1057 = n966 & n1056 ;
  assign n1058 = n1032 & n1050 ;
  assign n1059 = ~n966 & n1058 ;
  assign n1060 = ~n1057 & ~n1059 ;
  assign n1061 = n1055 & n1060 ;
  assign n1062 = ~n965 & ~n1061 ;
  assign n1063 = n944 & n1062 ;
  assign n1064 = ~n965 & n1061 ;
  assign n1065 = ~n944 & n1064 ;
  assign n1066 = ~n1063 & ~n1065 ;
  assign n1067 = n965 & ~n1061 ;
  assign n1068 = ~n944 & n1067 ;
  assign n1069 = n965 & n1061 ;
  assign n1070 = n944 & n1069 ;
  assign n1071 = ~n1068 & ~n1070 ;
  assign n1072 = n1066 & n1071 ;
  assign n1073 = ~n941 & n1072 ;
  assign n1074 = n931 & ~n1072 ;
  assign n1075 = ~n938 & n1074 ;
  assign n1076 = ~n1073 & ~n1075 ;
  assign n1077 = n931 & n1066 ;
  assign n1078 = ~n938 & n1077 ;
  assign n1079 = n1071 & ~n1078 ;
  assign n1080 = n944 & n1061 ;
  assign n1081 = n1055 & ~n1080 ;
  assign n1082 = ~n908 & ~n947 ;
  assign n1083 = ~n912 & n1082 ;
  assign n1084 = ~n946 & ~n1083 ;
  assign n1085 = ~\b[13]  & ~\b[14]  ;
  assign n1086 = \b[13]  & \b[14]  ;
  assign n1087 = ~n1085 & ~n1086 ;
  assign n1088 = n134 & n1087 ;
  assign n1089 = ~n1084 & n1088 ;
  assign n1090 = n134 & ~n1087 ;
  assign n1091 = ~n946 & n1090 ;
  assign n1092 = ~n1083 & n1091 ;
  assign n1093 = \a[0]  & \b[14]  ;
  assign n1094 = n133 & n1093 ;
  assign n1095 = ~\a[0]  & \b[12]  ;
  assign n1096 = n132 & n1095 ;
  assign n1097 = \b[13]  & n141 ;
  assign n1098 = ~n1096 & ~n1097 ;
  assign n1099 = ~n1094 & n1098 ;
  assign n1100 = ~n1092 & n1099 ;
  assign n1101 = ~n1089 & n1100 ;
  assign n1102 = ~\a[2]  & ~n1101 ;
  assign n1103 = \a[2]  & n1099 ;
  assign n1104 = ~n1092 & n1103 ;
  assign n1105 = ~n1089 & n1104 ;
  assign n1106 = ~n1102 & ~n1105 ;
  assign n1107 = n252 & ~n728 ;
  assign n1108 = ~n726 & n1107 ;
  assign n1109 = \b[9]  & n303 ;
  assign n1110 = n300 & n1109 ;
  assign n1111 = \b[11]  & n250 ;
  assign n1112 = \a[3]  & \b[10]  ;
  assign n1113 = n241 & n1112 ;
  assign n1114 = ~\a[3]  & \b[10]  ;
  assign n1115 = n244 & n1114 ;
  assign n1116 = ~n1113 & ~n1115 ;
  assign n1117 = ~n1111 & n1116 ;
  assign n1118 = ~n1110 & n1117 ;
  assign n1119 = ~\a[5]  & n1118 ;
  assign n1120 = ~n1108 & n1119 ;
  assign n1121 = ~n1108 & n1118 ;
  assign n1122 = \a[5]  & ~n1121 ;
  assign n1123 = ~n1120 & ~n1122 ;
  assign n1124 = ~n878 & ~n1030 ;
  assign n1125 = ~n882 & n1124 ;
  assign n1126 = ~n1031 & ~n1125 ;
  assign n1127 = n430 & ~n508 ;
  assign n1128 = ~n506 & n1127 ;
  assign n1129 = \b[6]  & n486 ;
  assign n1130 = n483 & n1129 ;
  assign n1131 = \b[8]  & n428 ;
  assign n1132 = \a[5]  & \b[7]  ;
  assign n1133 = n484 & n1132 ;
  assign n1134 = ~\a[6]  & \b[7]  ;
  assign n1135 = n422 & n1134 ;
  assign n1136 = ~n1133 & ~n1135 ;
  assign n1137 = ~n1131 & n1136 ;
  assign n1138 = ~n1130 & n1137 ;
  assign n1139 = ~n1128 & n1138 ;
  assign n1140 = ~\a[8]  & ~n1139 ;
  assign n1141 = \a[8]  & n1138 ;
  assign n1142 = ~n1128 & n1141 ;
  assign n1143 = ~n1140 & ~n1142 ;
  assign n1144 = ~n1008 & ~n1010 ;
  assign n1145 = ~n270 & n646 ;
  assign n1146 = ~n218 & n646 ;
  assign n1147 = ~n220 & n1146 ;
  assign n1148 = ~n1145 & ~n1147 ;
  assign n1149 = ~n273 & ~n1148 ;
  assign n1150 = \b[3]  & n796 ;
  assign n1151 = n793 & n1150 ;
  assign n1152 = \b[5]  & n644 ;
  assign n1153 = \a[9]  & \b[4]  ;
  assign n1154 = n635 & n1153 ;
  assign n1155 = ~\a[9]  & \b[4]  ;
  assign n1156 = n638 & n1155 ;
  assign n1157 = ~n1154 & ~n1156 ;
  assign n1158 = ~n1152 & n1157 ;
  assign n1159 = ~n1151 & n1158 ;
  assign n1160 = ~\a[11]  & n1159 ;
  assign n1161 = ~n1149 & n1160 ;
  assign n1162 = \a[11]  & ~n1159 ;
  assign n1163 = \a[11]  & ~n273 ;
  assign n1164 = ~n1148 & n1163 ;
  assign n1165 = ~n1162 & ~n1164 ;
  assign n1166 = ~n1161 & n1165 ;
  assign n1167 = \a[14]  & ~n848 ;
  assign n1168 = n993 & n1167 ;
  assign n1169 = n1001 & n1168 ;
  assign n1170 = \a[14]  & ~n1169 ;
  assign n1171 = \b[2]  & n997 ;
  assign n1172 = ~\a[12]  & \b[1]  ;
  assign n1173 = n991 & n1172 ;
  assign n1174 = \a[12]  & \b[1]  ;
  assign n1175 = n988 & n1174 ;
  assign n1176 = ~n1173 & ~n1175 ;
  assign n1177 = ~n1171 & n1176 ;
  assign n1178 = n157 & n999 ;
  assign n1179 = n847 & ~n996 ;
  assign n1180 = \a[12]  & ~\a[13]  ;
  assign n1181 = ~\a[12]  & \a[13]  ;
  assign n1182 = ~n1180 & ~n1181 ;
  assign n1183 = \b[0]  & n1182 ;
  assign n1184 = n1179 & n1183 ;
  assign n1185 = ~n1178 & ~n1184 ;
  assign n1186 = n1177 & n1185 ;
  assign n1187 = ~n1170 & ~n1186 ;
  assign n1188 = n1170 & n1186 ;
  assign n1189 = ~n1187 & ~n1188 ;
  assign n1190 = n1166 & ~n1189 ;
  assign n1191 = ~n1166 & n1189 ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1193 = ~n1144 & n1192 ;
  assign n1194 = ~n1008 & ~n1192 ;
  assign n1195 = ~n1010 & n1194 ;
  assign n1196 = ~n1193 & ~n1195 ;
  assign n1197 = n1143 & ~n1196 ;
  assign n1198 = ~n1143 & ~n1195 ;
  assign n1199 = ~n1193 & n1198 ;
  assign n1200 = ~n1197 & ~n1199 ;
  assign n1201 = n1126 & n1200 ;
  assign n1202 = ~n1126 & ~n1200 ;
  assign n1203 = ~n1201 & ~n1202 ;
  assign n1204 = ~n1123 & ~n1203 ;
  assign n1205 = n1123 & n1203 ;
  assign n1206 = ~n1204 & ~n1205 ;
  assign n1207 = ~n1106 & ~n1206 ;
  assign n1208 = ~n1081 & n1207 ;
  assign n1209 = ~n1106 & n1206 ;
  assign n1210 = n1081 & n1209 ;
  assign n1211 = ~n1208 & ~n1210 ;
  assign n1212 = n1106 & ~n1206 ;
  assign n1213 = n1081 & n1212 ;
  assign n1214 = n1106 & n1206 ;
  assign n1215 = ~n1081 & n1214 ;
  assign n1216 = ~n1213 & ~n1215 ;
  assign n1217 = n1211 & n1216 ;
  assign n1218 = n1079 & n1217 ;
  assign n1219 = ~n1079 & ~n1217 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = n1211 & ~n1218 ;
  assign n1222 = n1055 & ~n1205 ;
  assign n1223 = ~n1080 & n1222 ;
  assign n1224 = ~n1204 & ~n1223 ;
  assign n1225 = ~n946 & n1087 ;
  assign n1226 = ~n1083 & n1225 ;
  assign n1227 = ~n1086 & ~n1226 ;
  assign n1228 = ~\b[14]  & ~\b[15]  ;
  assign n1229 = \b[14]  & \b[15]  ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = ~n1227 & n1230 ;
  assign n1232 = ~n1086 & ~n1230 ;
  assign n1233 = ~n1226 & n1232 ;
  assign n1234 = n134 & ~n1233 ;
  assign n1235 = ~n1231 & n1234 ;
  assign n1236 = \a[0]  & \b[15]  ;
  assign n1237 = n133 & n1236 ;
  assign n1238 = ~\a[0]  & \b[13]  ;
  assign n1239 = n132 & n1238 ;
  assign n1240 = \b[14]  & n141 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = ~n1237 & n1241 ;
  assign n1243 = ~n1235 & n1242 ;
  assign n1244 = ~\a[2]  & ~n1243 ;
  assign n1245 = \a[2]  & n1242 ;
  assign n1246 = ~n1235 & n1245 ;
  assign n1247 = ~n1244 & ~n1246 ;
  assign n1248 = ~n1199 & ~n1201 ;
  assign n1249 = n252 & ~n912 ;
  assign n1250 = ~n910 & n1249 ;
  assign n1251 = \b[10]  & n303 ;
  assign n1252 = n300 & n1251 ;
  assign n1253 = \b[12]  & n250 ;
  assign n1254 = \a[3]  & \b[11]  ;
  assign n1255 = n241 & n1254 ;
  assign n1256 = ~\a[3]  & \b[11]  ;
  assign n1257 = n244 & n1256 ;
  assign n1258 = ~n1255 & ~n1257 ;
  assign n1259 = ~n1253 & n1258 ;
  assign n1260 = ~n1252 & n1259 ;
  assign n1261 = ~n1250 & n1260 ;
  assign n1262 = ~\a[5]  & ~n1261 ;
  assign n1263 = \a[5]  & n1260 ;
  assign n1264 = ~n1250 & n1263 ;
  assign n1265 = ~n1262 & ~n1264 ;
  assign n1266 = n430 & ~n589 ;
  assign n1267 = ~n587 & n1266 ;
  assign n1268 = \b[7]  & n486 ;
  assign n1269 = n483 & n1268 ;
  assign n1270 = \b[9]  & n428 ;
  assign n1271 = \a[5]  & \b[8]  ;
  assign n1272 = n484 & n1271 ;
  assign n1273 = ~\a[6]  & \b[8]  ;
  assign n1274 = n422 & n1273 ;
  assign n1275 = ~n1272 & ~n1274 ;
  assign n1276 = ~n1270 & n1275 ;
  assign n1277 = ~n1269 & n1276 ;
  assign n1278 = ~\a[8]  & n1277 ;
  assign n1279 = ~n1267 & n1278 ;
  assign n1280 = ~n1267 & n1277 ;
  assign n1281 = \a[8]  & ~n1280 ;
  assign n1282 = ~n1279 & ~n1281 ;
  assign n1283 = ~n1008 & ~n1190 ;
  assign n1284 = ~n1010 & n1283 ;
  assign n1285 = ~n1191 & ~n1284 ;
  assign n1286 = n177 & n999 ;
  assign n1287 = \b[3]  & n997 ;
  assign n1288 = \a[11]  & \b[2]  ;
  assign n1289 = n1180 & n1288 ;
  assign n1290 = ~\a[12]  & \b[2]  ;
  assign n1291 = n991 & n1290 ;
  assign n1292 = ~n1289 & ~n1291 ;
  assign n1293 = ~n1287 & n1292 ;
  assign n1294 = ~n1286 & n1293 ;
  assign n1295 = \b[1]  & n1182 ;
  assign n1296 = n1179 & n1295 ;
  assign n1297 = ~\a[14]  & ~n1296 ;
  assign n1298 = n1294 & n1297 ;
  assign n1299 = n1294 & ~n1296 ;
  assign n1300 = \a[14]  & ~n1299 ;
  assign n1301 = ~n1298 & ~n1300 ;
  assign n1302 = \a[14]  & ~\a[15]  ;
  assign n1303 = ~\a[14]  & \a[15]  ;
  assign n1304 = ~n1302 & ~n1303 ;
  assign n1305 = \b[0]  & ~n1304 ;
  assign n1306 = n1169 & n1186 ;
  assign n1307 = n1305 & n1306 ;
  assign n1308 = ~n1305 & ~n1306 ;
  assign n1309 = ~n1307 & ~n1308 ;
  assign n1310 = n1301 & n1309 ;
  assign n1311 = ~n1301 & ~n1309 ;
  assign n1312 = ~n1310 & ~n1311 ;
  assign n1313 = ~n323 & ~n551 ;
  assign n1314 = ~n643 & n1313 ;
  assign n1315 = n320 & n1314 ;
  assign n1316 = n323 & ~n551 ;
  assign n1317 = ~n643 & n1316 ;
  assign n1318 = ~n320 & n1317 ;
  assign n1319 = ~n1315 & ~n1318 ;
  assign n1320 = \b[4]  & n796 ;
  assign n1321 = n793 & n1320 ;
  assign n1322 = \b[6]  & n644 ;
  assign n1323 = \a[9]  & \b[5]  ;
  assign n1324 = n635 & n1323 ;
  assign n1325 = ~\a[9]  & \b[5]  ;
  assign n1326 = n638 & n1325 ;
  assign n1327 = ~n1324 & ~n1326 ;
  assign n1328 = ~n1322 & n1327 ;
  assign n1329 = ~n1321 & n1328 ;
  assign n1330 = n1319 & n1329 ;
  assign n1331 = ~\a[11]  & ~n1330 ;
  assign n1332 = \a[11]  & n1329 ;
  assign n1333 = n1319 & n1332 ;
  assign n1334 = ~n1331 & ~n1333 ;
  assign n1335 = n1312 & ~n1334 ;
  assign n1336 = ~n1312 & n1334 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = n1285 & n1337 ;
  assign n1339 = ~n1285 & ~n1337 ;
  assign n1340 = ~n1338 & ~n1339 ;
  assign n1341 = n1282 & n1340 ;
  assign n1342 = ~n1282 & ~n1340 ;
  assign n1343 = ~n1341 & ~n1342 ;
  assign n1344 = ~n1265 & ~n1343 ;
  assign n1345 = ~n1248 & n1344 ;
  assign n1346 = ~n1265 & n1343 ;
  assign n1347 = n1248 & n1346 ;
  assign n1348 = ~n1345 & ~n1347 ;
  assign n1349 = n1265 & ~n1343 ;
  assign n1350 = n1248 & n1349 ;
  assign n1351 = n1265 & n1343 ;
  assign n1352 = ~n1248 & n1351 ;
  assign n1353 = ~n1350 & ~n1352 ;
  assign n1354 = n1348 & n1353 ;
  assign n1355 = ~n1247 & ~n1354 ;
  assign n1356 = n1224 & n1355 ;
  assign n1357 = ~n1247 & n1354 ;
  assign n1358 = ~n1224 & n1357 ;
  assign n1359 = ~n1356 & ~n1358 ;
  assign n1360 = n1247 & ~n1354 ;
  assign n1361 = ~n1224 & n1360 ;
  assign n1362 = n1247 & n1354 ;
  assign n1363 = n1224 & n1362 ;
  assign n1364 = ~n1361 & ~n1363 ;
  assign n1365 = n1359 & n1364 ;
  assign n1366 = ~n1221 & n1365 ;
  assign n1367 = n1211 & ~n1365 ;
  assign n1368 = ~n1218 & n1367 ;
  assign n1369 = ~n1366 & ~n1368 ;
  assign n1370 = n1211 & n1359 ;
  assign n1371 = ~n1218 & n1370 ;
  assign n1372 = n1364 & ~n1371 ;
  assign n1373 = n1224 & n1354 ;
  assign n1374 = n1348 & ~n1373 ;
  assign n1375 = ~n1199 & ~n1341 ;
  assign n1376 = ~n1201 & n1375 ;
  assign n1377 = ~n1342 & ~n1376 ;
  assign n1378 = n252 & ~n951 ;
  assign n1379 = ~n949 & n1378 ;
  assign n1380 = \b[11]  & n303 ;
  assign n1381 = n300 & n1380 ;
  assign n1382 = \b[13]  & n250 ;
  assign n1383 = \a[3]  & \b[12]  ;
  assign n1384 = n241 & n1383 ;
  assign n1385 = ~\a[3]  & \b[12]  ;
  assign n1386 = n244 & n1385 ;
  assign n1387 = ~n1384 & ~n1386 ;
  assign n1388 = ~n1382 & n1387 ;
  assign n1389 = ~n1381 & n1388 ;
  assign n1390 = ~\a[5]  & n1389 ;
  assign n1391 = ~n1379 & n1390 ;
  assign n1392 = ~n1379 & n1389 ;
  assign n1393 = \a[5]  & ~n1392 ;
  assign n1394 = ~n1391 & ~n1393 ;
  assign n1395 = ~n1335 & ~n1338 ;
  assign n1396 = n430 & ~n721 ;
  assign n1397 = ~n1033 & n1396 ;
  assign n1398 = \b[8]  & n486 ;
  assign n1399 = n483 & n1398 ;
  assign n1400 = \b[10]  & n428 ;
  assign n1401 = \a[5]  & \b[9]  ;
  assign n1402 = n484 & n1401 ;
  assign n1403 = ~\a[6]  & \b[9]  ;
  assign n1404 = n422 & n1403 ;
  assign n1405 = ~n1402 & ~n1404 ;
  assign n1406 = ~n1400 & n1405 ;
  assign n1407 = ~n1399 & n1406 ;
  assign n1408 = ~n1397 & n1407 ;
  assign n1409 = ~\a[8]  & ~n1408 ;
  assign n1410 = \a[8]  & n1407 ;
  assign n1411 = ~n1397 & n1410 ;
  assign n1412 = ~n1409 & ~n1411 ;
  assign n1413 = ~n380 & n646 ;
  assign n1414 = ~n322 & n646 ;
  assign n1415 = ~n326 & n1414 ;
  assign n1416 = ~n1413 & ~n1415 ;
  assign n1417 = ~n383 & ~n1416 ;
  assign n1418 = \b[5]  & n796 ;
  assign n1419 = n793 & n1418 ;
  assign n1420 = \b[7]  & n644 ;
  assign n1421 = \a[9]  & \b[6]  ;
  assign n1422 = n635 & n1421 ;
  assign n1423 = ~\a[9]  & \b[6]  ;
  assign n1424 = n638 & n1423 ;
  assign n1425 = ~n1422 & ~n1424 ;
  assign n1426 = ~n1420 & n1425 ;
  assign n1427 = ~n1419 & n1426 ;
  assign n1428 = ~\a[11]  & n1427 ;
  assign n1429 = ~n1417 & n1428 ;
  assign n1430 = \a[11]  & ~n1427 ;
  assign n1431 = \a[11]  & ~n383 ;
  assign n1432 = ~n1416 & n1431 ;
  assign n1433 = ~n1430 & ~n1432 ;
  assign n1434 = ~n1429 & n1433 ;
  assign n1435 = ~n1307 & ~n1310 ;
  assign n1436 = n222 & n999 ;
  assign n1437 = \b[4]  & n997 ;
  assign n1438 = \a[11]  & \b[3]  ;
  assign n1439 = n1180 & n1438 ;
  assign n1440 = ~\a[12]  & \b[3]  ;
  assign n1441 = n991 & n1440 ;
  assign n1442 = ~n1439 & ~n1441 ;
  assign n1443 = ~n1437 & n1442 ;
  assign n1444 = \b[2]  & n1182 ;
  assign n1445 = n1179 & n1444 ;
  assign n1446 = \a[14]  & ~n1445 ;
  assign n1447 = n1443 & n1446 ;
  assign n1448 = ~n1436 & n1447 ;
  assign n1449 = n1443 & ~n1445 ;
  assign n1450 = ~n1436 & n1449 ;
  assign n1451 = ~\a[14]  & ~n1450 ;
  assign n1452 = ~n1448 & ~n1451 ;
  assign n1453 = \a[17]  & \b[0]  ;
  assign n1454 = ~n1304 & n1453 ;
  assign n1455 = \a[15]  & \b[0]  ;
  assign n1456 = \a[14]  & ~\a[16]  ;
  assign n1457 = n1455 & n1456 ;
  assign n1458 = ~\a[15]  & \b[0]  ;
  assign n1459 = ~\a[14]  & \a[16]  ;
  assign n1460 = n1458 & n1459 ;
  assign n1461 = ~n1457 & ~n1460 ;
  assign n1462 = \a[16]  & ~\a[17]  ;
  assign n1463 = ~\a[16]  & \a[17]  ;
  assign n1464 = ~n1462 & ~n1463 ;
  assign n1465 = ~n1304 & n1464 ;
  assign n1466 = \b[1]  & n1465 ;
  assign n1467 = ~n1304 & ~n1464 ;
  assign n1468 = ~n137 & n1467 ;
  assign n1469 = ~n1466 & ~n1468 ;
  assign n1470 = n1461 & n1469 ;
  assign n1471 = ~n1454 & ~n1470 ;
  assign n1472 = n1454 & n1461 ;
  assign n1473 = n1469 & n1472 ;
  assign n1474 = ~n1471 & ~n1473 ;
  assign n1475 = n1452 & n1474 ;
  assign n1476 = ~n1452 & ~n1474 ;
  assign n1477 = ~n1475 & ~n1476 ;
  assign n1478 = ~n1435 & n1477 ;
  assign n1479 = n1435 & ~n1477 ;
  assign n1480 = ~n1478 & ~n1479 ;
  assign n1481 = ~n1434 & ~n1480 ;
  assign n1482 = n1434 & n1480 ;
  assign n1483 = ~n1481 & ~n1482 ;
  assign n1484 = n1412 & ~n1483 ;
  assign n1485 = n1395 & n1484 ;
  assign n1486 = n1412 & n1483 ;
  assign n1487 = ~n1395 & n1486 ;
  assign n1488 = ~n1485 & ~n1487 ;
  assign n1489 = ~n1412 & ~n1483 ;
  assign n1490 = ~n1395 & n1489 ;
  assign n1491 = ~n1412 & n1483 ;
  assign n1492 = n1395 & n1491 ;
  assign n1493 = ~n1490 & ~n1492 ;
  assign n1494 = n1488 & n1493 ;
  assign n1495 = ~n1394 & ~n1494 ;
  assign n1496 = ~n1377 & n1495 ;
  assign n1497 = ~n1394 & n1494 ;
  assign n1498 = n1377 & n1497 ;
  assign n1499 = ~n1496 & ~n1498 ;
  assign n1500 = n1394 & ~n1494 ;
  assign n1501 = n1377 & n1500 ;
  assign n1502 = n1394 & n1494 ;
  assign n1503 = ~n1377 & n1502 ;
  assign n1504 = ~n1501 & ~n1503 ;
  assign n1505 = n1499 & n1504 ;
  assign n1506 = ~n1374 & n1505 ;
  assign n1507 = ~n1086 & ~n1229 ;
  assign n1508 = ~n1226 & n1507 ;
  assign n1509 = ~n1228 & ~n1508 ;
  assign n1510 = ~\b[15]  & ~\b[16]  ;
  assign n1511 = \b[15]  & \b[16]  ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = ~n1509 & ~n1512 ;
  assign n1514 = ~n1228 & n1512 ;
  assign n1515 = ~n1508 & n1514 ;
  assign n1516 = n134 & ~n1515 ;
  assign n1517 = ~n1513 & n1516 ;
  assign n1518 = \a[0]  & \b[16]  ;
  assign n1519 = n133 & n1518 ;
  assign n1520 = \b[15]  & n141 ;
  assign n1521 = ~\a[0]  & \a[2]  ;
  assign n1522 = ~\a[1]  & \b[14]  ;
  assign n1523 = n1521 & n1522 ;
  assign n1524 = ~n1520 & ~n1523 ;
  assign n1525 = ~n1519 & n1524 ;
  assign n1526 = \a[2]  & n1525 ;
  assign n1527 = ~n1517 & n1526 ;
  assign n1528 = ~n1517 & n1525 ;
  assign n1529 = ~\a[2]  & ~n1528 ;
  assign n1530 = ~n1527 & ~n1529 ;
  assign n1531 = n1348 & ~n1505 ;
  assign n1532 = ~n1373 & n1531 ;
  assign n1533 = ~n1530 & ~n1532 ;
  assign n1534 = ~n1506 & n1533 ;
  assign n1535 = ~n1505 & n1530 ;
  assign n1536 = n1374 & n1535 ;
  assign n1537 = n1505 & n1530 ;
  assign n1538 = ~n1374 & n1537 ;
  assign n1539 = ~n1536 & ~n1538 ;
  assign n1540 = ~n1534 & n1539 ;
  assign n1541 = n1372 & n1540 ;
  assign n1542 = ~n1372 & ~n1540 ;
  assign n1543 = ~n1541 & ~n1542 ;
  assign n1544 = ~n1534 & ~n1541 ;
  assign n1545 = n1348 & n1504 ;
  assign n1546 = ~n1373 & n1545 ;
  assign n1547 = n1499 & ~n1546 ;
  assign n1548 = n1377 & n1494 ;
  assign n1549 = n1493 & ~n1548 ;
  assign n1550 = n252 & n1087 ;
  assign n1551 = ~n1084 & n1550 ;
  assign n1552 = ~n946 & ~n1087 ;
  assign n1553 = n252 & n1552 ;
  assign n1554 = ~n1083 & n1553 ;
  assign n1555 = \b[12]  & n303 ;
  assign n1556 = n300 & n1555 ;
  assign n1557 = \b[14]  & n250 ;
  assign n1558 = \a[3]  & \b[13]  ;
  assign n1559 = n241 & n1558 ;
  assign n1560 = ~\a[3]  & \b[13]  ;
  assign n1561 = n244 & n1560 ;
  assign n1562 = ~n1559 & ~n1561 ;
  assign n1563 = ~n1557 & n1562 ;
  assign n1564 = ~n1556 & n1563 ;
  assign n1565 = ~n1554 & n1564 ;
  assign n1566 = ~n1551 & n1565 ;
  assign n1567 = ~\a[5]  & ~n1566 ;
  assign n1568 = \a[5]  & n1564 ;
  assign n1569 = ~n1554 & n1568 ;
  assign n1570 = ~n1551 & n1569 ;
  assign n1571 = ~n1567 & ~n1570 ;
  assign n1572 = n430 & ~n728 ;
  assign n1573 = ~n726 & n1572 ;
  assign n1574 = \b[9]  & n486 ;
  assign n1575 = n483 & n1574 ;
  assign n1576 = \b[11]  & n428 ;
  assign n1577 = \a[5]  & \b[10]  ;
  assign n1578 = n484 & n1577 ;
  assign n1579 = ~\a[6]  & \b[10]  ;
  assign n1580 = n422 & n1579 ;
  assign n1581 = ~n1578 & ~n1580 ;
  assign n1582 = ~n1576 & n1581 ;
  assign n1583 = ~n1575 & n1582 ;
  assign n1584 = ~\a[8]  & n1583 ;
  assign n1585 = ~n1573 & n1584 ;
  assign n1586 = ~n1573 & n1583 ;
  assign n1587 = \a[8]  & ~n1586 ;
  assign n1588 = ~n1585 & ~n1587 ;
  assign n1589 = ~n1335 & ~n1482 ;
  assign n1590 = ~n1338 & n1589 ;
  assign n1591 = ~n1481 & ~n1590 ;
  assign n1592 = ~n505 & ~n551 ;
  assign n1593 = ~n643 & n1592 ;
  assign n1594 = n502 & n1593 ;
  assign n1595 = n505 & ~n551 ;
  assign n1596 = ~n643 & n1595 ;
  assign n1597 = ~n502 & n1596 ;
  assign n1598 = ~n1594 & ~n1597 ;
  assign n1599 = \b[6]  & n796 ;
  assign n1600 = n793 & n1599 ;
  assign n1601 = \b[8]  & n644 ;
  assign n1602 = \a[9]  & \b[7]  ;
  assign n1603 = n635 & n1602 ;
  assign n1604 = ~\a[9]  & \b[7]  ;
  assign n1605 = n638 & n1604 ;
  assign n1606 = ~n1603 & ~n1605 ;
  assign n1607 = ~n1601 & n1606 ;
  assign n1608 = ~n1600 & n1607 ;
  assign n1609 = n1598 & n1608 ;
  assign n1610 = ~\a[11]  & ~n1609 ;
  assign n1611 = \a[11]  & n1608 ;
  assign n1612 = n1598 & n1611 ;
  assign n1613 = ~n1610 & ~n1612 ;
  assign n1614 = ~n1476 & ~n1478 ;
  assign n1615 = ~n270 & n999 ;
  assign n1616 = ~n218 & n999 ;
  assign n1617 = ~n220 & n1616 ;
  assign n1618 = ~n1615 & ~n1617 ;
  assign n1619 = ~n273 & ~n1618 ;
  assign n1620 = \b[3]  & n1182 ;
  assign n1621 = n1179 & n1620 ;
  assign n1622 = \b[5]  & n997 ;
  assign n1623 = \a[11]  & \b[4]  ;
  assign n1624 = n1180 & n1623 ;
  assign n1625 = ~\a[12]  & \b[4]  ;
  assign n1626 = n991 & n1625 ;
  assign n1627 = ~n1624 & ~n1626 ;
  assign n1628 = ~n1622 & n1627 ;
  assign n1629 = ~n1621 & n1628 ;
  assign n1630 = ~\a[14]  & n1629 ;
  assign n1631 = ~n1619 & n1630 ;
  assign n1632 = \a[14]  & ~n1629 ;
  assign n1633 = \a[14]  & ~n273 ;
  assign n1634 = ~n1618 & n1633 ;
  assign n1635 = ~n1632 & ~n1634 ;
  assign n1636 = ~n1631 & n1635 ;
  assign n1637 = \a[17]  & ~n1305 ;
  assign n1638 = n1461 & n1637 ;
  assign n1639 = n1469 & n1638 ;
  assign n1640 = \a[17]  & ~n1639 ;
  assign n1641 = \b[2]  & n1465 ;
  assign n1642 = ~\a[15]  & \b[1]  ;
  assign n1643 = n1459 & n1642 ;
  assign n1644 = \a[15]  & \b[1]  ;
  assign n1645 = n1456 & n1644 ;
  assign n1646 = ~n1643 & ~n1645 ;
  assign n1647 = ~n1641 & n1646 ;
  assign n1648 = n157 & n1467 ;
  assign n1649 = n1304 & ~n1464 ;
  assign n1650 = \a[15]  & ~\a[16]  ;
  assign n1651 = ~\a[15]  & \a[16]  ;
  assign n1652 = ~n1650 & ~n1651 ;
  assign n1653 = \b[0]  & n1652 ;
  assign n1654 = n1649 & n1653 ;
  assign n1655 = ~n1648 & ~n1654 ;
  assign n1656 = n1647 & n1655 ;
  assign n1657 = ~n1640 & ~n1656 ;
  assign n1658 = n1640 & n1656 ;
  assign n1659 = ~n1657 & ~n1658 ;
  assign n1660 = n1636 & ~n1659 ;
  assign n1661 = ~n1636 & n1659 ;
  assign n1662 = ~n1660 & ~n1661 ;
  assign n1663 = ~n1614 & n1662 ;
  assign n1664 = ~n1476 & ~n1662 ;
  assign n1665 = ~n1478 & n1664 ;
  assign n1666 = ~n1663 & ~n1665 ;
  assign n1667 = n1613 & ~n1666 ;
  assign n1668 = ~n1613 & ~n1665 ;
  assign n1669 = ~n1663 & n1668 ;
  assign n1670 = ~n1667 & ~n1669 ;
  assign n1671 = n1591 & n1670 ;
  assign n1672 = ~n1591 & ~n1670 ;
  assign n1673 = ~n1671 & ~n1672 ;
  assign n1674 = ~n1588 & ~n1673 ;
  assign n1675 = n1588 & n1673 ;
  assign n1676 = ~n1674 & ~n1675 ;
  assign n1677 = n1571 & ~n1676 ;
  assign n1678 = n1549 & n1677 ;
  assign n1679 = n1571 & n1676 ;
  assign n1680 = ~n1549 & n1679 ;
  assign n1681 = ~n1678 & ~n1680 ;
  assign n1682 = ~n1571 & ~n1676 ;
  assign n1683 = ~n1549 & n1682 ;
  assign n1684 = ~n1571 & n1676 ;
  assign n1685 = n1549 & n1684 ;
  assign n1686 = ~n1683 & ~n1685 ;
  assign n1687 = n1681 & n1686 ;
  assign n1688 = ~n1511 & ~n1515 ;
  assign n1689 = ~\b[16]  & ~\b[17]  ;
  assign n1690 = \b[16]  & \b[17]  ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = ~n1688 & n1691 ;
  assign n1693 = ~n1511 & ~n1691 ;
  assign n1694 = ~n1515 & n1693 ;
  assign n1695 = n134 & ~n1694 ;
  assign n1696 = ~n1692 & n1695 ;
  assign n1697 = \a[0]  & \b[17]  ;
  assign n1698 = n133 & n1697 ;
  assign n1699 = \b[16]  & n141 ;
  assign n1700 = ~\a[1]  & \b[15]  ;
  assign n1701 = n1521 & n1700 ;
  assign n1702 = ~n1699 & ~n1701 ;
  assign n1703 = ~n1698 & n1702 ;
  assign n1704 = ~n1696 & n1703 ;
  assign n1705 = ~\a[2]  & ~n1704 ;
  assign n1706 = \a[2]  & n1703 ;
  assign n1707 = ~n1696 & n1706 ;
  assign n1708 = ~n1705 & ~n1707 ;
  assign n1709 = ~n1687 & ~n1708 ;
  assign n1710 = n1547 & n1709 ;
  assign n1711 = n1687 & ~n1708 ;
  assign n1712 = ~n1547 & n1711 ;
  assign n1713 = ~n1710 & ~n1712 ;
  assign n1714 = ~n1687 & n1708 ;
  assign n1715 = ~n1547 & n1714 ;
  assign n1716 = n1687 & n1708 ;
  assign n1717 = n1547 & n1716 ;
  assign n1718 = ~n1715 & ~n1717 ;
  assign n1719 = n1713 & n1718 ;
  assign n1720 = ~n1544 & n1719 ;
  assign n1721 = ~n1534 & ~n1719 ;
  assign n1722 = ~n1541 & n1721 ;
  assign n1723 = ~n1720 & ~n1722 ;
  assign n1724 = ~n1534 & n1713 ;
  assign n1725 = ~n1541 & n1724 ;
  assign n1726 = n1718 & ~n1725 ;
  assign n1727 = n1547 & n1687 ;
  assign n1728 = n1686 & ~n1727 ;
  assign n1729 = n1493 & ~n1675 ;
  assign n1730 = ~n1548 & n1729 ;
  assign n1731 = ~n1674 & ~n1730 ;
  assign n1732 = n252 & ~n1233 ;
  assign n1733 = ~n1231 & n1732 ;
  assign n1734 = \b[13]  & n303 ;
  assign n1735 = n300 & n1734 ;
  assign n1736 = \b[15]  & n250 ;
  assign n1737 = \a[3]  & \b[14]  ;
  assign n1738 = n241 & n1737 ;
  assign n1739 = ~\a[3]  & \b[14]  ;
  assign n1740 = n244 & n1739 ;
  assign n1741 = ~n1738 & ~n1740 ;
  assign n1742 = ~n1736 & n1741 ;
  assign n1743 = ~n1735 & n1742 ;
  assign n1744 = ~n1733 & n1743 ;
  assign n1745 = ~\a[5]  & ~n1744 ;
  assign n1746 = \a[5]  & n1743 ;
  assign n1747 = ~n1733 & n1746 ;
  assign n1748 = ~n1745 & ~n1747 ;
  assign n1749 = ~n1669 & ~n1671 ;
  assign n1750 = n430 & ~n912 ;
  assign n1751 = ~n910 & n1750 ;
  assign n1752 = \b[10]  & n486 ;
  assign n1753 = n483 & n1752 ;
  assign n1754 = \b[12]  & n428 ;
  assign n1755 = \a[5]  & \b[11]  ;
  assign n1756 = n484 & n1755 ;
  assign n1757 = ~\a[6]  & \b[11]  ;
  assign n1758 = n422 & n1757 ;
  assign n1759 = ~n1756 & ~n1758 ;
  assign n1760 = ~n1754 & n1759 ;
  assign n1761 = ~n1753 & n1760 ;
  assign n1762 = ~n1751 & n1761 ;
  assign n1763 = ~\a[8]  & ~n1762 ;
  assign n1764 = \a[8]  & n1761 ;
  assign n1765 = ~n1751 & n1764 ;
  assign n1766 = ~n1763 & ~n1765 ;
  assign n1767 = ~n589 & n646 ;
  assign n1768 = ~n587 & n1767 ;
  assign n1769 = \b[7]  & n796 ;
  assign n1770 = n793 & n1769 ;
  assign n1771 = \b[9]  & n644 ;
  assign n1772 = \a[9]  & \b[8]  ;
  assign n1773 = n635 & n1772 ;
  assign n1774 = ~\a[9]  & \b[8]  ;
  assign n1775 = n638 & n1774 ;
  assign n1776 = ~n1773 & ~n1775 ;
  assign n1777 = ~n1771 & n1776 ;
  assign n1778 = ~n1770 & n1777 ;
  assign n1779 = ~n1768 & n1778 ;
  assign n1780 = ~\a[11]  & ~n1779 ;
  assign n1781 = \a[11]  & n1778 ;
  assign n1782 = ~n1768 & n1781 ;
  assign n1783 = ~n1780 & ~n1782 ;
  assign n1784 = ~n1476 & ~n1660 ;
  assign n1785 = ~n1478 & n1784 ;
  assign n1786 = ~n1661 & ~n1785 ;
  assign n1787 = n177 & n1467 ;
  assign n1788 = \b[3]  & n1465 ;
  assign n1789 = \a[14]  & \b[2]  ;
  assign n1790 = n1650 & n1789 ;
  assign n1791 = ~\a[15]  & \b[2]  ;
  assign n1792 = n1459 & n1791 ;
  assign n1793 = ~n1790 & ~n1792 ;
  assign n1794 = ~n1788 & n1793 ;
  assign n1795 = ~n1787 & n1794 ;
  assign n1796 = \b[1]  & n1652 ;
  assign n1797 = n1649 & n1796 ;
  assign n1798 = ~\a[17]  & ~n1797 ;
  assign n1799 = n1795 & n1798 ;
  assign n1800 = n1795 & ~n1797 ;
  assign n1801 = \a[17]  & ~n1800 ;
  assign n1802 = ~n1799 & ~n1801 ;
  assign n1803 = \a[17]  & ~\a[18]  ;
  assign n1804 = ~\a[17]  & \a[18]  ;
  assign n1805 = ~n1803 & ~n1804 ;
  assign n1806 = \b[0]  & ~n1805 ;
  assign n1807 = n1639 & n1656 ;
  assign n1808 = n1806 & n1807 ;
  assign n1809 = ~n1806 & ~n1807 ;
  assign n1810 = ~n1808 & ~n1809 ;
  assign n1811 = n1802 & n1810 ;
  assign n1812 = ~n1802 & ~n1810 ;
  assign n1813 = ~n1811 & ~n1812 ;
  assign n1814 = ~n323 & ~n847 ;
  assign n1815 = ~n996 & n1814 ;
  assign n1816 = n320 & n1815 ;
  assign n1817 = n323 & ~n847 ;
  assign n1818 = ~n996 & n1817 ;
  assign n1819 = ~n320 & n1818 ;
  assign n1820 = ~n1816 & ~n1819 ;
  assign n1821 = \b[4]  & n1182 ;
  assign n1822 = n1179 & n1821 ;
  assign n1823 = \b[6]  & n997 ;
  assign n1824 = \a[11]  & \b[5]  ;
  assign n1825 = n1180 & n1824 ;
  assign n1826 = ~\a[12]  & \b[5]  ;
  assign n1827 = n991 & n1826 ;
  assign n1828 = ~n1825 & ~n1827 ;
  assign n1829 = ~n1823 & n1828 ;
  assign n1830 = ~n1822 & n1829 ;
  assign n1831 = n1820 & n1830 ;
  assign n1832 = ~\a[14]  & ~n1831 ;
  assign n1833 = \a[14]  & n1830 ;
  assign n1834 = n1820 & n1833 ;
  assign n1835 = ~n1832 & ~n1834 ;
  assign n1836 = n1813 & ~n1835 ;
  assign n1837 = ~n1813 & n1835 ;
  assign n1838 = ~n1836 & ~n1837 ;
  assign n1839 = n1786 & n1838 ;
  assign n1840 = ~n1786 & ~n1838 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1842 = ~n1783 & n1841 ;
  assign n1843 = n1783 & ~n1841 ;
  assign n1844 = ~n1842 & ~n1843 ;
  assign n1845 = n1766 & ~n1844 ;
  assign n1846 = n1749 & n1845 ;
  assign n1847 = n1766 & n1844 ;
  assign n1848 = ~n1749 & n1847 ;
  assign n1849 = ~n1846 & ~n1848 ;
  assign n1850 = ~n1766 & ~n1844 ;
  assign n1851 = ~n1749 & n1850 ;
  assign n1852 = ~n1766 & n1844 ;
  assign n1853 = n1749 & n1852 ;
  assign n1854 = ~n1851 & ~n1853 ;
  assign n1855 = n1849 & n1854 ;
  assign n1856 = ~n1748 & ~n1855 ;
  assign n1857 = n1731 & n1856 ;
  assign n1858 = ~n1748 & n1855 ;
  assign n1859 = ~n1731 & n1858 ;
  assign n1860 = ~n1857 & ~n1859 ;
  assign n1861 = n1748 & ~n1855 ;
  assign n1862 = ~n1731 & n1861 ;
  assign n1863 = n1748 & n1855 ;
  assign n1864 = n1731 & n1863 ;
  assign n1865 = ~n1862 & ~n1864 ;
  assign n1866 = n1860 & n1865 ;
  assign n1867 = ~n1728 & n1866 ;
  assign n1868 = n1686 & ~n1866 ;
  assign n1869 = ~n1727 & n1868 ;
  assign n1870 = ~n1511 & ~n1690 ;
  assign n1871 = ~n1515 & n1870 ;
  assign n1872 = ~n1689 & ~n1871 ;
  assign n1873 = ~\b[17]  & ~\b[18]  ;
  assign n1874 = \b[17]  & \b[18]  ;
  assign n1875 = ~n1873 & ~n1874 ;
  assign n1876 = ~n1872 & ~n1875 ;
  assign n1877 = ~n1689 & n1875 ;
  assign n1878 = ~n1871 & n1877 ;
  assign n1879 = n134 & ~n1878 ;
  assign n1880 = ~n1876 & n1879 ;
  assign n1881 = \a[0]  & \b[18]  ;
  assign n1882 = n133 & n1881 ;
  assign n1883 = \b[17]  & n141 ;
  assign n1884 = ~\a[1]  & \b[16]  ;
  assign n1885 = n1521 & n1884 ;
  assign n1886 = ~n1883 & ~n1885 ;
  assign n1887 = ~n1882 & n1886 ;
  assign n1888 = \a[2]  & n1887 ;
  assign n1889 = ~n1880 & n1888 ;
  assign n1890 = ~n1880 & n1887 ;
  assign n1891 = ~\a[2]  & ~n1890 ;
  assign n1892 = ~n1889 & ~n1891 ;
  assign n1893 = ~n1869 & ~n1892 ;
  assign n1894 = ~n1867 & n1893 ;
  assign n1895 = ~n1866 & n1892 ;
  assign n1896 = n1728 & n1895 ;
  assign n1897 = n1866 & n1892 ;
  assign n1898 = ~n1728 & n1897 ;
  assign n1899 = ~n1896 & ~n1898 ;
  assign n1900 = ~n1894 & n1899 ;
  assign n1901 = n1726 & n1900 ;
  assign n1902 = ~n1726 & ~n1900 ;
  assign n1903 = ~n1901 & ~n1902 ;
  assign n1904 = ~n1894 & ~n1901 ;
  assign n1905 = n1686 & n1860 ;
  assign n1906 = ~n1727 & n1905 ;
  assign n1907 = n1865 & ~n1906 ;
  assign n1908 = ~n1669 & ~n1842 ;
  assign n1909 = ~n1671 & n1908 ;
  assign n1910 = ~n1843 & ~n1909 ;
  assign n1911 = ~n1836 & ~n1839 ;
  assign n1912 = ~n380 & n999 ;
  assign n1913 = ~n322 & n999 ;
  assign n1914 = ~n326 & n1913 ;
  assign n1915 = ~n1912 & ~n1914 ;
  assign n1916 = ~n383 & ~n1915 ;
  assign n1917 = \b[5]  & n1182 ;
  assign n1918 = n1179 & n1917 ;
  assign n1919 = \b[7]  & n997 ;
  assign n1920 = \a[11]  & \b[6]  ;
  assign n1921 = n1180 & n1920 ;
  assign n1922 = ~\a[12]  & \b[6]  ;
  assign n1923 = n991 & n1922 ;
  assign n1924 = ~n1921 & ~n1923 ;
  assign n1925 = ~n1919 & n1924 ;
  assign n1926 = ~n1918 & n1925 ;
  assign n1927 = ~\a[14]  & n1926 ;
  assign n1928 = ~n1916 & n1927 ;
  assign n1929 = \a[14]  & ~n1926 ;
  assign n1930 = \a[14]  & ~n383 ;
  assign n1931 = ~n1915 & n1930 ;
  assign n1932 = ~n1929 & ~n1931 ;
  assign n1933 = ~n1928 & n1932 ;
  assign n1934 = ~n1808 & ~n1811 ;
  assign n1935 = n222 & n1467 ;
  assign n1936 = \b[4]  & n1465 ;
  assign n1937 = ~\a[15]  & \b[3]  ;
  assign n1938 = n1459 & n1937 ;
  assign n1939 = \a[15]  & \b[3]  ;
  assign n1940 = n1456 & n1939 ;
  assign n1941 = ~n1938 & ~n1940 ;
  assign n1942 = ~n1936 & n1941 ;
  assign n1943 = \b[2]  & n1652 ;
  assign n1944 = n1649 & n1943 ;
  assign n1945 = \a[17]  & ~n1944 ;
  assign n1946 = n1942 & n1945 ;
  assign n1947 = ~n1935 & n1946 ;
  assign n1948 = n1942 & ~n1944 ;
  assign n1949 = ~n1935 & n1948 ;
  assign n1950 = ~\a[17]  & ~n1949 ;
  assign n1951 = ~n1947 & ~n1950 ;
  assign n1952 = \a[20]  & \b[0]  ;
  assign n1953 = ~n1805 & n1952 ;
  assign n1954 = \a[18]  & ~\a[19]  ;
  assign n1955 = n1453 & n1954 ;
  assign n1956 = ~\a[18]  & \b[0]  ;
  assign n1957 = ~\a[17]  & \a[19]  ;
  assign n1958 = n1956 & n1957 ;
  assign n1959 = ~n1955 & ~n1958 ;
  assign n1960 = \a[19]  & ~\a[20]  ;
  assign n1961 = ~\a[19]  & \a[20]  ;
  assign n1962 = ~n1960 & ~n1961 ;
  assign n1963 = ~n1805 & n1962 ;
  assign n1964 = \b[1]  & n1963 ;
  assign n1965 = ~n1805 & ~n1962 ;
  assign n1966 = ~n137 & n1965 ;
  assign n1967 = ~n1964 & ~n1966 ;
  assign n1968 = n1959 & n1967 ;
  assign n1969 = n1953 & ~n1968 ;
  assign n1970 = ~n1953 & n1959 ;
  assign n1971 = n1967 & n1970 ;
  assign n1972 = ~n1969 & ~n1971 ;
  assign n1973 = ~n1951 & n1972 ;
  assign n1974 = n1951 & ~n1972 ;
  assign n1975 = ~n1973 & ~n1974 ;
  assign n1976 = ~n1934 & n1975 ;
  assign n1977 = n1934 & ~n1975 ;
  assign n1978 = ~n1976 & ~n1977 ;
  assign n1979 = n1933 & n1978 ;
  assign n1980 = ~n1933 & ~n1978 ;
  assign n1981 = ~n1979 & ~n1980 ;
  assign n1982 = n646 & ~n721 ;
  assign n1983 = ~n1033 & n1982 ;
  assign n1984 = \b[8]  & n796 ;
  assign n1985 = n793 & n1984 ;
  assign n1986 = \b[10]  & n644 ;
  assign n1987 = \a[9]  & \b[9]  ;
  assign n1988 = n635 & n1987 ;
  assign n1989 = ~\a[9]  & \b[9]  ;
  assign n1990 = n638 & n1989 ;
  assign n1991 = ~n1988 & ~n1990 ;
  assign n1992 = ~n1986 & n1991 ;
  assign n1993 = ~n1985 & n1992 ;
  assign n1994 = ~n1983 & n1993 ;
  assign n1995 = ~\a[11]  & ~n1994 ;
  assign n1996 = \a[11]  & n1993 ;
  assign n1997 = ~n1983 & n1996 ;
  assign n1998 = ~n1995 & ~n1997 ;
  assign n1999 = ~n1981 & ~n1998 ;
  assign n2000 = ~n1911 & n1999 ;
  assign n2001 = n1981 & ~n1998 ;
  assign n2002 = n1911 & n2001 ;
  assign n2003 = ~n2000 & ~n2002 ;
  assign n2004 = ~n1981 & n1998 ;
  assign n2005 = n1911 & n2004 ;
  assign n2006 = n1981 & n1998 ;
  assign n2007 = ~n1911 & n2006 ;
  assign n2008 = ~n2005 & ~n2007 ;
  assign n2009 = n2003 & n2008 ;
  assign n2010 = n430 & ~n951 ;
  assign n2011 = ~n949 & n2010 ;
  assign n2012 = \b[11]  & n486 ;
  assign n2013 = n483 & n2012 ;
  assign n2014 = \b[13]  & n428 ;
  assign n2015 = \a[5]  & \b[12]  ;
  assign n2016 = n484 & n2015 ;
  assign n2017 = ~\a[6]  & \b[12]  ;
  assign n2018 = n422 & n2017 ;
  assign n2019 = ~n2016 & ~n2018 ;
  assign n2020 = ~n2014 & n2019 ;
  assign n2021 = ~n2013 & n2020 ;
  assign n2022 = ~n2011 & n2021 ;
  assign n2023 = ~\a[8]  & ~n2022 ;
  assign n2024 = \a[8]  & n2021 ;
  assign n2025 = ~n2011 & n2024 ;
  assign n2026 = ~n2023 & ~n2025 ;
  assign n2027 = ~n2009 & n2026 ;
  assign n2028 = ~n1910 & n2027 ;
  assign n2029 = n2009 & n2026 ;
  assign n2030 = n1910 & n2029 ;
  assign n2031 = ~n2028 & ~n2030 ;
  assign n2032 = ~n2009 & ~n2026 ;
  assign n2033 = n1910 & n2032 ;
  assign n2034 = n2009 & ~n2026 ;
  assign n2035 = ~n1910 & n2034 ;
  assign n2036 = ~n2033 & ~n2035 ;
  assign n2037 = n2031 & n2036 ;
  assign n2038 = n1731 & n1855 ;
  assign n2039 = n1854 & ~n2038 ;
  assign n2040 = n2037 & ~n2039 ;
  assign n2041 = n1854 & ~n2037 ;
  assign n2042 = ~n2038 & n2041 ;
  assign n2043 = n252 & n1512 ;
  assign n2044 = ~n1509 & n2043 ;
  assign n2045 = n252 & ~n1512 ;
  assign n2046 = ~n1228 & n2045 ;
  assign n2047 = ~n1508 & n2046 ;
  assign n2048 = \b[14]  & n303 ;
  assign n2049 = n300 & n2048 ;
  assign n2050 = \b[16]  & n250 ;
  assign n2051 = \a[3]  & \b[15]  ;
  assign n2052 = n241 & n2051 ;
  assign n2053 = ~\a[3]  & \b[15]  ;
  assign n2054 = n244 & n2053 ;
  assign n2055 = ~n2052 & ~n2054 ;
  assign n2056 = ~n2050 & n2055 ;
  assign n2057 = ~n2049 & n2056 ;
  assign n2058 = ~n2047 & n2057 ;
  assign n2059 = ~n2044 & n2058 ;
  assign n2060 = ~\a[5]  & ~n2059 ;
  assign n2061 = \a[5]  & n2057 ;
  assign n2062 = ~n2047 & n2061 ;
  assign n2063 = ~n2044 & n2062 ;
  assign n2064 = ~n2060 & ~n2063 ;
  assign n2065 = ~n2042 & ~n2064 ;
  assign n2066 = ~n2040 & n2065 ;
  assign n2067 = n2037 & n2064 ;
  assign n2068 = ~n2039 & n2067 ;
  assign n2069 = ~n2037 & n2064 ;
  assign n2070 = n2039 & n2069 ;
  assign n2071 = ~n2068 & ~n2070 ;
  assign n2072 = ~n2066 & n2071 ;
  assign n2073 = ~n1874 & ~n1878 ;
  assign n2074 = ~\b[18]  & ~\b[19]  ;
  assign n2075 = \b[18]  & \b[19]  ;
  assign n2076 = ~n2074 & ~n2075 ;
  assign n2077 = ~n2073 & n2076 ;
  assign n2078 = ~n1874 & ~n2076 ;
  assign n2079 = ~n1878 & n2078 ;
  assign n2080 = n134 & ~n2079 ;
  assign n2081 = ~n2077 & n2080 ;
  assign n2082 = \a[0]  & \b[19]  ;
  assign n2083 = n133 & n2082 ;
  assign n2084 = \b[18]  & n141 ;
  assign n2085 = ~\a[1]  & \b[17]  ;
  assign n2086 = n1521 & n2085 ;
  assign n2087 = ~n2084 & ~n2086 ;
  assign n2088 = ~n2083 & n2087 ;
  assign n2089 = ~n2081 & n2088 ;
  assign n2090 = ~\a[2]  & ~n2089 ;
  assign n2091 = \a[2]  & n2088 ;
  assign n2092 = ~n2081 & n2091 ;
  assign n2093 = ~n2090 & ~n2092 ;
  assign n2094 = ~n2072 & ~n2093 ;
  assign n2095 = n1907 & n2094 ;
  assign n2096 = n2072 & ~n2093 ;
  assign n2097 = ~n1907 & n2096 ;
  assign n2098 = ~n2095 & ~n2097 ;
  assign n2099 = ~n2072 & n2093 ;
  assign n2100 = ~n1907 & n2099 ;
  assign n2101 = n2072 & n2093 ;
  assign n2102 = n1907 & n2101 ;
  assign n2103 = ~n2100 & ~n2102 ;
  assign n2104 = n2098 & n2103 ;
  assign n2105 = ~n1904 & n2104 ;
  assign n2106 = ~n1894 & ~n2104 ;
  assign n2107 = ~n1901 & n2106 ;
  assign n2108 = ~n2105 & ~n2107 ;
  assign n2109 = ~n1894 & n2098 ;
  assign n2110 = ~n1901 & n2109 ;
  assign n2111 = n2103 & ~n2110 ;
  assign n2112 = n1907 & n2072 ;
  assign n2113 = ~n2066 & ~n2112 ;
  assign n2114 = n1854 & n2036 ;
  assign n2115 = ~n2038 & n2114 ;
  assign n2116 = n2031 & ~n2115 ;
  assign n2117 = n252 & ~n1694 ;
  assign n2118 = ~n1692 & n2117 ;
  assign n2119 = \b[15]  & n303 ;
  assign n2120 = n300 & n2119 ;
  assign n2121 = \b[17]  & n250 ;
  assign n2122 = \a[3]  & \b[16]  ;
  assign n2123 = n241 & n2122 ;
  assign n2124 = ~\a[3]  & \b[16]  ;
  assign n2125 = n244 & n2124 ;
  assign n2126 = ~n2123 & ~n2125 ;
  assign n2127 = ~n2121 & n2126 ;
  assign n2128 = ~n2120 & n2127 ;
  assign n2129 = ~n2118 & n2128 ;
  assign n2130 = ~\a[5]  & ~n2129 ;
  assign n2131 = \a[5]  & n2128 ;
  assign n2132 = ~n2118 & n2131 ;
  assign n2133 = ~n2130 & ~n2132 ;
  assign n2134 = n1910 & n2009 ;
  assign n2135 = n2003 & ~n2134 ;
  assign n2136 = n646 & ~n728 ;
  assign n2137 = ~n726 & n2136 ;
  assign n2138 = \b[9]  & n796 ;
  assign n2139 = n793 & n2138 ;
  assign n2140 = \b[11]  & n644 ;
  assign n2141 = \a[9]  & \b[10]  ;
  assign n2142 = n635 & n2141 ;
  assign n2143 = ~\a[9]  & \b[10]  ;
  assign n2144 = n638 & n2143 ;
  assign n2145 = ~n2142 & ~n2144 ;
  assign n2146 = ~n2140 & n2145 ;
  assign n2147 = ~n2139 & n2146 ;
  assign n2148 = ~\a[11]  & n2147 ;
  assign n2149 = ~n2137 & n2148 ;
  assign n2150 = ~n2137 & n2147 ;
  assign n2151 = \a[11]  & ~n2150 ;
  assign n2152 = ~n2149 & ~n2151 ;
  assign n2153 = ~n1836 & ~n1979 ;
  assign n2154 = ~n1839 & n2153 ;
  assign n2155 = ~n1980 & ~n2154 ;
  assign n2156 = ~n505 & ~n847 ;
  assign n2157 = ~n996 & n2156 ;
  assign n2158 = n502 & n2157 ;
  assign n2159 = n505 & ~n847 ;
  assign n2160 = ~n996 & n2159 ;
  assign n2161 = ~n502 & n2160 ;
  assign n2162 = ~n2158 & ~n2161 ;
  assign n2163 = \b[6]  & n1182 ;
  assign n2164 = n1179 & n2163 ;
  assign n2165 = \b[8]  & n997 ;
  assign n2166 = \a[11]  & \b[7]  ;
  assign n2167 = n1180 & n2166 ;
  assign n2168 = ~\a[12]  & \b[7]  ;
  assign n2169 = n991 & n2168 ;
  assign n2170 = ~n2167 & ~n2169 ;
  assign n2171 = ~n2165 & n2170 ;
  assign n2172 = ~n2164 & n2171 ;
  assign n2173 = n2162 & n2172 ;
  assign n2174 = ~\a[14]  & ~n2173 ;
  assign n2175 = \a[14]  & n2172 ;
  assign n2176 = n2162 & n2175 ;
  assign n2177 = ~n2174 & ~n2176 ;
  assign n2178 = ~n1973 & ~n1976 ;
  assign n2179 = ~n270 & n1467 ;
  assign n2180 = ~n218 & n1467 ;
  assign n2181 = ~n220 & n2180 ;
  assign n2182 = ~n2179 & ~n2181 ;
  assign n2183 = ~n273 & ~n2182 ;
  assign n2184 = \b[3]  & n1652 ;
  assign n2185 = n1649 & n2184 ;
  assign n2186 = ~\a[15]  & \b[4]  ;
  assign n2187 = n1459 & n2186 ;
  assign n2188 = ~n2185 & ~n2187 ;
  assign n2189 = \b[5]  & n1465 ;
  assign n2190 = \a[15]  & \b[4]  ;
  assign n2191 = n1456 & n2190 ;
  assign n2192 = \a[17]  & ~n2191 ;
  assign n2193 = ~n2189 & n2192 ;
  assign n2194 = n2188 & n2193 ;
  assign n2195 = ~n2183 & n2194 ;
  assign n2196 = ~n2189 & ~n2191 ;
  assign n2197 = n2188 & n2196 ;
  assign n2198 = ~\a[17]  & ~n2197 ;
  assign n2199 = ~\a[17]  & ~n273 ;
  assign n2200 = ~n2182 & n2199 ;
  assign n2201 = ~n2198 & ~n2200 ;
  assign n2202 = ~n2195 & n2201 ;
  assign n2203 = \a[20]  & ~n1806 ;
  assign n2204 = n1959 & n2203 ;
  assign n2205 = n1967 & n2204 ;
  assign n2206 = \a[20]  & ~n2205 ;
  assign n2207 = \b[2]  & n1963 ;
  assign n2208 = ~\a[18]  & \b[1]  ;
  assign n2209 = n1957 & n2208 ;
  assign n2210 = \a[17]  & ~\a[19]  ;
  assign n2211 = \a[18]  & \b[1]  ;
  assign n2212 = n2210 & n2211 ;
  assign n2213 = ~n2209 & ~n2212 ;
  assign n2214 = ~n2207 & n2213 ;
  assign n2215 = n157 & n1965 ;
  assign n2216 = n1805 & ~n1962 ;
  assign n2217 = ~\a[18]  & \a[19]  ;
  assign n2218 = ~n1954 & ~n2217 ;
  assign n2219 = \b[0]  & n2218 ;
  assign n2220 = n2216 & n2219 ;
  assign n2221 = ~n2215 & ~n2220 ;
  assign n2222 = n2214 & n2221 ;
  assign n2223 = ~n2206 & ~n2222 ;
  assign n2224 = n2206 & n2222 ;
  assign n2225 = ~n2223 & ~n2224 ;
  assign n2226 = ~n2202 & ~n2225 ;
  assign n2227 = n2202 & n2225 ;
  assign n2228 = ~n2226 & ~n2227 ;
  assign n2229 = ~n2178 & n2228 ;
  assign n2230 = ~n1973 & ~n2228 ;
  assign n2231 = ~n1976 & n2230 ;
  assign n2232 = ~n2229 & ~n2231 ;
  assign n2233 = n2177 & ~n2232 ;
  assign n2234 = ~n2177 & ~n2231 ;
  assign n2235 = ~n2229 & n2234 ;
  assign n2236 = ~n2233 & ~n2235 ;
  assign n2237 = n2155 & n2236 ;
  assign n2238 = ~n2155 & ~n2236 ;
  assign n2239 = ~n2237 & ~n2238 ;
  assign n2240 = ~n2152 & ~n2239 ;
  assign n2241 = n2152 & n2239 ;
  assign n2242 = ~n2240 & ~n2241 ;
  assign n2243 = ~n359 & ~n946 ;
  assign n2244 = ~n1087 & n2243 ;
  assign n2245 = ~n1083 & n2244 ;
  assign n2246 = ~n427 & n2245 ;
  assign n2247 = n430 & n1087 ;
  assign n2248 = ~n1084 & n2247 ;
  assign n2249 = ~n2246 & ~n2248 ;
  assign n2250 = \b[12]  & n486 ;
  assign n2251 = n483 & n2250 ;
  assign n2252 = \b[14]  & n428 ;
  assign n2253 = \a[5]  & \b[13]  ;
  assign n2254 = n484 & n2253 ;
  assign n2255 = ~\a[6]  & \b[13]  ;
  assign n2256 = n422 & n2255 ;
  assign n2257 = ~n2254 & ~n2256 ;
  assign n2258 = ~n2252 & n2257 ;
  assign n2259 = ~n2251 & n2258 ;
  assign n2260 = n2249 & n2259 ;
  assign n2261 = ~\a[8]  & ~n2260 ;
  assign n2262 = \a[8]  & n2259 ;
  assign n2263 = n2249 & n2262 ;
  assign n2264 = ~n2261 & ~n2263 ;
  assign n2265 = ~n2242 & ~n2264 ;
  assign n2266 = ~n2135 & n2265 ;
  assign n2267 = n2242 & ~n2264 ;
  assign n2268 = n2135 & n2267 ;
  assign n2269 = ~n2266 & ~n2268 ;
  assign n2270 = ~n2242 & n2264 ;
  assign n2271 = n2135 & n2270 ;
  assign n2272 = n2242 & n2264 ;
  assign n2273 = ~n2135 & n2272 ;
  assign n2274 = ~n2271 & ~n2273 ;
  assign n2275 = n2269 & n2274 ;
  assign n2276 = ~n2133 & ~n2275 ;
  assign n2277 = n2116 & n2276 ;
  assign n2278 = ~n2133 & n2275 ;
  assign n2279 = ~n2116 & n2278 ;
  assign n2280 = ~n2277 & ~n2279 ;
  assign n2281 = n2133 & ~n2275 ;
  assign n2282 = ~n2116 & n2281 ;
  assign n2283 = n2133 & n2275 ;
  assign n2284 = n2116 & n2283 ;
  assign n2285 = ~n2282 & ~n2284 ;
  assign n2286 = n2280 & n2285 ;
  assign n2287 = ~n2113 & n2286 ;
  assign n2288 = ~n1874 & ~n2075 ;
  assign n2289 = ~n1878 & n2288 ;
  assign n2290 = ~n2074 & ~n2289 ;
  assign n2291 = ~\b[19]  & ~\b[20]  ;
  assign n2292 = \b[19]  & \b[20]  ;
  assign n2293 = ~n2291 & ~n2292 ;
  assign n2294 = n134 & n2293 ;
  assign n2295 = ~n2290 & n2294 ;
  assign n2296 = n134 & ~n2293 ;
  assign n2297 = ~n2074 & n2296 ;
  assign n2298 = ~n2289 & n2297 ;
  assign n2299 = \a[0]  & \b[20]  ;
  assign n2300 = n133 & n2299 ;
  assign n2301 = \b[19]  & n141 ;
  assign n2302 = ~\a[1]  & \b[18]  ;
  assign n2303 = n1521 & n2302 ;
  assign n2304 = ~n2301 & ~n2303 ;
  assign n2305 = ~n2300 & n2304 ;
  assign n2306 = \a[2]  & n2305 ;
  assign n2307 = ~n2298 & n2306 ;
  assign n2308 = ~n2295 & n2307 ;
  assign n2309 = ~n2298 & n2305 ;
  assign n2310 = ~n2295 & n2309 ;
  assign n2311 = ~\a[2]  & ~n2310 ;
  assign n2312 = ~n2308 & ~n2311 ;
  assign n2313 = ~n2066 & ~n2286 ;
  assign n2314 = ~n2112 & n2313 ;
  assign n2315 = ~n2312 & ~n2314 ;
  assign n2316 = ~n2287 & n2315 ;
  assign n2317 = ~n2286 & n2312 ;
  assign n2318 = n2113 & n2317 ;
  assign n2319 = n2286 & n2312 ;
  assign n2320 = ~n2113 & n2319 ;
  assign n2321 = ~n2318 & ~n2320 ;
  assign n2322 = ~n2316 & n2321 ;
  assign n2323 = n2111 & n2322 ;
  assign n2324 = ~n2111 & ~n2322 ;
  assign n2325 = ~n2323 & ~n2324 ;
  assign n2326 = ~n2316 & ~n2323 ;
  assign n2327 = ~n2066 & n2280 ;
  assign n2328 = ~n2112 & n2327 ;
  assign n2329 = n2285 & ~n2328 ;
  assign n2330 = n2116 & n2275 ;
  assign n2331 = n2269 & ~n2330 ;
  assign n2332 = n2003 & ~n2241 ;
  assign n2333 = ~n2134 & n2332 ;
  assign n2334 = ~n2240 & ~n2333 ;
  assign n2335 = n430 & ~n1233 ;
  assign n2336 = ~n1231 & n2335 ;
  assign n2337 = \b[13]  & n486 ;
  assign n2338 = n483 & n2337 ;
  assign n2339 = \b[15]  & n428 ;
  assign n2340 = \a[5]  & \b[14]  ;
  assign n2341 = n484 & n2340 ;
  assign n2342 = ~\a[6]  & \b[14]  ;
  assign n2343 = n422 & n2342 ;
  assign n2344 = ~n2341 & ~n2343 ;
  assign n2345 = ~n2339 & n2344 ;
  assign n2346 = ~n2338 & n2345 ;
  assign n2347 = ~n2336 & n2346 ;
  assign n2348 = ~\a[8]  & ~n2347 ;
  assign n2349 = \a[8]  & n2346 ;
  assign n2350 = ~n2336 & n2349 ;
  assign n2351 = ~n2348 & ~n2350 ;
  assign n2352 = ~n2235 & ~n2237 ;
  assign n2353 = n646 & ~n912 ;
  assign n2354 = ~n910 & n2353 ;
  assign n2355 = \b[10]  & n796 ;
  assign n2356 = n793 & n2355 ;
  assign n2357 = \b[12]  & n644 ;
  assign n2358 = \a[9]  & \b[11]  ;
  assign n2359 = n635 & n2358 ;
  assign n2360 = ~\a[9]  & \b[11]  ;
  assign n2361 = n638 & n2360 ;
  assign n2362 = ~n2359 & ~n2361 ;
  assign n2363 = ~n2357 & n2362 ;
  assign n2364 = ~n2356 & n2363 ;
  assign n2365 = ~n2354 & n2364 ;
  assign n2366 = ~\a[11]  & ~n2365 ;
  assign n2367 = \a[11]  & n2364 ;
  assign n2368 = ~n2354 & n2367 ;
  assign n2369 = ~n2366 & ~n2368 ;
  assign n2370 = ~n1973 & ~n2226 ;
  assign n2371 = ~n1976 & n2370 ;
  assign n2372 = ~n2227 & ~n2371 ;
  assign n2373 = ~n586 & n999 ;
  assign n2374 = ~n504 & n999 ;
  assign n2375 = ~n508 & n2374 ;
  assign n2376 = ~n2373 & ~n2375 ;
  assign n2377 = ~n589 & ~n2376 ;
  assign n2378 = \b[7]  & n1182 ;
  assign n2379 = n1179 & n2378 ;
  assign n2380 = \b[9]  & n997 ;
  assign n2381 = \a[12]  & \b[8]  ;
  assign n2382 = n988 & n2381 ;
  assign n2383 = ~\a[12]  & \b[8]  ;
  assign n2384 = n991 & n2383 ;
  assign n2385 = ~n2382 & ~n2384 ;
  assign n2386 = ~n2380 & n2385 ;
  assign n2387 = ~n2379 & n2386 ;
  assign n2388 = ~\a[14]  & n2387 ;
  assign n2389 = ~n2377 & n2388 ;
  assign n2390 = \a[14]  & ~n2387 ;
  assign n2391 = \a[14]  & ~n589 ;
  assign n2392 = ~n2376 & n2391 ;
  assign n2393 = ~n2390 & ~n2392 ;
  assign n2394 = ~n2389 & n2393 ;
  assign n2395 = n177 & n1965 ;
  assign n2396 = \b[3]  & n1963 ;
  assign n2397 = \a[17]  & \b[2]  ;
  assign n2398 = n1954 & n2397 ;
  assign n2399 = ~\a[18]  & \b[2]  ;
  assign n2400 = n1957 & n2399 ;
  assign n2401 = ~n2398 & ~n2400 ;
  assign n2402 = ~n2396 & n2401 ;
  assign n2403 = ~n2395 & n2402 ;
  assign n2404 = \b[1]  & n2218 ;
  assign n2405 = n2216 & n2404 ;
  assign n2406 = ~\a[20]  & ~n2405 ;
  assign n2407 = n2403 & n2406 ;
  assign n2408 = n2403 & ~n2405 ;
  assign n2409 = \a[20]  & ~n2408 ;
  assign n2410 = ~n2407 & ~n2409 ;
  assign n2411 = \a[20]  & ~\a[21]  ;
  assign n2412 = ~\a[20]  & \a[21]  ;
  assign n2413 = ~n2411 & ~n2412 ;
  assign n2414 = \b[0]  & ~n2413 ;
  assign n2415 = n2205 & n2222 ;
  assign n2416 = n2414 & n2415 ;
  assign n2417 = ~n2414 & ~n2415 ;
  assign n2418 = ~n2416 & ~n2417 ;
  assign n2419 = n2410 & n2418 ;
  assign n2420 = ~n2410 & ~n2418 ;
  assign n2421 = ~n2419 & ~n2420 ;
  assign n2422 = ~n323 & ~n1304 ;
  assign n2423 = ~n1464 & n2422 ;
  assign n2424 = n320 & n2423 ;
  assign n2425 = n323 & ~n1304 ;
  assign n2426 = ~n1464 & n2425 ;
  assign n2427 = ~n320 & n2426 ;
  assign n2428 = ~n2424 & ~n2427 ;
  assign n2429 = \b[4]  & n1652 ;
  assign n2430 = n1649 & n2429 ;
  assign n2431 = ~\a[15]  & \b[5]  ;
  assign n2432 = n1459 & n2431 ;
  assign n2433 = ~n2430 & ~n2432 ;
  assign n2434 = \b[6]  & n1465 ;
  assign n2435 = \a[15]  & \b[5]  ;
  assign n2436 = n1456 & n2435 ;
  assign n2437 = \a[17]  & ~n2436 ;
  assign n2438 = ~n2434 & n2437 ;
  assign n2439 = n2433 & n2438 ;
  assign n2440 = n2428 & n2439 ;
  assign n2441 = ~n2434 & ~n2436 ;
  assign n2442 = n2433 & n2441 ;
  assign n2443 = n2428 & n2442 ;
  assign n2444 = ~\a[17]  & ~n2443 ;
  assign n2445 = ~n2440 & ~n2444 ;
  assign n2446 = n2421 & ~n2445 ;
  assign n2447 = ~n2421 & n2445 ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2449 = n2394 & ~n2448 ;
  assign n2450 = n2372 & n2449 ;
  assign n2451 = n2394 & n2448 ;
  assign n2452 = ~n2372 & n2451 ;
  assign n2453 = ~n2450 & ~n2452 ;
  assign n2454 = ~n2394 & ~n2448 ;
  assign n2455 = ~n2372 & n2454 ;
  assign n2456 = ~n2394 & n2448 ;
  assign n2457 = n2372 & n2456 ;
  assign n2458 = ~n2455 & ~n2457 ;
  assign n2459 = n2453 & n2458 ;
  assign n2460 = n2369 & ~n2459 ;
  assign n2461 = n2352 & n2460 ;
  assign n2462 = n2369 & n2459 ;
  assign n2463 = ~n2352 & n2462 ;
  assign n2464 = ~n2461 & ~n2463 ;
  assign n2465 = ~n2352 & n2459 ;
  assign n2466 = ~n2235 & ~n2459 ;
  assign n2467 = ~n2237 & n2466 ;
  assign n2468 = ~n2369 & ~n2467 ;
  assign n2469 = ~n2465 & n2468 ;
  assign n2470 = n2464 & ~n2469 ;
  assign n2471 = ~n2351 & ~n2470 ;
  assign n2472 = n2334 & n2471 ;
  assign n2473 = ~n2351 & n2470 ;
  assign n2474 = ~n2334 & n2473 ;
  assign n2475 = ~n2472 & ~n2474 ;
  assign n2476 = n2351 & ~n2470 ;
  assign n2477 = ~n2334 & n2476 ;
  assign n2478 = n2351 & n2470 ;
  assign n2479 = n2334 & n2478 ;
  assign n2480 = ~n2477 & ~n2479 ;
  assign n2481 = n2475 & n2480 ;
  assign n2482 = ~n2331 & n2481 ;
  assign n2483 = n2269 & ~n2481 ;
  assign n2484 = ~n2330 & n2483 ;
  assign n2485 = n252 & n1875 ;
  assign n2486 = ~n1872 & n2485 ;
  assign n2487 = n252 & ~n1875 ;
  assign n2488 = ~n1689 & n2487 ;
  assign n2489 = ~n1871 & n2488 ;
  assign n2490 = \b[16]  & n303 ;
  assign n2491 = n300 & n2490 ;
  assign n2492 = \b[18]  & n250 ;
  assign n2493 = \a[3]  & \b[17]  ;
  assign n2494 = n241 & n2493 ;
  assign n2495 = ~\a[3]  & \b[17]  ;
  assign n2496 = n244 & n2495 ;
  assign n2497 = ~n2494 & ~n2496 ;
  assign n2498 = ~n2492 & n2497 ;
  assign n2499 = ~n2491 & n2498 ;
  assign n2500 = ~n2489 & n2499 ;
  assign n2501 = ~n2486 & n2500 ;
  assign n2502 = ~\a[5]  & ~n2501 ;
  assign n2503 = \a[5]  & n2499 ;
  assign n2504 = ~n2489 & n2503 ;
  assign n2505 = ~n2486 & n2504 ;
  assign n2506 = ~n2502 & ~n2505 ;
  assign n2507 = ~n2484 & ~n2506 ;
  assign n2508 = ~n2482 & n2507 ;
  assign n2509 = ~n2481 & n2506 ;
  assign n2510 = n2331 & n2509 ;
  assign n2511 = n2481 & n2506 ;
  assign n2512 = ~n2331 & n2511 ;
  assign n2513 = ~n2510 & ~n2512 ;
  assign n2514 = ~n2508 & n2513 ;
  assign n2515 = ~n2074 & n2293 ;
  assign n2516 = ~n2289 & n2515 ;
  assign n2517 = ~n2292 & ~n2516 ;
  assign n2518 = ~\b[20]  & ~\b[21]  ;
  assign n2519 = \b[20]  & \b[21]  ;
  assign n2520 = ~n2518 & ~n2519 ;
  assign n2521 = ~n2517 & n2520 ;
  assign n2522 = ~n2292 & ~n2520 ;
  assign n2523 = ~n2516 & n2522 ;
  assign n2524 = n134 & ~n2523 ;
  assign n2525 = ~n2521 & n2524 ;
  assign n2526 = \a[0]  & \b[21]  ;
  assign n2527 = n133 & n2526 ;
  assign n2528 = \b[20]  & n141 ;
  assign n2529 = ~\a[1]  & \b[19]  ;
  assign n2530 = n1521 & n2529 ;
  assign n2531 = ~n2528 & ~n2530 ;
  assign n2532 = ~n2527 & n2531 ;
  assign n2533 = ~n2525 & n2532 ;
  assign n2534 = ~\a[2]  & ~n2533 ;
  assign n2535 = \a[2]  & n2532 ;
  assign n2536 = ~n2525 & n2535 ;
  assign n2537 = ~n2534 & ~n2536 ;
  assign n2538 = ~n2514 & ~n2537 ;
  assign n2539 = n2329 & n2538 ;
  assign n2540 = n2514 & ~n2537 ;
  assign n2541 = ~n2329 & n2540 ;
  assign n2542 = ~n2539 & ~n2541 ;
  assign n2543 = ~n2514 & n2537 ;
  assign n2544 = ~n2329 & n2543 ;
  assign n2545 = n2514 & n2537 ;
  assign n2546 = n2329 & n2545 ;
  assign n2547 = ~n2544 & ~n2546 ;
  assign n2548 = n2542 & n2547 ;
  assign n2549 = ~n2326 & n2548 ;
  assign n2550 = ~n2316 & ~n2548 ;
  assign n2551 = ~n2323 & n2550 ;
  assign n2552 = ~n2549 & ~n2551 ;
  assign n2553 = ~n2316 & n2542 ;
  assign n2554 = ~n2323 & n2553 ;
  assign n2555 = n2547 & ~n2554 ;
  assign n2556 = n2329 & n2514 ;
  assign n2557 = ~n2508 & ~n2556 ;
  assign n2558 = n2269 & n2475 ;
  assign n2559 = ~n2330 & n2558 ;
  assign n2560 = n2480 & ~n2559 ;
  assign n2561 = n2334 & n2470 ;
  assign n2562 = ~n2469 & ~n2561 ;
  assign n2563 = ~n2235 & n2453 ;
  assign n2564 = ~n2237 & n2563 ;
  assign n2565 = n2458 & ~n2564 ;
  assign n2566 = n2372 & n2448 ;
  assign n2567 = ~n2446 & ~n2566 ;
  assign n2568 = ~n380 & n1467 ;
  assign n2569 = ~n322 & n1467 ;
  assign n2570 = ~n326 & n2569 ;
  assign n2571 = ~n2568 & ~n2570 ;
  assign n2572 = ~n383 & ~n2571 ;
  assign n2573 = \b[5]  & n1652 ;
  assign n2574 = n1649 & n2573 ;
  assign n2575 = \b[7]  & n1465 ;
  assign n2576 = \a[15]  & \b[6]  ;
  assign n2577 = n1456 & n2576 ;
  assign n2578 = ~\a[15]  & \b[6]  ;
  assign n2579 = n1459 & n2578 ;
  assign n2580 = ~n2577 & ~n2579 ;
  assign n2581 = ~n2575 & n2580 ;
  assign n2582 = ~n2574 & n2581 ;
  assign n2583 = ~\a[17]  & n2582 ;
  assign n2584 = ~n2572 & n2583 ;
  assign n2585 = \a[17]  & ~n2582 ;
  assign n2586 = \a[17]  & ~n383 ;
  assign n2587 = ~n2571 & n2586 ;
  assign n2588 = ~n2585 & ~n2587 ;
  assign n2589 = ~n2584 & n2588 ;
  assign n2590 = ~n2416 & ~n2419 ;
  assign n2591 = n222 & n1965 ;
  assign n2592 = \b[4]  & n1963 ;
  assign n2593 = \a[17]  & \b[3]  ;
  assign n2594 = n1954 & n2593 ;
  assign n2595 = ~\a[18]  & \b[3]  ;
  assign n2596 = n1957 & n2595 ;
  assign n2597 = ~n2594 & ~n2596 ;
  assign n2598 = ~n2592 & n2597 ;
  assign n2599 = \b[2]  & n2218 ;
  assign n2600 = n2216 & n2599 ;
  assign n2601 = \a[20]  & ~n2600 ;
  assign n2602 = n2598 & n2601 ;
  assign n2603 = ~n2591 & n2602 ;
  assign n2604 = n2598 & ~n2600 ;
  assign n2605 = ~n2591 & n2604 ;
  assign n2606 = ~\a[20]  & ~n2605 ;
  assign n2607 = ~n2603 & ~n2606 ;
  assign n2608 = \a[23]  & \b[0]  ;
  assign n2609 = ~n2413 & n2608 ;
  assign n2610 = \a[21]  & \b[0]  ;
  assign n2611 = \a[20]  & ~\a[22]  ;
  assign n2612 = n2610 & n2611 ;
  assign n2613 = ~\a[21]  & \b[0]  ;
  assign n2614 = ~\a[20]  & \a[22]  ;
  assign n2615 = n2613 & n2614 ;
  assign n2616 = ~n2612 & ~n2615 ;
  assign n2617 = \a[22]  & ~\a[23]  ;
  assign n2618 = ~\a[22]  & \a[23]  ;
  assign n2619 = ~n2617 & ~n2618 ;
  assign n2620 = ~n2413 & n2619 ;
  assign n2621 = \b[1]  & n2620 ;
  assign n2622 = ~n2413 & ~n2619 ;
  assign n2623 = ~n137 & n2622 ;
  assign n2624 = ~n2621 & ~n2623 ;
  assign n2625 = n2616 & n2624 ;
  assign n2626 = n2609 & ~n2625 ;
  assign n2627 = ~n2609 & n2616 ;
  assign n2628 = n2624 & n2627 ;
  assign n2629 = ~n2626 & ~n2628 ;
  assign n2630 = ~n2607 & n2629 ;
  assign n2631 = n2607 & ~n2629 ;
  assign n2632 = ~n2630 & ~n2631 ;
  assign n2633 = ~n2590 & n2632 ;
  assign n2634 = n2590 & ~n2632 ;
  assign n2635 = ~n2633 & ~n2634 ;
  assign n2636 = n2589 & n2635 ;
  assign n2637 = ~n2589 & ~n2635 ;
  assign n2638 = ~n2636 & ~n2637 ;
  assign n2639 = ~n685 & ~n847 ;
  assign n2640 = ~n996 & n2639 ;
  assign n2641 = n682 & n2640 ;
  assign n2642 = n685 & ~n847 ;
  assign n2643 = ~n996 & n2642 ;
  assign n2644 = ~n682 & n2643 ;
  assign n2645 = ~n2641 & ~n2644 ;
  assign n2646 = \b[8]  & n1182 ;
  assign n2647 = n1179 & n2646 ;
  assign n2648 = ~\a[11]  & \b[9]  ;
  assign n2649 = n1181 & n2648 ;
  assign n2650 = ~n2647 & ~n2649 ;
  assign n2651 = \b[10]  & n997 ;
  assign n2652 = \a[12]  & \b[9]  ;
  assign n2653 = n988 & n2652 ;
  assign n2654 = \a[14]  & ~n2653 ;
  assign n2655 = ~n2651 & n2654 ;
  assign n2656 = n2650 & n2655 ;
  assign n2657 = n2645 & n2656 ;
  assign n2658 = ~n2651 & ~n2653 ;
  assign n2659 = n2650 & n2658 ;
  assign n2660 = n2645 & n2659 ;
  assign n2661 = ~\a[14]  & ~n2660 ;
  assign n2662 = ~n2657 & ~n2661 ;
  assign n2663 = ~n2638 & ~n2662 ;
  assign n2664 = ~n2567 & n2663 ;
  assign n2665 = n2638 & ~n2662 ;
  assign n2666 = n2567 & n2665 ;
  assign n2667 = ~n2664 & ~n2666 ;
  assign n2668 = ~n2638 & n2662 ;
  assign n2669 = n2567 & n2668 ;
  assign n2670 = n2638 & n2662 ;
  assign n2671 = ~n2567 & n2670 ;
  assign n2672 = ~n2669 & ~n2671 ;
  assign n2673 = n2667 & n2672 ;
  assign n2674 = n646 & ~n951 ;
  assign n2675 = ~n949 & n2674 ;
  assign n2676 = \b[11]  & n796 ;
  assign n2677 = n793 & n2676 ;
  assign n2678 = \b[13]  & n644 ;
  assign n2679 = \a[9]  & \b[12]  ;
  assign n2680 = n635 & n2679 ;
  assign n2681 = ~\a[9]  & \b[12]  ;
  assign n2682 = n638 & n2681 ;
  assign n2683 = ~n2680 & ~n2682 ;
  assign n2684 = ~n2678 & n2683 ;
  assign n2685 = ~n2677 & n2684 ;
  assign n2686 = ~\a[11]  & n2685 ;
  assign n2687 = ~n2675 & n2686 ;
  assign n2688 = ~n2675 & n2685 ;
  assign n2689 = \a[11]  & ~n2688 ;
  assign n2690 = ~n2687 & ~n2689 ;
  assign n2691 = ~n2673 & ~n2690 ;
  assign n2692 = ~n2565 & n2691 ;
  assign n2693 = n2673 & ~n2690 ;
  assign n2694 = n2565 & n2693 ;
  assign n2695 = ~n2692 & ~n2694 ;
  assign n2696 = ~n2673 & n2690 ;
  assign n2697 = n2565 & n2696 ;
  assign n2698 = n2673 & n2690 ;
  assign n2699 = ~n2565 & n2698 ;
  assign n2700 = ~n2697 & ~n2699 ;
  assign n2701 = n2695 & n2700 ;
  assign n2702 = ~n2562 & n2701 ;
  assign n2703 = n430 & n1512 ;
  assign n2704 = ~n1509 & n2703 ;
  assign n2705 = n430 & ~n1512 ;
  assign n2706 = ~n1228 & n2705 ;
  assign n2707 = ~n1508 & n2706 ;
  assign n2708 = \b[14]  & n486 ;
  assign n2709 = n483 & n2708 ;
  assign n2710 = \b[16]  & n428 ;
  assign n2711 = \a[5]  & \b[15]  ;
  assign n2712 = n484 & n2711 ;
  assign n2713 = ~\a[6]  & \b[15]  ;
  assign n2714 = n422 & n2713 ;
  assign n2715 = ~n2712 & ~n2714 ;
  assign n2716 = ~n2710 & n2715 ;
  assign n2717 = ~n2709 & n2716 ;
  assign n2718 = ~n2707 & n2717 ;
  assign n2719 = ~n2704 & n2718 ;
  assign n2720 = ~\a[8]  & ~n2719 ;
  assign n2721 = \a[8]  & n2717 ;
  assign n2722 = ~n2707 & n2721 ;
  assign n2723 = ~n2704 & n2722 ;
  assign n2724 = ~n2720 & ~n2723 ;
  assign n2725 = ~n2469 & ~n2701 ;
  assign n2726 = ~n2561 & n2725 ;
  assign n2727 = ~n2724 & ~n2726 ;
  assign n2728 = ~n2702 & n2727 ;
  assign n2729 = ~n2701 & n2724 ;
  assign n2730 = n2562 & n2729 ;
  assign n2731 = n2701 & n2724 ;
  assign n2732 = ~n2562 & n2731 ;
  assign n2733 = ~n2730 & ~n2732 ;
  assign n2734 = ~n2728 & n2733 ;
  assign n2735 = n252 & ~n2079 ;
  assign n2736 = ~n2077 & n2735 ;
  assign n2737 = \b[17]  & n303 ;
  assign n2738 = n300 & n2737 ;
  assign n2739 = \b[19]  & n250 ;
  assign n2740 = \a[3]  & \b[18]  ;
  assign n2741 = n241 & n2740 ;
  assign n2742 = ~\a[3]  & \b[18]  ;
  assign n2743 = n244 & n2742 ;
  assign n2744 = ~n2741 & ~n2743 ;
  assign n2745 = ~n2739 & n2744 ;
  assign n2746 = ~n2738 & n2745 ;
  assign n2747 = ~n2736 & n2746 ;
  assign n2748 = ~\a[5]  & ~n2747 ;
  assign n2749 = \a[5]  & n2746 ;
  assign n2750 = ~n2736 & n2749 ;
  assign n2751 = ~n2748 & ~n2750 ;
  assign n2752 = ~n2734 & ~n2751 ;
  assign n2753 = n2560 & n2752 ;
  assign n2754 = n2734 & ~n2751 ;
  assign n2755 = ~n2560 & n2754 ;
  assign n2756 = ~n2753 & ~n2755 ;
  assign n2757 = ~n2734 & n2751 ;
  assign n2758 = ~n2560 & n2757 ;
  assign n2759 = n2734 & n2751 ;
  assign n2760 = n2560 & n2759 ;
  assign n2761 = ~n2758 & ~n2760 ;
  assign n2762 = n2756 & n2761 ;
  assign n2763 = ~n2292 & ~n2519 ;
  assign n2764 = ~n2516 & n2763 ;
  assign n2765 = ~n2518 & ~n2764 ;
  assign n2766 = ~\b[21]  & ~\b[22]  ;
  assign n2767 = \b[21]  & \b[22]  ;
  assign n2768 = ~n2766 & ~n2767 ;
  assign n2769 = ~n2765 & ~n2768 ;
  assign n2770 = ~n2518 & n2768 ;
  assign n2771 = ~n2764 & n2770 ;
  assign n2772 = n134 & ~n2771 ;
  assign n2773 = ~n2769 & n2772 ;
  assign n2774 = \a[0]  & \b[22]  ;
  assign n2775 = n133 & n2774 ;
  assign n2776 = \b[21]  & n141 ;
  assign n2777 = ~\a[1]  & \b[20]  ;
  assign n2778 = n1521 & n2777 ;
  assign n2779 = ~n2776 & ~n2778 ;
  assign n2780 = ~n2775 & n2779 ;
  assign n2781 = \a[2]  & n2780 ;
  assign n2782 = ~n2773 & n2781 ;
  assign n2783 = ~n2773 & n2780 ;
  assign n2784 = ~\a[2]  & ~n2783 ;
  assign n2785 = ~n2782 & ~n2784 ;
  assign n2786 = ~n2762 & n2785 ;
  assign n2787 = n2557 & n2786 ;
  assign n2788 = n2762 & n2785 ;
  assign n2789 = ~n2557 & n2788 ;
  assign n2790 = ~n2787 & ~n2789 ;
  assign n2791 = ~n2557 & n2762 ;
  assign n2792 = ~n2508 & ~n2762 ;
  assign n2793 = ~n2556 & n2792 ;
  assign n2794 = ~n2785 & ~n2793 ;
  assign n2795 = ~n2791 & n2794 ;
  assign n2796 = n2790 & ~n2795 ;
  assign n2797 = n2555 & n2796 ;
  assign n2798 = ~n2555 & ~n2796 ;
  assign n2799 = ~n2797 & ~n2798 ;
  assign n2800 = ~n2795 & ~n2797 ;
  assign n2801 = ~n2508 & n2756 ;
  assign n2802 = ~n2556 & n2801 ;
  assign n2803 = n2761 & ~n2802 ;
  assign n2804 = n2560 & n2734 ;
  assign n2805 = ~n2728 & ~n2804 ;
  assign n2806 = ~n2469 & n2700 ;
  assign n2807 = ~n2561 & n2806 ;
  assign n2808 = n2695 & ~n2807 ;
  assign n2809 = n430 & ~n1694 ;
  assign n2810 = ~n1692 & n2809 ;
  assign n2811 = \b[15]  & n486 ;
  assign n2812 = n483 & n2811 ;
  assign n2813 = \b[17]  & n428 ;
  assign n2814 = \a[5]  & \b[16]  ;
  assign n2815 = n484 & n2814 ;
  assign n2816 = ~\a[6]  & \b[16]  ;
  assign n2817 = n422 & n2816 ;
  assign n2818 = ~n2815 & ~n2817 ;
  assign n2819 = ~n2813 & n2818 ;
  assign n2820 = ~n2812 & n2819 ;
  assign n2821 = ~n2810 & n2820 ;
  assign n2822 = ~\a[8]  & ~n2821 ;
  assign n2823 = \a[8]  & n2820 ;
  assign n2824 = ~n2810 & n2823 ;
  assign n2825 = ~n2822 & ~n2824 ;
  assign n2826 = n2565 & n2673 ;
  assign n2827 = n2667 & ~n2826 ;
  assign n2828 = ~n728 & n999 ;
  assign n2829 = ~n726 & n2828 ;
  assign n2830 = \b[9]  & n1182 ;
  assign n2831 = n1179 & n2830 ;
  assign n2832 = ~\a[11]  & \b[10]  ;
  assign n2833 = n1181 & n2832 ;
  assign n2834 = ~n2831 & ~n2833 ;
  assign n2835 = \b[11]  & n997 ;
  assign n2836 = \a[12]  & \b[10]  ;
  assign n2837 = n988 & n2836 ;
  assign n2838 = \a[14]  & ~n2837 ;
  assign n2839 = ~n2835 & n2838 ;
  assign n2840 = n2834 & n2839 ;
  assign n2841 = ~n2829 & n2840 ;
  assign n2842 = ~n2835 & ~n2837 ;
  assign n2843 = n2834 & n2842 ;
  assign n2844 = ~n2829 & n2843 ;
  assign n2845 = ~\a[14]  & ~n2844 ;
  assign n2846 = ~n2841 & ~n2845 ;
  assign n2847 = ~n2446 & ~n2636 ;
  assign n2848 = ~n2566 & n2847 ;
  assign n2849 = ~n2637 & ~n2848 ;
  assign n2850 = ~n505 & ~n1304 ;
  assign n2851 = ~n1464 & n2850 ;
  assign n2852 = n502 & n2851 ;
  assign n2853 = n505 & ~n1304 ;
  assign n2854 = ~n1464 & n2853 ;
  assign n2855 = ~n502 & n2854 ;
  assign n2856 = ~n2852 & ~n2855 ;
  assign n2857 = \b[6]  & n1652 ;
  assign n2858 = n1649 & n2857 ;
  assign n2859 = ~\a[15]  & \b[7]  ;
  assign n2860 = n1459 & n2859 ;
  assign n2861 = ~n2858 & ~n2860 ;
  assign n2862 = \b[8]  & n1465 ;
  assign n2863 = \a[15]  & \b[7]  ;
  assign n2864 = n1456 & n2863 ;
  assign n2865 = \a[17]  & ~n2864 ;
  assign n2866 = ~n2862 & n2865 ;
  assign n2867 = n2861 & n2866 ;
  assign n2868 = n2856 & n2867 ;
  assign n2869 = ~n2862 & ~n2864 ;
  assign n2870 = n2861 & n2869 ;
  assign n2871 = n2856 & n2870 ;
  assign n2872 = ~\a[17]  & ~n2871 ;
  assign n2873 = ~n2868 & ~n2872 ;
  assign n2874 = ~n2630 & ~n2633 ;
  assign n2875 = ~n270 & n1965 ;
  assign n2876 = ~n218 & n1965 ;
  assign n2877 = ~n220 & n2876 ;
  assign n2878 = ~n2875 & ~n2877 ;
  assign n2879 = ~n273 & ~n2878 ;
  assign n2880 = \b[3]  & n2218 ;
  assign n2881 = n2216 & n2880 ;
  assign n2882 = \b[5]  & n1963 ;
  assign n2883 = \a[17]  & \b[4]  ;
  assign n2884 = n1954 & n2883 ;
  assign n2885 = ~\a[18]  & \b[4]  ;
  assign n2886 = n1957 & n2885 ;
  assign n2887 = ~n2884 & ~n2886 ;
  assign n2888 = ~n2882 & n2887 ;
  assign n2889 = ~n2881 & n2888 ;
  assign n2890 = ~\a[20]  & n2889 ;
  assign n2891 = ~n2879 & n2890 ;
  assign n2892 = \a[20]  & ~n2889 ;
  assign n2893 = \a[20]  & ~n273 ;
  assign n2894 = ~n2878 & n2893 ;
  assign n2895 = ~n2892 & ~n2894 ;
  assign n2896 = ~n2891 & n2895 ;
  assign n2897 = \a[23]  & ~n2414 ;
  assign n2898 = n2616 & n2897 ;
  assign n2899 = n2624 & n2898 ;
  assign n2900 = \a[23]  & ~n2899 ;
  assign n2901 = \b[2]  & n2620 ;
  assign n2902 = ~\a[21]  & \b[1]  ;
  assign n2903 = n2614 & n2902 ;
  assign n2904 = \a[21]  & \b[1]  ;
  assign n2905 = n2611 & n2904 ;
  assign n2906 = ~n2903 & ~n2905 ;
  assign n2907 = ~n2901 & n2906 ;
  assign n2908 = n157 & n2622 ;
  assign n2909 = n2413 & ~n2619 ;
  assign n2910 = \a[21]  & ~\a[22]  ;
  assign n2911 = ~\a[21]  & \a[22]  ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = \b[0]  & n2912 ;
  assign n2914 = n2909 & n2913 ;
  assign n2915 = ~n2908 & ~n2914 ;
  assign n2916 = n2907 & n2915 ;
  assign n2917 = ~n2900 & ~n2916 ;
  assign n2918 = n2900 & n2916 ;
  assign n2919 = ~n2917 & ~n2918 ;
  assign n2920 = n2896 & ~n2919 ;
  assign n2921 = ~n2896 & n2919 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = ~n2874 & n2922 ;
  assign n2924 = ~n2630 & ~n2922 ;
  assign n2925 = ~n2633 & n2924 ;
  assign n2926 = ~n2923 & ~n2925 ;
  assign n2927 = n2873 & ~n2926 ;
  assign n2928 = ~n2873 & ~n2925 ;
  assign n2929 = ~n2923 & n2928 ;
  assign n2930 = ~n2927 & ~n2929 ;
  assign n2931 = n2849 & n2930 ;
  assign n2932 = ~n2849 & ~n2930 ;
  assign n2933 = ~n2931 & ~n2932 ;
  assign n2934 = n2846 & ~n2933 ;
  assign n2935 = ~n2846 & n2933 ;
  assign n2936 = ~n2934 & ~n2935 ;
  assign n2937 = ~n551 & ~n946 ;
  assign n2938 = ~n1087 & n2937 ;
  assign n2939 = ~n1083 & n2938 ;
  assign n2940 = ~n643 & n2939 ;
  assign n2941 = n646 & n1087 ;
  assign n2942 = ~n1084 & n2941 ;
  assign n2943 = ~n2940 & ~n2942 ;
  assign n2944 = \b[12]  & n796 ;
  assign n2945 = n793 & n2944 ;
  assign n2946 = ~\a[9]  & \b[13]  ;
  assign n2947 = n638 & n2946 ;
  assign n2948 = ~n2945 & ~n2947 ;
  assign n2949 = \b[14]  & n644 ;
  assign n2950 = \a[9]  & \b[13]  ;
  assign n2951 = n635 & n2950 ;
  assign n2952 = \a[11]  & ~n2951 ;
  assign n2953 = ~n2949 & n2952 ;
  assign n2954 = n2948 & n2953 ;
  assign n2955 = n2943 & n2954 ;
  assign n2956 = ~n2949 & ~n2951 ;
  assign n2957 = n2948 & n2956 ;
  assign n2958 = n2943 & n2957 ;
  assign n2959 = ~\a[11]  & ~n2958 ;
  assign n2960 = ~n2955 & ~n2959 ;
  assign n2961 = ~n2936 & ~n2960 ;
  assign n2962 = ~n2827 & n2961 ;
  assign n2963 = n2936 & ~n2960 ;
  assign n2964 = n2827 & n2963 ;
  assign n2965 = ~n2962 & ~n2964 ;
  assign n2966 = ~n2936 & n2960 ;
  assign n2967 = n2827 & n2966 ;
  assign n2968 = n2936 & n2960 ;
  assign n2969 = ~n2827 & n2968 ;
  assign n2970 = ~n2967 & ~n2969 ;
  assign n2971 = n2965 & n2970 ;
  assign n2972 = ~n2825 & ~n2971 ;
  assign n2973 = n2808 & n2972 ;
  assign n2974 = ~n2825 & n2971 ;
  assign n2975 = ~n2808 & n2974 ;
  assign n2976 = ~n2973 & ~n2975 ;
  assign n2977 = n2825 & ~n2971 ;
  assign n2978 = ~n2808 & n2977 ;
  assign n2979 = n2825 & n2971 ;
  assign n2980 = n2808 & n2979 ;
  assign n2981 = ~n2978 & ~n2980 ;
  assign n2982 = n2976 & n2981 ;
  assign n2983 = ~n2805 & n2982 ;
  assign n2984 = n252 & n2293 ;
  assign n2985 = ~n2290 & n2984 ;
  assign n2986 = n252 & ~n2293 ;
  assign n2987 = ~n2074 & n2986 ;
  assign n2988 = ~n2289 & n2987 ;
  assign n2989 = \b[18]  & n303 ;
  assign n2990 = n300 & n2989 ;
  assign n2991 = \b[20]  & n250 ;
  assign n2992 = \a[3]  & \b[19]  ;
  assign n2993 = n241 & n2992 ;
  assign n2994 = ~\a[3]  & \b[19]  ;
  assign n2995 = n244 & n2994 ;
  assign n2996 = ~n2993 & ~n2995 ;
  assign n2997 = ~n2991 & n2996 ;
  assign n2998 = ~n2990 & n2997 ;
  assign n2999 = ~n2988 & n2998 ;
  assign n3000 = ~n2985 & n2999 ;
  assign n3001 = ~\a[5]  & ~n3000 ;
  assign n3002 = \a[5]  & n2998 ;
  assign n3003 = ~n2988 & n3002 ;
  assign n3004 = ~n2985 & n3003 ;
  assign n3005 = ~n3001 & ~n3004 ;
  assign n3006 = ~n2728 & ~n2982 ;
  assign n3007 = ~n2804 & n3006 ;
  assign n3008 = ~n3005 & ~n3007 ;
  assign n3009 = ~n2983 & n3008 ;
  assign n3010 = ~n2982 & n3005 ;
  assign n3011 = n2805 & n3010 ;
  assign n3012 = n2982 & n3005 ;
  assign n3013 = ~n2805 & n3012 ;
  assign n3014 = ~n3011 & ~n3013 ;
  assign n3015 = ~n3009 & n3014 ;
  assign n3016 = ~n2767 & ~n2771 ;
  assign n3017 = ~\b[22]  & ~\b[23]  ;
  assign n3018 = \b[22]  & \b[23]  ;
  assign n3019 = ~n3017 & ~n3018 ;
  assign n3020 = ~n3016 & n3019 ;
  assign n3021 = ~n2767 & ~n3019 ;
  assign n3022 = ~n2771 & n3021 ;
  assign n3023 = n134 & ~n3022 ;
  assign n3024 = ~n3020 & n3023 ;
  assign n3025 = \a[0]  & \b[23]  ;
  assign n3026 = n133 & n3025 ;
  assign n3027 = \b[22]  & n141 ;
  assign n3028 = ~\a[1]  & \b[21]  ;
  assign n3029 = n1521 & n3028 ;
  assign n3030 = ~n3027 & ~n3029 ;
  assign n3031 = ~n3026 & n3030 ;
  assign n3032 = ~n3024 & n3031 ;
  assign n3033 = ~\a[2]  & ~n3032 ;
  assign n3034 = \a[2]  & n3031 ;
  assign n3035 = ~n3024 & n3034 ;
  assign n3036 = ~n3033 & ~n3035 ;
  assign n3037 = ~n3015 & ~n3036 ;
  assign n3038 = n2803 & n3037 ;
  assign n3039 = n3015 & ~n3036 ;
  assign n3040 = ~n2803 & n3039 ;
  assign n3041 = ~n3038 & ~n3040 ;
  assign n3042 = ~n3015 & n3036 ;
  assign n3043 = ~n2803 & n3042 ;
  assign n3044 = n3015 & n3036 ;
  assign n3045 = n2803 & n3044 ;
  assign n3046 = ~n3043 & ~n3045 ;
  assign n3047 = n3041 & n3046 ;
  assign n3048 = ~n2800 & n3047 ;
  assign n3049 = ~n2795 & ~n3047 ;
  assign n3050 = ~n2797 & n3049 ;
  assign n3051 = ~n3048 & ~n3050 ;
  assign n3052 = ~n2795 & n3041 ;
  assign n3053 = ~n2797 & n3052 ;
  assign n3054 = n3046 & ~n3053 ;
  assign n3055 = n2803 & n3015 ;
  assign n3056 = ~n3009 & ~n3055 ;
  assign n3057 = n252 & ~n2523 ;
  assign n3058 = ~n2521 & n3057 ;
  assign n3059 = \b[19]  & n303 ;
  assign n3060 = n300 & n3059 ;
  assign n3061 = \b[21]  & n250 ;
  assign n3062 = \a[3]  & \b[20]  ;
  assign n3063 = n241 & n3062 ;
  assign n3064 = ~\a[3]  & \b[20]  ;
  assign n3065 = n244 & n3064 ;
  assign n3066 = ~n3063 & ~n3065 ;
  assign n3067 = ~n3061 & n3066 ;
  assign n3068 = ~n3060 & n3067 ;
  assign n3069 = ~n3058 & n3068 ;
  assign n3070 = ~\a[5]  & ~n3069 ;
  assign n3071 = \a[5]  & n3068 ;
  assign n3072 = ~n3058 & n3071 ;
  assign n3073 = ~n3070 & ~n3072 ;
  assign n3074 = ~n2728 & n2976 ;
  assign n3075 = n2981 & ~n3074 ;
  assign n3076 = n2734 & n2981 ;
  assign n3077 = n2560 & n3076 ;
  assign n3078 = ~n3075 & ~n3077 ;
  assign n3079 = n2808 & n2971 ;
  assign n3080 = n2965 & ~n3079 ;
  assign n3081 = n2667 & ~n2935 ;
  assign n3082 = ~n2826 & n3081 ;
  assign n3083 = ~n2934 & ~n3082 ;
  assign n3084 = ~n2929 & ~n2931 ;
  assign n3085 = ~n847 & ~n909 ;
  assign n3086 = ~n996 & n3085 ;
  assign n3087 = n906 & n3086 ;
  assign n3088 = ~n847 & n909 ;
  assign n3089 = ~n996 & n3088 ;
  assign n3090 = ~n906 & n3089 ;
  assign n3091 = ~n3087 & ~n3090 ;
  assign n3092 = \b[10]  & n1182 ;
  assign n3093 = n1179 & n3092 ;
  assign n3094 = ~\a[11]  & \b[11]  ;
  assign n3095 = n1181 & n3094 ;
  assign n3096 = ~n3093 & ~n3095 ;
  assign n3097 = \b[12]  & n997 ;
  assign n3098 = \a[12]  & \b[11]  ;
  assign n3099 = n988 & n3098 ;
  assign n3100 = \a[14]  & ~n3099 ;
  assign n3101 = ~n3097 & n3100 ;
  assign n3102 = n3096 & n3101 ;
  assign n3103 = n3091 & n3102 ;
  assign n3104 = ~n3097 & ~n3099 ;
  assign n3105 = n3096 & n3104 ;
  assign n3106 = n3091 & n3105 ;
  assign n3107 = ~\a[14]  & ~n3106 ;
  assign n3108 = ~n3103 & ~n3107 ;
  assign n3109 = ~n2630 & ~n2920 ;
  assign n3110 = ~n2633 & n3109 ;
  assign n3111 = ~n2921 & ~n3110 ;
  assign n3112 = ~n586 & n1467 ;
  assign n3113 = ~n504 & n1467 ;
  assign n3114 = ~n508 & n3113 ;
  assign n3115 = ~n3112 & ~n3114 ;
  assign n3116 = ~n589 & ~n3115 ;
  assign n3117 = \b[7]  & n1652 ;
  assign n3118 = n1649 & n3117 ;
  assign n3119 = ~\a[15]  & \b[8]  ;
  assign n3120 = n1459 & n3119 ;
  assign n3121 = ~n3118 & ~n3120 ;
  assign n3122 = \b[9]  & n1465 ;
  assign n3123 = \a[15]  & \b[8]  ;
  assign n3124 = n1456 & n3123 ;
  assign n3125 = \a[17]  & ~n3124 ;
  assign n3126 = ~n3122 & n3125 ;
  assign n3127 = n3121 & n3126 ;
  assign n3128 = ~n3116 & n3127 ;
  assign n3129 = ~n3122 & ~n3124 ;
  assign n3130 = n3121 & n3129 ;
  assign n3131 = ~\a[17]  & ~n3130 ;
  assign n3132 = ~\a[17]  & ~n589 ;
  assign n3133 = ~n3115 & n3132 ;
  assign n3134 = ~n3131 & ~n3133 ;
  assign n3135 = ~n3128 & n3134 ;
  assign n3136 = n177 & n2622 ;
  assign n3137 = \b[3]  & n2620 ;
  assign n3138 = \a[20]  & \b[2]  ;
  assign n3139 = n2910 & n3138 ;
  assign n3140 = ~\a[21]  & \b[2]  ;
  assign n3141 = n2614 & n3140 ;
  assign n3142 = ~n3139 & ~n3141 ;
  assign n3143 = ~n3137 & n3142 ;
  assign n3144 = ~n3136 & n3143 ;
  assign n3145 = \b[1]  & n2912 ;
  assign n3146 = n2909 & n3145 ;
  assign n3147 = ~\a[23]  & ~n3146 ;
  assign n3148 = n3144 & n3147 ;
  assign n3149 = n3144 & ~n3146 ;
  assign n3150 = \a[23]  & ~n3149 ;
  assign n3151 = ~n3148 & ~n3150 ;
  assign n3152 = \a[23]  & ~\a[24]  ;
  assign n3153 = ~\a[23]  & \a[24]  ;
  assign n3154 = ~n3152 & ~n3153 ;
  assign n3155 = \b[0]  & ~n3154 ;
  assign n3156 = n2899 & n2916 ;
  assign n3157 = n3155 & n3156 ;
  assign n3158 = ~n3155 & ~n3156 ;
  assign n3159 = ~n3157 & ~n3158 ;
  assign n3160 = n3151 & n3159 ;
  assign n3161 = ~n3151 & ~n3159 ;
  assign n3162 = ~n3160 & ~n3161 ;
  assign n3163 = ~n323 & ~n1805 ;
  assign n3164 = ~n1962 & n3163 ;
  assign n3165 = n320 & n3164 ;
  assign n3166 = n323 & ~n1805 ;
  assign n3167 = ~n1962 & n3166 ;
  assign n3168 = ~n320 & n3167 ;
  assign n3169 = ~n3165 & ~n3168 ;
  assign n3170 = \b[4]  & n2218 ;
  assign n3171 = n2216 & n3170 ;
  assign n3172 = \b[6]  & n1963 ;
  assign n3173 = \a[17]  & \b[5]  ;
  assign n3174 = n1954 & n3173 ;
  assign n3175 = ~\a[18]  & \b[5]  ;
  assign n3176 = n1957 & n3175 ;
  assign n3177 = ~n3174 & ~n3176 ;
  assign n3178 = ~n3172 & n3177 ;
  assign n3179 = ~n3171 & n3178 ;
  assign n3180 = n3169 & n3179 ;
  assign n3181 = ~\a[20]  & ~n3180 ;
  assign n3182 = \a[20]  & n3179 ;
  assign n3183 = n3169 & n3182 ;
  assign n3184 = ~n3181 & ~n3183 ;
  assign n3185 = n3162 & ~n3184 ;
  assign n3186 = ~n3162 & n3184 ;
  assign n3187 = ~n3185 & ~n3186 ;
  assign n3188 = ~n3135 & ~n3187 ;
  assign n3189 = n3111 & n3188 ;
  assign n3190 = ~n3135 & n3187 ;
  assign n3191 = ~n3111 & n3190 ;
  assign n3192 = ~n3189 & ~n3191 ;
  assign n3193 = n3135 & ~n3187 ;
  assign n3194 = ~n3111 & n3193 ;
  assign n3195 = n3135 & n3187 ;
  assign n3196 = n3111 & n3195 ;
  assign n3197 = ~n3194 & ~n3196 ;
  assign n3198 = n3192 & n3197 ;
  assign n3199 = n3108 & ~n3198 ;
  assign n3200 = n3084 & n3199 ;
  assign n3201 = n3108 & n3198 ;
  assign n3202 = ~n3084 & n3201 ;
  assign n3203 = ~n3200 & ~n3202 ;
  assign n3204 = ~n3084 & n3198 ;
  assign n3205 = ~n2929 & ~n3198 ;
  assign n3206 = ~n2931 & n3205 ;
  assign n3207 = ~n3108 & ~n3206 ;
  assign n3208 = ~n3204 & n3207 ;
  assign n3209 = n3203 & ~n3208 ;
  assign n3210 = n646 & ~n1233 ;
  assign n3211 = ~n1231 & n3210 ;
  assign n3212 = \b[15]  & n644 ;
  assign n3213 = \a[9]  & \b[14]  ;
  assign n3214 = n635 & n3213 ;
  assign n3215 = ~n3212 & ~n3214 ;
  assign n3216 = \b[13]  & n796 ;
  assign n3217 = n793 & n3216 ;
  assign n3218 = ~\a[9]  & \b[14]  ;
  assign n3219 = n638 & n3218 ;
  assign n3220 = ~n3217 & ~n3219 ;
  assign n3221 = n3215 & n3220 ;
  assign n3222 = ~n3211 & n3221 ;
  assign n3223 = ~\a[11]  & ~n3222 ;
  assign n3224 = \a[11]  & n3221 ;
  assign n3225 = ~n3211 & n3224 ;
  assign n3226 = ~n3223 & ~n3225 ;
  assign n3227 = ~n3209 & ~n3226 ;
  assign n3228 = n3083 & n3227 ;
  assign n3229 = n3209 & ~n3226 ;
  assign n3230 = ~n3083 & n3229 ;
  assign n3231 = ~n3228 & ~n3230 ;
  assign n3232 = ~n3209 & n3226 ;
  assign n3233 = ~n3083 & n3232 ;
  assign n3234 = n3209 & n3226 ;
  assign n3235 = n3083 & n3234 ;
  assign n3236 = ~n3233 & ~n3235 ;
  assign n3237 = n3231 & n3236 ;
  assign n3238 = n430 & n1875 ;
  assign n3239 = ~n1872 & n3238 ;
  assign n3240 = n430 & ~n1875 ;
  assign n3241 = ~n1689 & n3240 ;
  assign n3242 = ~n1871 & n3241 ;
  assign n3243 = \b[16]  & n486 ;
  assign n3244 = n483 & n3243 ;
  assign n3245 = \b[18]  & n428 ;
  assign n3246 = \a[6]  & \b[17]  ;
  assign n3247 = n419 & n3246 ;
  assign n3248 = ~\a[6]  & \b[17]  ;
  assign n3249 = n422 & n3248 ;
  assign n3250 = ~n3247 & ~n3249 ;
  assign n3251 = ~n3245 & n3250 ;
  assign n3252 = ~n3244 & n3251 ;
  assign n3253 = ~n3242 & n3252 ;
  assign n3254 = ~n3239 & n3253 ;
  assign n3255 = ~\a[8]  & ~n3254 ;
  assign n3256 = \a[8]  & n3252 ;
  assign n3257 = ~n3242 & n3256 ;
  assign n3258 = ~n3239 & n3257 ;
  assign n3259 = ~n3255 & ~n3258 ;
  assign n3260 = ~n3237 & n3259 ;
  assign n3261 = n3080 & n3260 ;
  assign n3262 = n3237 & n3259 ;
  assign n3263 = ~n3080 & n3262 ;
  assign n3264 = ~n3261 & ~n3263 ;
  assign n3265 = ~n3080 & n3237 ;
  assign n3266 = n2965 & ~n3237 ;
  assign n3267 = ~n3079 & n3266 ;
  assign n3268 = ~n3259 & ~n3267 ;
  assign n3269 = ~n3265 & n3268 ;
  assign n3270 = n3264 & ~n3269 ;
  assign n3271 = ~n3078 & n3270 ;
  assign n3272 = n3078 & ~n3270 ;
  assign n3273 = ~n3271 & ~n3272 ;
  assign n3274 = ~n3073 & n3273 ;
  assign n3275 = n3073 & ~n3273 ;
  assign n3276 = ~n3274 & ~n3275 ;
  assign n3277 = ~n3056 & n3276 ;
  assign n3278 = ~n2767 & ~n3018 ;
  assign n3279 = ~n2771 & n3278 ;
  assign n3280 = ~n3017 & ~n3279 ;
  assign n3281 = ~\b[23]  & ~\b[24]  ;
  assign n3282 = \b[23]  & \b[24]  ;
  assign n3283 = ~n3281 & ~n3282 ;
  assign n3284 = n134 & n3283 ;
  assign n3285 = ~n3280 & n3284 ;
  assign n3286 = n134 & ~n3283 ;
  assign n3287 = ~n3017 & n3286 ;
  assign n3288 = ~n3279 & n3287 ;
  assign n3289 = \a[0]  & \b[24]  ;
  assign n3290 = n133 & n3289 ;
  assign n3291 = \b[23]  & n141 ;
  assign n3292 = ~\a[1]  & \b[22]  ;
  assign n3293 = n1521 & n3292 ;
  assign n3294 = ~n3291 & ~n3293 ;
  assign n3295 = ~n3290 & n3294 ;
  assign n3296 = \a[2]  & n3295 ;
  assign n3297 = ~n3288 & n3296 ;
  assign n3298 = ~n3285 & n3297 ;
  assign n3299 = ~n3288 & n3295 ;
  assign n3300 = ~n3285 & n3299 ;
  assign n3301 = ~\a[2]  & ~n3300 ;
  assign n3302 = ~n3298 & ~n3301 ;
  assign n3303 = ~n3009 & ~n3276 ;
  assign n3304 = ~n3055 & n3303 ;
  assign n3305 = ~n3302 & ~n3304 ;
  assign n3306 = ~n3277 & n3305 ;
  assign n3307 = ~n3276 & n3302 ;
  assign n3308 = n3056 & n3307 ;
  assign n3309 = n3276 & n3302 ;
  assign n3310 = ~n3056 & n3309 ;
  assign n3311 = ~n3308 & ~n3310 ;
  assign n3312 = ~n3306 & n3311 ;
  assign n3313 = n3054 & n3312 ;
  assign n3314 = ~n3054 & ~n3312 ;
  assign n3315 = ~n3313 & ~n3314 ;
  assign n3316 = ~n3306 & ~n3313 ;
  assign n3317 = ~n3009 & ~n3274 ;
  assign n3318 = ~n3055 & n3317 ;
  assign n3319 = ~n3275 & ~n3318 ;
  assign n3320 = ~n3269 & ~n3271 ;
  assign n3321 = n252 & ~n2771 ;
  assign n3322 = ~n2769 & n3321 ;
  assign n3323 = \b[20]  & n303 ;
  assign n3324 = n300 & n3323 ;
  assign n3325 = \b[22]  & n250 ;
  assign n3326 = \a[3]  & \b[21]  ;
  assign n3327 = n241 & n3326 ;
  assign n3328 = ~\a[3]  & \b[21]  ;
  assign n3329 = n244 & n3328 ;
  assign n3330 = ~n3327 & ~n3329 ;
  assign n3331 = ~n3325 & n3330 ;
  assign n3332 = ~n3324 & n3331 ;
  assign n3333 = ~n3322 & n3332 ;
  assign n3334 = ~\a[5]  & ~n3333 ;
  assign n3335 = \a[5]  & n3332 ;
  assign n3336 = ~n3322 & n3335 ;
  assign n3337 = ~n3334 & ~n3336 ;
  assign n3338 = n2965 & n3231 ;
  assign n3339 = ~n3079 & n3338 ;
  assign n3340 = n3236 & ~n3339 ;
  assign n3341 = n3083 & n3209 ;
  assign n3342 = ~n3208 & ~n3341 ;
  assign n3343 = ~n2929 & n3192 ;
  assign n3344 = ~n2931 & n3343 ;
  assign n3345 = n3197 & ~n3344 ;
  assign n3346 = n3111 & n3187 ;
  assign n3347 = ~n3185 & ~n3346 ;
  assign n3348 = ~n380 & n1965 ;
  assign n3349 = ~n322 & n1965 ;
  assign n3350 = ~n326 & n3349 ;
  assign n3351 = ~n3348 & ~n3350 ;
  assign n3352 = ~n383 & ~n3351 ;
  assign n3353 = \b[5]  & n2218 ;
  assign n3354 = n2216 & n3353 ;
  assign n3355 = \b[7]  & n1963 ;
  assign n3356 = \a[17]  & \b[6]  ;
  assign n3357 = n1954 & n3356 ;
  assign n3358 = ~\a[18]  & \b[6]  ;
  assign n3359 = n1957 & n3358 ;
  assign n3360 = ~n3357 & ~n3359 ;
  assign n3361 = ~n3355 & n3360 ;
  assign n3362 = ~n3354 & n3361 ;
  assign n3363 = ~\a[20]  & n3362 ;
  assign n3364 = ~n3352 & n3363 ;
  assign n3365 = \a[20]  & ~n3362 ;
  assign n3366 = \a[20]  & ~n383 ;
  assign n3367 = ~n3351 & n3366 ;
  assign n3368 = ~n3365 & ~n3367 ;
  assign n3369 = ~n3364 & n3368 ;
  assign n3370 = ~n3157 & ~n3160 ;
  assign n3371 = n222 & n2622 ;
  assign n3372 = \b[4]  & n2620 ;
  assign n3373 = \a[20]  & \b[3]  ;
  assign n3374 = n2910 & n3373 ;
  assign n3375 = ~\a[21]  & \b[3]  ;
  assign n3376 = n2614 & n3375 ;
  assign n3377 = ~n3374 & ~n3376 ;
  assign n3378 = ~n3372 & n3377 ;
  assign n3379 = \b[2]  & n2912 ;
  assign n3380 = n2909 & n3379 ;
  assign n3381 = \a[23]  & ~n3380 ;
  assign n3382 = n3378 & n3381 ;
  assign n3383 = ~n3371 & n3382 ;
  assign n3384 = n3378 & ~n3380 ;
  assign n3385 = ~n3371 & n3384 ;
  assign n3386 = ~\a[23]  & ~n3385 ;
  assign n3387 = ~n3383 & ~n3386 ;
  assign n3388 = \a[26]  & \b[0]  ;
  assign n3389 = ~n3154 & n3388 ;
  assign n3390 = \a[24]  & \b[0]  ;
  assign n3391 = \a[23]  & ~\a[25]  ;
  assign n3392 = n3390 & n3391 ;
  assign n3393 = ~\a[24]  & \b[0]  ;
  assign n3394 = ~\a[23]  & \a[25]  ;
  assign n3395 = n3393 & n3394 ;
  assign n3396 = ~n3392 & ~n3395 ;
  assign n3397 = \a[25]  & ~\a[26]  ;
  assign n3398 = ~\a[25]  & \a[26]  ;
  assign n3399 = ~n3397 & ~n3398 ;
  assign n3400 = ~n3154 & n3399 ;
  assign n3401 = \b[1]  & n3400 ;
  assign n3402 = ~n3154 & ~n3399 ;
  assign n3403 = ~n137 & n3402 ;
  assign n3404 = ~n3401 & ~n3403 ;
  assign n3405 = n3396 & n3404 ;
  assign n3406 = n3389 & ~n3405 ;
  assign n3407 = ~n3389 & n3396 ;
  assign n3408 = n3404 & n3407 ;
  assign n3409 = ~n3406 & ~n3408 ;
  assign n3410 = ~n3387 & n3409 ;
  assign n3411 = n3387 & ~n3409 ;
  assign n3412 = ~n3410 & ~n3411 ;
  assign n3413 = ~n3370 & n3412 ;
  assign n3414 = n3370 & ~n3412 ;
  assign n3415 = ~n3413 & ~n3414 ;
  assign n3416 = n3369 & n3415 ;
  assign n3417 = ~n3369 & ~n3415 ;
  assign n3418 = ~n3416 & ~n3417 ;
  assign n3419 = ~n685 & ~n1304 ;
  assign n3420 = ~n1464 & n3419 ;
  assign n3421 = n682 & n3420 ;
  assign n3422 = n685 & ~n1304 ;
  assign n3423 = ~n1464 & n3422 ;
  assign n3424 = ~n682 & n3423 ;
  assign n3425 = ~n3421 & ~n3424 ;
  assign n3426 = \b[8]  & n1652 ;
  assign n3427 = n1649 & n3426 ;
  assign n3428 = ~\a[15]  & \b[9]  ;
  assign n3429 = n1459 & n3428 ;
  assign n3430 = ~n3427 & ~n3429 ;
  assign n3431 = \b[10]  & n1465 ;
  assign n3432 = \a[15]  & \b[9]  ;
  assign n3433 = n1456 & n3432 ;
  assign n3434 = \a[17]  & ~n3433 ;
  assign n3435 = ~n3431 & n3434 ;
  assign n3436 = n3430 & n3435 ;
  assign n3437 = n3425 & n3436 ;
  assign n3438 = ~n3431 & ~n3433 ;
  assign n3439 = n3430 & n3438 ;
  assign n3440 = n3425 & n3439 ;
  assign n3441 = ~\a[17]  & ~n3440 ;
  assign n3442 = ~n3437 & ~n3441 ;
  assign n3443 = ~n3418 & ~n3442 ;
  assign n3444 = ~n3347 & n3443 ;
  assign n3445 = n3418 & ~n3442 ;
  assign n3446 = n3347 & n3445 ;
  assign n3447 = ~n3444 & ~n3446 ;
  assign n3448 = ~n3418 & n3442 ;
  assign n3449 = n3347 & n3448 ;
  assign n3450 = n3418 & n3442 ;
  assign n3451 = ~n3347 & n3450 ;
  assign n3452 = ~n3449 & ~n3451 ;
  assign n3453 = n3447 & n3452 ;
  assign n3454 = ~n951 & n999 ;
  assign n3455 = ~n949 & n3454 ;
  assign n3456 = \b[11]  & n1182 ;
  assign n3457 = n1179 & n3456 ;
  assign n3458 = ~\a[11]  & \b[12]  ;
  assign n3459 = n1181 & n3458 ;
  assign n3460 = ~n3457 & ~n3459 ;
  assign n3461 = \b[13]  & n997 ;
  assign n3462 = \a[12]  & \b[12]  ;
  assign n3463 = n988 & n3462 ;
  assign n3464 = \a[14]  & ~n3463 ;
  assign n3465 = ~n3461 & n3464 ;
  assign n3466 = n3460 & n3465 ;
  assign n3467 = ~n3455 & n3466 ;
  assign n3468 = ~n3461 & ~n3463 ;
  assign n3469 = n3460 & n3468 ;
  assign n3470 = ~n3455 & n3469 ;
  assign n3471 = ~\a[14]  & ~n3470 ;
  assign n3472 = ~n3467 & ~n3471 ;
  assign n3473 = ~n3453 & n3472 ;
  assign n3474 = ~n3345 & n3473 ;
  assign n3475 = n3453 & n3472 ;
  assign n3476 = n3345 & n3475 ;
  assign n3477 = ~n3474 & ~n3476 ;
  assign n3478 = ~n3453 & ~n3472 ;
  assign n3479 = n3345 & n3478 ;
  assign n3480 = n3453 & ~n3472 ;
  assign n3481 = ~n3345 & n3480 ;
  assign n3482 = ~n3479 & ~n3481 ;
  assign n3483 = n3477 & n3482 ;
  assign n3484 = n646 & n1512 ;
  assign n3485 = ~n1509 & n3484 ;
  assign n3486 = n646 & ~n1512 ;
  assign n3487 = ~n1228 & n3486 ;
  assign n3488 = ~n1508 & n3487 ;
  assign n3489 = \b[14]  & n796 ;
  assign n3490 = n793 & n3489 ;
  assign n3491 = ~\a[9]  & \b[15]  ;
  assign n3492 = n638 & n3491 ;
  assign n3493 = ~n3490 & ~n3492 ;
  assign n3494 = \b[16]  & n644 ;
  assign n3495 = \a[9]  & \b[15]  ;
  assign n3496 = n635 & n3495 ;
  assign n3497 = \a[11]  & ~n3496 ;
  assign n3498 = ~n3494 & n3497 ;
  assign n3499 = n3493 & n3498 ;
  assign n3500 = ~n3488 & n3499 ;
  assign n3501 = ~n3485 & n3500 ;
  assign n3502 = ~n3494 & ~n3496 ;
  assign n3503 = n3493 & n3502 ;
  assign n3504 = ~n3488 & n3503 ;
  assign n3505 = ~n3485 & n3504 ;
  assign n3506 = ~\a[11]  & ~n3505 ;
  assign n3507 = ~n3501 & ~n3506 ;
  assign n3508 = ~n3483 & ~n3507 ;
  assign n3509 = ~n3342 & n3508 ;
  assign n3510 = n3483 & ~n3507 ;
  assign n3511 = n3342 & n3510 ;
  assign n3512 = ~n3509 & ~n3511 ;
  assign n3513 = ~n3342 & ~n3483 ;
  assign n3514 = ~n3208 & n3483 ;
  assign n3515 = ~n3341 & n3514 ;
  assign n3516 = n3507 & ~n3515 ;
  assign n3517 = ~n3513 & n3516 ;
  assign n3518 = n3512 & ~n3517 ;
  assign n3519 = n430 & ~n2079 ;
  assign n3520 = ~n2077 & n3519 ;
  assign n3521 = \b[17]  & n486 ;
  assign n3522 = n483 & n3521 ;
  assign n3523 = \b[19]  & n428 ;
  assign n3524 = \a[6]  & \b[18]  ;
  assign n3525 = n419 & n3524 ;
  assign n3526 = ~\a[6]  & \b[18]  ;
  assign n3527 = n422 & n3526 ;
  assign n3528 = ~n3525 & ~n3527 ;
  assign n3529 = ~n3523 & n3528 ;
  assign n3530 = ~n3522 & n3529 ;
  assign n3531 = ~n3520 & n3530 ;
  assign n3532 = ~\a[8]  & ~n3531 ;
  assign n3533 = \a[8]  & n3530 ;
  assign n3534 = ~n3520 & n3533 ;
  assign n3535 = ~n3532 & ~n3534 ;
  assign n3536 = ~n3518 & ~n3535 ;
  assign n3537 = n3340 & n3536 ;
  assign n3538 = n3518 & ~n3535 ;
  assign n3539 = ~n3340 & n3538 ;
  assign n3540 = ~n3537 & ~n3539 ;
  assign n3541 = ~n3518 & n3535 ;
  assign n3542 = ~n3340 & n3541 ;
  assign n3543 = n3518 & n3535 ;
  assign n3544 = n3340 & n3543 ;
  assign n3545 = ~n3542 & ~n3544 ;
  assign n3546 = n3540 & n3545 ;
  assign n3547 = ~n3337 & ~n3546 ;
  assign n3548 = ~n3320 & n3547 ;
  assign n3549 = ~n3337 & n3546 ;
  assign n3550 = n3320 & n3549 ;
  assign n3551 = ~n3548 & ~n3550 ;
  assign n3552 = n3337 & ~n3546 ;
  assign n3553 = n3320 & n3552 ;
  assign n3554 = n3337 & n3546 ;
  assign n3555 = ~n3320 & n3554 ;
  assign n3556 = ~n3553 & ~n3555 ;
  assign n3557 = n3551 & n3556 ;
  assign n3558 = ~n3319 & ~n3557 ;
  assign n3559 = ~n3017 & n3283 ;
  assign n3560 = ~n3279 & n3559 ;
  assign n3561 = ~n3282 & ~n3560 ;
  assign n3562 = ~\b[24]  & ~\b[25]  ;
  assign n3563 = \b[24]  & \b[25]  ;
  assign n3564 = ~n3562 & ~n3563 ;
  assign n3565 = ~n3561 & n3564 ;
  assign n3566 = ~n3282 & ~n3564 ;
  assign n3567 = ~n3560 & n3566 ;
  assign n3568 = n134 & ~n3567 ;
  assign n3569 = ~n3565 & n3568 ;
  assign n3570 = \a[0]  & \b[25]  ;
  assign n3571 = n133 & n3570 ;
  assign n3572 = \b[24]  & n141 ;
  assign n3573 = ~\a[1]  & \b[23]  ;
  assign n3574 = n1521 & n3573 ;
  assign n3575 = ~n3572 & ~n3574 ;
  assign n3576 = ~n3571 & n3575 ;
  assign n3577 = ~n3569 & n3576 ;
  assign n3578 = ~\a[2]  & ~n3577 ;
  assign n3579 = \a[2]  & n3576 ;
  assign n3580 = ~n3569 & n3579 ;
  assign n3581 = ~n3578 & ~n3580 ;
  assign n3582 = ~n3275 & n3557 ;
  assign n3583 = ~n3318 & n3582 ;
  assign n3584 = ~n3581 & ~n3583 ;
  assign n3585 = ~n3558 & n3584 ;
  assign n3586 = ~n3557 & n3581 ;
  assign n3587 = ~n3319 & n3586 ;
  assign n3588 = n3557 & n3581 ;
  assign n3589 = n3319 & n3588 ;
  assign n3590 = ~n3587 & ~n3589 ;
  assign n3591 = ~n3585 & n3590 ;
  assign n3592 = ~n3316 & n3591 ;
  assign n3593 = ~n3306 & ~n3591 ;
  assign n3594 = ~n3313 & n3593 ;
  assign n3595 = ~n3592 & ~n3594 ;
  assign n3596 = ~n3306 & ~n3585 ;
  assign n3597 = ~n3313 & n3596 ;
  assign n3598 = n3551 & ~n3583 ;
  assign n3599 = ~n3282 & ~n3563 ;
  assign n3600 = ~n3560 & n3599 ;
  assign n3601 = ~n3562 & ~n3600 ;
  assign n3602 = ~\b[25]  & ~\b[26]  ;
  assign n3603 = \b[25]  & \b[26]  ;
  assign n3604 = ~n3602 & ~n3603 ;
  assign n3605 = n134 & n3604 ;
  assign n3606 = ~n3601 & n3605 ;
  assign n3607 = n134 & ~n3604 ;
  assign n3608 = ~n3562 & n3607 ;
  assign n3609 = ~n3600 & n3608 ;
  assign n3610 = \a[0]  & \b[26]  ;
  assign n3611 = n133 & n3610 ;
  assign n3612 = \b[25]  & n141 ;
  assign n3613 = ~\a[1]  & \b[24]  ;
  assign n3614 = n1521 & n3613 ;
  assign n3615 = ~n3612 & ~n3614 ;
  assign n3616 = ~n3611 & n3615 ;
  assign n3617 = \a[2]  & n3616 ;
  assign n3618 = ~n3609 & n3617 ;
  assign n3619 = ~n3606 & n3618 ;
  assign n3620 = ~n3609 & n3616 ;
  assign n3621 = ~n3606 & n3620 ;
  assign n3622 = ~\a[2]  & ~n3621 ;
  assign n3623 = ~n3619 & ~n3622 ;
  assign n3624 = ~n3269 & n3540 ;
  assign n3625 = ~n3271 & n3624 ;
  assign n3626 = n3545 & ~n3625 ;
  assign n3627 = n3340 & n3518 ;
  assign n3628 = n3512 & ~n3627 ;
  assign n3629 = ~n3208 & n3482 ;
  assign n3630 = ~n3341 & n3629 ;
  assign n3631 = n3477 & ~n3630 ;
  assign n3632 = n646 & ~n1694 ;
  assign n3633 = ~n1692 & n3632 ;
  assign n3634 = \b[17]  & n644 ;
  assign n3635 = \a[9]  & \b[16]  ;
  assign n3636 = n635 & n3635 ;
  assign n3637 = ~n3634 & ~n3636 ;
  assign n3638 = \b[15]  & n796 ;
  assign n3639 = n793 & n3638 ;
  assign n3640 = ~\a[9]  & \b[16]  ;
  assign n3641 = n638 & n3640 ;
  assign n3642 = ~n3639 & ~n3641 ;
  assign n3643 = n3637 & n3642 ;
  assign n3644 = ~n3633 & n3643 ;
  assign n3645 = ~\a[11]  & ~n3644 ;
  assign n3646 = \a[11]  & n3643 ;
  assign n3647 = ~n3633 & n3646 ;
  assign n3648 = ~n3645 & ~n3647 ;
  assign n3649 = n3345 & n3453 ;
  assign n3650 = n3447 & ~n3649 ;
  assign n3651 = ~n728 & n1467 ;
  assign n3652 = ~n726 & n3651 ;
  assign n3653 = \b[9]  & n1652 ;
  assign n3654 = n1649 & n3653 ;
  assign n3655 = ~\a[15]  & \b[10]  ;
  assign n3656 = n1459 & n3655 ;
  assign n3657 = ~n3654 & ~n3656 ;
  assign n3658 = \b[11]  & n1465 ;
  assign n3659 = \a[15]  & \b[10]  ;
  assign n3660 = n1456 & n3659 ;
  assign n3661 = \a[17]  & ~n3660 ;
  assign n3662 = ~n3658 & n3661 ;
  assign n3663 = n3657 & n3662 ;
  assign n3664 = ~n3652 & n3663 ;
  assign n3665 = ~n3658 & ~n3660 ;
  assign n3666 = n3657 & n3665 ;
  assign n3667 = ~n3652 & n3666 ;
  assign n3668 = ~\a[17]  & ~n3667 ;
  assign n3669 = ~n3664 & ~n3668 ;
  assign n3670 = ~n3185 & ~n3416 ;
  assign n3671 = ~n3346 & n3670 ;
  assign n3672 = ~n3417 & ~n3671 ;
  assign n3673 = ~n505 & ~n1805 ;
  assign n3674 = ~n1962 & n3673 ;
  assign n3675 = n502 & n3674 ;
  assign n3676 = n505 & ~n1805 ;
  assign n3677 = ~n1962 & n3676 ;
  assign n3678 = ~n502 & n3677 ;
  assign n3679 = ~n3675 & ~n3678 ;
  assign n3680 = \b[6]  & n2218 ;
  assign n3681 = n2216 & n3680 ;
  assign n3682 = \b[8]  & n1963 ;
  assign n3683 = \a[17]  & \b[7]  ;
  assign n3684 = n1954 & n3683 ;
  assign n3685 = ~\a[18]  & \b[7]  ;
  assign n3686 = n1957 & n3685 ;
  assign n3687 = ~n3684 & ~n3686 ;
  assign n3688 = ~n3682 & n3687 ;
  assign n3689 = ~n3681 & n3688 ;
  assign n3690 = n3679 & n3689 ;
  assign n3691 = ~\a[20]  & ~n3690 ;
  assign n3692 = \a[20]  & n3689 ;
  assign n3693 = n3679 & n3692 ;
  assign n3694 = ~n3691 & ~n3693 ;
  assign n3695 = ~n3410 & ~n3413 ;
  assign n3696 = ~n270 & n2622 ;
  assign n3697 = ~n218 & n2622 ;
  assign n3698 = ~n220 & n3697 ;
  assign n3699 = ~n3696 & ~n3698 ;
  assign n3700 = ~n273 & ~n3699 ;
  assign n3701 = \b[3]  & n2912 ;
  assign n3702 = n2909 & n3701 ;
  assign n3703 = \b[5]  & n2620 ;
  assign n3704 = \a[20]  & \b[4]  ;
  assign n3705 = n2910 & n3704 ;
  assign n3706 = ~\a[21]  & \b[4]  ;
  assign n3707 = n2614 & n3706 ;
  assign n3708 = ~n3705 & ~n3707 ;
  assign n3709 = ~n3703 & n3708 ;
  assign n3710 = ~n3702 & n3709 ;
  assign n3711 = ~\a[23]  & n3710 ;
  assign n3712 = ~n3700 & n3711 ;
  assign n3713 = \a[23]  & ~n3710 ;
  assign n3714 = \a[23]  & ~n273 ;
  assign n3715 = ~n3699 & n3714 ;
  assign n3716 = ~n3713 & ~n3715 ;
  assign n3717 = ~n3712 & n3716 ;
  assign n3718 = \a[26]  & ~n3155 ;
  assign n3719 = n3396 & n3718 ;
  assign n3720 = n3404 & n3719 ;
  assign n3721 = \a[26]  & ~n3720 ;
  assign n3722 = \b[2]  & n3400 ;
  assign n3723 = ~\a[24]  & \b[1]  ;
  assign n3724 = n3394 & n3723 ;
  assign n3725 = \a[24]  & \b[1]  ;
  assign n3726 = n3391 & n3725 ;
  assign n3727 = ~n3724 & ~n3726 ;
  assign n3728 = ~n3722 & n3727 ;
  assign n3729 = n157 & n3402 ;
  assign n3730 = n3154 & ~n3399 ;
  assign n3731 = \a[24]  & ~\a[25]  ;
  assign n3732 = ~\a[24]  & \a[25]  ;
  assign n3733 = ~n3731 & ~n3732 ;
  assign n3734 = \b[0]  & n3733 ;
  assign n3735 = n3730 & n3734 ;
  assign n3736 = ~n3729 & ~n3735 ;
  assign n3737 = n3728 & n3736 ;
  assign n3738 = ~n3721 & ~n3737 ;
  assign n3739 = n3721 & n3737 ;
  assign n3740 = ~n3738 & ~n3739 ;
  assign n3741 = n3717 & ~n3740 ;
  assign n3742 = ~n3717 & n3740 ;
  assign n3743 = ~n3741 & ~n3742 ;
  assign n3744 = ~n3695 & n3743 ;
  assign n3745 = ~n3410 & ~n3743 ;
  assign n3746 = ~n3413 & n3745 ;
  assign n3747 = ~n3744 & ~n3746 ;
  assign n3748 = n3694 & ~n3747 ;
  assign n3749 = ~n3694 & ~n3746 ;
  assign n3750 = ~n3744 & n3749 ;
  assign n3751 = ~n3748 & ~n3750 ;
  assign n3752 = n3672 & n3751 ;
  assign n3753 = ~n3672 & ~n3751 ;
  assign n3754 = ~n3752 & ~n3753 ;
  assign n3755 = n3669 & ~n3754 ;
  assign n3756 = ~n3669 & n3754 ;
  assign n3757 = ~n3755 & ~n3756 ;
  assign n3758 = n999 & n1087 ;
  assign n3759 = ~n1084 & n3758 ;
  assign n3760 = n999 & n1552 ;
  assign n3761 = ~n1083 & n3760 ;
  assign n3762 = \b[12]  & n1182 ;
  assign n3763 = n1179 & n3762 ;
  assign n3764 = ~\a[11]  & \b[13]  ;
  assign n3765 = n1181 & n3764 ;
  assign n3766 = ~n3763 & ~n3765 ;
  assign n3767 = \b[14]  & n997 ;
  assign n3768 = \a[12]  & \b[13]  ;
  assign n3769 = n988 & n3768 ;
  assign n3770 = \a[14]  & ~n3769 ;
  assign n3771 = ~n3767 & n3770 ;
  assign n3772 = n3766 & n3771 ;
  assign n3773 = ~n3761 & n3772 ;
  assign n3774 = ~n3759 & n3773 ;
  assign n3775 = ~n3767 & ~n3769 ;
  assign n3776 = n3766 & n3775 ;
  assign n3777 = ~n3761 & n3776 ;
  assign n3778 = ~n3759 & n3777 ;
  assign n3779 = ~\a[14]  & ~n3778 ;
  assign n3780 = ~n3774 & ~n3779 ;
  assign n3781 = ~n3757 & ~n3780 ;
  assign n3782 = ~n3650 & n3781 ;
  assign n3783 = n3757 & ~n3780 ;
  assign n3784 = n3650 & n3783 ;
  assign n3785 = ~n3782 & ~n3784 ;
  assign n3786 = ~n3757 & n3780 ;
  assign n3787 = n3650 & n3786 ;
  assign n3788 = n3757 & n3780 ;
  assign n3789 = ~n3650 & n3788 ;
  assign n3790 = ~n3787 & ~n3789 ;
  assign n3791 = n3785 & n3790 ;
  assign n3792 = ~n3648 & ~n3791 ;
  assign n3793 = n3631 & n3792 ;
  assign n3794 = ~n3648 & n3791 ;
  assign n3795 = ~n3631 & n3794 ;
  assign n3796 = ~n3793 & ~n3795 ;
  assign n3797 = n3648 & ~n3791 ;
  assign n3798 = ~n3631 & n3797 ;
  assign n3799 = n3648 & n3791 ;
  assign n3800 = n3631 & n3799 ;
  assign n3801 = ~n3798 & ~n3800 ;
  assign n3802 = n3796 & n3801 ;
  assign n3803 = ~n3628 & n3802 ;
  assign n3804 = n3512 & ~n3802 ;
  assign n3805 = ~n3627 & n3804 ;
  assign n3806 = n430 & n2293 ;
  assign n3807 = ~n2290 & n3806 ;
  assign n3808 = n430 & ~n2293 ;
  assign n3809 = ~n2074 & n3808 ;
  assign n3810 = ~n2289 & n3809 ;
  assign n3811 = \b[18]  & n486 ;
  assign n3812 = n483 & n3811 ;
  assign n3813 = \b[20]  & n428 ;
  assign n3814 = \a[6]  & \b[19]  ;
  assign n3815 = n419 & n3814 ;
  assign n3816 = ~\a[6]  & \b[19]  ;
  assign n3817 = n422 & n3816 ;
  assign n3818 = ~n3815 & ~n3817 ;
  assign n3819 = ~n3813 & n3818 ;
  assign n3820 = ~n3812 & n3819 ;
  assign n3821 = ~n3810 & n3820 ;
  assign n3822 = ~n3807 & n3821 ;
  assign n3823 = ~\a[8]  & ~n3822 ;
  assign n3824 = \a[8]  & n3820 ;
  assign n3825 = ~n3810 & n3824 ;
  assign n3826 = ~n3807 & n3825 ;
  assign n3827 = ~n3823 & ~n3826 ;
  assign n3828 = ~n3805 & ~n3827 ;
  assign n3829 = ~n3803 & n3828 ;
  assign n3830 = ~n3802 & n3827 ;
  assign n3831 = n3628 & n3830 ;
  assign n3832 = n3802 & n3827 ;
  assign n3833 = ~n3628 & n3832 ;
  assign n3834 = ~n3831 & ~n3833 ;
  assign n3835 = ~n3829 & n3834 ;
  assign n3836 = ~n3626 & ~n3835 ;
  assign n3837 = n3626 & n3835 ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = n252 & ~n3022 ;
  assign n3840 = ~n3020 & n3839 ;
  assign n3841 = \b[23]  & n250 ;
  assign n3842 = \a[3]  & \b[22]  ;
  assign n3843 = n241 & n3842 ;
  assign n3844 = ~n3841 & ~n3843 ;
  assign n3845 = \b[21]  & n303 ;
  assign n3846 = n300 & n3845 ;
  assign n3847 = ~\a[3]  & \b[22]  ;
  assign n3848 = n244 & n3847 ;
  assign n3849 = ~n3846 & ~n3848 ;
  assign n3850 = n3844 & n3849 ;
  assign n3851 = ~n3840 & n3850 ;
  assign n3852 = ~\a[5]  & ~n3851 ;
  assign n3853 = \a[5]  & n3850 ;
  assign n3854 = ~n3840 & n3853 ;
  assign n3855 = ~n3852 & ~n3854 ;
  assign n3856 = n3838 & ~n3855 ;
  assign n3857 = ~n3838 & n3855 ;
  assign n3858 = ~n3856 & ~n3857 ;
  assign n3859 = ~n3623 & ~n3858 ;
  assign n3860 = ~n3598 & n3859 ;
  assign n3861 = ~n3623 & n3858 ;
  assign n3862 = n3598 & n3861 ;
  assign n3863 = ~n3860 & ~n3862 ;
  assign n3864 = n3623 & ~n3858 ;
  assign n3865 = n3598 & n3864 ;
  assign n3866 = n3623 & n3858 ;
  assign n3867 = ~n3598 & n3866 ;
  assign n3868 = ~n3865 & ~n3867 ;
  assign n3869 = n3863 & n3868 ;
  assign n3870 = n3590 & n3869 ;
  assign n3871 = ~n3597 & n3870 ;
  assign n3872 = n3590 & ~n3597 ;
  assign n3873 = ~n3869 & ~n3872 ;
  assign n3874 = ~n3871 & ~n3873 ;
  assign n3875 = n3863 & ~n3871 ;
  assign n3876 = n3551 & ~n3856 ;
  assign n3877 = ~n3583 & n3876 ;
  assign n3878 = ~n3857 & ~n3877 ;
  assign n3879 = ~n3829 & ~n3837 ;
  assign n3880 = n3512 & n3796 ;
  assign n3881 = ~n3627 & n3880 ;
  assign n3882 = n3801 & ~n3881 ;
  assign n3883 = n3631 & n3791 ;
  assign n3884 = n3785 & ~n3883 ;
  assign n3885 = n3447 & ~n3756 ;
  assign n3886 = ~n3649 & n3885 ;
  assign n3887 = ~n3755 & ~n3886 ;
  assign n3888 = ~n3750 & ~n3752 ;
  assign n3889 = ~n909 & ~n1304 ;
  assign n3890 = ~n1464 & n3889 ;
  assign n3891 = n906 & n3890 ;
  assign n3892 = n909 & ~n1304 ;
  assign n3893 = ~n1464 & n3892 ;
  assign n3894 = ~n906 & n3893 ;
  assign n3895 = ~n3891 & ~n3894 ;
  assign n3896 = \b[10]  & n1652 ;
  assign n3897 = n1649 & n3896 ;
  assign n3898 = ~\a[15]  & \b[11]  ;
  assign n3899 = n1459 & n3898 ;
  assign n3900 = ~n3897 & ~n3899 ;
  assign n3901 = \b[12]  & n1465 ;
  assign n3902 = \a[15]  & \b[11]  ;
  assign n3903 = n1456 & n3902 ;
  assign n3904 = \a[17]  & ~n3903 ;
  assign n3905 = ~n3901 & n3904 ;
  assign n3906 = n3900 & n3905 ;
  assign n3907 = n3895 & n3906 ;
  assign n3908 = ~n3901 & ~n3903 ;
  assign n3909 = n3900 & n3908 ;
  assign n3910 = n3895 & n3909 ;
  assign n3911 = ~\a[17]  & ~n3910 ;
  assign n3912 = ~n3907 & ~n3911 ;
  assign n3913 = ~n3410 & ~n3741 ;
  assign n3914 = ~n3413 & n3913 ;
  assign n3915 = ~n3742 & ~n3914 ;
  assign n3916 = ~n586 & n1965 ;
  assign n3917 = ~n504 & n1965 ;
  assign n3918 = ~n508 & n3917 ;
  assign n3919 = ~n3916 & ~n3918 ;
  assign n3920 = ~n589 & ~n3919 ;
  assign n3921 = \b[7]  & n2218 ;
  assign n3922 = n2216 & n3921 ;
  assign n3923 = \b[9]  & n1963 ;
  assign n3924 = \a[17]  & \b[8]  ;
  assign n3925 = n1954 & n3924 ;
  assign n3926 = ~\a[18]  & \b[8]  ;
  assign n3927 = n1957 & n3926 ;
  assign n3928 = ~n3925 & ~n3927 ;
  assign n3929 = ~n3923 & n3928 ;
  assign n3930 = ~n3922 & n3929 ;
  assign n3931 = ~\a[20]  & n3930 ;
  assign n3932 = ~n3920 & n3931 ;
  assign n3933 = \a[20]  & ~n3930 ;
  assign n3934 = \a[20]  & ~n589 ;
  assign n3935 = ~n3919 & n3934 ;
  assign n3936 = ~n3933 & ~n3935 ;
  assign n3937 = ~n3932 & n3936 ;
  assign n3938 = n177 & n3402 ;
  assign n3939 = \b[3]  & n3400 ;
  assign n3940 = \a[23]  & \b[2]  ;
  assign n3941 = n3731 & n3940 ;
  assign n3942 = ~\a[24]  & \b[2]  ;
  assign n3943 = n3394 & n3942 ;
  assign n3944 = ~n3941 & ~n3943 ;
  assign n3945 = ~n3939 & n3944 ;
  assign n3946 = ~n3938 & n3945 ;
  assign n3947 = \b[1]  & n3733 ;
  assign n3948 = n3730 & n3947 ;
  assign n3949 = ~\a[26]  & ~n3948 ;
  assign n3950 = n3946 & n3949 ;
  assign n3951 = n3946 & ~n3948 ;
  assign n3952 = \a[26]  & ~n3951 ;
  assign n3953 = ~n3950 & ~n3952 ;
  assign n3954 = \a[26]  & ~\a[27]  ;
  assign n3955 = ~\a[26]  & \a[27]  ;
  assign n3956 = ~n3954 & ~n3955 ;
  assign n3957 = \b[0]  & ~n3956 ;
  assign n3958 = n3720 & n3737 ;
  assign n3959 = n3957 & n3958 ;
  assign n3960 = ~n3957 & ~n3958 ;
  assign n3961 = ~n3959 & ~n3960 ;
  assign n3962 = n3953 & n3961 ;
  assign n3963 = ~n3953 & ~n3961 ;
  assign n3964 = ~n3962 & ~n3963 ;
  assign n3965 = ~n323 & ~n2413 ;
  assign n3966 = ~n2619 & n3965 ;
  assign n3967 = n320 & n3966 ;
  assign n3968 = n323 & ~n2413 ;
  assign n3969 = ~n2619 & n3968 ;
  assign n3970 = ~n320 & n3969 ;
  assign n3971 = ~n3967 & ~n3970 ;
  assign n3972 = \b[4]  & n2912 ;
  assign n3973 = n2909 & n3972 ;
  assign n3974 = \b[6]  & n2620 ;
  assign n3975 = \a[20]  & \b[5]  ;
  assign n3976 = n2910 & n3975 ;
  assign n3977 = ~\a[21]  & \b[5]  ;
  assign n3978 = n2614 & n3977 ;
  assign n3979 = ~n3976 & ~n3978 ;
  assign n3980 = ~n3974 & n3979 ;
  assign n3981 = ~n3973 & n3980 ;
  assign n3982 = n3971 & n3981 ;
  assign n3983 = ~\a[23]  & ~n3982 ;
  assign n3984 = \a[23]  & n3981 ;
  assign n3985 = n3971 & n3984 ;
  assign n3986 = ~n3983 & ~n3985 ;
  assign n3987 = n3964 & ~n3986 ;
  assign n3988 = ~n3964 & n3986 ;
  assign n3989 = ~n3987 & ~n3988 ;
  assign n3990 = n3937 & ~n3989 ;
  assign n3991 = n3915 & n3990 ;
  assign n3992 = n3937 & n3989 ;
  assign n3993 = ~n3915 & n3992 ;
  assign n3994 = ~n3991 & ~n3993 ;
  assign n3995 = ~n3937 & ~n3989 ;
  assign n3996 = ~n3915 & n3995 ;
  assign n3997 = ~n3937 & n3989 ;
  assign n3998 = n3915 & n3997 ;
  assign n3999 = ~n3996 & ~n3998 ;
  assign n4000 = n3994 & n3999 ;
  assign n4001 = n3912 & ~n4000 ;
  assign n4002 = n3888 & n4001 ;
  assign n4003 = n3912 & n4000 ;
  assign n4004 = ~n3888 & n4003 ;
  assign n4005 = ~n4002 & ~n4004 ;
  assign n4006 = ~n3888 & n4000 ;
  assign n4007 = ~n3750 & ~n4000 ;
  assign n4008 = ~n3752 & n4007 ;
  assign n4009 = ~n3912 & ~n4008 ;
  assign n4010 = ~n4006 & n4009 ;
  assign n4011 = n4005 & ~n4010 ;
  assign n4012 = n999 & ~n1233 ;
  assign n4013 = ~n1231 & n4012 ;
  assign n4014 = \b[13]  & n1182 ;
  assign n4015 = n1179 & n4014 ;
  assign n4016 = ~\a[11]  & \b[14]  ;
  assign n4017 = n1181 & n4016 ;
  assign n4018 = ~n4015 & ~n4017 ;
  assign n4019 = \b[15]  & n997 ;
  assign n4020 = \a[12]  & \b[14]  ;
  assign n4021 = n988 & n4020 ;
  assign n4022 = \a[14]  & ~n4021 ;
  assign n4023 = ~n4019 & n4022 ;
  assign n4024 = n4018 & n4023 ;
  assign n4025 = ~n4013 & n4024 ;
  assign n4026 = ~n4019 & ~n4021 ;
  assign n4027 = n4018 & n4026 ;
  assign n4028 = ~n4013 & n4027 ;
  assign n4029 = ~\a[14]  & ~n4028 ;
  assign n4030 = ~n4025 & ~n4029 ;
  assign n4031 = ~n4011 & ~n4030 ;
  assign n4032 = n3887 & n4031 ;
  assign n4033 = n4011 & ~n4030 ;
  assign n4034 = ~n3887 & n4033 ;
  assign n4035 = ~n4032 & ~n4034 ;
  assign n4036 = ~n4011 & n4030 ;
  assign n4037 = ~n3887 & n4036 ;
  assign n4038 = n4011 & n4030 ;
  assign n4039 = n3887 & n4038 ;
  assign n4040 = ~n4037 & ~n4039 ;
  assign n4041 = n4035 & n4040 ;
  assign n4042 = ~n3884 & n4041 ;
  assign n4043 = n3785 & ~n4041 ;
  assign n4044 = ~n3883 & n4043 ;
  assign n4045 = n646 & n1875 ;
  assign n4046 = ~n1872 & n4045 ;
  assign n4047 = n646 & ~n1875 ;
  assign n4048 = ~n1689 & n4047 ;
  assign n4049 = ~n1871 & n4048 ;
  assign n4050 = \b[16]  & n796 ;
  assign n4051 = n793 & n4050 ;
  assign n4052 = ~\a[9]  & \b[17]  ;
  assign n4053 = n638 & n4052 ;
  assign n4054 = ~n4051 & ~n4053 ;
  assign n4055 = \b[18]  & n644 ;
  assign n4056 = \a[9]  & \b[17]  ;
  assign n4057 = n635 & n4056 ;
  assign n4058 = \a[11]  & ~n4057 ;
  assign n4059 = ~n4055 & n4058 ;
  assign n4060 = n4054 & n4059 ;
  assign n4061 = ~n4049 & n4060 ;
  assign n4062 = ~n4046 & n4061 ;
  assign n4063 = ~n4055 & ~n4057 ;
  assign n4064 = n4054 & n4063 ;
  assign n4065 = ~n4049 & n4064 ;
  assign n4066 = ~n4046 & n4065 ;
  assign n4067 = ~\a[11]  & ~n4066 ;
  assign n4068 = ~n4062 & ~n4067 ;
  assign n4069 = ~n4044 & ~n4068 ;
  assign n4070 = ~n4042 & n4069 ;
  assign n4071 = ~n4041 & n4068 ;
  assign n4072 = n3884 & n4071 ;
  assign n4073 = n4041 & n4068 ;
  assign n4074 = ~n3884 & n4073 ;
  assign n4075 = ~n4072 & ~n4074 ;
  assign n4076 = ~n4070 & n4075 ;
  assign n4077 = n430 & ~n2523 ;
  assign n4078 = ~n2521 & n4077 ;
  assign n4079 = \b[19]  & n486 ;
  assign n4080 = n483 & n4079 ;
  assign n4081 = \b[21]  & n428 ;
  assign n4082 = \a[6]  & \b[20]  ;
  assign n4083 = n419 & n4082 ;
  assign n4084 = ~\a[6]  & \b[20]  ;
  assign n4085 = n422 & n4084 ;
  assign n4086 = ~n4083 & ~n4085 ;
  assign n4087 = ~n4081 & n4086 ;
  assign n4088 = ~n4080 & n4087 ;
  assign n4089 = ~n4078 & n4088 ;
  assign n4090 = ~\a[8]  & ~n4089 ;
  assign n4091 = \a[8]  & n4088 ;
  assign n4092 = ~n4078 & n4091 ;
  assign n4093 = ~n4090 & ~n4092 ;
  assign n4094 = ~n4076 & n4093 ;
  assign n4095 = ~n3882 & n4094 ;
  assign n4096 = n4076 & n4093 ;
  assign n4097 = n3882 & n4096 ;
  assign n4098 = ~n4095 & ~n4097 ;
  assign n4099 = ~n4076 & ~n4093 ;
  assign n4100 = n3882 & n4099 ;
  assign n4101 = n4076 & ~n4093 ;
  assign n4102 = ~n3882 & n4101 ;
  assign n4103 = ~n4100 & ~n4102 ;
  assign n4104 = n4098 & n4103 ;
  assign n4105 = n252 & n3283 ;
  assign n4106 = ~n3280 & n4105 ;
  assign n4107 = ~n3017 & ~n3283 ;
  assign n4108 = n252 & n4107 ;
  assign n4109 = ~n3279 & n4108 ;
  assign n4110 = \b[22]  & n303 ;
  assign n4111 = n300 & n4110 ;
  assign n4112 = ~\a[3]  & \b[23]  ;
  assign n4113 = n244 & n4112 ;
  assign n4114 = ~n4111 & ~n4113 ;
  assign n4115 = \b[24]  & n250 ;
  assign n4116 = \a[3]  & \b[23]  ;
  assign n4117 = n241 & n4116 ;
  assign n4118 = \a[5]  & ~n4117 ;
  assign n4119 = ~n4115 & n4118 ;
  assign n4120 = n4114 & n4119 ;
  assign n4121 = ~n4109 & n4120 ;
  assign n4122 = ~n4106 & n4121 ;
  assign n4123 = ~n4115 & ~n4117 ;
  assign n4124 = n4114 & n4123 ;
  assign n4125 = ~n4109 & n4124 ;
  assign n4126 = ~n4106 & n4125 ;
  assign n4127 = ~\a[5]  & ~n4126 ;
  assign n4128 = ~n4122 & ~n4127 ;
  assign n4129 = ~n4104 & ~n4128 ;
  assign n4130 = ~n3879 & n4129 ;
  assign n4131 = n4104 & ~n4128 ;
  assign n4132 = n3879 & n4131 ;
  assign n4133 = ~n4130 & ~n4132 ;
  assign n4134 = n4104 & n4128 ;
  assign n4135 = ~n3879 & n4134 ;
  assign n4136 = ~n4104 & n4128 ;
  assign n4137 = n3879 & n4136 ;
  assign n4138 = ~n4135 & ~n4137 ;
  assign n4139 = n4133 & n4138 ;
  assign n4140 = ~n3562 & n3604 ;
  assign n4141 = ~n3600 & n4140 ;
  assign n4142 = ~n3603 & ~n4141 ;
  assign n4143 = ~\b[26]  & ~\b[27]  ;
  assign n4144 = \b[26]  & \b[27]  ;
  assign n4145 = ~n4143 & ~n4144 ;
  assign n4146 = ~n4142 & n4145 ;
  assign n4147 = ~n3603 & ~n4145 ;
  assign n4148 = ~n4141 & n4147 ;
  assign n4149 = n134 & ~n4148 ;
  assign n4150 = ~n4146 & n4149 ;
  assign n4151 = \a[0]  & \b[27]  ;
  assign n4152 = n133 & n4151 ;
  assign n4153 = \b[26]  & n141 ;
  assign n4154 = ~\a[1]  & \b[25]  ;
  assign n4155 = n1521 & n4154 ;
  assign n4156 = ~n4153 & ~n4155 ;
  assign n4157 = ~n4152 & n4156 ;
  assign n4158 = ~n4150 & n4157 ;
  assign n4159 = ~\a[2]  & ~n4158 ;
  assign n4160 = \a[2]  & n4157 ;
  assign n4161 = ~n4150 & n4160 ;
  assign n4162 = ~n4159 & ~n4161 ;
  assign n4163 = ~n4139 & n4162 ;
  assign n4164 = ~n3878 & n4163 ;
  assign n4165 = n4139 & n4162 ;
  assign n4166 = n3878 & n4165 ;
  assign n4167 = ~n4164 & ~n4166 ;
  assign n4168 = ~n4139 & ~n4162 ;
  assign n4169 = n3878 & n4168 ;
  assign n4170 = n4139 & ~n4162 ;
  assign n4171 = ~n3878 & n4170 ;
  assign n4172 = ~n4169 & ~n4171 ;
  assign n4173 = n4167 & n4172 ;
  assign n4174 = ~n3875 & n4173 ;
  assign n4175 = n3863 & ~n4173 ;
  assign n4176 = ~n3871 & n4175 ;
  assign n4177 = ~n4174 & ~n4176 ;
  assign n4178 = n3863 & n4172 ;
  assign n4179 = ~n3871 & n4178 ;
  assign n4180 = n4167 & ~n4179 ;
  assign n4181 = n3878 & n4139 ;
  assign n4182 = n4133 & ~n4181 ;
  assign n4183 = n3882 & n4076 ;
  assign n4184 = ~n4070 & ~n4183 ;
  assign n4185 = n3785 & n4035 ;
  assign n4186 = ~n3883 & n4185 ;
  assign n4187 = n4040 & ~n4186 ;
  assign n4188 = n3887 & n4011 ;
  assign n4189 = ~n4010 & ~n4188 ;
  assign n4190 = ~n3750 & n3994 ;
  assign n4191 = ~n3752 & n4190 ;
  assign n4192 = n3999 & ~n4191 ;
  assign n4193 = n3915 & n3989 ;
  assign n4194 = ~n3987 & ~n4193 ;
  assign n4195 = ~n380 & n2622 ;
  assign n4196 = ~n322 & n2622 ;
  assign n4197 = ~n326 & n4196 ;
  assign n4198 = ~n4195 & ~n4197 ;
  assign n4199 = ~n383 & ~n4198 ;
  assign n4200 = \b[5]  & n2912 ;
  assign n4201 = n2909 & n4200 ;
  assign n4202 = \b[7]  & n2620 ;
  assign n4203 = \a[20]  & \b[6]  ;
  assign n4204 = n2910 & n4203 ;
  assign n4205 = ~\a[21]  & \b[6]  ;
  assign n4206 = n2614 & n4205 ;
  assign n4207 = ~n4204 & ~n4206 ;
  assign n4208 = ~n4202 & n4207 ;
  assign n4209 = ~n4201 & n4208 ;
  assign n4210 = ~\a[23]  & n4209 ;
  assign n4211 = ~n4199 & n4210 ;
  assign n4212 = \a[23]  & ~n4209 ;
  assign n4213 = \a[23]  & ~n383 ;
  assign n4214 = ~n4198 & n4213 ;
  assign n4215 = ~n4212 & ~n4214 ;
  assign n4216 = ~n4211 & n4215 ;
  assign n4217 = ~n3959 & ~n3962 ;
  assign n4218 = n222 & n3402 ;
  assign n4219 = \b[4]  & n3400 ;
  assign n4220 = \a[23]  & \b[3]  ;
  assign n4221 = n3731 & n4220 ;
  assign n4222 = ~\a[24]  & \b[3]  ;
  assign n4223 = n3394 & n4222 ;
  assign n4224 = ~n4221 & ~n4223 ;
  assign n4225 = ~n4219 & n4224 ;
  assign n4226 = \b[2]  & n3733 ;
  assign n4227 = n3730 & n4226 ;
  assign n4228 = \a[26]  & ~n4227 ;
  assign n4229 = n4225 & n4228 ;
  assign n4230 = ~n4218 & n4229 ;
  assign n4231 = n4225 & ~n4227 ;
  assign n4232 = ~n4218 & n4231 ;
  assign n4233 = ~\a[26]  & ~n4232 ;
  assign n4234 = ~n4230 & ~n4233 ;
  assign n4235 = \a[29]  & \b[0]  ;
  assign n4236 = ~n3956 & n4235 ;
  assign n4237 = \a[27]  & \b[0]  ;
  assign n4238 = \a[26]  & ~\a[28]  ;
  assign n4239 = n4237 & n4238 ;
  assign n4240 = ~\a[27]  & \b[0]  ;
  assign n4241 = ~\a[26]  & \a[28]  ;
  assign n4242 = n4240 & n4241 ;
  assign n4243 = ~n4239 & ~n4242 ;
  assign n4244 = \a[28]  & ~\a[29]  ;
  assign n4245 = ~\a[28]  & \a[29]  ;
  assign n4246 = ~n4244 & ~n4245 ;
  assign n4247 = ~n3956 & n4246 ;
  assign n4248 = \b[1]  & n4247 ;
  assign n4249 = ~n3956 & ~n4246 ;
  assign n4250 = ~n137 & n4249 ;
  assign n4251 = ~n4248 & ~n4250 ;
  assign n4252 = n4243 & n4251 ;
  assign n4253 = n4236 & ~n4252 ;
  assign n4254 = ~n4236 & n4243 ;
  assign n4255 = n4251 & n4254 ;
  assign n4256 = ~n4253 & ~n4255 ;
  assign n4257 = ~n4234 & n4256 ;
  assign n4258 = n4234 & ~n4256 ;
  assign n4259 = ~n4257 & ~n4258 ;
  assign n4260 = ~n4217 & n4259 ;
  assign n4261 = n4217 & ~n4259 ;
  assign n4262 = ~n4260 & ~n4261 ;
  assign n4263 = n4216 & n4262 ;
  assign n4264 = ~n4216 & ~n4262 ;
  assign n4265 = ~n4263 & ~n4264 ;
  assign n4266 = ~n685 & ~n1805 ;
  assign n4267 = ~n1962 & n4266 ;
  assign n4268 = n682 & n4267 ;
  assign n4269 = n685 & ~n1805 ;
  assign n4270 = ~n1962 & n4269 ;
  assign n4271 = ~n682 & n4270 ;
  assign n4272 = ~n4268 & ~n4271 ;
  assign n4273 = \b[8]  & n2218 ;
  assign n4274 = n2216 & n4273 ;
  assign n4275 = \b[10]  & n1963 ;
  assign n4276 = \a[17]  & \b[9]  ;
  assign n4277 = n1954 & n4276 ;
  assign n4278 = ~\a[18]  & \b[9]  ;
  assign n4279 = n1957 & n4278 ;
  assign n4280 = ~n4277 & ~n4279 ;
  assign n4281 = ~n4275 & n4280 ;
  assign n4282 = ~n4274 & n4281 ;
  assign n4283 = n4272 & n4282 ;
  assign n4284 = ~\a[20]  & ~n4283 ;
  assign n4285 = \a[20]  & n4282 ;
  assign n4286 = n4272 & n4285 ;
  assign n4287 = ~n4284 & ~n4286 ;
  assign n4288 = ~n4265 & ~n4287 ;
  assign n4289 = ~n4194 & n4288 ;
  assign n4290 = n4265 & ~n4287 ;
  assign n4291 = n4194 & n4290 ;
  assign n4292 = ~n4289 & ~n4291 ;
  assign n4293 = ~n4265 & n4287 ;
  assign n4294 = n4194 & n4293 ;
  assign n4295 = n4265 & n4287 ;
  assign n4296 = ~n4194 & n4295 ;
  assign n4297 = ~n4294 & ~n4296 ;
  assign n4298 = n4292 & n4297 ;
  assign n4299 = ~n948 & n1467 ;
  assign n4300 = ~n908 & n1467 ;
  assign n4301 = ~n912 & n4300 ;
  assign n4302 = ~n4299 & ~n4301 ;
  assign n4303 = ~n951 & ~n4302 ;
  assign n4304 = \b[11]  & n1652 ;
  assign n4305 = n1649 & n4304 ;
  assign n4306 = ~\a[15]  & \b[12]  ;
  assign n4307 = n1459 & n4306 ;
  assign n4308 = ~n4305 & ~n4307 ;
  assign n4309 = \b[13]  & n1465 ;
  assign n4310 = \a[15]  & \b[12]  ;
  assign n4311 = n1456 & n4310 ;
  assign n4312 = \a[17]  & ~n4311 ;
  assign n4313 = ~n4309 & n4312 ;
  assign n4314 = n4308 & n4313 ;
  assign n4315 = ~n4303 & n4314 ;
  assign n4316 = ~n4309 & ~n4311 ;
  assign n4317 = n4308 & n4316 ;
  assign n4318 = ~\a[17]  & ~n4317 ;
  assign n4319 = ~\a[17]  & ~n951 ;
  assign n4320 = ~n4302 & n4319 ;
  assign n4321 = ~n4318 & ~n4320 ;
  assign n4322 = ~n4315 & n4321 ;
  assign n4323 = ~n4298 & ~n4322 ;
  assign n4324 = n4192 & n4323 ;
  assign n4325 = n4298 & ~n4322 ;
  assign n4326 = ~n4192 & n4325 ;
  assign n4327 = ~n4324 & ~n4326 ;
  assign n4328 = ~n4298 & n4322 ;
  assign n4329 = ~n4192 & n4328 ;
  assign n4330 = n4298 & n4322 ;
  assign n4331 = n4192 & n4330 ;
  assign n4332 = ~n4329 & ~n4331 ;
  assign n4333 = n4327 & n4332 ;
  assign n4334 = ~n4189 & n4333 ;
  assign n4335 = n999 & n1512 ;
  assign n4336 = ~n1509 & n4335 ;
  assign n4337 = ~n1228 & ~n1512 ;
  assign n4338 = n999 & n4337 ;
  assign n4339 = ~n1508 & n4338 ;
  assign n4340 = \b[14]  & n1182 ;
  assign n4341 = n1179 & n4340 ;
  assign n4342 = ~\a[11]  & \b[15]  ;
  assign n4343 = n1181 & n4342 ;
  assign n4344 = ~n4341 & ~n4343 ;
  assign n4345 = \b[16]  & n997 ;
  assign n4346 = \a[12]  & \b[15]  ;
  assign n4347 = n988 & n4346 ;
  assign n4348 = \a[14]  & ~n4347 ;
  assign n4349 = ~n4345 & n4348 ;
  assign n4350 = n4344 & n4349 ;
  assign n4351 = ~n4339 & n4350 ;
  assign n4352 = ~n4336 & n4351 ;
  assign n4353 = ~n4345 & ~n4347 ;
  assign n4354 = n4344 & n4353 ;
  assign n4355 = ~n4339 & n4354 ;
  assign n4356 = ~n4336 & n4355 ;
  assign n4357 = ~\a[14]  & ~n4356 ;
  assign n4358 = ~n4352 & ~n4357 ;
  assign n4359 = ~n4010 & ~n4333 ;
  assign n4360 = ~n4188 & n4359 ;
  assign n4361 = ~n4358 & ~n4360 ;
  assign n4362 = ~n4334 & n4361 ;
  assign n4363 = ~n4333 & n4358 ;
  assign n4364 = n4189 & n4363 ;
  assign n4365 = n4333 & n4358 ;
  assign n4366 = ~n4189 & n4365 ;
  assign n4367 = ~n4364 & ~n4366 ;
  assign n4368 = ~n4362 & n4367 ;
  assign n4369 = n646 & ~n2079 ;
  assign n4370 = ~n2077 & n4369 ;
  assign n4371 = \b[19]  & n644 ;
  assign n4372 = \a[9]  & \b[18]  ;
  assign n4373 = n635 & n4372 ;
  assign n4374 = ~n4371 & ~n4373 ;
  assign n4375 = \b[17]  & n796 ;
  assign n4376 = n793 & n4375 ;
  assign n4377 = ~\a[9]  & \b[18]  ;
  assign n4378 = n638 & n4377 ;
  assign n4379 = ~n4376 & ~n4378 ;
  assign n4380 = n4374 & n4379 ;
  assign n4381 = ~n4370 & n4380 ;
  assign n4382 = ~\a[11]  & ~n4381 ;
  assign n4383 = \a[11]  & n4380 ;
  assign n4384 = ~n4370 & n4383 ;
  assign n4385 = ~n4382 & ~n4384 ;
  assign n4386 = ~n4368 & ~n4385 ;
  assign n4387 = n4187 & n4386 ;
  assign n4388 = n4368 & ~n4385 ;
  assign n4389 = ~n4187 & n4388 ;
  assign n4390 = ~n4387 & ~n4389 ;
  assign n4391 = ~n4368 & n4385 ;
  assign n4392 = ~n4187 & n4391 ;
  assign n4393 = n4368 & n4385 ;
  assign n4394 = n4187 & n4393 ;
  assign n4395 = ~n4392 & ~n4394 ;
  assign n4396 = n4390 & n4395 ;
  assign n4397 = n430 & ~n2771 ;
  assign n4398 = ~n2769 & n4397 ;
  assign n4399 = \b[20]  & n486 ;
  assign n4400 = n483 & n4399 ;
  assign n4401 = \b[22]  & n428 ;
  assign n4402 = \a[6]  & \b[21]  ;
  assign n4403 = n419 & n4402 ;
  assign n4404 = ~\a[6]  & \b[21]  ;
  assign n4405 = n422 & n4404 ;
  assign n4406 = ~n4403 & ~n4405 ;
  assign n4407 = ~n4401 & n4406 ;
  assign n4408 = ~n4400 & n4407 ;
  assign n4409 = ~n4398 & n4408 ;
  assign n4410 = ~\a[8]  & ~n4409 ;
  assign n4411 = \a[8]  & n4408 ;
  assign n4412 = ~n4398 & n4411 ;
  assign n4413 = ~n4410 & ~n4412 ;
  assign n4414 = ~n4396 & n4413 ;
  assign n4415 = n4184 & n4414 ;
  assign n4416 = n4396 & n4413 ;
  assign n4417 = ~n4184 & n4416 ;
  assign n4418 = ~n4415 & ~n4417 ;
  assign n4419 = ~n4184 & n4396 ;
  assign n4420 = ~n4070 & ~n4396 ;
  assign n4421 = ~n4183 & n4420 ;
  assign n4422 = ~n4413 & ~n4421 ;
  assign n4423 = ~n4419 & n4422 ;
  assign n4424 = n4418 & ~n4423 ;
  assign n4425 = ~n3829 & n4103 ;
  assign n4426 = ~n3837 & n4425 ;
  assign n4427 = n4098 & ~n4426 ;
  assign n4428 = n4424 & n4427 ;
  assign n4429 = ~n4424 & ~n4427 ;
  assign n4430 = ~n4428 & ~n4429 ;
  assign n4431 = n252 & ~n3567 ;
  assign n4432 = ~n3565 & n4431 ;
  assign n4433 = \b[25]  & n250 ;
  assign n4434 = \a[3]  & \b[24]  ;
  assign n4435 = n241 & n4434 ;
  assign n4436 = ~n4433 & ~n4435 ;
  assign n4437 = \b[23]  & n303 ;
  assign n4438 = n300 & n4437 ;
  assign n4439 = ~\a[3]  & \b[24]  ;
  assign n4440 = n244 & n4439 ;
  assign n4441 = ~n4438 & ~n4440 ;
  assign n4442 = n4436 & n4441 ;
  assign n4443 = ~n4432 & n4442 ;
  assign n4444 = ~\a[5]  & ~n4443 ;
  assign n4445 = \a[5]  & n4442 ;
  assign n4446 = ~n4432 & n4445 ;
  assign n4447 = ~n4444 & ~n4446 ;
  assign n4448 = n4430 & ~n4447 ;
  assign n4449 = ~n4430 & n4447 ;
  assign n4450 = ~n4448 & ~n4449 ;
  assign n4451 = ~n3603 & ~n4144 ;
  assign n4452 = ~n4141 & n4451 ;
  assign n4453 = ~n4143 & ~n4452 ;
  assign n4454 = ~\b[27]  & ~\b[28]  ;
  assign n4455 = \b[27]  & \b[28]  ;
  assign n4456 = ~n4454 & ~n4455 ;
  assign n4457 = n134 & n4456 ;
  assign n4458 = ~n4453 & n4457 ;
  assign n4459 = n134 & ~n4456 ;
  assign n4460 = ~n4143 & n4459 ;
  assign n4461 = ~n4452 & n4460 ;
  assign n4462 = \a[0]  & \b[28]  ;
  assign n4463 = n133 & n4462 ;
  assign n4464 = \b[27]  & n141 ;
  assign n4465 = ~\a[1]  & \b[26]  ;
  assign n4466 = n1521 & n4465 ;
  assign n4467 = ~n4464 & ~n4466 ;
  assign n4468 = ~n4463 & n4467 ;
  assign n4469 = \a[2]  & n4468 ;
  assign n4470 = ~n4461 & n4469 ;
  assign n4471 = ~n4458 & n4470 ;
  assign n4472 = ~n4461 & n4468 ;
  assign n4473 = ~n4458 & n4472 ;
  assign n4474 = ~\a[2]  & ~n4473 ;
  assign n4475 = ~n4471 & ~n4474 ;
  assign n4476 = ~n4450 & n4475 ;
  assign n4477 = n4182 & n4476 ;
  assign n4478 = n4450 & n4475 ;
  assign n4479 = ~n4182 & n4478 ;
  assign n4480 = ~n4477 & ~n4479 ;
  assign n4481 = ~n4450 & ~n4475 ;
  assign n4482 = ~n4182 & n4481 ;
  assign n4483 = n4450 & ~n4475 ;
  assign n4484 = n4182 & n4483 ;
  assign n4485 = ~n4482 & ~n4484 ;
  assign n4486 = n4480 & n4485 ;
  assign n4487 = n4180 & n4486 ;
  assign n4488 = ~n4180 & ~n4486 ;
  assign n4489 = ~n4487 & ~n4488 ;
  assign n4490 = n4485 & ~n4487 ;
  assign n4491 = n4133 & ~n4448 ;
  assign n4492 = ~n4181 & n4491 ;
  assign n4493 = ~n4449 & ~n4492 ;
  assign n4494 = ~n4143 & n4456 ;
  assign n4495 = ~n4452 & n4494 ;
  assign n4496 = ~n4455 & ~n4495 ;
  assign n4497 = ~\b[28]  & ~\b[29]  ;
  assign n4498 = \b[28]  & \b[29]  ;
  assign n4499 = ~n4497 & ~n4498 ;
  assign n4500 = ~n4496 & n4499 ;
  assign n4501 = ~n4455 & ~n4499 ;
  assign n4502 = ~n4495 & n4501 ;
  assign n4503 = n134 & ~n4502 ;
  assign n4504 = ~n4500 & n4503 ;
  assign n4505 = \a[0]  & \b[29]  ;
  assign n4506 = n133 & n4505 ;
  assign n4507 = \b[28]  & n141 ;
  assign n4508 = ~\a[1]  & \b[27]  ;
  assign n4509 = n1521 & n4508 ;
  assign n4510 = ~n4507 & ~n4509 ;
  assign n4511 = ~n4506 & n4510 ;
  assign n4512 = ~n4504 & n4511 ;
  assign n4513 = ~\a[2]  & ~n4512 ;
  assign n4514 = \a[2]  & n4511 ;
  assign n4515 = ~n4504 & n4514 ;
  assign n4516 = ~n4513 & ~n4515 ;
  assign n4517 = ~n4423 & ~n4428 ;
  assign n4518 = ~n3601 & ~n3604 ;
  assign n4519 = n252 & ~n4141 ;
  assign n4520 = ~n4518 & n4519 ;
  assign n4521 = \b[24]  & n303 ;
  assign n4522 = n300 & n4521 ;
  assign n4523 = ~\a[3]  & \b[25]  ;
  assign n4524 = n244 & n4523 ;
  assign n4525 = ~n4522 & ~n4524 ;
  assign n4526 = \b[26]  & n250 ;
  assign n4527 = \a[3]  & \b[25]  ;
  assign n4528 = n241 & n4527 ;
  assign n4529 = \a[5]  & ~n4528 ;
  assign n4530 = ~n4526 & n4529 ;
  assign n4531 = n4525 & n4530 ;
  assign n4532 = ~n4520 & n4531 ;
  assign n4533 = ~n4526 & ~n4528 ;
  assign n4534 = n4525 & n4533 ;
  assign n4535 = ~n4520 & n4534 ;
  assign n4536 = ~\a[5]  & ~n4535 ;
  assign n4537 = ~n4532 & ~n4536 ;
  assign n4538 = n430 & ~n3022 ;
  assign n4539 = ~n3020 & n4538 ;
  assign n4540 = \b[21]  & n486 ;
  assign n4541 = n483 & n4540 ;
  assign n4542 = \b[23]  & n428 ;
  assign n4543 = \a[6]  & \b[22]  ;
  assign n4544 = n419 & n4543 ;
  assign n4545 = ~\a[6]  & \b[22]  ;
  assign n4546 = n422 & n4545 ;
  assign n4547 = ~n4544 & ~n4546 ;
  assign n4548 = ~n4542 & n4547 ;
  assign n4549 = ~n4541 & n4548 ;
  assign n4550 = ~n4539 & n4549 ;
  assign n4551 = ~\a[8]  & ~n4550 ;
  assign n4552 = \a[8]  & n4549 ;
  assign n4553 = ~n4539 & n4552 ;
  assign n4554 = ~n4551 & ~n4553 ;
  assign n4555 = ~n4070 & n4390 ;
  assign n4556 = n4395 & ~n4555 ;
  assign n4557 = n4076 & n4395 ;
  assign n4558 = n3882 & n4557 ;
  assign n4559 = ~n4556 & ~n4558 ;
  assign n4560 = n4187 & n4368 ;
  assign n4561 = ~n4362 & ~n4560 ;
  assign n4562 = ~n4010 & n4327 ;
  assign n4563 = ~n4188 & n4562 ;
  assign n4564 = n4332 & ~n4563 ;
  assign n4565 = n4192 & n4298 ;
  assign n4566 = n4292 & ~n4565 ;
  assign n4567 = ~n728 & n1965 ;
  assign n4568 = ~n726 & n4567 ;
  assign n4569 = \b[9]  & n2218 ;
  assign n4570 = n2216 & n4569 ;
  assign n4571 = \b[11]  & n1963 ;
  assign n4572 = \a[17]  & \b[10]  ;
  assign n4573 = n1954 & n4572 ;
  assign n4574 = ~\a[18]  & \b[10]  ;
  assign n4575 = n1957 & n4574 ;
  assign n4576 = ~n4573 & ~n4575 ;
  assign n4577 = ~n4571 & n4576 ;
  assign n4578 = ~n4570 & n4577 ;
  assign n4579 = ~\a[20]  & n4578 ;
  assign n4580 = ~n4568 & n4579 ;
  assign n4581 = ~n4568 & n4578 ;
  assign n4582 = \a[20]  & ~n4581 ;
  assign n4583 = ~n4580 & ~n4582 ;
  assign n4584 = ~n3987 & ~n4263 ;
  assign n4585 = ~n4193 & n4584 ;
  assign n4586 = ~n4264 & ~n4585 ;
  assign n4587 = ~n505 & ~n2413 ;
  assign n4588 = ~n2619 & n4587 ;
  assign n4589 = n502 & n4588 ;
  assign n4590 = n505 & ~n2413 ;
  assign n4591 = ~n2619 & n4590 ;
  assign n4592 = ~n502 & n4591 ;
  assign n4593 = ~n4589 & ~n4592 ;
  assign n4594 = \b[6]  & n2912 ;
  assign n4595 = n2909 & n4594 ;
  assign n4596 = \b[8]  & n2620 ;
  assign n4597 = \a[20]  & \b[7]  ;
  assign n4598 = n2910 & n4597 ;
  assign n4599 = ~\a[21]  & \b[7]  ;
  assign n4600 = n2614 & n4599 ;
  assign n4601 = ~n4598 & ~n4600 ;
  assign n4602 = ~n4596 & n4601 ;
  assign n4603 = ~n4595 & n4602 ;
  assign n4604 = n4593 & n4603 ;
  assign n4605 = ~\a[23]  & ~n4604 ;
  assign n4606 = \a[23]  & n4603 ;
  assign n4607 = n4593 & n4606 ;
  assign n4608 = ~n4605 & ~n4607 ;
  assign n4609 = ~n4257 & ~n4260 ;
  assign n4610 = ~n270 & n3402 ;
  assign n4611 = ~n218 & n3402 ;
  assign n4612 = ~n220 & n4611 ;
  assign n4613 = ~n4610 & ~n4612 ;
  assign n4614 = ~n273 & ~n4613 ;
  assign n4615 = \b[3]  & n3733 ;
  assign n4616 = n3730 & n4615 ;
  assign n4617 = \b[5]  & n3400 ;
  assign n4618 = \a[23]  & \b[4]  ;
  assign n4619 = n3731 & n4618 ;
  assign n4620 = ~\a[24]  & \b[4]  ;
  assign n4621 = n3394 & n4620 ;
  assign n4622 = ~n4619 & ~n4621 ;
  assign n4623 = ~n4617 & n4622 ;
  assign n4624 = ~n4616 & n4623 ;
  assign n4625 = ~\a[26]  & n4624 ;
  assign n4626 = ~n4614 & n4625 ;
  assign n4627 = \a[26]  & ~n4624 ;
  assign n4628 = \a[26]  & ~n273 ;
  assign n4629 = ~n4613 & n4628 ;
  assign n4630 = ~n4627 & ~n4629 ;
  assign n4631 = ~n4626 & n4630 ;
  assign n4632 = \a[29]  & ~n3957 ;
  assign n4633 = n4243 & n4632 ;
  assign n4634 = n4251 & n4633 ;
  assign n4635 = \a[29]  & ~n4634 ;
  assign n4636 = \b[2]  & n4247 ;
  assign n4637 = ~\a[27]  & \b[1]  ;
  assign n4638 = n4241 & n4637 ;
  assign n4639 = \a[27]  & \b[1]  ;
  assign n4640 = n4238 & n4639 ;
  assign n4641 = ~n4638 & ~n4640 ;
  assign n4642 = ~n4636 & n4641 ;
  assign n4643 = n157 & n4249 ;
  assign n4644 = n3956 & ~n4246 ;
  assign n4645 = \a[27]  & ~\a[28]  ;
  assign n4646 = ~\a[27]  & \a[28]  ;
  assign n4647 = ~n4645 & ~n4646 ;
  assign n4648 = \b[0]  & n4647 ;
  assign n4649 = n4644 & n4648 ;
  assign n4650 = ~n4643 & ~n4649 ;
  assign n4651 = n4642 & n4650 ;
  assign n4652 = ~n4635 & ~n4651 ;
  assign n4653 = n4635 & n4651 ;
  assign n4654 = ~n4652 & ~n4653 ;
  assign n4655 = n4631 & ~n4654 ;
  assign n4656 = ~n4631 & n4654 ;
  assign n4657 = ~n4655 & ~n4656 ;
  assign n4658 = ~n4609 & n4657 ;
  assign n4659 = ~n4257 & ~n4657 ;
  assign n4660 = ~n4260 & n4659 ;
  assign n4661 = ~n4658 & ~n4660 ;
  assign n4662 = n4608 & ~n4661 ;
  assign n4663 = ~n4608 & ~n4660 ;
  assign n4664 = ~n4658 & n4663 ;
  assign n4665 = ~n4662 & ~n4664 ;
  assign n4666 = n4586 & n4665 ;
  assign n4667 = ~n4586 & ~n4665 ;
  assign n4668 = ~n4666 & ~n4667 ;
  assign n4669 = ~n4583 & ~n4668 ;
  assign n4670 = n4583 & n4668 ;
  assign n4671 = ~n4669 & ~n4670 ;
  assign n4672 = n1087 & n1467 ;
  assign n4673 = ~n1084 & n4672 ;
  assign n4674 = n1467 & n1552 ;
  assign n4675 = ~n1083 & n4674 ;
  assign n4676 = \b[12]  & n1652 ;
  assign n4677 = n1649 & n4676 ;
  assign n4678 = ~\a[15]  & \b[13]  ;
  assign n4679 = n1459 & n4678 ;
  assign n4680 = ~n4677 & ~n4679 ;
  assign n4681 = \b[14]  & n1465 ;
  assign n4682 = \a[15]  & \b[13]  ;
  assign n4683 = n1456 & n4682 ;
  assign n4684 = \a[17]  & ~n4683 ;
  assign n4685 = ~n4681 & n4684 ;
  assign n4686 = n4680 & n4685 ;
  assign n4687 = ~n4675 & n4686 ;
  assign n4688 = ~n4673 & n4687 ;
  assign n4689 = ~n4681 & ~n4683 ;
  assign n4690 = n4680 & n4689 ;
  assign n4691 = ~n4675 & n4690 ;
  assign n4692 = ~n4673 & n4691 ;
  assign n4693 = ~\a[17]  & ~n4692 ;
  assign n4694 = ~n4688 & ~n4693 ;
  assign n4695 = ~n4671 & ~n4694 ;
  assign n4696 = ~n4566 & n4695 ;
  assign n4697 = n4671 & ~n4694 ;
  assign n4698 = n4566 & n4697 ;
  assign n4699 = ~n4696 & ~n4698 ;
  assign n4700 = ~n4671 & n4694 ;
  assign n4701 = n4566 & n4700 ;
  assign n4702 = n4671 & n4694 ;
  assign n4703 = ~n4566 & n4702 ;
  assign n4704 = ~n4701 & ~n4703 ;
  assign n4705 = n4699 & n4704 ;
  assign n4706 = n999 & ~n1694 ;
  assign n4707 = ~n1692 & n4706 ;
  assign n4708 = \b[15]  & n1182 ;
  assign n4709 = n1179 & n4708 ;
  assign n4710 = ~\a[11]  & \b[16]  ;
  assign n4711 = n1181 & n4710 ;
  assign n4712 = ~n4709 & ~n4711 ;
  assign n4713 = \b[17]  & n997 ;
  assign n4714 = \a[12]  & \b[16]  ;
  assign n4715 = n988 & n4714 ;
  assign n4716 = \a[14]  & ~n4715 ;
  assign n4717 = ~n4713 & n4716 ;
  assign n4718 = n4712 & n4717 ;
  assign n4719 = ~n4707 & n4718 ;
  assign n4720 = ~n4713 & ~n4715 ;
  assign n4721 = n4712 & n4720 ;
  assign n4722 = ~n4707 & n4721 ;
  assign n4723 = ~\a[14]  & ~n4722 ;
  assign n4724 = ~n4719 & ~n4723 ;
  assign n4725 = ~n4705 & ~n4724 ;
  assign n4726 = n4564 & n4725 ;
  assign n4727 = n4705 & ~n4724 ;
  assign n4728 = ~n4564 & n4727 ;
  assign n4729 = ~n4726 & ~n4728 ;
  assign n4730 = ~n4705 & n4724 ;
  assign n4731 = ~n4564 & n4730 ;
  assign n4732 = n4705 & n4724 ;
  assign n4733 = n4564 & n4732 ;
  assign n4734 = ~n4731 & ~n4733 ;
  assign n4735 = n4729 & n4734 ;
  assign n4736 = ~n4561 & n4735 ;
  assign n4737 = ~n4362 & ~n4735 ;
  assign n4738 = ~n4560 & n4737 ;
  assign n4739 = n646 & n2293 ;
  assign n4740 = ~n2290 & n4739 ;
  assign n4741 = n646 & ~n2293 ;
  assign n4742 = ~n2074 & n4741 ;
  assign n4743 = ~n2289 & n4742 ;
  assign n4744 = \b[18]  & n796 ;
  assign n4745 = n793 & n4744 ;
  assign n4746 = ~\a[9]  & \b[19]  ;
  assign n4747 = n638 & n4746 ;
  assign n4748 = ~n4745 & ~n4747 ;
  assign n4749 = \b[20]  & n644 ;
  assign n4750 = \a[9]  & \b[19]  ;
  assign n4751 = n635 & n4750 ;
  assign n4752 = \a[11]  & ~n4751 ;
  assign n4753 = ~n4749 & n4752 ;
  assign n4754 = n4748 & n4753 ;
  assign n4755 = ~n4743 & n4754 ;
  assign n4756 = ~n4740 & n4755 ;
  assign n4757 = ~n4749 & ~n4751 ;
  assign n4758 = n4748 & n4757 ;
  assign n4759 = ~n4743 & n4758 ;
  assign n4760 = ~n4740 & n4759 ;
  assign n4761 = ~\a[11]  & ~n4760 ;
  assign n4762 = ~n4756 & ~n4761 ;
  assign n4763 = ~n4738 & ~n4762 ;
  assign n4764 = ~n4736 & n4763 ;
  assign n4765 = ~n4735 & n4762 ;
  assign n4766 = n4561 & n4765 ;
  assign n4767 = n4735 & n4762 ;
  assign n4768 = ~n4561 & n4767 ;
  assign n4769 = ~n4766 & ~n4768 ;
  assign n4770 = ~n4764 & n4769 ;
  assign n4771 = ~n4559 & n4770 ;
  assign n4772 = n4559 & ~n4770 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4774 = ~n4554 & n4773 ;
  assign n4775 = n4554 & ~n4773 ;
  assign n4776 = ~n4774 & ~n4775 ;
  assign n4777 = ~n4537 & ~n4776 ;
  assign n4778 = ~n4517 & n4777 ;
  assign n4779 = ~n4537 & n4776 ;
  assign n4780 = n4517 & n4779 ;
  assign n4781 = ~n4778 & ~n4780 ;
  assign n4782 = n4537 & ~n4776 ;
  assign n4783 = n4517 & n4782 ;
  assign n4784 = n4537 & n4776 ;
  assign n4785 = ~n4517 & n4784 ;
  assign n4786 = ~n4783 & ~n4785 ;
  assign n4787 = n4781 & n4786 ;
  assign n4788 = ~n4516 & ~n4787 ;
  assign n4789 = n4493 & n4788 ;
  assign n4790 = ~n4516 & n4787 ;
  assign n4791 = ~n4493 & n4790 ;
  assign n4792 = ~n4789 & ~n4791 ;
  assign n4793 = n4516 & ~n4787 ;
  assign n4794 = ~n4493 & n4793 ;
  assign n4795 = n4516 & n4787 ;
  assign n4796 = n4493 & n4795 ;
  assign n4797 = ~n4794 & ~n4796 ;
  assign n4798 = n4792 & n4797 ;
  assign n4799 = ~n4490 & n4798 ;
  assign n4800 = n4485 & ~n4798 ;
  assign n4801 = ~n4487 & n4800 ;
  assign n4802 = ~n4799 & ~n4801 ;
  assign n4803 = n4485 & n4792 ;
  assign n4804 = ~n4487 & n4803 ;
  assign n4805 = n4797 & ~n4804 ;
  assign n4806 = n4493 & n4787 ;
  assign n4807 = n4781 & ~n4806 ;
  assign n4808 = ~n4423 & ~n4774 ;
  assign n4809 = ~n4428 & n4808 ;
  assign n4810 = ~n4775 & ~n4809 ;
  assign n4811 = ~n4764 & ~n4771 ;
  assign n4812 = n430 & n3283 ;
  assign n4813 = ~n3280 & n4812 ;
  assign n4814 = n430 & n4107 ;
  assign n4815 = ~n3279 & n4814 ;
  assign n4816 = \b[22]  & n486 ;
  assign n4817 = n483 & n4816 ;
  assign n4818 = \b[24]  & n428 ;
  assign n4819 = \a[6]  & \b[23]  ;
  assign n4820 = n419 & n4819 ;
  assign n4821 = ~\a[6]  & \b[23]  ;
  assign n4822 = n422 & n4821 ;
  assign n4823 = ~n4820 & ~n4822 ;
  assign n4824 = ~n4818 & n4823 ;
  assign n4825 = ~n4817 & n4824 ;
  assign n4826 = ~n4815 & n4825 ;
  assign n4827 = ~n4813 & n4826 ;
  assign n4828 = ~\a[8]  & ~n4827 ;
  assign n4829 = \a[8]  & n4825 ;
  assign n4830 = ~n4815 & n4829 ;
  assign n4831 = ~n4813 & n4830 ;
  assign n4832 = ~n4828 & ~n4831 ;
  assign n4833 = ~n4362 & n4729 ;
  assign n4834 = ~n4560 & n4833 ;
  assign n4835 = n4734 & ~n4834 ;
  assign n4836 = n4564 & n4705 ;
  assign n4837 = n4699 & ~n4836 ;
  assign n4838 = n4292 & ~n4670 ;
  assign n4839 = ~n4565 & n4838 ;
  assign n4840 = ~n4669 & ~n4839 ;
  assign n4841 = ~n4664 & ~n4666 ;
  assign n4842 = ~n909 & ~n1805 ;
  assign n4843 = ~n1962 & n4842 ;
  assign n4844 = n906 & n4843 ;
  assign n4845 = n909 & ~n1805 ;
  assign n4846 = ~n1962 & n4845 ;
  assign n4847 = ~n906 & n4846 ;
  assign n4848 = ~n4844 & ~n4847 ;
  assign n4849 = \b[10]  & n2218 ;
  assign n4850 = n2216 & n4849 ;
  assign n4851 = ~\a[18]  & \b[11]  ;
  assign n4852 = n1957 & n4851 ;
  assign n4853 = ~n4850 & ~n4852 ;
  assign n4854 = \b[12]  & n1963 ;
  assign n4855 = \a[18]  & \b[11]  ;
  assign n4856 = n2210 & n4855 ;
  assign n4857 = \a[20]  & ~n4856 ;
  assign n4858 = ~n4854 & n4857 ;
  assign n4859 = n4853 & n4858 ;
  assign n4860 = n4848 & n4859 ;
  assign n4861 = ~n4854 & ~n4856 ;
  assign n4862 = n4853 & n4861 ;
  assign n4863 = n4848 & n4862 ;
  assign n4864 = ~\a[20]  & ~n4863 ;
  assign n4865 = ~n4860 & ~n4864 ;
  assign n4866 = ~n4257 & ~n4655 ;
  assign n4867 = ~n4260 & n4866 ;
  assign n4868 = ~n4656 & ~n4867 ;
  assign n4869 = ~n586 & n2622 ;
  assign n4870 = ~n504 & n2622 ;
  assign n4871 = ~n508 & n4870 ;
  assign n4872 = ~n4869 & ~n4871 ;
  assign n4873 = ~n589 & ~n4872 ;
  assign n4874 = \b[7]  & n2912 ;
  assign n4875 = n2909 & n4874 ;
  assign n4876 = \b[9]  & n2620 ;
  assign n4877 = \a[20]  & \b[8]  ;
  assign n4878 = n2910 & n4877 ;
  assign n4879 = ~\a[21]  & \b[8]  ;
  assign n4880 = n2614 & n4879 ;
  assign n4881 = ~n4878 & ~n4880 ;
  assign n4882 = ~n4876 & n4881 ;
  assign n4883 = ~n4875 & n4882 ;
  assign n4884 = ~\a[23]  & n4883 ;
  assign n4885 = ~n4873 & n4884 ;
  assign n4886 = \a[23]  & ~n4883 ;
  assign n4887 = \a[23]  & ~n589 ;
  assign n4888 = ~n4872 & n4887 ;
  assign n4889 = ~n4886 & ~n4888 ;
  assign n4890 = ~n4885 & n4889 ;
  assign n4891 = n177 & n4249 ;
  assign n4892 = \b[3]  & n4247 ;
  assign n4893 = \a[26]  & \b[2]  ;
  assign n4894 = n4645 & n4893 ;
  assign n4895 = ~\a[27]  & \b[2]  ;
  assign n4896 = n4241 & n4895 ;
  assign n4897 = ~n4894 & ~n4896 ;
  assign n4898 = ~n4892 & n4897 ;
  assign n4899 = ~n4891 & n4898 ;
  assign n4900 = \b[1]  & n4647 ;
  assign n4901 = n4644 & n4900 ;
  assign n4902 = ~\a[29]  & ~n4901 ;
  assign n4903 = n4899 & n4902 ;
  assign n4904 = n4899 & ~n4901 ;
  assign n4905 = \a[29]  & ~n4904 ;
  assign n4906 = ~n4903 & ~n4905 ;
  assign n4907 = \a[29]  & ~\a[30]  ;
  assign n4908 = ~\a[29]  & \a[30]  ;
  assign n4909 = ~n4907 & ~n4908 ;
  assign n4910 = \b[0]  & ~n4909 ;
  assign n4911 = n4634 & n4651 ;
  assign n4912 = n4910 & n4911 ;
  assign n4913 = ~n4910 & ~n4911 ;
  assign n4914 = ~n4912 & ~n4913 ;
  assign n4915 = n4906 & n4914 ;
  assign n4916 = ~n4906 & ~n4914 ;
  assign n4917 = ~n4915 & ~n4916 ;
  assign n4918 = ~n323 & ~n3154 ;
  assign n4919 = ~n3399 & n4918 ;
  assign n4920 = n320 & n4919 ;
  assign n4921 = n323 & ~n3154 ;
  assign n4922 = ~n3399 & n4921 ;
  assign n4923 = ~n320 & n4922 ;
  assign n4924 = ~n4920 & ~n4923 ;
  assign n4925 = \b[4]  & n3733 ;
  assign n4926 = n3730 & n4925 ;
  assign n4927 = \b[6]  & n3400 ;
  assign n4928 = \a[23]  & \b[5]  ;
  assign n4929 = n3731 & n4928 ;
  assign n4930 = ~\a[24]  & \b[5]  ;
  assign n4931 = n3394 & n4930 ;
  assign n4932 = ~n4929 & ~n4931 ;
  assign n4933 = ~n4927 & n4932 ;
  assign n4934 = ~n4926 & n4933 ;
  assign n4935 = n4924 & n4934 ;
  assign n4936 = ~\a[26]  & ~n4935 ;
  assign n4937 = \a[26]  & n4934 ;
  assign n4938 = n4924 & n4937 ;
  assign n4939 = ~n4936 & ~n4938 ;
  assign n4940 = n4917 & ~n4939 ;
  assign n4941 = ~n4917 & n4939 ;
  assign n4942 = ~n4940 & ~n4941 ;
  assign n4943 = n4890 & ~n4942 ;
  assign n4944 = n4868 & n4943 ;
  assign n4945 = n4890 & n4942 ;
  assign n4946 = ~n4868 & n4945 ;
  assign n4947 = ~n4944 & ~n4946 ;
  assign n4948 = ~n4890 & ~n4942 ;
  assign n4949 = ~n4868 & n4948 ;
  assign n4950 = ~n4890 & n4942 ;
  assign n4951 = n4868 & n4950 ;
  assign n4952 = ~n4949 & ~n4951 ;
  assign n4953 = n4947 & n4952 ;
  assign n4954 = n4865 & ~n4953 ;
  assign n4955 = n4841 & n4954 ;
  assign n4956 = n4865 & n4953 ;
  assign n4957 = ~n4841 & n4956 ;
  assign n4958 = ~n4955 & ~n4957 ;
  assign n4959 = ~n4841 & n4953 ;
  assign n4960 = ~n4664 & ~n4953 ;
  assign n4961 = ~n4666 & n4960 ;
  assign n4962 = ~n4865 & ~n4961 ;
  assign n4963 = ~n4959 & n4962 ;
  assign n4964 = n4958 & ~n4963 ;
  assign n4965 = ~n1233 & n1467 ;
  assign n4966 = ~n1231 & n4965 ;
  assign n4967 = \b[13]  & n1652 ;
  assign n4968 = n1649 & n4967 ;
  assign n4969 = ~\a[15]  & \b[14]  ;
  assign n4970 = n1459 & n4969 ;
  assign n4971 = ~n4968 & ~n4970 ;
  assign n4972 = \b[15]  & n1465 ;
  assign n4973 = \a[15]  & \b[14]  ;
  assign n4974 = n1456 & n4973 ;
  assign n4975 = \a[17]  & ~n4974 ;
  assign n4976 = ~n4972 & n4975 ;
  assign n4977 = n4971 & n4976 ;
  assign n4978 = ~n4966 & n4977 ;
  assign n4979 = ~n4972 & ~n4974 ;
  assign n4980 = n4971 & n4979 ;
  assign n4981 = ~n4966 & n4980 ;
  assign n4982 = ~\a[17]  & ~n4981 ;
  assign n4983 = ~n4978 & ~n4982 ;
  assign n4984 = ~n4964 & ~n4983 ;
  assign n4985 = n4840 & n4984 ;
  assign n4986 = n4964 & ~n4983 ;
  assign n4987 = ~n4840 & n4986 ;
  assign n4988 = ~n4985 & ~n4987 ;
  assign n4989 = ~n4964 & n4983 ;
  assign n4990 = ~n4840 & n4989 ;
  assign n4991 = n4964 & n4983 ;
  assign n4992 = n4840 & n4991 ;
  assign n4993 = ~n4990 & ~n4992 ;
  assign n4994 = n4988 & n4993 ;
  assign n4995 = ~n4837 & n4994 ;
  assign n4996 = n4699 & ~n4994 ;
  assign n4997 = ~n4836 & n4996 ;
  assign n4998 = n999 & n1875 ;
  assign n4999 = ~n1872 & n4998 ;
  assign n5000 = ~n1689 & ~n1875 ;
  assign n5001 = n999 & n5000 ;
  assign n5002 = ~n1871 & n5001 ;
  assign n5003 = \b[16]  & n1182 ;
  assign n5004 = n1179 & n5003 ;
  assign n5005 = ~\a[11]  & \b[17]  ;
  assign n5006 = n1181 & n5005 ;
  assign n5007 = ~n5004 & ~n5006 ;
  assign n5008 = \b[18]  & n997 ;
  assign n5009 = \a[12]  & \b[17]  ;
  assign n5010 = n988 & n5009 ;
  assign n5011 = \a[14]  & ~n5010 ;
  assign n5012 = ~n5008 & n5011 ;
  assign n5013 = n5007 & n5012 ;
  assign n5014 = ~n5002 & n5013 ;
  assign n5015 = ~n4999 & n5014 ;
  assign n5016 = ~n5008 & ~n5010 ;
  assign n5017 = n5007 & n5016 ;
  assign n5018 = ~n5002 & n5017 ;
  assign n5019 = ~n4999 & n5018 ;
  assign n5020 = ~\a[14]  & ~n5019 ;
  assign n5021 = ~n5015 & ~n5020 ;
  assign n5022 = ~n4997 & ~n5021 ;
  assign n5023 = ~n4995 & n5022 ;
  assign n5024 = ~n4994 & n5021 ;
  assign n5025 = n4837 & n5024 ;
  assign n5026 = n4994 & n5021 ;
  assign n5027 = ~n4837 & n5026 ;
  assign n5028 = ~n5025 & ~n5027 ;
  assign n5029 = ~n5023 & n5028 ;
  assign n5030 = n646 & ~n2523 ;
  assign n5031 = ~n2521 & n5030 ;
  assign n5032 = \b[21]  & n644 ;
  assign n5033 = \a[9]  & \b[20]  ;
  assign n5034 = n635 & n5033 ;
  assign n5035 = ~n5032 & ~n5034 ;
  assign n5036 = \b[19]  & n796 ;
  assign n5037 = n793 & n5036 ;
  assign n5038 = ~\a[9]  & \b[20]  ;
  assign n5039 = n638 & n5038 ;
  assign n5040 = ~n5037 & ~n5039 ;
  assign n5041 = n5035 & n5040 ;
  assign n5042 = ~n5031 & n5041 ;
  assign n5043 = ~\a[11]  & ~n5042 ;
  assign n5044 = \a[11]  & n5041 ;
  assign n5045 = ~n5031 & n5044 ;
  assign n5046 = ~n5043 & ~n5045 ;
  assign n5047 = ~n5029 & ~n5046 ;
  assign n5048 = n4835 & n5047 ;
  assign n5049 = n5029 & ~n5046 ;
  assign n5050 = ~n4835 & n5049 ;
  assign n5051 = ~n5048 & ~n5050 ;
  assign n5052 = ~n5029 & n5046 ;
  assign n5053 = ~n4835 & n5052 ;
  assign n5054 = n5029 & n5046 ;
  assign n5055 = n4835 & n5054 ;
  assign n5056 = ~n5053 & ~n5055 ;
  assign n5057 = n5051 & n5056 ;
  assign n5058 = ~n4832 & ~n5057 ;
  assign n5059 = ~n4811 & n5058 ;
  assign n5060 = ~n4832 & n5057 ;
  assign n5061 = n4811 & n5060 ;
  assign n5062 = ~n5059 & ~n5061 ;
  assign n5063 = n4832 & ~n5057 ;
  assign n5064 = n4811 & n5063 ;
  assign n5065 = n4832 & n5057 ;
  assign n5066 = ~n4811 & n5065 ;
  assign n5067 = ~n5064 & ~n5066 ;
  assign n5068 = n5062 & n5067 ;
  assign n5069 = n252 & ~n4148 ;
  assign n5070 = ~n4146 & n5069 ;
  assign n5071 = \b[27]  & n250 ;
  assign n5072 = \a[3]  & \b[26]  ;
  assign n5073 = n241 & n5072 ;
  assign n5074 = ~n5071 & ~n5073 ;
  assign n5075 = \b[25]  & n303 ;
  assign n5076 = n300 & n5075 ;
  assign n5077 = ~\a[3]  & \b[26]  ;
  assign n5078 = n244 & n5077 ;
  assign n5079 = ~n5076 & ~n5078 ;
  assign n5080 = n5074 & n5079 ;
  assign n5081 = ~n5070 & n5080 ;
  assign n5082 = ~\a[5]  & ~n5081 ;
  assign n5083 = \a[5]  & n5080 ;
  assign n5084 = ~n5070 & n5083 ;
  assign n5085 = ~n5082 & ~n5084 ;
  assign n5086 = ~n5068 & ~n5085 ;
  assign n5087 = n4810 & n5086 ;
  assign n5088 = n5068 & ~n5085 ;
  assign n5089 = ~n4810 & n5088 ;
  assign n5090 = ~n5087 & ~n5089 ;
  assign n5091 = ~n5068 & n5085 ;
  assign n5092 = ~n4810 & n5091 ;
  assign n5093 = n5068 & n5085 ;
  assign n5094 = n4810 & n5093 ;
  assign n5095 = ~n5092 & ~n5094 ;
  assign n5096 = n5090 & n5095 ;
  assign n5097 = ~n4807 & n5096 ;
  assign n5098 = n4781 & ~n5096 ;
  assign n5099 = ~n4806 & n5098 ;
  assign n5100 = ~n4455 & ~n4498 ;
  assign n5101 = ~n4495 & n5100 ;
  assign n5102 = ~n4497 & ~n5101 ;
  assign n5103 = ~\b[29]  & ~\b[30]  ;
  assign n5104 = \b[29]  & \b[30]  ;
  assign n5105 = ~n5103 & ~n5104 ;
  assign n5106 = n134 & n5105 ;
  assign n5107 = ~n5102 & n5106 ;
  assign n5108 = n134 & ~n5105 ;
  assign n5109 = ~n4497 & n5108 ;
  assign n5110 = ~n5101 & n5109 ;
  assign n5111 = \a[0]  & \b[30]  ;
  assign n5112 = n133 & n5111 ;
  assign n5113 = \b[29]  & n141 ;
  assign n5114 = ~\a[1]  & \b[28]  ;
  assign n5115 = n1521 & n5114 ;
  assign n5116 = ~n5113 & ~n5115 ;
  assign n5117 = ~n5112 & n5116 ;
  assign n5118 = \a[2]  & n5117 ;
  assign n5119 = ~n5110 & n5118 ;
  assign n5120 = ~n5107 & n5119 ;
  assign n5121 = ~n5110 & n5117 ;
  assign n5122 = ~n5107 & n5121 ;
  assign n5123 = ~\a[2]  & ~n5122 ;
  assign n5124 = ~n5120 & ~n5123 ;
  assign n5125 = ~n5099 & ~n5124 ;
  assign n5126 = ~n5097 & n5125 ;
  assign n5127 = ~n5096 & n5124 ;
  assign n5128 = n4807 & n5127 ;
  assign n5129 = n5096 & n5124 ;
  assign n5130 = ~n4807 & n5129 ;
  assign n5131 = ~n5128 & ~n5130 ;
  assign n5132 = ~n5126 & n5131 ;
  assign n5133 = n4805 & n5132 ;
  assign n5134 = ~n4805 & ~n5132 ;
  assign n5135 = ~n5133 & ~n5134 ;
  assign n5136 = ~n5126 & ~n5133 ;
  assign n5137 = n4781 & n5090 ;
  assign n5138 = ~n4806 & n5137 ;
  assign n5139 = n5095 & ~n5138 ;
  assign n5140 = n4810 & n5068 ;
  assign n5141 = n5062 & ~n5140 ;
  assign n5142 = ~n4764 & n5051 ;
  assign n5143 = ~n4771 & n5142 ;
  assign n5144 = n5056 & ~n5143 ;
  assign n5145 = n4835 & n5029 ;
  assign n5146 = ~n5023 & ~n5145 ;
  assign n5147 = n4699 & n4988 ;
  assign n5148 = ~n4836 & n5147 ;
  assign n5149 = n4993 & ~n5148 ;
  assign n5150 = n4840 & n4964 ;
  assign n5151 = ~n4963 & ~n5150 ;
  assign n5152 = ~n4664 & n4947 ;
  assign n5153 = ~n4666 & n5152 ;
  assign n5154 = n4952 & ~n5153 ;
  assign n5155 = n4868 & n4942 ;
  assign n5156 = ~n4940 & ~n5155 ;
  assign n5157 = ~n380 & n3402 ;
  assign n5158 = ~n322 & n3402 ;
  assign n5159 = ~n326 & n5158 ;
  assign n5160 = ~n5157 & ~n5159 ;
  assign n5161 = ~n383 & ~n5160 ;
  assign n5162 = \b[5]  & n3733 ;
  assign n5163 = n3730 & n5162 ;
  assign n5164 = \b[7]  & n3400 ;
  assign n5165 = \a[23]  & \b[6]  ;
  assign n5166 = n3731 & n5165 ;
  assign n5167 = ~\a[24]  & \b[6]  ;
  assign n5168 = n3394 & n5167 ;
  assign n5169 = ~n5166 & ~n5168 ;
  assign n5170 = ~n5164 & n5169 ;
  assign n5171 = ~n5163 & n5170 ;
  assign n5172 = ~\a[26]  & n5171 ;
  assign n5173 = ~n5161 & n5172 ;
  assign n5174 = \a[26]  & ~n5171 ;
  assign n5175 = \a[26]  & ~n383 ;
  assign n5176 = ~n5160 & n5175 ;
  assign n5177 = ~n5174 & ~n5176 ;
  assign n5178 = ~n5173 & n5177 ;
  assign n5179 = ~n4912 & ~n4915 ;
  assign n5180 = n222 & n4249 ;
  assign n5181 = \b[4]  & n4247 ;
  assign n5182 = \a[26]  & \b[3]  ;
  assign n5183 = n4645 & n5182 ;
  assign n5184 = ~\a[27]  & \b[3]  ;
  assign n5185 = n4241 & n5184 ;
  assign n5186 = ~n5183 & ~n5185 ;
  assign n5187 = ~n5181 & n5186 ;
  assign n5188 = \b[2]  & n4647 ;
  assign n5189 = n4644 & n5188 ;
  assign n5190 = \a[29]  & ~n5189 ;
  assign n5191 = n5187 & n5190 ;
  assign n5192 = ~n5180 & n5191 ;
  assign n5193 = n5187 & ~n5189 ;
  assign n5194 = ~n5180 & n5193 ;
  assign n5195 = ~\a[29]  & ~n5194 ;
  assign n5196 = ~n5192 & ~n5195 ;
  assign n5197 = \a[32]  & \b[0]  ;
  assign n5198 = ~n4909 & n5197 ;
  assign n5199 = \a[30]  & \b[0]  ;
  assign n5200 = \a[29]  & ~\a[31]  ;
  assign n5201 = n5199 & n5200 ;
  assign n5202 = ~\a[30]  & \b[0]  ;
  assign n5203 = ~\a[29]  & \a[31]  ;
  assign n5204 = n5202 & n5203 ;
  assign n5205 = ~n5201 & ~n5204 ;
  assign n5206 = \a[31]  & ~\a[32]  ;
  assign n5207 = ~\a[31]  & \a[32]  ;
  assign n5208 = ~n5206 & ~n5207 ;
  assign n5209 = ~n4909 & n5208 ;
  assign n5210 = \b[1]  & n5209 ;
  assign n5211 = ~n4909 & ~n5208 ;
  assign n5212 = ~n137 & n5211 ;
  assign n5213 = ~n5210 & ~n5212 ;
  assign n5214 = n5205 & n5213 ;
  assign n5215 = n5198 & ~n5214 ;
  assign n5216 = ~n5198 & n5205 ;
  assign n5217 = n5213 & n5216 ;
  assign n5218 = ~n5215 & ~n5217 ;
  assign n5219 = ~n5196 & n5218 ;
  assign n5220 = n5196 & ~n5218 ;
  assign n5221 = ~n5219 & ~n5220 ;
  assign n5222 = ~n5179 & n5221 ;
  assign n5223 = n5179 & ~n5221 ;
  assign n5224 = ~n5222 & ~n5223 ;
  assign n5225 = n5178 & n5224 ;
  assign n5226 = ~n5178 & ~n5224 ;
  assign n5227 = ~n5225 & ~n5226 ;
  assign n5228 = ~n685 & ~n2413 ;
  assign n5229 = ~n2619 & n5228 ;
  assign n5230 = n682 & n5229 ;
  assign n5231 = n685 & ~n2413 ;
  assign n5232 = ~n2619 & n5231 ;
  assign n5233 = ~n682 & n5232 ;
  assign n5234 = ~n5230 & ~n5233 ;
  assign n5235 = \b[8]  & n2912 ;
  assign n5236 = n2909 & n5235 ;
  assign n5237 = \b[10]  & n2620 ;
  assign n5238 = \a[20]  & \b[9]  ;
  assign n5239 = n2910 & n5238 ;
  assign n5240 = ~\a[21]  & \b[9]  ;
  assign n5241 = n2614 & n5240 ;
  assign n5242 = ~n5239 & ~n5241 ;
  assign n5243 = ~n5237 & n5242 ;
  assign n5244 = ~n5236 & n5243 ;
  assign n5245 = n5234 & n5244 ;
  assign n5246 = ~\a[23]  & ~n5245 ;
  assign n5247 = \a[23]  & n5244 ;
  assign n5248 = n5234 & n5247 ;
  assign n5249 = ~n5246 & ~n5248 ;
  assign n5250 = ~n5227 & ~n5249 ;
  assign n5251 = ~n5156 & n5250 ;
  assign n5252 = n5227 & ~n5249 ;
  assign n5253 = n5156 & n5252 ;
  assign n5254 = ~n5251 & ~n5253 ;
  assign n5255 = ~n5227 & n5249 ;
  assign n5256 = n5156 & n5255 ;
  assign n5257 = n5227 & n5249 ;
  assign n5258 = ~n5156 & n5257 ;
  assign n5259 = ~n5256 & ~n5258 ;
  assign n5260 = n5254 & n5259 ;
  assign n5261 = ~n948 & n1965 ;
  assign n5262 = ~n908 & n1965 ;
  assign n5263 = ~n912 & n5262 ;
  assign n5264 = ~n5261 & ~n5263 ;
  assign n5265 = ~n951 & ~n5264 ;
  assign n5266 = \b[11]  & n2218 ;
  assign n5267 = n2216 & n5266 ;
  assign n5268 = ~\a[18]  & \b[12]  ;
  assign n5269 = n1957 & n5268 ;
  assign n5270 = ~n5267 & ~n5269 ;
  assign n5271 = \b[13]  & n1963 ;
  assign n5272 = \a[18]  & \b[12]  ;
  assign n5273 = n2210 & n5272 ;
  assign n5274 = \a[20]  & ~n5273 ;
  assign n5275 = ~n5271 & n5274 ;
  assign n5276 = n5270 & n5275 ;
  assign n5277 = ~n5265 & n5276 ;
  assign n5278 = ~n5271 & ~n5273 ;
  assign n5279 = n5270 & n5278 ;
  assign n5280 = ~\a[20]  & ~n5279 ;
  assign n5281 = ~\a[20]  & ~n951 ;
  assign n5282 = ~n5264 & n5281 ;
  assign n5283 = ~n5280 & ~n5282 ;
  assign n5284 = ~n5277 & n5283 ;
  assign n5285 = ~n5260 & n5284 ;
  assign n5286 = ~n5154 & n5285 ;
  assign n5287 = n5260 & n5284 ;
  assign n5288 = n5154 & n5287 ;
  assign n5289 = ~n5286 & ~n5288 ;
  assign n5290 = ~n5260 & ~n5284 ;
  assign n5291 = n5154 & n5290 ;
  assign n5292 = n5260 & ~n5284 ;
  assign n5293 = ~n5154 & n5292 ;
  assign n5294 = ~n5291 & ~n5293 ;
  assign n5295 = n5289 & n5294 ;
  assign n5296 = ~n1304 & ~n1512 ;
  assign n5297 = ~n1464 & n5296 ;
  assign n5298 = n1509 & n5297 ;
  assign n5299 = ~n1304 & n1512 ;
  assign n5300 = ~n1464 & n5299 ;
  assign n5301 = ~n1509 & n5300 ;
  assign n5302 = ~n5298 & ~n5301 ;
  assign n5303 = \b[14]  & n1652 ;
  assign n5304 = n1649 & n5303 ;
  assign n5305 = ~\a[15]  & \b[15]  ;
  assign n5306 = n1459 & n5305 ;
  assign n5307 = ~n5304 & ~n5306 ;
  assign n5308 = \b[16]  & n1465 ;
  assign n5309 = \a[15]  & \b[15]  ;
  assign n5310 = n1456 & n5309 ;
  assign n5311 = \a[17]  & ~n5310 ;
  assign n5312 = ~n5308 & n5311 ;
  assign n5313 = n5307 & n5312 ;
  assign n5314 = n5302 & n5313 ;
  assign n5315 = ~n5308 & ~n5310 ;
  assign n5316 = n5307 & n5315 ;
  assign n5317 = n5302 & n5316 ;
  assign n5318 = ~\a[17]  & ~n5317 ;
  assign n5319 = ~n5314 & ~n5318 ;
  assign n5320 = ~n5295 & ~n5319 ;
  assign n5321 = ~n5151 & n5320 ;
  assign n5322 = n5295 & ~n5319 ;
  assign n5323 = n5151 & n5322 ;
  assign n5324 = ~n5321 & ~n5323 ;
  assign n5325 = ~n5151 & ~n5295 ;
  assign n5326 = ~n4963 & n5295 ;
  assign n5327 = ~n5150 & n5326 ;
  assign n5328 = n5319 & ~n5327 ;
  assign n5329 = ~n5325 & n5328 ;
  assign n5330 = n5324 & ~n5329 ;
  assign n5331 = n999 & ~n2079 ;
  assign n5332 = ~n2077 & n5331 ;
  assign n5333 = \b[17]  & n1182 ;
  assign n5334 = n1179 & n5333 ;
  assign n5335 = ~\a[11]  & \b[18]  ;
  assign n5336 = n1181 & n5335 ;
  assign n5337 = ~n5334 & ~n5336 ;
  assign n5338 = \b[19]  & n997 ;
  assign n5339 = \a[12]  & \b[18]  ;
  assign n5340 = n988 & n5339 ;
  assign n5341 = \a[14]  & ~n5340 ;
  assign n5342 = ~n5338 & n5341 ;
  assign n5343 = n5337 & n5342 ;
  assign n5344 = ~n5332 & n5343 ;
  assign n5345 = ~n5338 & ~n5340 ;
  assign n5346 = n5337 & n5345 ;
  assign n5347 = ~n5332 & n5346 ;
  assign n5348 = ~\a[14]  & ~n5347 ;
  assign n5349 = ~n5344 & ~n5348 ;
  assign n5350 = ~n5330 & ~n5349 ;
  assign n5351 = n5149 & n5350 ;
  assign n5352 = n5330 & ~n5349 ;
  assign n5353 = ~n5149 & n5352 ;
  assign n5354 = ~n5351 & ~n5353 ;
  assign n5355 = ~n5330 & n5349 ;
  assign n5356 = ~n5149 & n5355 ;
  assign n5357 = n5330 & n5349 ;
  assign n5358 = n5149 & n5357 ;
  assign n5359 = ~n5356 & ~n5358 ;
  assign n5360 = n5354 & n5359 ;
  assign n5361 = ~n5146 & n5360 ;
  assign n5362 = ~n5023 & ~n5360 ;
  assign n5363 = ~n5145 & n5362 ;
  assign n5364 = n646 & n2768 ;
  assign n5365 = ~n2765 & n5364 ;
  assign n5366 = n646 & ~n2768 ;
  assign n5367 = ~n2518 & n5366 ;
  assign n5368 = ~n2764 & n5367 ;
  assign n5369 = \b[20]  & n796 ;
  assign n5370 = n793 & n5369 ;
  assign n5371 = ~\a[9]  & \b[21]  ;
  assign n5372 = n638 & n5371 ;
  assign n5373 = ~n5370 & ~n5372 ;
  assign n5374 = \b[22]  & n644 ;
  assign n5375 = \a[9]  & \b[21]  ;
  assign n5376 = n635 & n5375 ;
  assign n5377 = \a[11]  & ~n5376 ;
  assign n5378 = ~n5374 & n5377 ;
  assign n5379 = n5373 & n5378 ;
  assign n5380 = ~n5368 & n5379 ;
  assign n5381 = ~n5365 & n5380 ;
  assign n5382 = ~n5374 & ~n5376 ;
  assign n5383 = n5373 & n5382 ;
  assign n5384 = ~n5368 & n5383 ;
  assign n5385 = ~n5365 & n5384 ;
  assign n5386 = ~\a[11]  & ~n5385 ;
  assign n5387 = ~n5381 & ~n5386 ;
  assign n5388 = ~n5363 & ~n5387 ;
  assign n5389 = ~n5361 & n5388 ;
  assign n5390 = ~n5360 & n5387 ;
  assign n5391 = n5146 & n5390 ;
  assign n5392 = n5360 & n5387 ;
  assign n5393 = ~n5146 & n5392 ;
  assign n5394 = ~n5391 & ~n5393 ;
  assign n5395 = ~n5389 & n5394 ;
  assign n5396 = ~n5144 & ~n5395 ;
  assign n5397 = n5144 & n5395 ;
  assign n5398 = ~n5396 & ~n5397 ;
  assign n5399 = n430 & ~n3567 ;
  assign n5400 = ~n3565 & n5399 ;
  assign n5401 = \b[25]  & n428 ;
  assign n5402 = \a[6]  & \b[24]  ;
  assign n5403 = n419 & n5402 ;
  assign n5404 = ~n5401 & ~n5403 ;
  assign n5405 = \b[23]  & n486 ;
  assign n5406 = n483 & n5405 ;
  assign n5407 = ~\a[6]  & \b[24]  ;
  assign n5408 = n422 & n5407 ;
  assign n5409 = ~n5406 & ~n5408 ;
  assign n5410 = n5404 & n5409 ;
  assign n5411 = ~n5400 & n5410 ;
  assign n5412 = ~\a[8]  & ~n5411 ;
  assign n5413 = \a[8]  & n5410 ;
  assign n5414 = ~n5400 & n5413 ;
  assign n5415 = ~n5412 & ~n5414 ;
  assign n5416 = n5398 & ~n5415 ;
  assign n5417 = ~n5398 & n5415 ;
  assign n5418 = ~n5416 & ~n5417 ;
  assign n5419 = n252 & n4456 ;
  assign n5420 = ~n4453 & n5419 ;
  assign n5421 = ~n4143 & ~n4456 ;
  assign n5422 = n252 & n5421 ;
  assign n5423 = ~n4452 & n5422 ;
  assign n5424 = \b[26]  & n303 ;
  assign n5425 = n300 & n5424 ;
  assign n5426 = ~\a[3]  & \b[27]  ;
  assign n5427 = n244 & n5426 ;
  assign n5428 = ~n5425 & ~n5427 ;
  assign n5429 = \b[28]  & n250 ;
  assign n5430 = \a[3]  & \b[27]  ;
  assign n5431 = n241 & n5430 ;
  assign n5432 = \a[5]  & ~n5431 ;
  assign n5433 = ~n5429 & n5432 ;
  assign n5434 = n5428 & n5433 ;
  assign n5435 = ~n5423 & n5434 ;
  assign n5436 = ~n5420 & n5435 ;
  assign n5437 = ~n5429 & ~n5431 ;
  assign n5438 = n5428 & n5437 ;
  assign n5439 = ~n5423 & n5438 ;
  assign n5440 = ~n5420 & n5439 ;
  assign n5441 = ~\a[5]  & ~n5440 ;
  assign n5442 = ~n5436 & ~n5441 ;
  assign n5443 = ~n5418 & ~n5442 ;
  assign n5444 = ~n5141 & n5443 ;
  assign n5445 = n5418 & ~n5442 ;
  assign n5446 = n5141 & n5445 ;
  assign n5447 = ~n5444 & ~n5446 ;
  assign n5448 = ~n5418 & n5442 ;
  assign n5449 = n5141 & n5448 ;
  assign n5450 = n5418 & n5442 ;
  assign n5451 = ~n5141 & n5450 ;
  assign n5452 = ~n5449 & ~n5451 ;
  assign n5453 = n5447 & n5452 ;
  assign n5454 = ~n4497 & n5105 ;
  assign n5455 = ~n5101 & n5454 ;
  assign n5456 = ~n5104 & ~n5455 ;
  assign n5457 = ~\b[30]  & ~\b[31]  ;
  assign n5458 = \b[30]  & \b[31]  ;
  assign n5459 = ~n5457 & ~n5458 ;
  assign n5460 = ~n5456 & n5459 ;
  assign n5461 = ~n5104 & ~n5459 ;
  assign n5462 = ~n5455 & n5461 ;
  assign n5463 = n134 & ~n5462 ;
  assign n5464 = ~n5460 & n5463 ;
  assign n5465 = \a[0]  & \b[31]  ;
  assign n5466 = n133 & n5465 ;
  assign n5467 = \b[30]  & n141 ;
  assign n5468 = ~\a[1]  & \b[29]  ;
  assign n5469 = n1521 & n5468 ;
  assign n5470 = ~n5467 & ~n5469 ;
  assign n5471 = ~n5466 & n5470 ;
  assign n5472 = ~n5464 & n5471 ;
  assign n5473 = ~\a[2]  & ~n5472 ;
  assign n5474 = \a[2]  & n5471 ;
  assign n5475 = ~n5464 & n5474 ;
  assign n5476 = ~n5473 & ~n5475 ;
  assign n5477 = ~n5453 & ~n5476 ;
  assign n5478 = n5139 & n5477 ;
  assign n5479 = n5453 & ~n5476 ;
  assign n5480 = ~n5139 & n5479 ;
  assign n5481 = ~n5478 & ~n5480 ;
  assign n5482 = ~n5453 & n5476 ;
  assign n5483 = ~n5139 & n5482 ;
  assign n5484 = n5453 & n5476 ;
  assign n5485 = n5139 & n5484 ;
  assign n5486 = ~n5483 & ~n5485 ;
  assign n5487 = n5481 & n5486 ;
  assign n5488 = ~n5136 & n5487 ;
  assign n5489 = ~n5126 & ~n5487 ;
  assign n5490 = ~n5133 & n5489 ;
  assign n5491 = ~n5488 & ~n5490 ;
  assign n5492 = ~n5126 & n5481 ;
  assign n5493 = ~n5133 & n5492 ;
  assign n5494 = n5486 & ~n5493 ;
  assign n5495 = n5139 & n5453 ;
  assign n5496 = n5447 & ~n5495 ;
  assign n5497 = n5062 & ~n5416 ;
  assign n5498 = ~n5140 & n5497 ;
  assign n5499 = ~n5417 & ~n5498 ;
  assign n5500 = ~n5389 & ~n5397 ;
  assign n5501 = ~n5023 & n5354 ;
  assign n5502 = ~n5145 & n5501 ;
  assign n5503 = n5359 & ~n5502 ;
  assign n5504 = n646 & ~n3022 ;
  assign n5505 = ~n3020 & n5504 ;
  assign n5506 = \b[23]  & n644 ;
  assign n5507 = \a[9]  & \b[22]  ;
  assign n5508 = n635 & n5507 ;
  assign n5509 = ~n5506 & ~n5508 ;
  assign n5510 = \b[21]  & n796 ;
  assign n5511 = n793 & n5510 ;
  assign n5512 = ~\a[9]  & \b[22]  ;
  assign n5513 = n638 & n5512 ;
  assign n5514 = ~n5511 & ~n5513 ;
  assign n5515 = n5509 & n5514 ;
  assign n5516 = ~n5505 & n5515 ;
  assign n5517 = ~\a[11]  & ~n5516 ;
  assign n5518 = \a[11]  & n5515 ;
  assign n5519 = ~n5505 & n5518 ;
  assign n5520 = ~n5517 & ~n5519 ;
  assign n5521 = n5149 & n5330 ;
  assign n5522 = n5324 & ~n5521 ;
  assign n5523 = ~n4963 & n5294 ;
  assign n5524 = ~n5150 & n5523 ;
  assign n5525 = n5289 & ~n5524 ;
  assign n5526 = n5154 & n5260 ;
  assign n5527 = n5254 & ~n5526 ;
  assign n5528 = n1087 & n1965 ;
  assign n5529 = ~n1084 & n5528 ;
  assign n5530 = ~n1087 & n1965 ;
  assign n5531 = ~n946 & n5530 ;
  assign n5532 = ~n1083 & n5531 ;
  assign n5533 = \b[12]  & n2218 ;
  assign n5534 = n2216 & n5533 ;
  assign n5535 = ~\a[18]  & \b[13]  ;
  assign n5536 = n1957 & n5535 ;
  assign n5537 = ~n5534 & ~n5536 ;
  assign n5538 = \b[14]  & n1963 ;
  assign n5539 = \a[18]  & \b[13]  ;
  assign n5540 = n2210 & n5539 ;
  assign n5541 = \a[20]  & ~n5540 ;
  assign n5542 = ~n5538 & n5541 ;
  assign n5543 = n5537 & n5542 ;
  assign n5544 = ~n5532 & n5543 ;
  assign n5545 = ~n5529 & n5544 ;
  assign n5546 = ~n5538 & ~n5540 ;
  assign n5547 = n5537 & n5546 ;
  assign n5548 = ~n5532 & n5547 ;
  assign n5549 = ~n5529 & n5548 ;
  assign n5550 = ~\a[20]  & ~n5549 ;
  assign n5551 = ~n5545 & ~n5550 ;
  assign n5552 = ~n4940 & ~n5225 ;
  assign n5553 = ~n5155 & n5552 ;
  assign n5554 = ~n5226 & ~n5553 ;
  assign n5555 = ~n5219 & ~n5222 ;
  assign n5556 = ~n270 & n4249 ;
  assign n5557 = ~n218 & n4249 ;
  assign n5558 = ~n220 & n5557 ;
  assign n5559 = ~n5556 & ~n5558 ;
  assign n5560 = ~n273 & ~n5559 ;
  assign n5561 = \b[3]  & n4647 ;
  assign n5562 = n4644 & n5561 ;
  assign n5563 = ~\a[26]  & \b[4]  ;
  assign n5564 = n4646 & n5563 ;
  assign n5565 = ~n5562 & ~n5564 ;
  assign n5566 = \b[5]  & n4247 ;
  assign n5567 = \a[27]  & \b[4]  ;
  assign n5568 = n4238 & n5567 ;
  assign n5569 = \a[29]  & ~n5568 ;
  assign n5570 = ~n5566 & n5569 ;
  assign n5571 = n5565 & n5570 ;
  assign n5572 = ~n5560 & n5571 ;
  assign n5573 = ~n5566 & ~n5568 ;
  assign n5574 = n5565 & n5573 ;
  assign n5575 = ~\a[29]  & ~n5574 ;
  assign n5576 = ~\a[29]  & ~n273 ;
  assign n5577 = ~n5559 & n5576 ;
  assign n5578 = ~n5575 & ~n5577 ;
  assign n5579 = ~n5572 & n5578 ;
  assign n5580 = \a[32]  & ~n4910 ;
  assign n5581 = n5205 & n5580 ;
  assign n5582 = n5213 & n5581 ;
  assign n5583 = \a[32]  & ~n5582 ;
  assign n5584 = \b[2]  & n5209 ;
  assign n5585 = ~\a[30]  & \b[1]  ;
  assign n5586 = n5203 & n5585 ;
  assign n5587 = \a[30]  & \b[1]  ;
  assign n5588 = n5200 & n5587 ;
  assign n5589 = ~n5586 & ~n5588 ;
  assign n5590 = ~n5584 & n5589 ;
  assign n5591 = n157 & n5211 ;
  assign n5592 = n4909 & ~n5208 ;
  assign n5593 = \a[30]  & ~\a[31]  ;
  assign n5594 = ~\a[30]  & \a[31]  ;
  assign n5595 = ~n5593 & ~n5594 ;
  assign n5596 = \b[0]  & n5595 ;
  assign n5597 = n5592 & n5596 ;
  assign n5598 = ~n5591 & ~n5597 ;
  assign n5599 = n5590 & n5598 ;
  assign n5600 = ~n5583 & ~n5599 ;
  assign n5601 = n5583 & n5599 ;
  assign n5602 = ~n5600 & ~n5601 ;
  assign n5603 = ~n5579 & ~n5602 ;
  assign n5604 = n5579 & n5602 ;
  assign n5605 = ~n5603 & ~n5604 ;
  assign n5606 = ~n5555 & n5605 ;
  assign n5607 = ~n505 & ~n3154 ;
  assign n5608 = ~n3399 & n5607 ;
  assign n5609 = n502 & n5608 ;
  assign n5610 = n505 & ~n3154 ;
  assign n5611 = ~n3399 & n5610 ;
  assign n5612 = ~n502 & n5611 ;
  assign n5613 = ~n5609 & ~n5612 ;
  assign n5614 = \b[6]  & n3733 ;
  assign n5615 = n3730 & n5614 ;
  assign n5616 = \b[8]  & n3400 ;
  assign n5617 = \a[24]  & \b[7]  ;
  assign n5618 = n3391 & n5617 ;
  assign n5619 = ~\a[24]  & \b[7]  ;
  assign n5620 = n3394 & n5619 ;
  assign n5621 = ~n5618 & ~n5620 ;
  assign n5622 = ~n5616 & n5621 ;
  assign n5623 = ~n5615 & n5622 ;
  assign n5624 = n5613 & n5623 ;
  assign n5625 = ~\a[26]  & ~n5624 ;
  assign n5626 = \a[26]  & n5623 ;
  assign n5627 = n5613 & n5626 ;
  assign n5628 = ~n5625 & ~n5627 ;
  assign n5629 = ~n5219 & ~n5605 ;
  assign n5630 = ~n5222 & n5629 ;
  assign n5631 = ~n5628 & ~n5630 ;
  assign n5632 = ~n5606 & n5631 ;
  assign n5633 = ~n5606 & ~n5630 ;
  assign n5634 = n5628 & ~n5633 ;
  assign n5635 = ~n5632 & ~n5634 ;
  assign n5636 = ~n5554 & ~n5635 ;
  assign n5637 = n5554 & n5635 ;
  assign n5638 = ~n5636 & ~n5637 ;
  assign n5639 = ~n728 & n2622 ;
  assign n5640 = ~n726 & n5639 ;
  assign n5641 = \b[9]  & n2912 ;
  assign n5642 = n2909 & n5641 ;
  assign n5643 = \b[11]  & n2620 ;
  assign n5644 = \a[20]  & \b[10]  ;
  assign n5645 = n2910 & n5644 ;
  assign n5646 = ~\a[21]  & \b[10]  ;
  assign n5647 = n2614 & n5646 ;
  assign n5648 = ~n5645 & ~n5647 ;
  assign n5649 = ~n5643 & n5648 ;
  assign n5650 = ~n5642 & n5649 ;
  assign n5651 = ~\a[23]  & n5650 ;
  assign n5652 = ~n5640 & n5651 ;
  assign n5653 = ~n5640 & n5650 ;
  assign n5654 = \a[23]  & ~n5653 ;
  assign n5655 = ~n5652 & ~n5654 ;
  assign n5656 = n5638 & n5655 ;
  assign n5657 = ~n5638 & ~n5655 ;
  assign n5658 = ~n5656 & ~n5657 ;
  assign n5659 = n5551 & ~n5658 ;
  assign n5660 = n5527 & n5659 ;
  assign n5661 = n5551 & n5658 ;
  assign n5662 = ~n5527 & n5661 ;
  assign n5663 = ~n5660 & ~n5662 ;
  assign n5664 = ~n5551 & ~n5658 ;
  assign n5665 = ~n5527 & n5664 ;
  assign n5666 = ~n5551 & n5658 ;
  assign n5667 = n5527 & n5666 ;
  assign n5668 = ~n5665 & ~n5667 ;
  assign n5669 = n5663 & n5668 ;
  assign n5670 = n1467 & ~n1694 ;
  assign n5671 = ~n1692 & n5670 ;
  assign n5672 = \b[15]  & n1652 ;
  assign n5673 = n1649 & n5672 ;
  assign n5674 = ~\a[15]  & \b[16]  ;
  assign n5675 = n1459 & n5674 ;
  assign n5676 = ~n5673 & ~n5675 ;
  assign n5677 = \b[17]  & n1465 ;
  assign n5678 = \a[15]  & \b[16]  ;
  assign n5679 = n1456 & n5678 ;
  assign n5680 = \a[17]  & ~n5679 ;
  assign n5681 = ~n5677 & n5680 ;
  assign n5682 = n5676 & n5681 ;
  assign n5683 = ~n5671 & n5682 ;
  assign n5684 = ~n5677 & ~n5679 ;
  assign n5685 = n5676 & n5684 ;
  assign n5686 = ~n5671 & n5685 ;
  assign n5687 = ~\a[17]  & ~n5686 ;
  assign n5688 = ~n5683 & ~n5687 ;
  assign n5689 = ~n5669 & ~n5688 ;
  assign n5690 = n5525 & n5689 ;
  assign n5691 = n5669 & ~n5688 ;
  assign n5692 = ~n5525 & n5691 ;
  assign n5693 = ~n5690 & ~n5692 ;
  assign n5694 = ~n5669 & n5688 ;
  assign n5695 = ~n5525 & n5694 ;
  assign n5696 = n5669 & n5688 ;
  assign n5697 = n5525 & n5696 ;
  assign n5698 = ~n5695 & ~n5697 ;
  assign n5699 = n5693 & n5698 ;
  assign n5700 = ~n5522 & n5699 ;
  assign n5701 = n5324 & ~n5699 ;
  assign n5702 = ~n5521 & n5701 ;
  assign n5703 = n999 & n2293 ;
  assign n5704 = ~n2290 & n5703 ;
  assign n5705 = ~n2074 & ~n2293 ;
  assign n5706 = n999 & n5705 ;
  assign n5707 = ~n2289 & n5706 ;
  assign n5708 = \b[18]  & n1182 ;
  assign n5709 = n1179 & n5708 ;
  assign n5710 = ~\a[11]  & \b[19]  ;
  assign n5711 = n1181 & n5710 ;
  assign n5712 = ~n5709 & ~n5711 ;
  assign n5713 = \b[20]  & n997 ;
  assign n5714 = \a[12]  & \b[19]  ;
  assign n5715 = n988 & n5714 ;
  assign n5716 = \a[14]  & ~n5715 ;
  assign n5717 = ~n5713 & n5716 ;
  assign n5718 = n5712 & n5717 ;
  assign n5719 = ~n5707 & n5718 ;
  assign n5720 = ~n5704 & n5719 ;
  assign n5721 = ~n5713 & ~n5715 ;
  assign n5722 = n5712 & n5721 ;
  assign n5723 = ~n5707 & n5722 ;
  assign n5724 = ~n5704 & n5723 ;
  assign n5725 = ~\a[14]  & ~n5724 ;
  assign n5726 = ~n5720 & ~n5725 ;
  assign n5727 = ~n5702 & ~n5726 ;
  assign n5728 = ~n5700 & n5727 ;
  assign n5729 = ~n5699 & n5726 ;
  assign n5730 = n5522 & n5729 ;
  assign n5731 = n5699 & n5726 ;
  assign n5732 = ~n5522 & n5731 ;
  assign n5733 = ~n5730 & ~n5732 ;
  assign n5734 = ~n5728 & n5733 ;
  assign n5735 = n5520 & ~n5734 ;
  assign n5736 = ~n5503 & n5735 ;
  assign n5737 = n5520 & n5734 ;
  assign n5738 = n5503 & n5737 ;
  assign n5739 = ~n5736 & ~n5738 ;
  assign n5740 = ~n5520 & ~n5734 ;
  assign n5741 = n5503 & n5740 ;
  assign n5742 = ~n5520 & n5734 ;
  assign n5743 = ~n5503 & n5742 ;
  assign n5744 = ~n5741 & ~n5743 ;
  assign n5745 = n5739 & n5744 ;
  assign n5746 = n430 & ~n4141 ;
  assign n5747 = ~n4518 & n5746 ;
  assign n5748 = \b[24]  & n486 ;
  assign n5749 = n483 & n5748 ;
  assign n5750 = ~\a[6]  & \b[25]  ;
  assign n5751 = n422 & n5750 ;
  assign n5752 = ~n5749 & ~n5751 ;
  assign n5753 = \b[26]  & n428 ;
  assign n5754 = \a[6]  & \b[25]  ;
  assign n5755 = n419 & n5754 ;
  assign n5756 = \a[8]  & ~n5755 ;
  assign n5757 = ~n5753 & n5756 ;
  assign n5758 = n5752 & n5757 ;
  assign n5759 = ~n5747 & n5758 ;
  assign n5760 = ~n5753 & ~n5755 ;
  assign n5761 = n5752 & n5760 ;
  assign n5762 = ~n5747 & n5761 ;
  assign n5763 = ~\a[8]  & ~n5762 ;
  assign n5764 = ~n5759 & ~n5763 ;
  assign n5765 = ~n5745 & ~n5764 ;
  assign n5766 = ~n5500 & n5765 ;
  assign n5767 = n5745 & ~n5764 ;
  assign n5768 = n5500 & n5767 ;
  assign n5769 = ~n5766 & ~n5768 ;
  assign n5770 = ~n5745 & n5764 ;
  assign n5771 = n5500 & n5770 ;
  assign n5772 = n5745 & n5764 ;
  assign n5773 = ~n5500 & n5772 ;
  assign n5774 = ~n5771 & ~n5773 ;
  assign n5775 = n5769 & n5774 ;
  assign n5776 = n252 & ~n4502 ;
  assign n5777 = ~n4500 & n5776 ;
  assign n5778 = \b[29]  & n250 ;
  assign n5779 = \a[3]  & \b[28]  ;
  assign n5780 = n241 & n5779 ;
  assign n5781 = ~n5778 & ~n5780 ;
  assign n5782 = \b[27]  & n303 ;
  assign n5783 = n300 & n5782 ;
  assign n5784 = ~\a[3]  & \b[28]  ;
  assign n5785 = n244 & n5784 ;
  assign n5786 = ~n5783 & ~n5785 ;
  assign n5787 = n5781 & n5786 ;
  assign n5788 = ~n5777 & n5787 ;
  assign n5789 = ~\a[5]  & ~n5788 ;
  assign n5790 = \a[5]  & n5787 ;
  assign n5791 = ~n5777 & n5790 ;
  assign n5792 = ~n5789 & ~n5791 ;
  assign n5793 = ~n5775 & ~n5792 ;
  assign n5794 = n5499 & n5793 ;
  assign n5795 = n5775 & ~n5792 ;
  assign n5796 = ~n5499 & n5795 ;
  assign n5797 = ~n5794 & ~n5796 ;
  assign n5798 = ~n5775 & n5792 ;
  assign n5799 = ~n5499 & n5798 ;
  assign n5800 = n5775 & n5792 ;
  assign n5801 = n5499 & n5800 ;
  assign n5802 = ~n5799 & ~n5801 ;
  assign n5803 = n5797 & n5802 ;
  assign n5804 = ~n5496 & n5803 ;
  assign n5805 = ~n5104 & ~n5458 ;
  assign n5806 = ~n5455 & n5805 ;
  assign n5807 = ~n5457 & ~n5806 ;
  assign n5808 = ~\b[31]  & ~\b[32]  ;
  assign n5809 = \b[31]  & \b[32]  ;
  assign n5810 = ~n5808 & ~n5809 ;
  assign n5811 = n134 & n5810 ;
  assign n5812 = ~n5807 & n5811 ;
  assign n5813 = n134 & ~n5810 ;
  assign n5814 = ~n5457 & n5813 ;
  assign n5815 = ~n5806 & n5814 ;
  assign n5816 = \a[0]  & \b[32]  ;
  assign n5817 = n133 & n5816 ;
  assign n5818 = \b[31]  & n141 ;
  assign n5819 = ~\a[1]  & \b[30]  ;
  assign n5820 = n1521 & n5819 ;
  assign n5821 = ~n5818 & ~n5820 ;
  assign n5822 = ~n5817 & n5821 ;
  assign n5823 = \a[2]  & n5822 ;
  assign n5824 = ~n5815 & n5823 ;
  assign n5825 = ~n5812 & n5824 ;
  assign n5826 = ~n5815 & n5822 ;
  assign n5827 = ~n5812 & n5826 ;
  assign n5828 = ~\a[2]  & ~n5827 ;
  assign n5829 = ~n5825 & ~n5828 ;
  assign n5830 = n5447 & ~n5803 ;
  assign n5831 = ~n5495 & n5830 ;
  assign n5832 = ~n5829 & ~n5831 ;
  assign n5833 = ~n5804 & n5832 ;
  assign n5834 = ~n5803 & n5829 ;
  assign n5835 = n5496 & n5834 ;
  assign n5836 = n5803 & n5829 ;
  assign n5837 = ~n5496 & n5836 ;
  assign n5838 = ~n5835 & ~n5837 ;
  assign n5839 = ~n5833 & n5838 ;
  assign n5840 = n5494 & n5839 ;
  assign n5841 = ~n5494 & ~n5839 ;
  assign n5842 = ~n5840 & ~n5841 ;
  assign n5843 = ~n5833 & ~n5840 ;
  assign n5844 = n5447 & n5797 ;
  assign n5845 = ~n5495 & n5844 ;
  assign n5846 = n5802 & ~n5845 ;
  assign n5847 = ~n5457 & n5810 ;
  assign n5848 = ~n5806 & n5847 ;
  assign n5849 = ~n5809 & ~n5848 ;
  assign n5850 = ~\b[32]  & ~\b[33]  ;
  assign n5851 = \b[32]  & \b[33]  ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = ~n5849 & n5852 ;
  assign n5854 = ~n5809 & ~n5852 ;
  assign n5855 = ~n5848 & n5854 ;
  assign n5856 = n134 & ~n5855 ;
  assign n5857 = ~n5853 & n5856 ;
  assign n5858 = \a[0]  & \b[33]  ;
  assign n5859 = n133 & n5858 ;
  assign n5860 = \b[32]  & n141 ;
  assign n5861 = ~\a[1]  & \b[31]  ;
  assign n5862 = n1521 & n5861 ;
  assign n5863 = ~n5860 & ~n5862 ;
  assign n5864 = ~n5859 & n5863 ;
  assign n5865 = ~n5857 & n5864 ;
  assign n5866 = ~\a[2]  & ~n5865 ;
  assign n5867 = \a[2]  & n5864 ;
  assign n5868 = ~n5857 & n5867 ;
  assign n5869 = ~n5866 & ~n5868 ;
  assign n5870 = n5499 & n5775 ;
  assign n5871 = n5769 & ~n5870 ;
  assign n5872 = ~n5389 & n5744 ;
  assign n5873 = ~n5397 & n5872 ;
  assign n5874 = n5739 & ~n5873 ;
  assign n5875 = n5503 & n5734 ;
  assign n5876 = ~n5728 & ~n5875 ;
  assign n5877 = n646 & n3283 ;
  assign n5878 = ~n3280 & n5877 ;
  assign n5879 = n646 & n4107 ;
  assign n5880 = ~n3279 & n5879 ;
  assign n5881 = \b[22]  & n796 ;
  assign n5882 = n793 & n5881 ;
  assign n5883 = ~\a[9]  & \b[23]  ;
  assign n5884 = n638 & n5883 ;
  assign n5885 = ~n5882 & ~n5884 ;
  assign n5886 = \b[24]  & n644 ;
  assign n5887 = \a[9]  & \b[23]  ;
  assign n5888 = n635 & n5887 ;
  assign n5889 = \a[11]  & ~n5888 ;
  assign n5890 = ~n5886 & n5889 ;
  assign n5891 = n5885 & n5890 ;
  assign n5892 = ~n5880 & n5891 ;
  assign n5893 = ~n5878 & n5892 ;
  assign n5894 = ~n5886 & ~n5888 ;
  assign n5895 = n5885 & n5894 ;
  assign n5896 = ~n5880 & n5895 ;
  assign n5897 = ~n5878 & n5896 ;
  assign n5898 = ~\a[11]  & ~n5897 ;
  assign n5899 = ~n5893 & ~n5898 ;
  assign n5900 = n5324 & n5693 ;
  assign n5901 = ~n5521 & n5900 ;
  assign n5902 = n5698 & ~n5901 ;
  assign n5903 = n5525 & n5669 ;
  assign n5904 = n5668 & ~n5903 ;
  assign n5905 = n5254 & ~n5656 ;
  assign n5906 = ~n5526 & n5905 ;
  assign n5907 = ~n5657 & ~n5906 ;
  assign n5908 = ~n5632 & ~n5637 ;
  assign n5909 = ~n5219 & ~n5603 ;
  assign n5910 = ~n5222 & n5909 ;
  assign n5911 = ~n5604 & ~n5910 ;
  assign n5912 = ~n586 & n3402 ;
  assign n5913 = ~n504 & n3402 ;
  assign n5914 = ~n508 & n5913 ;
  assign n5915 = ~n5912 & ~n5914 ;
  assign n5916 = ~n589 & ~n5915 ;
  assign n5917 = \b[7]  & n3733 ;
  assign n5918 = n3730 & n5917 ;
  assign n5919 = \b[9]  & n3400 ;
  assign n5920 = \a[24]  & \b[8]  ;
  assign n5921 = n3391 & n5920 ;
  assign n5922 = ~\a[24]  & \b[8]  ;
  assign n5923 = n3394 & n5922 ;
  assign n5924 = ~n5921 & ~n5923 ;
  assign n5925 = ~n5919 & n5924 ;
  assign n5926 = ~n5918 & n5925 ;
  assign n5927 = ~\a[26]  & n5926 ;
  assign n5928 = ~n5916 & n5927 ;
  assign n5929 = \a[26]  & ~n5926 ;
  assign n5930 = \a[26]  & ~n589 ;
  assign n5931 = ~n5915 & n5930 ;
  assign n5932 = ~n5929 & ~n5931 ;
  assign n5933 = ~n5928 & n5932 ;
  assign n5934 = n177 & n5211 ;
  assign n5935 = \b[3]  & n5209 ;
  assign n5936 = \a[29]  & \b[2]  ;
  assign n5937 = n5593 & n5936 ;
  assign n5938 = ~\a[30]  & \b[2]  ;
  assign n5939 = n5203 & n5938 ;
  assign n5940 = ~n5937 & ~n5939 ;
  assign n5941 = ~n5935 & n5940 ;
  assign n5942 = ~n5934 & n5941 ;
  assign n5943 = \b[1]  & n5595 ;
  assign n5944 = n5592 & n5943 ;
  assign n5945 = ~\a[32]  & ~n5944 ;
  assign n5946 = n5942 & n5945 ;
  assign n5947 = n5942 & ~n5944 ;
  assign n5948 = \a[32]  & ~n5947 ;
  assign n5949 = ~n5946 & ~n5948 ;
  assign n5950 = \a[32]  & ~\a[33]  ;
  assign n5951 = ~\a[32]  & \a[33]  ;
  assign n5952 = ~n5950 & ~n5951 ;
  assign n5953 = \b[0]  & ~n5952 ;
  assign n5954 = n5582 & n5599 ;
  assign n5955 = n5953 & n5954 ;
  assign n5956 = ~n5953 & ~n5954 ;
  assign n5957 = ~n5955 & ~n5956 ;
  assign n5958 = n5949 & n5957 ;
  assign n5959 = ~n5949 & ~n5957 ;
  assign n5960 = ~n5958 & ~n5959 ;
  assign n5961 = ~n323 & ~n3956 ;
  assign n5962 = ~n4246 & n5961 ;
  assign n5963 = n320 & n5962 ;
  assign n5964 = n323 & ~n3956 ;
  assign n5965 = ~n4246 & n5964 ;
  assign n5966 = ~n320 & n5965 ;
  assign n5967 = ~n5963 & ~n5966 ;
  assign n5968 = \b[4]  & n4647 ;
  assign n5969 = n4644 & n5968 ;
  assign n5970 = ~\a[26]  & \b[5]  ;
  assign n5971 = n4646 & n5970 ;
  assign n5972 = ~n5969 & ~n5971 ;
  assign n5973 = \b[6]  & n4247 ;
  assign n5974 = \a[27]  & \b[5]  ;
  assign n5975 = n4238 & n5974 ;
  assign n5976 = \a[29]  & ~n5975 ;
  assign n5977 = ~n5973 & n5976 ;
  assign n5978 = n5972 & n5977 ;
  assign n5979 = n5967 & n5978 ;
  assign n5980 = ~n5973 & ~n5975 ;
  assign n5981 = n5972 & n5980 ;
  assign n5982 = n5967 & n5981 ;
  assign n5983 = ~\a[29]  & ~n5982 ;
  assign n5984 = ~n5979 & ~n5983 ;
  assign n5985 = n5960 & ~n5984 ;
  assign n5986 = ~n5960 & n5984 ;
  assign n5987 = ~n5985 & ~n5986 ;
  assign n5988 = n5933 & ~n5987 ;
  assign n5989 = n5911 & n5988 ;
  assign n5990 = n5933 & n5987 ;
  assign n5991 = ~n5911 & n5990 ;
  assign n5992 = ~n5989 & ~n5991 ;
  assign n5993 = ~n5933 & ~n5987 ;
  assign n5994 = ~n5911 & n5993 ;
  assign n5995 = ~n5933 & n5987 ;
  assign n5996 = n5911 & n5995 ;
  assign n5997 = ~n5994 & ~n5996 ;
  assign n5998 = n5992 & n5997 ;
  assign n5999 = ~n909 & ~n2413 ;
  assign n6000 = ~n2619 & n5999 ;
  assign n6001 = n906 & n6000 ;
  assign n6002 = n909 & ~n2413 ;
  assign n6003 = ~n2619 & n6002 ;
  assign n6004 = ~n906 & n6003 ;
  assign n6005 = ~n6001 & ~n6004 ;
  assign n6006 = \b[10]  & n2912 ;
  assign n6007 = n2909 & n6006 ;
  assign n6008 = \b[12]  & n2620 ;
  assign n6009 = \a[20]  & \b[11]  ;
  assign n6010 = n2910 & n6009 ;
  assign n6011 = ~\a[21]  & \b[11]  ;
  assign n6012 = n2614 & n6011 ;
  assign n6013 = ~n6010 & ~n6012 ;
  assign n6014 = ~n6008 & n6013 ;
  assign n6015 = ~n6007 & n6014 ;
  assign n6016 = n6005 & n6015 ;
  assign n6017 = ~\a[23]  & ~n6016 ;
  assign n6018 = \a[23]  & n6015 ;
  assign n6019 = n6005 & n6018 ;
  assign n6020 = ~n6017 & ~n6019 ;
  assign n6021 = ~n5998 & n6020 ;
  assign n6022 = n5908 & n6021 ;
  assign n6023 = n5998 & n6020 ;
  assign n6024 = ~n5908 & n6023 ;
  assign n6025 = ~n6022 & ~n6024 ;
  assign n6026 = ~n5908 & n5998 ;
  assign n6027 = ~n5632 & ~n5998 ;
  assign n6028 = ~n5637 & n6027 ;
  assign n6029 = ~n6020 & ~n6028 ;
  assign n6030 = ~n6026 & n6029 ;
  assign n6031 = n6025 & ~n6030 ;
  assign n6032 = ~n1233 & n1965 ;
  assign n6033 = ~n1231 & n6032 ;
  assign n6034 = \b[13]  & n2218 ;
  assign n6035 = n2216 & n6034 ;
  assign n6036 = ~\a[18]  & \b[14]  ;
  assign n6037 = n1957 & n6036 ;
  assign n6038 = ~n6035 & ~n6037 ;
  assign n6039 = \b[15]  & n1963 ;
  assign n6040 = \a[18]  & \b[14]  ;
  assign n6041 = n2210 & n6040 ;
  assign n6042 = \a[20]  & ~n6041 ;
  assign n6043 = ~n6039 & n6042 ;
  assign n6044 = n6038 & n6043 ;
  assign n6045 = ~n6033 & n6044 ;
  assign n6046 = ~n6039 & ~n6041 ;
  assign n6047 = n6038 & n6046 ;
  assign n6048 = ~n6033 & n6047 ;
  assign n6049 = ~\a[20]  & ~n6048 ;
  assign n6050 = ~n6045 & ~n6049 ;
  assign n6051 = ~n6031 & ~n6050 ;
  assign n6052 = n5907 & n6051 ;
  assign n6053 = n6031 & ~n6050 ;
  assign n6054 = ~n5907 & n6053 ;
  assign n6055 = ~n6052 & ~n6054 ;
  assign n6056 = ~n6031 & n6050 ;
  assign n6057 = ~n5907 & n6056 ;
  assign n6058 = n6031 & n6050 ;
  assign n6059 = n5907 & n6058 ;
  assign n6060 = ~n6057 & ~n6059 ;
  assign n6061 = n6055 & n6060 ;
  assign n6062 = ~n5904 & n6061 ;
  assign n6063 = n1467 & n1875 ;
  assign n6064 = ~n1872 & n6063 ;
  assign n6065 = n1467 & n5000 ;
  assign n6066 = ~n1871 & n6065 ;
  assign n6067 = \b[16]  & n1652 ;
  assign n6068 = n1649 & n6067 ;
  assign n6069 = ~\a[15]  & \b[17]  ;
  assign n6070 = n1459 & n6069 ;
  assign n6071 = ~n6068 & ~n6070 ;
  assign n6072 = \b[18]  & n1465 ;
  assign n6073 = \a[15]  & \b[17]  ;
  assign n6074 = n1456 & n6073 ;
  assign n6075 = \a[17]  & ~n6074 ;
  assign n6076 = ~n6072 & n6075 ;
  assign n6077 = n6071 & n6076 ;
  assign n6078 = ~n6066 & n6077 ;
  assign n6079 = ~n6064 & n6078 ;
  assign n6080 = ~n6072 & ~n6074 ;
  assign n6081 = n6071 & n6080 ;
  assign n6082 = ~n6066 & n6081 ;
  assign n6083 = ~n6064 & n6082 ;
  assign n6084 = ~\a[17]  & ~n6083 ;
  assign n6085 = ~n6079 & ~n6084 ;
  assign n6086 = n5668 & ~n6061 ;
  assign n6087 = ~n5903 & n6086 ;
  assign n6088 = ~n6085 & ~n6087 ;
  assign n6089 = ~n6062 & n6088 ;
  assign n6090 = ~n6061 & n6085 ;
  assign n6091 = n5904 & n6090 ;
  assign n6092 = n6061 & n6085 ;
  assign n6093 = ~n5904 & n6092 ;
  assign n6094 = ~n6091 & ~n6093 ;
  assign n6095 = ~n6089 & n6094 ;
  assign n6096 = n999 & ~n2523 ;
  assign n6097 = ~n2521 & n6096 ;
  assign n6098 = \b[19]  & n1182 ;
  assign n6099 = n1179 & n6098 ;
  assign n6100 = ~\a[11]  & \b[20]  ;
  assign n6101 = n1181 & n6100 ;
  assign n6102 = ~n6099 & ~n6101 ;
  assign n6103 = \b[21]  & n997 ;
  assign n6104 = \a[12]  & \b[20]  ;
  assign n6105 = n988 & n6104 ;
  assign n6106 = \a[14]  & ~n6105 ;
  assign n6107 = ~n6103 & n6106 ;
  assign n6108 = n6102 & n6107 ;
  assign n6109 = ~n6097 & n6108 ;
  assign n6110 = ~n6103 & ~n6105 ;
  assign n6111 = n6102 & n6110 ;
  assign n6112 = ~n6097 & n6111 ;
  assign n6113 = ~\a[14]  & ~n6112 ;
  assign n6114 = ~n6109 & ~n6113 ;
  assign n6115 = ~n6095 & ~n6114 ;
  assign n6116 = n5902 & n6115 ;
  assign n6117 = n6095 & ~n6114 ;
  assign n6118 = ~n5902 & n6117 ;
  assign n6119 = ~n6116 & ~n6118 ;
  assign n6120 = ~n6095 & n6114 ;
  assign n6121 = ~n5902 & n6120 ;
  assign n6122 = n6095 & n6114 ;
  assign n6123 = n5902 & n6122 ;
  assign n6124 = ~n6121 & ~n6123 ;
  assign n6125 = n6119 & n6124 ;
  assign n6126 = n5899 & ~n6125 ;
  assign n6127 = n5876 & n6126 ;
  assign n6128 = n5899 & n6125 ;
  assign n6129 = ~n5876 & n6128 ;
  assign n6130 = ~n6127 & ~n6129 ;
  assign n6131 = ~n5876 & n6125 ;
  assign n6132 = ~n5728 & ~n6125 ;
  assign n6133 = ~n5875 & n6132 ;
  assign n6134 = ~n5899 & ~n6133 ;
  assign n6135 = ~n6131 & n6134 ;
  assign n6136 = n6130 & ~n6135 ;
  assign n6137 = n5874 & n6136 ;
  assign n6138 = ~n5874 & ~n6136 ;
  assign n6139 = ~n6137 & ~n6138 ;
  assign n6140 = n430 & ~n4148 ;
  assign n6141 = ~n4146 & n6140 ;
  assign n6142 = \b[27]  & n428 ;
  assign n6143 = \a[6]  & \b[26]  ;
  assign n6144 = n419 & n6143 ;
  assign n6145 = ~n6142 & ~n6144 ;
  assign n6146 = \b[25]  & n486 ;
  assign n6147 = n483 & n6146 ;
  assign n6148 = ~\a[6]  & \b[26]  ;
  assign n6149 = n422 & n6148 ;
  assign n6150 = ~n6147 & ~n6149 ;
  assign n6151 = n6145 & n6150 ;
  assign n6152 = ~n6141 & n6151 ;
  assign n6153 = ~\a[8]  & ~n6152 ;
  assign n6154 = \a[8]  & n6151 ;
  assign n6155 = ~n6141 & n6154 ;
  assign n6156 = ~n6153 & ~n6155 ;
  assign n6157 = n6139 & ~n6156 ;
  assign n6158 = ~n6139 & n6156 ;
  assign n6159 = ~n6157 & ~n6158 ;
  assign n6160 = ~n5102 & ~n5105 ;
  assign n6161 = n252 & ~n5455 ;
  assign n6162 = ~n6160 & n6161 ;
  assign n6163 = \b[28]  & n303 ;
  assign n6164 = n300 & n6163 ;
  assign n6165 = ~\a[3]  & \b[29]  ;
  assign n6166 = n244 & n6165 ;
  assign n6167 = ~n6164 & ~n6166 ;
  assign n6168 = \b[30]  & n250 ;
  assign n6169 = \a[3]  & \b[29]  ;
  assign n6170 = n241 & n6169 ;
  assign n6171 = \a[5]  & ~n6170 ;
  assign n6172 = ~n6168 & n6171 ;
  assign n6173 = n6167 & n6172 ;
  assign n6174 = ~n6162 & n6173 ;
  assign n6175 = ~n6168 & ~n6170 ;
  assign n6176 = n6167 & n6175 ;
  assign n6177 = ~n6162 & n6176 ;
  assign n6178 = ~\a[5]  & ~n6177 ;
  assign n6179 = ~n6174 & ~n6178 ;
  assign n6180 = ~n6159 & ~n6179 ;
  assign n6181 = ~n5871 & n6180 ;
  assign n6182 = n6159 & ~n6179 ;
  assign n6183 = n5871 & n6182 ;
  assign n6184 = ~n6181 & ~n6183 ;
  assign n6185 = ~n6159 & n6179 ;
  assign n6186 = n5871 & n6185 ;
  assign n6187 = n6159 & n6179 ;
  assign n6188 = ~n5871 & n6187 ;
  assign n6189 = ~n6186 & ~n6188 ;
  assign n6190 = n6184 & n6189 ;
  assign n6191 = ~n5869 & ~n6190 ;
  assign n6192 = n5846 & n6191 ;
  assign n6193 = ~n5869 & n6190 ;
  assign n6194 = ~n5846 & n6193 ;
  assign n6195 = ~n6192 & ~n6194 ;
  assign n6196 = n5869 & ~n6190 ;
  assign n6197 = ~n5846 & n6196 ;
  assign n6198 = n5869 & n6190 ;
  assign n6199 = n5846 & n6198 ;
  assign n6200 = ~n6197 & ~n6199 ;
  assign n6201 = n6195 & n6200 ;
  assign n6202 = ~n5843 & n6201 ;
  assign n6203 = ~n5833 & ~n6201 ;
  assign n6204 = ~n5840 & n6203 ;
  assign n6205 = ~n6202 & ~n6204 ;
  assign n6206 = ~n5833 & n6195 ;
  assign n6207 = ~n5840 & n6206 ;
  assign n6208 = n6200 & ~n6207 ;
  assign n6209 = n5846 & n6190 ;
  assign n6210 = n6184 & ~n6209 ;
  assign n6211 = n5769 & ~n6157 ;
  assign n6212 = ~n5870 & n6211 ;
  assign n6213 = ~n6158 & ~n6212 ;
  assign n6214 = ~n6135 & ~n6137 ;
  assign n6215 = n430 & n4456 ;
  assign n6216 = ~n4453 & n6215 ;
  assign n6217 = n430 & n5421 ;
  assign n6218 = ~n4452 & n6217 ;
  assign n6219 = \b[26]  & n486 ;
  assign n6220 = n483 & n6219 ;
  assign n6221 = ~\a[6]  & \b[27]  ;
  assign n6222 = n422 & n6221 ;
  assign n6223 = ~n6220 & ~n6222 ;
  assign n6224 = \b[28]  & n428 ;
  assign n6225 = \a[6]  & \b[27]  ;
  assign n6226 = n419 & n6225 ;
  assign n6227 = \a[8]  & ~n6226 ;
  assign n6228 = ~n6224 & n6227 ;
  assign n6229 = n6223 & n6228 ;
  assign n6230 = ~n6218 & n6229 ;
  assign n6231 = ~n6216 & n6230 ;
  assign n6232 = ~n6224 & ~n6226 ;
  assign n6233 = n6223 & n6232 ;
  assign n6234 = ~n6218 & n6233 ;
  assign n6235 = ~n6216 & n6234 ;
  assign n6236 = ~\a[8]  & ~n6235 ;
  assign n6237 = ~n6231 & ~n6236 ;
  assign n6238 = ~n5728 & n6119 ;
  assign n6239 = ~n5875 & n6238 ;
  assign n6240 = n6124 & ~n6239 ;
  assign n6241 = n5902 & n6095 ;
  assign n6242 = ~n6089 & ~n6241 ;
  assign n6243 = n5668 & n6055 ;
  assign n6244 = ~n5903 & n6243 ;
  assign n6245 = n6060 & ~n6244 ;
  assign n6246 = n5907 & n6031 ;
  assign n6247 = ~n6030 & ~n6246 ;
  assign n6248 = ~n5632 & n5992 ;
  assign n6249 = ~n5637 & n6248 ;
  assign n6250 = n5997 & ~n6249 ;
  assign n6251 = n5911 & n5987 ;
  assign n6252 = ~n5985 & ~n6251 ;
  assign n6253 = ~n380 & n4249 ;
  assign n6254 = ~n322 & n4249 ;
  assign n6255 = ~n326 & n6254 ;
  assign n6256 = ~n6253 & ~n6255 ;
  assign n6257 = ~n383 & ~n6256 ;
  assign n6258 = \b[5]  & n4647 ;
  assign n6259 = n4644 & n6258 ;
  assign n6260 = ~\a[26]  & \b[6]  ;
  assign n6261 = n4646 & n6260 ;
  assign n6262 = ~n6259 & ~n6261 ;
  assign n6263 = \b[7]  & n4247 ;
  assign n6264 = \a[27]  & \b[6]  ;
  assign n6265 = n4238 & n6264 ;
  assign n6266 = \a[29]  & ~n6265 ;
  assign n6267 = ~n6263 & n6266 ;
  assign n6268 = n6262 & n6267 ;
  assign n6269 = ~n6257 & n6268 ;
  assign n6270 = ~n6263 & ~n6265 ;
  assign n6271 = n6262 & n6270 ;
  assign n6272 = ~\a[29]  & ~n6271 ;
  assign n6273 = ~\a[29]  & ~n383 ;
  assign n6274 = ~n6256 & n6273 ;
  assign n6275 = ~n6272 & ~n6274 ;
  assign n6276 = ~n6269 & n6275 ;
  assign n6277 = ~n5955 & ~n5958 ;
  assign n6278 = n222 & n5211 ;
  assign n6279 = \b[4]  & n5209 ;
  assign n6280 = \a[29]  & \b[3]  ;
  assign n6281 = n5593 & n6280 ;
  assign n6282 = ~\a[30]  & \b[3]  ;
  assign n6283 = n5203 & n6282 ;
  assign n6284 = ~n6281 & ~n6283 ;
  assign n6285 = ~n6279 & n6284 ;
  assign n6286 = \b[2]  & n5595 ;
  assign n6287 = n5592 & n6286 ;
  assign n6288 = \a[32]  & ~n6287 ;
  assign n6289 = n6285 & n6288 ;
  assign n6290 = ~n6278 & n6289 ;
  assign n6291 = n6285 & ~n6287 ;
  assign n6292 = ~n6278 & n6291 ;
  assign n6293 = ~\a[32]  & ~n6292 ;
  assign n6294 = ~n6290 & ~n6293 ;
  assign n6295 = \a[35]  & \b[0]  ;
  assign n6296 = ~n5952 & n6295 ;
  assign n6297 = \a[33]  & \b[0]  ;
  assign n6298 = \a[32]  & ~\a[34]  ;
  assign n6299 = n6297 & n6298 ;
  assign n6300 = ~\a[33]  & \b[0]  ;
  assign n6301 = ~\a[32]  & \a[34]  ;
  assign n6302 = n6300 & n6301 ;
  assign n6303 = ~n6299 & ~n6302 ;
  assign n6304 = \a[34]  & ~\a[35]  ;
  assign n6305 = ~\a[34]  & \a[35]  ;
  assign n6306 = ~n6304 & ~n6305 ;
  assign n6307 = ~n5952 & n6306 ;
  assign n6308 = \b[1]  & n6307 ;
  assign n6309 = ~n5952 & ~n6306 ;
  assign n6310 = ~n137 & n6309 ;
  assign n6311 = ~n6308 & ~n6310 ;
  assign n6312 = n6303 & n6311 ;
  assign n6313 = n6296 & ~n6312 ;
  assign n6314 = ~n6296 & n6303 ;
  assign n6315 = n6311 & n6314 ;
  assign n6316 = ~n6313 & ~n6315 ;
  assign n6317 = n6294 & ~n6316 ;
  assign n6318 = ~n6294 & n6316 ;
  assign n6319 = ~n6317 & ~n6318 ;
  assign n6320 = ~n6277 & n6319 ;
  assign n6321 = n6277 & ~n6319 ;
  assign n6322 = ~n6320 & ~n6321 ;
  assign n6323 = n6276 & ~n6322 ;
  assign n6324 = ~n6276 & n6322 ;
  assign n6325 = ~n6323 & ~n6324 ;
  assign n6326 = ~n685 & ~n3154 ;
  assign n6327 = ~n3399 & n6326 ;
  assign n6328 = n682 & n6327 ;
  assign n6329 = n685 & ~n3154 ;
  assign n6330 = ~n3399 & n6329 ;
  assign n6331 = ~n682 & n6330 ;
  assign n6332 = ~n6328 & ~n6331 ;
  assign n6333 = \b[8]  & n3733 ;
  assign n6334 = n3730 & n6333 ;
  assign n6335 = \b[10]  & n3400 ;
  assign n6336 = \a[24]  & \b[9]  ;
  assign n6337 = n3391 & n6336 ;
  assign n6338 = ~\a[24]  & \b[9]  ;
  assign n6339 = n3394 & n6338 ;
  assign n6340 = ~n6337 & ~n6339 ;
  assign n6341 = ~n6335 & n6340 ;
  assign n6342 = ~n6334 & n6341 ;
  assign n6343 = n6332 & n6342 ;
  assign n6344 = ~\a[26]  & ~n6343 ;
  assign n6345 = \a[26]  & n6342 ;
  assign n6346 = n6332 & n6345 ;
  assign n6347 = ~n6344 & ~n6346 ;
  assign n6348 = ~n6325 & ~n6347 ;
  assign n6349 = ~n6252 & n6348 ;
  assign n6350 = n6325 & ~n6347 ;
  assign n6351 = n6252 & n6350 ;
  assign n6352 = ~n6349 & ~n6351 ;
  assign n6353 = ~n6325 & n6347 ;
  assign n6354 = n6252 & n6353 ;
  assign n6355 = n6325 & n6347 ;
  assign n6356 = ~n6252 & n6355 ;
  assign n6357 = ~n6354 & ~n6356 ;
  assign n6358 = n6352 & n6357 ;
  assign n6359 = ~n948 & n2622 ;
  assign n6360 = ~n908 & n2622 ;
  assign n6361 = ~n912 & n6360 ;
  assign n6362 = ~n6359 & ~n6361 ;
  assign n6363 = ~n951 & ~n6362 ;
  assign n6364 = \b[11]  & n2912 ;
  assign n6365 = n2909 & n6364 ;
  assign n6366 = \b[13]  & n2620 ;
  assign n6367 = \a[20]  & \b[12]  ;
  assign n6368 = n2910 & n6367 ;
  assign n6369 = ~\a[21]  & \b[12]  ;
  assign n6370 = n2614 & n6369 ;
  assign n6371 = ~n6368 & ~n6370 ;
  assign n6372 = ~n6366 & n6371 ;
  assign n6373 = ~n6365 & n6372 ;
  assign n6374 = ~\a[23]  & n6373 ;
  assign n6375 = ~n6363 & n6374 ;
  assign n6376 = \a[23]  & ~n6373 ;
  assign n6377 = \a[23]  & ~n951 ;
  assign n6378 = ~n6362 & n6377 ;
  assign n6379 = ~n6376 & ~n6378 ;
  assign n6380 = ~n6375 & n6379 ;
  assign n6381 = ~n6358 & n6380 ;
  assign n6382 = n6250 & n6381 ;
  assign n6383 = n6358 & n6380 ;
  assign n6384 = ~n6250 & n6383 ;
  assign n6385 = ~n6382 & ~n6384 ;
  assign n6386 = ~n6358 & ~n6380 ;
  assign n6387 = ~n6250 & n6386 ;
  assign n6388 = n6358 & ~n6380 ;
  assign n6389 = n6250 & n6388 ;
  assign n6390 = ~n6387 & ~n6389 ;
  assign n6391 = n6385 & n6390 ;
  assign n6392 = ~n6247 & n6391 ;
  assign n6393 = ~n1512 & ~n1805 ;
  assign n6394 = ~n1962 & n6393 ;
  assign n6395 = n1509 & n6394 ;
  assign n6396 = n1512 & ~n1805 ;
  assign n6397 = ~n1962 & n6396 ;
  assign n6398 = ~n1509 & n6397 ;
  assign n6399 = ~n6395 & ~n6398 ;
  assign n6400 = \b[14]  & n2218 ;
  assign n6401 = n2216 & n6400 ;
  assign n6402 = ~\a[18]  & \b[15]  ;
  assign n6403 = n1957 & n6402 ;
  assign n6404 = ~n6401 & ~n6403 ;
  assign n6405 = \b[16]  & n1963 ;
  assign n6406 = \a[18]  & \b[15]  ;
  assign n6407 = n2210 & n6406 ;
  assign n6408 = \a[20]  & ~n6407 ;
  assign n6409 = ~n6405 & n6408 ;
  assign n6410 = n6404 & n6409 ;
  assign n6411 = n6399 & n6410 ;
  assign n6412 = ~n6405 & ~n6407 ;
  assign n6413 = n6404 & n6412 ;
  assign n6414 = n6399 & n6413 ;
  assign n6415 = ~\a[20]  & ~n6414 ;
  assign n6416 = ~n6411 & ~n6415 ;
  assign n6417 = ~n6030 & ~n6391 ;
  assign n6418 = ~n6246 & n6417 ;
  assign n6419 = ~n6416 & ~n6418 ;
  assign n6420 = ~n6392 & n6419 ;
  assign n6421 = ~n6391 & n6416 ;
  assign n6422 = n6247 & n6421 ;
  assign n6423 = n6391 & n6416 ;
  assign n6424 = ~n6247 & n6423 ;
  assign n6425 = ~n6422 & ~n6424 ;
  assign n6426 = ~n6420 & n6425 ;
  assign n6427 = n1467 & ~n2079 ;
  assign n6428 = ~n2077 & n6427 ;
  assign n6429 = \b[17]  & n1652 ;
  assign n6430 = n1649 & n6429 ;
  assign n6431 = ~\a[15]  & \b[18]  ;
  assign n6432 = n1459 & n6431 ;
  assign n6433 = ~n6430 & ~n6432 ;
  assign n6434 = \b[19]  & n1465 ;
  assign n6435 = \a[15]  & \b[18]  ;
  assign n6436 = n1456 & n6435 ;
  assign n6437 = \a[17]  & ~n6436 ;
  assign n6438 = ~n6434 & n6437 ;
  assign n6439 = n6433 & n6438 ;
  assign n6440 = ~n6428 & n6439 ;
  assign n6441 = ~n6434 & ~n6436 ;
  assign n6442 = n6433 & n6441 ;
  assign n6443 = ~n6428 & n6442 ;
  assign n6444 = ~\a[17]  & ~n6443 ;
  assign n6445 = ~n6440 & ~n6444 ;
  assign n6446 = ~n6426 & ~n6445 ;
  assign n6447 = n6245 & n6446 ;
  assign n6448 = n6426 & ~n6445 ;
  assign n6449 = ~n6245 & n6448 ;
  assign n6450 = ~n6447 & ~n6449 ;
  assign n6451 = ~n6426 & n6445 ;
  assign n6452 = ~n6245 & n6451 ;
  assign n6453 = n6426 & n6445 ;
  assign n6454 = n6245 & n6453 ;
  assign n6455 = ~n6452 & ~n6454 ;
  assign n6456 = n6450 & n6455 ;
  assign n6457 = ~n6242 & n6456 ;
  assign n6458 = ~n6089 & ~n6456 ;
  assign n6459 = ~n6241 & n6458 ;
  assign n6460 = n999 & n2768 ;
  assign n6461 = ~n2765 & n6460 ;
  assign n6462 = ~n2518 & ~n2768 ;
  assign n6463 = n999 & n6462 ;
  assign n6464 = ~n2764 & n6463 ;
  assign n6465 = \b[20]  & n1182 ;
  assign n6466 = n1179 & n6465 ;
  assign n6467 = ~\a[11]  & \b[21]  ;
  assign n6468 = n1181 & n6467 ;
  assign n6469 = ~n6466 & ~n6468 ;
  assign n6470 = \b[22]  & n997 ;
  assign n6471 = \a[12]  & \b[21]  ;
  assign n6472 = n988 & n6471 ;
  assign n6473 = \a[14]  & ~n6472 ;
  assign n6474 = ~n6470 & n6473 ;
  assign n6475 = n6469 & n6474 ;
  assign n6476 = ~n6464 & n6475 ;
  assign n6477 = ~n6461 & n6476 ;
  assign n6478 = ~n6470 & ~n6472 ;
  assign n6479 = n6469 & n6478 ;
  assign n6480 = ~n6464 & n6479 ;
  assign n6481 = ~n6461 & n6480 ;
  assign n6482 = ~\a[14]  & ~n6481 ;
  assign n6483 = ~n6477 & ~n6482 ;
  assign n6484 = ~n6459 & ~n6483 ;
  assign n6485 = ~n6457 & n6484 ;
  assign n6486 = ~n6456 & n6483 ;
  assign n6487 = n6242 & n6486 ;
  assign n6488 = n6456 & n6483 ;
  assign n6489 = ~n6242 & n6488 ;
  assign n6490 = ~n6487 & ~n6489 ;
  assign n6491 = ~n6485 & n6490 ;
  assign n6492 = n646 & ~n3567 ;
  assign n6493 = ~n3565 & n6492 ;
  assign n6494 = \b[25]  & n644 ;
  assign n6495 = \a[9]  & \b[24]  ;
  assign n6496 = n635 & n6495 ;
  assign n6497 = ~n6494 & ~n6496 ;
  assign n6498 = \b[23]  & n796 ;
  assign n6499 = n793 & n6498 ;
  assign n6500 = ~\a[9]  & \b[24]  ;
  assign n6501 = n638 & n6500 ;
  assign n6502 = ~n6499 & ~n6501 ;
  assign n6503 = n6497 & n6502 ;
  assign n6504 = ~n6493 & n6503 ;
  assign n6505 = ~\a[11]  & ~n6504 ;
  assign n6506 = \a[11]  & n6503 ;
  assign n6507 = ~n6493 & n6506 ;
  assign n6508 = ~n6505 & ~n6507 ;
  assign n6509 = ~n6491 & ~n6508 ;
  assign n6510 = n6240 & n6509 ;
  assign n6511 = n6491 & ~n6508 ;
  assign n6512 = ~n6240 & n6511 ;
  assign n6513 = ~n6510 & ~n6512 ;
  assign n6514 = ~n6491 & n6508 ;
  assign n6515 = ~n6240 & n6514 ;
  assign n6516 = n6491 & n6508 ;
  assign n6517 = n6240 & n6516 ;
  assign n6518 = ~n6515 & ~n6517 ;
  assign n6519 = n6513 & n6518 ;
  assign n6520 = ~n6237 & ~n6519 ;
  assign n6521 = ~n6214 & n6520 ;
  assign n6522 = ~n6237 & n6519 ;
  assign n6523 = n6214 & n6522 ;
  assign n6524 = ~n6521 & ~n6523 ;
  assign n6525 = n6237 & ~n6519 ;
  assign n6526 = n6214 & n6525 ;
  assign n6527 = n6237 & n6519 ;
  assign n6528 = ~n6214 & n6527 ;
  assign n6529 = ~n6526 & ~n6528 ;
  assign n6530 = n6524 & n6529 ;
  assign n6531 = n252 & ~n5462 ;
  assign n6532 = ~n5460 & n6531 ;
  assign n6533 = \b[31]  & n250 ;
  assign n6534 = \a[3]  & \b[30]  ;
  assign n6535 = n241 & n6534 ;
  assign n6536 = ~n6533 & ~n6535 ;
  assign n6537 = \b[29]  & n303 ;
  assign n6538 = n300 & n6537 ;
  assign n6539 = ~\a[3]  & \b[30]  ;
  assign n6540 = n244 & n6539 ;
  assign n6541 = ~n6538 & ~n6540 ;
  assign n6542 = n6536 & n6541 ;
  assign n6543 = ~n6532 & n6542 ;
  assign n6544 = ~\a[5]  & ~n6543 ;
  assign n6545 = \a[5]  & n6542 ;
  assign n6546 = ~n6532 & n6545 ;
  assign n6547 = ~n6544 & ~n6546 ;
  assign n6548 = ~n6530 & ~n6547 ;
  assign n6549 = n6213 & n6548 ;
  assign n6550 = n6530 & ~n6547 ;
  assign n6551 = ~n6213 & n6550 ;
  assign n6552 = ~n6549 & ~n6551 ;
  assign n6553 = ~n6530 & n6547 ;
  assign n6554 = ~n6213 & n6553 ;
  assign n6555 = n6530 & n6547 ;
  assign n6556 = n6213 & n6555 ;
  assign n6557 = ~n6554 & ~n6556 ;
  assign n6558 = n6552 & n6557 ;
  assign n6559 = ~n6210 & n6558 ;
  assign n6560 = ~n5809 & ~n5851 ;
  assign n6561 = ~n5848 & n6560 ;
  assign n6562 = ~n5850 & ~n6561 ;
  assign n6563 = ~\b[33]  & ~\b[34]  ;
  assign n6564 = \b[33]  & \b[34]  ;
  assign n6565 = ~n6563 & ~n6564 ;
  assign n6566 = n134 & n6565 ;
  assign n6567 = ~n6562 & n6566 ;
  assign n6568 = n134 & ~n6565 ;
  assign n6569 = ~n5850 & n6568 ;
  assign n6570 = ~n6561 & n6569 ;
  assign n6571 = \a[0]  & \b[34]  ;
  assign n6572 = n133 & n6571 ;
  assign n6573 = \b[33]  & n141 ;
  assign n6574 = ~\a[1]  & \b[32]  ;
  assign n6575 = n1521 & n6574 ;
  assign n6576 = ~n6573 & ~n6575 ;
  assign n6577 = ~n6572 & n6576 ;
  assign n6578 = \a[2]  & n6577 ;
  assign n6579 = ~n6570 & n6578 ;
  assign n6580 = ~n6567 & n6579 ;
  assign n6581 = ~n6570 & n6577 ;
  assign n6582 = ~n6567 & n6581 ;
  assign n6583 = ~\a[2]  & ~n6582 ;
  assign n6584 = ~n6580 & ~n6583 ;
  assign n6585 = n6184 & ~n6558 ;
  assign n6586 = ~n6209 & n6585 ;
  assign n6587 = ~n6584 & ~n6586 ;
  assign n6588 = ~n6559 & n6587 ;
  assign n6589 = ~n6558 & n6584 ;
  assign n6590 = n6210 & n6589 ;
  assign n6591 = n6558 & n6584 ;
  assign n6592 = ~n6210 & n6591 ;
  assign n6593 = ~n6590 & ~n6592 ;
  assign n6594 = ~n6588 & n6593 ;
  assign n6595 = n6208 & n6594 ;
  assign n6596 = ~n6208 & ~n6594 ;
  assign n6597 = ~n6595 & ~n6596 ;
  assign n6598 = ~n6588 & ~n6595 ;
  assign n6599 = n6184 & n6552 ;
  assign n6600 = ~n6209 & n6599 ;
  assign n6601 = n6557 & ~n6600 ;
  assign n6602 = ~n5850 & n6565 ;
  assign n6603 = ~n6561 & n6602 ;
  assign n6604 = ~n6564 & ~n6603 ;
  assign n6605 = ~\b[34]  & ~\b[35]  ;
  assign n6606 = \b[34]  & \b[35]  ;
  assign n6607 = ~n6605 & ~n6606 ;
  assign n6608 = ~n6604 & n6607 ;
  assign n6609 = ~n6564 & ~n6607 ;
  assign n6610 = ~n6603 & n6609 ;
  assign n6611 = n134 & ~n6610 ;
  assign n6612 = ~n6608 & n6611 ;
  assign n6613 = \a[0]  & \b[35]  ;
  assign n6614 = n133 & n6613 ;
  assign n6615 = \b[34]  & n141 ;
  assign n6616 = ~\a[1]  & \b[33]  ;
  assign n6617 = n1521 & n6616 ;
  assign n6618 = ~n6615 & ~n6617 ;
  assign n6619 = ~n6614 & n6618 ;
  assign n6620 = ~n6612 & n6619 ;
  assign n6621 = ~\a[2]  & ~n6620 ;
  assign n6622 = \a[2]  & n6619 ;
  assign n6623 = ~n6612 & n6622 ;
  assign n6624 = ~n6621 & ~n6623 ;
  assign n6625 = n6213 & n6530 ;
  assign n6626 = n6524 & ~n6625 ;
  assign n6627 = ~n6135 & n6513 ;
  assign n6628 = ~n6137 & n6627 ;
  assign n6629 = n6518 & ~n6628 ;
  assign n6630 = n6240 & n6491 ;
  assign n6631 = ~n6485 & ~n6630 ;
  assign n6632 = n646 & ~n4141 ;
  assign n6633 = ~n4518 & n6632 ;
  assign n6634 = \b[24]  & n796 ;
  assign n6635 = n793 & n6634 ;
  assign n6636 = ~\a[9]  & \b[25]  ;
  assign n6637 = n638 & n6636 ;
  assign n6638 = ~n6635 & ~n6637 ;
  assign n6639 = \b[26]  & n644 ;
  assign n6640 = \a[9]  & \b[25]  ;
  assign n6641 = n635 & n6640 ;
  assign n6642 = \a[11]  & ~n6641 ;
  assign n6643 = ~n6639 & n6642 ;
  assign n6644 = n6638 & n6643 ;
  assign n6645 = ~n6633 & n6644 ;
  assign n6646 = ~n6639 & ~n6641 ;
  assign n6647 = n6638 & n6646 ;
  assign n6648 = ~n6633 & n6647 ;
  assign n6649 = ~\a[11]  & ~n6648 ;
  assign n6650 = ~n6645 & ~n6649 ;
  assign n6651 = ~n6089 & n6450 ;
  assign n6652 = ~n6241 & n6651 ;
  assign n6653 = n6455 & ~n6652 ;
  assign n6654 = n999 & ~n3022 ;
  assign n6655 = ~n3020 & n6654 ;
  assign n6656 = \b[21]  & n1182 ;
  assign n6657 = n1179 & n6656 ;
  assign n6658 = ~\a[11]  & \b[22]  ;
  assign n6659 = n1181 & n6658 ;
  assign n6660 = ~n6657 & ~n6659 ;
  assign n6661 = \b[23]  & n997 ;
  assign n6662 = \a[12]  & \b[22]  ;
  assign n6663 = n988 & n6662 ;
  assign n6664 = \a[14]  & ~n6663 ;
  assign n6665 = ~n6661 & n6664 ;
  assign n6666 = n6660 & n6665 ;
  assign n6667 = ~n6655 & n6666 ;
  assign n6668 = ~n6661 & ~n6663 ;
  assign n6669 = n6660 & n6668 ;
  assign n6670 = ~n6655 & n6669 ;
  assign n6671 = ~\a[14]  & ~n6670 ;
  assign n6672 = ~n6667 & ~n6671 ;
  assign n6673 = n6245 & n6426 ;
  assign n6674 = ~n6420 & ~n6673 ;
  assign n6675 = ~n6030 & n6385 ;
  assign n6676 = ~n6246 & n6675 ;
  assign n6677 = n6390 & ~n6676 ;
  assign n6678 = n6250 & n6358 ;
  assign n6679 = n6352 & ~n6678 ;
  assign n6680 = n1087 & n2622 ;
  assign n6681 = ~n1084 & n6680 ;
  assign n6682 = n1552 & n2622 ;
  assign n6683 = ~n1083 & n6682 ;
  assign n6684 = \b[12]  & n2912 ;
  assign n6685 = n2909 & n6684 ;
  assign n6686 = \b[14]  & n2620 ;
  assign n6687 = \a[20]  & \b[13]  ;
  assign n6688 = n2910 & n6687 ;
  assign n6689 = ~\a[21]  & \b[13]  ;
  assign n6690 = n2614 & n6689 ;
  assign n6691 = ~n6688 & ~n6690 ;
  assign n6692 = ~n6686 & n6691 ;
  assign n6693 = ~n6685 & n6692 ;
  assign n6694 = ~n6683 & n6693 ;
  assign n6695 = ~n6681 & n6694 ;
  assign n6696 = ~\a[23]  & ~n6695 ;
  assign n6697 = \a[23]  & n6693 ;
  assign n6698 = ~n6683 & n6697 ;
  assign n6699 = ~n6681 & n6698 ;
  assign n6700 = ~n6696 & ~n6699 ;
  assign n6701 = ~n728 & n3402 ;
  assign n6702 = ~n726 & n6701 ;
  assign n6703 = \b[9]  & n3733 ;
  assign n6704 = n3730 & n6703 ;
  assign n6705 = \b[11]  & n3400 ;
  assign n6706 = \a[24]  & \b[10]  ;
  assign n6707 = n3391 & n6706 ;
  assign n6708 = ~\a[24]  & \b[10]  ;
  assign n6709 = n3394 & n6708 ;
  assign n6710 = ~n6707 & ~n6709 ;
  assign n6711 = ~n6705 & n6710 ;
  assign n6712 = ~n6704 & n6711 ;
  assign n6713 = ~\a[26]  & n6712 ;
  assign n6714 = ~n6702 & n6713 ;
  assign n6715 = ~n6702 & n6712 ;
  assign n6716 = \a[26]  & ~n6715 ;
  assign n6717 = ~n6714 & ~n6716 ;
  assign n6718 = ~n5985 & ~n6324 ;
  assign n6719 = ~n6251 & n6718 ;
  assign n6720 = ~n6323 & ~n6719 ;
  assign n6721 = ~n505 & ~n3956 ;
  assign n6722 = ~n4246 & n6721 ;
  assign n6723 = n502 & n6722 ;
  assign n6724 = n505 & ~n3956 ;
  assign n6725 = ~n4246 & n6724 ;
  assign n6726 = ~n502 & n6725 ;
  assign n6727 = ~n6723 & ~n6726 ;
  assign n6728 = \b[6]  & n4647 ;
  assign n6729 = n4644 & n6728 ;
  assign n6730 = ~\a[26]  & \b[7]  ;
  assign n6731 = n4646 & n6730 ;
  assign n6732 = ~n6729 & ~n6731 ;
  assign n6733 = \b[8]  & n4247 ;
  assign n6734 = \a[27]  & \b[7]  ;
  assign n6735 = n4238 & n6734 ;
  assign n6736 = \a[29]  & ~n6735 ;
  assign n6737 = ~n6733 & n6736 ;
  assign n6738 = n6732 & n6737 ;
  assign n6739 = n6727 & n6738 ;
  assign n6740 = ~n6733 & ~n6735 ;
  assign n6741 = n6732 & n6740 ;
  assign n6742 = n6727 & n6741 ;
  assign n6743 = ~\a[29]  & ~n6742 ;
  assign n6744 = ~n6739 & ~n6743 ;
  assign n6745 = ~n6318 & ~n6320 ;
  assign n6746 = ~n273 & n5211 ;
  assign n6747 = ~n271 & n6746 ;
  assign n6748 = \b[3]  & n5595 ;
  assign n6749 = n5592 & n6748 ;
  assign n6750 = \b[5]  & n5209 ;
  assign n6751 = \a[29]  & \b[4]  ;
  assign n6752 = n5593 & n6751 ;
  assign n6753 = ~\a[30]  & \b[4]  ;
  assign n6754 = n5203 & n6753 ;
  assign n6755 = ~n6752 & ~n6754 ;
  assign n6756 = ~n6750 & n6755 ;
  assign n6757 = ~n6749 & n6756 ;
  assign n6758 = ~n6747 & n6757 ;
  assign n6759 = ~\a[32]  & ~n6758 ;
  assign n6760 = \a[32]  & n6757 ;
  assign n6761 = ~n6747 & n6760 ;
  assign n6762 = ~n6759 & ~n6761 ;
  assign n6763 = \a[35]  & ~n5953 ;
  assign n6764 = n6303 & n6763 ;
  assign n6765 = n6311 & n6764 ;
  assign n6766 = \a[35]  & ~n6765 ;
  assign n6767 = \b[2]  & n6307 ;
  assign n6768 = ~\a[33]  & \b[1]  ;
  assign n6769 = n6301 & n6768 ;
  assign n6770 = \a[33]  & \b[1]  ;
  assign n6771 = n6298 & n6770 ;
  assign n6772 = ~n6769 & ~n6771 ;
  assign n6773 = ~n6767 & n6772 ;
  assign n6774 = n157 & n6309 ;
  assign n6775 = n5952 & ~n6306 ;
  assign n6776 = \a[33]  & ~\a[34]  ;
  assign n6777 = ~\a[33]  & \a[34]  ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = \b[0]  & n6778 ;
  assign n6780 = n6775 & n6779 ;
  assign n6781 = ~n6774 & ~n6780 ;
  assign n6782 = n6773 & n6781 ;
  assign n6783 = ~n6766 & ~n6782 ;
  assign n6784 = n6766 & n6782 ;
  assign n6785 = ~n6783 & ~n6784 ;
  assign n6786 = ~n6762 & ~n6785 ;
  assign n6787 = n6762 & n6785 ;
  assign n6788 = ~n6786 & ~n6787 ;
  assign n6789 = ~n6745 & n6788 ;
  assign n6790 = n6745 & ~n6788 ;
  assign n6791 = ~n6789 & ~n6790 ;
  assign n6792 = ~n6744 & n6791 ;
  assign n6793 = n6744 & ~n6791 ;
  assign n6794 = ~n6792 & ~n6793 ;
  assign n6795 = n6720 & n6794 ;
  assign n6796 = ~n6720 & ~n6794 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6798 = n6717 & n6797 ;
  assign n6799 = ~n6717 & ~n6797 ;
  assign n6800 = ~n6798 & ~n6799 ;
  assign n6801 = n6700 & ~n6800 ;
  assign n6802 = n6679 & n6801 ;
  assign n6803 = n6700 & n6800 ;
  assign n6804 = ~n6679 & n6803 ;
  assign n6805 = ~n6802 & ~n6804 ;
  assign n6806 = ~n6700 & ~n6800 ;
  assign n6807 = ~n6679 & n6806 ;
  assign n6808 = ~n6700 & n6800 ;
  assign n6809 = n6679 & n6808 ;
  assign n6810 = ~n6807 & ~n6809 ;
  assign n6811 = n6805 & n6810 ;
  assign n6812 = ~n1694 & n1965 ;
  assign n6813 = ~n1692 & n6812 ;
  assign n6814 = \b[15]  & n2218 ;
  assign n6815 = n2216 & n6814 ;
  assign n6816 = ~\a[18]  & \b[16]  ;
  assign n6817 = n1957 & n6816 ;
  assign n6818 = ~n6815 & ~n6817 ;
  assign n6819 = \b[17]  & n1963 ;
  assign n6820 = \a[18]  & \b[16]  ;
  assign n6821 = n2210 & n6820 ;
  assign n6822 = \a[20]  & ~n6821 ;
  assign n6823 = ~n6819 & n6822 ;
  assign n6824 = n6818 & n6823 ;
  assign n6825 = ~n6813 & n6824 ;
  assign n6826 = ~n6819 & ~n6821 ;
  assign n6827 = n6818 & n6826 ;
  assign n6828 = ~n6813 & n6827 ;
  assign n6829 = ~\a[20]  & ~n6828 ;
  assign n6830 = ~n6825 & ~n6829 ;
  assign n6831 = ~n6811 & ~n6830 ;
  assign n6832 = n6677 & n6831 ;
  assign n6833 = n6811 & ~n6830 ;
  assign n6834 = ~n6677 & n6833 ;
  assign n6835 = ~n6832 & ~n6834 ;
  assign n6836 = ~n6811 & n6830 ;
  assign n6837 = ~n6677 & n6836 ;
  assign n6838 = n6811 & n6830 ;
  assign n6839 = n6677 & n6838 ;
  assign n6840 = ~n6837 & ~n6839 ;
  assign n6841 = n6835 & n6840 ;
  assign n6842 = ~n6674 & n6841 ;
  assign n6843 = ~n6420 & ~n6841 ;
  assign n6844 = ~n6673 & n6843 ;
  assign n6845 = n1467 & n2293 ;
  assign n6846 = ~n2290 & n6845 ;
  assign n6847 = n1467 & n5705 ;
  assign n6848 = ~n2289 & n6847 ;
  assign n6849 = \b[18]  & n1652 ;
  assign n6850 = n1649 & n6849 ;
  assign n6851 = ~\a[15]  & \b[19]  ;
  assign n6852 = n1459 & n6851 ;
  assign n6853 = ~n6850 & ~n6852 ;
  assign n6854 = \b[20]  & n1465 ;
  assign n6855 = \a[15]  & \b[19]  ;
  assign n6856 = n1456 & n6855 ;
  assign n6857 = \a[17]  & ~n6856 ;
  assign n6858 = ~n6854 & n6857 ;
  assign n6859 = n6853 & n6858 ;
  assign n6860 = ~n6848 & n6859 ;
  assign n6861 = ~n6846 & n6860 ;
  assign n6862 = ~n6854 & ~n6856 ;
  assign n6863 = n6853 & n6862 ;
  assign n6864 = ~n6848 & n6863 ;
  assign n6865 = ~n6846 & n6864 ;
  assign n6866 = ~\a[17]  & ~n6865 ;
  assign n6867 = ~n6861 & ~n6866 ;
  assign n6868 = ~n6844 & ~n6867 ;
  assign n6869 = ~n6842 & n6868 ;
  assign n6870 = ~n6841 & n6867 ;
  assign n6871 = n6674 & n6870 ;
  assign n6872 = n6841 & n6867 ;
  assign n6873 = ~n6674 & n6872 ;
  assign n6874 = ~n6871 & ~n6873 ;
  assign n6875 = ~n6869 & n6874 ;
  assign n6876 = n6672 & ~n6875 ;
  assign n6877 = ~n6653 & n6876 ;
  assign n6878 = n6672 & n6875 ;
  assign n6879 = n6653 & n6878 ;
  assign n6880 = ~n6877 & ~n6879 ;
  assign n6881 = ~n6672 & ~n6875 ;
  assign n6882 = n6653 & n6881 ;
  assign n6883 = ~n6672 & n6875 ;
  assign n6884 = ~n6653 & n6883 ;
  assign n6885 = ~n6882 & ~n6884 ;
  assign n6886 = n6880 & n6885 ;
  assign n6887 = n6650 & ~n6886 ;
  assign n6888 = n6631 & n6887 ;
  assign n6889 = n6650 & n6886 ;
  assign n6890 = ~n6631 & n6889 ;
  assign n6891 = ~n6888 & ~n6890 ;
  assign n6892 = ~n6631 & n6886 ;
  assign n6893 = ~n6485 & ~n6886 ;
  assign n6894 = ~n6630 & n6893 ;
  assign n6895 = ~n6650 & ~n6894 ;
  assign n6896 = ~n6892 & n6895 ;
  assign n6897 = n6891 & ~n6896 ;
  assign n6898 = n6629 & n6897 ;
  assign n6899 = ~n6629 & ~n6897 ;
  assign n6900 = ~n6898 & ~n6899 ;
  assign n6901 = n430 & ~n4502 ;
  assign n6902 = ~n4500 & n6901 ;
  assign n6903 = \b[29]  & n428 ;
  assign n6904 = \a[6]  & \b[28]  ;
  assign n6905 = n419 & n6904 ;
  assign n6906 = ~n6903 & ~n6905 ;
  assign n6907 = \b[27]  & n486 ;
  assign n6908 = n483 & n6907 ;
  assign n6909 = ~\a[6]  & \b[28]  ;
  assign n6910 = n422 & n6909 ;
  assign n6911 = ~n6908 & ~n6910 ;
  assign n6912 = n6906 & n6911 ;
  assign n6913 = ~n6902 & n6912 ;
  assign n6914 = ~\a[8]  & ~n6913 ;
  assign n6915 = \a[8]  & n6912 ;
  assign n6916 = ~n6902 & n6915 ;
  assign n6917 = ~n6914 & ~n6916 ;
  assign n6918 = n6900 & ~n6917 ;
  assign n6919 = ~n6900 & n6917 ;
  assign n6920 = ~n6918 & ~n6919 ;
  assign n6921 = n252 & n5810 ;
  assign n6922 = ~n5807 & n6921 ;
  assign n6923 = n252 & ~n5810 ;
  assign n6924 = ~n5457 & n6923 ;
  assign n6925 = ~n5806 & n6924 ;
  assign n6926 = \b[30]  & n303 ;
  assign n6927 = n300 & n6926 ;
  assign n6928 = ~\a[3]  & \b[31]  ;
  assign n6929 = n244 & n6928 ;
  assign n6930 = ~n6927 & ~n6929 ;
  assign n6931 = \b[32]  & n250 ;
  assign n6932 = \a[3]  & \b[31]  ;
  assign n6933 = n241 & n6932 ;
  assign n6934 = \a[5]  & ~n6933 ;
  assign n6935 = ~n6931 & n6934 ;
  assign n6936 = n6930 & n6935 ;
  assign n6937 = ~n6925 & n6936 ;
  assign n6938 = ~n6922 & n6937 ;
  assign n6939 = ~n6931 & ~n6933 ;
  assign n6940 = n6930 & n6939 ;
  assign n6941 = ~n6925 & n6940 ;
  assign n6942 = ~n6922 & n6941 ;
  assign n6943 = ~\a[5]  & ~n6942 ;
  assign n6944 = ~n6938 & ~n6943 ;
  assign n6945 = ~n6920 & ~n6944 ;
  assign n6946 = ~n6626 & n6945 ;
  assign n6947 = n6920 & ~n6944 ;
  assign n6948 = n6626 & n6947 ;
  assign n6949 = ~n6946 & ~n6948 ;
  assign n6950 = ~n6920 & n6944 ;
  assign n6951 = n6626 & n6950 ;
  assign n6952 = n6920 & n6944 ;
  assign n6953 = ~n6626 & n6952 ;
  assign n6954 = ~n6951 & ~n6953 ;
  assign n6955 = n6949 & n6954 ;
  assign n6956 = ~n6624 & ~n6955 ;
  assign n6957 = n6601 & n6956 ;
  assign n6958 = ~n6624 & n6955 ;
  assign n6959 = ~n6601 & n6958 ;
  assign n6960 = ~n6957 & ~n6959 ;
  assign n6961 = n6624 & ~n6955 ;
  assign n6962 = ~n6601 & n6961 ;
  assign n6963 = n6624 & n6955 ;
  assign n6964 = n6601 & n6963 ;
  assign n6965 = ~n6962 & ~n6964 ;
  assign n6966 = n6960 & n6965 ;
  assign n6967 = ~n6598 & n6966 ;
  assign n6968 = ~n6588 & ~n6966 ;
  assign n6969 = ~n6595 & n6968 ;
  assign n6970 = ~n6967 & ~n6969 ;
  assign n6971 = ~n6588 & n6960 ;
  assign n6972 = ~n6595 & n6971 ;
  assign n6973 = n6965 & ~n6972 ;
  assign n6974 = n6601 & n6955 ;
  assign n6975 = n6949 & ~n6974 ;
  assign n6976 = n6524 & ~n6918 ;
  assign n6977 = ~n6625 & n6976 ;
  assign n6978 = ~n6919 & ~n6977 ;
  assign n6979 = n252 & ~n5855 ;
  assign n6980 = ~n5853 & n6979 ;
  assign n6981 = \b[33]  & n250 ;
  assign n6982 = \a[3]  & \b[32]  ;
  assign n6983 = n241 & n6982 ;
  assign n6984 = ~n6981 & ~n6983 ;
  assign n6985 = \b[31]  & n303 ;
  assign n6986 = n300 & n6985 ;
  assign n6987 = ~\a[3]  & \b[32]  ;
  assign n6988 = n244 & n6987 ;
  assign n6989 = ~n6986 & ~n6988 ;
  assign n6990 = n6984 & n6989 ;
  assign n6991 = ~n6980 & n6990 ;
  assign n6992 = ~\a[5]  & ~n6991 ;
  assign n6993 = \a[5]  & n6990 ;
  assign n6994 = ~n6980 & n6993 ;
  assign n6995 = ~n6992 & ~n6994 ;
  assign n6996 = ~n6896 & ~n6898 ;
  assign n6997 = n430 & ~n5455 ;
  assign n6998 = ~n6160 & n6997 ;
  assign n6999 = \b[28]  & n486 ;
  assign n7000 = n483 & n6999 ;
  assign n7001 = ~\a[6]  & \b[29]  ;
  assign n7002 = n422 & n7001 ;
  assign n7003 = ~n7000 & ~n7002 ;
  assign n7004 = \b[30]  & n428 ;
  assign n7005 = \a[6]  & \b[29]  ;
  assign n7006 = n419 & n7005 ;
  assign n7007 = \a[8]  & ~n7006 ;
  assign n7008 = ~n7004 & n7007 ;
  assign n7009 = n7003 & n7008 ;
  assign n7010 = ~n6998 & n7009 ;
  assign n7011 = ~n7004 & ~n7006 ;
  assign n7012 = n7003 & n7011 ;
  assign n7013 = ~n6998 & n7012 ;
  assign n7014 = ~\a[8]  & ~n7013 ;
  assign n7015 = ~n7010 & ~n7014 ;
  assign n7016 = ~n6485 & n6885 ;
  assign n7017 = ~n6630 & n7016 ;
  assign n7018 = n6880 & ~n7017 ;
  assign n7019 = n6653 & n6875 ;
  assign n7020 = ~n6869 & ~n7019 ;
  assign n7021 = n999 & n3283 ;
  assign n7022 = ~n3280 & n7021 ;
  assign n7023 = n999 & n4107 ;
  assign n7024 = ~n3279 & n7023 ;
  assign n7025 = \b[22]  & n1182 ;
  assign n7026 = n1179 & n7025 ;
  assign n7027 = ~\a[11]  & \b[23]  ;
  assign n7028 = n1181 & n7027 ;
  assign n7029 = ~n7026 & ~n7028 ;
  assign n7030 = \b[24]  & n997 ;
  assign n7031 = \a[12]  & \b[23]  ;
  assign n7032 = n988 & n7031 ;
  assign n7033 = \a[14]  & ~n7032 ;
  assign n7034 = ~n7030 & n7033 ;
  assign n7035 = n7029 & n7034 ;
  assign n7036 = ~n7024 & n7035 ;
  assign n7037 = ~n7022 & n7036 ;
  assign n7038 = ~n7030 & ~n7032 ;
  assign n7039 = n7029 & n7038 ;
  assign n7040 = ~n7024 & n7039 ;
  assign n7041 = ~n7022 & n7040 ;
  assign n7042 = ~\a[14]  & ~n7041 ;
  assign n7043 = ~n7037 & ~n7042 ;
  assign n7044 = ~n6420 & n6835 ;
  assign n7045 = ~n6673 & n7044 ;
  assign n7046 = n6840 & ~n7045 ;
  assign n7047 = n6677 & n6811 ;
  assign n7048 = n6810 & ~n7047 ;
  assign n7049 = n6352 & ~n6798 ;
  assign n7050 = ~n6678 & n7049 ;
  assign n7051 = ~n6799 & ~n7050 ;
  assign n7052 = ~n6792 & ~n6795 ;
  assign n7053 = ~n6318 & ~n6786 ;
  assign n7054 = ~n6320 & n7053 ;
  assign n7055 = ~n6787 & ~n7054 ;
  assign n7056 = ~n586 & n4249 ;
  assign n7057 = ~n504 & n4249 ;
  assign n7058 = ~n508 & n7057 ;
  assign n7059 = ~n7056 & ~n7058 ;
  assign n7060 = ~n589 & ~n7059 ;
  assign n7061 = \b[7]  & n4647 ;
  assign n7062 = n4644 & n7061 ;
  assign n7063 = ~\a[26]  & \b[8]  ;
  assign n7064 = n4646 & n7063 ;
  assign n7065 = ~n7062 & ~n7064 ;
  assign n7066 = \b[9]  & n4247 ;
  assign n7067 = \a[27]  & \b[8]  ;
  assign n7068 = n4238 & n7067 ;
  assign n7069 = \a[29]  & ~n7068 ;
  assign n7070 = ~n7066 & n7069 ;
  assign n7071 = n7065 & n7070 ;
  assign n7072 = ~n7060 & n7071 ;
  assign n7073 = ~n7066 & ~n7068 ;
  assign n7074 = n7065 & n7073 ;
  assign n7075 = ~\a[29]  & ~n7074 ;
  assign n7076 = ~\a[29]  & ~n589 ;
  assign n7077 = ~n7059 & n7076 ;
  assign n7078 = ~n7075 & ~n7077 ;
  assign n7079 = ~n7072 & n7078 ;
  assign n7080 = n177 & n6309 ;
  assign n7081 = \b[3]  & n6307 ;
  assign n7082 = \a[32]  & \b[2]  ;
  assign n7083 = n6776 & n7082 ;
  assign n7084 = ~\a[33]  & \b[2]  ;
  assign n7085 = n6301 & n7084 ;
  assign n7086 = ~n7083 & ~n7085 ;
  assign n7087 = ~n7081 & n7086 ;
  assign n7088 = ~n7080 & n7087 ;
  assign n7089 = \b[1]  & n6778 ;
  assign n7090 = n6775 & n7089 ;
  assign n7091 = ~\a[35]  & ~n7090 ;
  assign n7092 = n7088 & n7091 ;
  assign n7093 = n7088 & ~n7090 ;
  assign n7094 = \a[35]  & ~n7093 ;
  assign n7095 = ~n7092 & ~n7094 ;
  assign n7096 = \a[35]  & ~\a[36]  ;
  assign n7097 = ~\a[35]  & \a[36]  ;
  assign n7098 = ~n7096 & ~n7097 ;
  assign n7099 = \b[0]  & ~n7098 ;
  assign n7100 = n6765 & n6782 ;
  assign n7101 = n7099 & n7100 ;
  assign n7102 = ~n7099 & ~n7100 ;
  assign n7103 = ~n7101 & ~n7102 ;
  assign n7104 = n7095 & n7103 ;
  assign n7105 = ~n7095 & ~n7103 ;
  assign n7106 = ~n7104 & ~n7105 ;
  assign n7107 = ~n323 & ~n4909 ;
  assign n7108 = ~n5208 & n7107 ;
  assign n7109 = n320 & n7108 ;
  assign n7110 = n323 & ~n4909 ;
  assign n7111 = ~n5208 & n7110 ;
  assign n7112 = ~n320 & n7111 ;
  assign n7113 = ~n7109 & ~n7112 ;
  assign n7114 = \b[4]  & n5595 ;
  assign n7115 = n5592 & n7114 ;
  assign n7116 = \b[6]  & n5209 ;
  assign n7117 = \a[29]  & \b[5]  ;
  assign n7118 = n5593 & n7117 ;
  assign n7119 = ~\a[30]  & \b[5]  ;
  assign n7120 = n5203 & n7119 ;
  assign n7121 = ~n7118 & ~n7120 ;
  assign n7122 = ~n7116 & n7121 ;
  assign n7123 = ~n7115 & n7122 ;
  assign n7124 = n7113 & n7123 ;
  assign n7125 = ~\a[32]  & ~n7124 ;
  assign n7126 = \a[32]  & n7123 ;
  assign n7127 = n7113 & n7126 ;
  assign n7128 = ~n7125 & ~n7127 ;
  assign n7129 = n7106 & ~n7128 ;
  assign n7130 = ~n7106 & n7128 ;
  assign n7131 = ~n7129 & ~n7130 ;
  assign n7132 = ~n7079 & ~n7131 ;
  assign n7133 = n7055 & n7132 ;
  assign n7134 = ~n7079 & n7131 ;
  assign n7135 = ~n7055 & n7134 ;
  assign n7136 = ~n7133 & ~n7135 ;
  assign n7137 = n7079 & ~n7131 ;
  assign n7138 = ~n7055 & n7137 ;
  assign n7139 = n7079 & n7131 ;
  assign n7140 = n7055 & n7139 ;
  assign n7141 = ~n7138 & ~n7140 ;
  assign n7142 = n7136 & n7141 ;
  assign n7143 = ~n909 & ~n3154 ;
  assign n7144 = ~n3399 & n7143 ;
  assign n7145 = n906 & n7144 ;
  assign n7146 = n909 & ~n3154 ;
  assign n7147 = ~n3399 & n7146 ;
  assign n7148 = ~n906 & n7147 ;
  assign n7149 = ~n7145 & ~n7148 ;
  assign n7150 = \b[10]  & n3733 ;
  assign n7151 = n3730 & n7150 ;
  assign n7152 = \b[12]  & n3400 ;
  assign n7153 = \a[24]  & \b[11]  ;
  assign n7154 = n3391 & n7153 ;
  assign n7155 = ~\a[24]  & \b[11]  ;
  assign n7156 = n3394 & n7155 ;
  assign n7157 = ~n7154 & ~n7156 ;
  assign n7158 = ~n7152 & n7157 ;
  assign n7159 = ~n7151 & n7158 ;
  assign n7160 = n7149 & n7159 ;
  assign n7161 = ~\a[26]  & ~n7160 ;
  assign n7162 = \a[26]  & n7159 ;
  assign n7163 = n7149 & n7162 ;
  assign n7164 = ~n7161 & ~n7163 ;
  assign n7165 = ~n7142 & n7164 ;
  assign n7166 = n7052 & n7165 ;
  assign n7167 = n7142 & n7164 ;
  assign n7168 = ~n7052 & n7167 ;
  assign n7169 = ~n7166 & ~n7168 ;
  assign n7170 = ~n7052 & n7142 ;
  assign n7171 = ~n6792 & ~n7142 ;
  assign n7172 = ~n6795 & n7171 ;
  assign n7173 = ~n7164 & ~n7172 ;
  assign n7174 = ~n7170 & n7173 ;
  assign n7175 = n7169 & ~n7174 ;
  assign n7176 = ~n1233 & n2622 ;
  assign n7177 = ~n1231 & n7176 ;
  assign n7178 = \b[13]  & n2912 ;
  assign n7179 = n2909 & n7178 ;
  assign n7180 = \b[15]  & n2620 ;
  assign n7181 = \a[21]  & \b[14]  ;
  assign n7182 = n2611 & n7181 ;
  assign n7183 = ~\a[21]  & \b[14]  ;
  assign n7184 = n2614 & n7183 ;
  assign n7185 = ~n7182 & ~n7184 ;
  assign n7186 = ~n7180 & n7185 ;
  assign n7187 = ~n7179 & n7186 ;
  assign n7188 = ~\a[23]  & n7187 ;
  assign n7189 = ~n7177 & n7188 ;
  assign n7190 = ~n7177 & n7187 ;
  assign n7191 = \a[23]  & ~n7190 ;
  assign n7192 = ~n7189 & ~n7191 ;
  assign n7193 = n7175 & n7192 ;
  assign n7194 = ~n7051 & n7193 ;
  assign n7195 = ~n7175 & n7192 ;
  assign n7196 = n7051 & n7195 ;
  assign n7197 = ~n7194 & ~n7196 ;
  assign n7198 = ~n7175 & ~n7192 ;
  assign n7199 = ~n7051 & n7198 ;
  assign n7200 = n7175 & ~n7192 ;
  assign n7201 = n7051 & n7200 ;
  assign n7202 = ~n7199 & ~n7201 ;
  assign n7203 = n7197 & n7202 ;
  assign n7204 = ~n7048 & n7203 ;
  assign n7205 = n1875 & n1965 ;
  assign n7206 = ~n1872 & n7205 ;
  assign n7207 = n1965 & n5000 ;
  assign n7208 = ~n1871 & n7207 ;
  assign n7209 = \b[16]  & n2218 ;
  assign n7210 = n2216 & n7209 ;
  assign n7211 = ~\a[18]  & \b[17]  ;
  assign n7212 = n1957 & n7211 ;
  assign n7213 = ~n7210 & ~n7212 ;
  assign n7214 = \b[18]  & n1963 ;
  assign n7215 = \a[18]  & \b[17]  ;
  assign n7216 = n2210 & n7215 ;
  assign n7217 = \a[20]  & ~n7216 ;
  assign n7218 = ~n7214 & n7217 ;
  assign n7219 = n7213 & n7218 ;
  assign n7220 = ~n7208 & n7219 ;
  assign n7221 = ~n7206 & n7220 ;
  assign n7222 = ~n7214 & ~n7216 ;
  assign n7223 = n7213 & n7222 ;
  assign n7224 = ~n7208 & n7223 ;
  assign n7225 = ~n7206 & n7224 ;
  assign n7226 = ~\a[20]  & ~n7225 ;
  assign n7227 = ~n7221 & ~n7226 ;
  assign n7228 = n6810 & ~n7203 ;
  assign n7229 = ~n7047 & n7228 ;
  assign n7230 = ~n7227 & ~n7229 ;
  assign n7231 = ~n7204 & n7230 ;
  assign n7232 = ~n7203 & n7227 ;
  assign n7233 = n7048 & n7232 ;
  assign n7234 = n7203 & n7227 ;
  assign n7235 = ~n7048 & n7234 ;
  assign n7236 = ~n7233 & ~n7235 ;
  assign n7237 = ~n7231 & n7236 ;
  assign n7238 = n1467 & ~n2523 ;
  assign n7239 = ~n2521 & n7238 ;
  assign n7240 = \b[19]  & n1652 ;
  assign n7241 = n1649 & n7240 ;
  assign n7242 = ~\a[15]  & \b[20]  ;
  assign n7243 = n1459 & n7242 ;
  assign n7244 = ~n7241 & ~n7243 ;
  assign n7245 = \b[21]  & n1465 ;
  assign n7246 = \a[15]  & \b[20]  ;
  assign n7247 = n1456 & n7246 ;
  assign n7248 = \a[17]  & ~n7247 ;
  assign n7249 = ~n7245 & n7248 ;
  assign n7250 = n7244 & n7249 ;
  assign n7251 = ~n7239 & n7250 ;
  assign n7252 = ~n7245 & ~n7247 ;
  assign n7253 = n7244 & n7252 ;
  assign n7254 = ~n7239 & n7253 ;
  assign n7255 = ~\a[17]  & ~n7254 ;
  assign n7256 = ~n7251 & ~n7255 ;
  assign n7257 = ~n7237 & ~n7256 ;
  assign n7258 = n7046 & n7257 ;
  assign n7259 = n7237 & ~n7256 ;
  assign n7260 = ~n7046 & n7259 ;
  assign n7261 = ~n7258 & ~n7260 ;
  assign n7262 = ~n7237 & n7256 ;
  assign n7263 = ~n7046 & n7262 ;
  assign n7264 = n7237 & n7256 ;
  assign n7265 = n7046 & n7264 ;
  assign n7266 = ~n7263 & ~n7265 ;
  assign n7267 = n7261 & n7266 ;
  assign n7268 = n7043 & ~n7267 ;
  assign n7269 = n7020 & n7268 ;
  assign n7270 = n7043 & n7267 ;
  assign n7271 = ~n7020 & n7270 ;
  assign n7272 = ~n7269 & ~n7271 ;
  assign n7273 = ~n7020 & n7267 ;
  assign n7274 = ~n6869 & ~n7267 ;
  assign n7275 = ~n7019 & n7274 ;
  assign n7276 = ~n7043 & ~n7275 ;
  assign n7277 = ~n7273 & n7276 ;
  assign n7278 = n7272 & ~n7277 ;
  assign n7279 = n646 & ~n4148 ;
  assign n7280 = ~n4146 & n7279 ;
  assign n7281 = \b[27]  & n644 ;
  assign n7282 = \a[9]  & \b[26]  ;
  assign n7283 = n635 & n7282 ;
  assign n7284 = ~n7281 & ~n7283 ;
  assign n7285 = \b[25]  & n796 ;
  assign n7286 = n793 & n7285 ;
  assign n7287 = ~\a[9]  & \b[26]  ;
  assign n7288 = n638 & n7287 ;
  assign n7289 = ~n7286 & ~n7288 ;
  assign n7290 = n7284 & n7289 ;
  assign n7291 = ~n7280 & n7290 ;
  assign n7292 = ~\a[11]  & ~n7291 ;
  assign n7293 = \a[11]  & n7290 ;
  assign n7294 = ~n7280 & n7293 ;
  assign n7295 = ~n7292 & ~n7294 ;
  assign n7296 = ~n7278 & ~n7295 ;
  assign n7297 = n7018 & n7296 ;
  assign n7298 = n7278 & ~n7295 ;
  assign n7299 = ~n7018 & n7298 ;
  assign n7300 = ~n7297 & ~n7299 ;
  assign n7301 = ~n7278 & n7295 ;
  assign n7302 = ~n7018 & n7301 ;
  assign n7303 = n7278 & n7295 ;
  assign n7304 = n7018 & n7303 ;
  assign n7305 = ~n7302 & ~n7304 ;
  assign n7306 = n7300 & n7305 ;
  assign n7307 = n7015 & ~n7306 ;
  assign n7308 = n6996 & n7307 ;
  assign n7309 = n7015 & n7306 ;
  assign n7310 = ~n6996 & n7309 ;
  assign n7311 = ~n7308 & ~n7310 ;
  assign n7312 = ~n7015 & ~n7306 ;
  assign n7313 = ~n6996 & n7312 ;
  assign n7314 = ~n7015 & n7306 ;
  assign n7315 = n6996 & n7314 ;
  assign n7316 = ~n7313 & ~n7315 ;
  assign n7317 = n7311 & n7316 ;
  assign n7318 = ~n6995 & ~n7317 ;
  assign n7319 = n6978 & n7318 ;
  assign n7320 = ~n6995 & n7317 ;
  assign n7321 = ~n6978 & n7320 ;
  assign n7322 = ~n7319 & ~n7321 ;
  assign n7323 = n6995 & ~n7317 ;
  assign n7324 = ~n6978 & n7323 ;
  assign n7325 = n6995 & n7317 ;
  assign n7326 = n6978 & n7325 ;
  assign n7327 = ~n7324 & ~n7326 ;
  assign n7328 = n7322 & n7327 ;
  assign n7329 = ~n6975 & n7328 ;
  assign n7330 = n6949 & ~n7328 ;
  assign n7331 = ~n6974 & n7330 ;
  assign n7332 = ~n6564 & ~n6606 ;
  assign n7333 = ~n6603 & n7332 ;
  assign n7334 = ~n6605 & ~n7333 ;
  assign n7335 = ~\b[35]  & ~\b[36]  ;
  assign n7336 = \b[35]  & \b[36]  ;
  assign n7337 = ~n7335 & ~n7336 ;
  assign n7338 = n134 & n7337 ;
  assign n7339 = ~n7334 & n7338 ;
  assign n7340 = n134 & ~n7337 ;
  assign n7341 = ~n6605 & n7340 ;
  assign n7342 = ~n7333 & n7341 ;
  assign n7343 = \a[0]  & \b[36]  ;
  assign n7344 = n133 & n7343 ;
  assign n7345 = \b[35]  & n141 ;
  assign n7346 = ~\a[1]  & \b[34]  ;
  assign n7347 = n1521 & n7346 ;
  assign n7348 = ~n7345 & ~n7347 ;
  assign n7349 = ~n7344 & n7348 ;
  assign n7350 = \a[2]  & n7349 ;
  assign n7351 = ~n7342 & n7350 ;
  assign n7352 = ~n7339 & n7351 ;
  assign n7353 = ~n7342 & n7349 ;
  assign n7354 = ~n7339 & n7353 ;
  assign n7355 = ~\a[2]  & ~n7354 ;
  assign n7356 = ~n7352 & ~n7355 ;
  assign n7357 = ~n7331 & ~n7356 ;
  assign n7358 = ~n7329 & n7357 ;
  assign n7359 = ~n7328 & n7356 ;
  assign n7360 = n6975 & n7359 ;
  assign n7361 = n7328 & n7356 ;
  assign n7362 = ~n6975 & n7361 ;
  assign n7363 = ~n7360 & ~n7362 ;
  assign n7364 = ~n7358 & n7363 ;
  assign n7365 = n6973 & n7364 ;
  assign n7366 = ~n6973 & ~n7364 ;
  assign n7367 = ~n7365 & ~n7366 ;
  assign n7368 = ~n7358 & ~n7365 ;
  assign n7369 = n6949 & n7322 ;
  assign n7370 = ~n6974 & n7369 ;
  assign n7371 = n7327 & ~n7370 ;
  assign n7372 = n6978 & n7317 ;
  assign n7373 = n7316 & ~n7372 ;
  assign n7374 = n430 & ~n5462 ;
  assign n7375 = ~n5460 & n7374 ;
  assign n7376 = \b[31]  & n428 ;
  assign n7377 = \a[6]  & \b[30]  ;
  assign n7378 = n419 & n7377 ;
  assign n7379 = ~n7376 & ~n7378 ;
  assign n7380 = \b[29]  & n486 ;
  assign n7381 = n483 & n7380 ;
  assign n7382 = ~\a[6]  & \b[30]  ;
  assign n7383 = n422 & n7382 ;
  assign n7384 = ~n7381 & ~n7383 ;
  assign n7385 = n7379 & n7384 ;
  assign n7386 = ~n7375 & n7385 ;
  assign n7387 = ~\a[8]  & ~n7386 ;
  assign n7388 = \a[8]  & n7385 ;
  assign n7389 = ~n7375 & n7388 ;
  assign n7390 = ~n7387 & ~n7389 ;
  assign n7391 = ~n6896 & n7300 ;
  assign n7392 = ~n6898 & n7391 ;
  assign n7393 = n7305 & ~n7392 ;
  assign n7394 = n7018 & n7278 ;
  assign n7395 = ~n7277 & ~n7394 ;
  assign n7396 = n646 & n4456 ;
  assign n7397 = ~n4453 & n7396 ;
  assign n7398 = n646 & n5421 ;
  assign n7399 = ~n4452 & n7398 ;
  assign n7400 = \b[26]  & n796 ;
  assign n7401 = n793 & n7400 ;
  assign n7402 = ~\a[9]  & \b[27]  ;
  assign n7403 = n638 & n7402 ;
  assign n7404 = ~n7401 & ~n7403 ;
  assign n7405 = \b[28]  & n644 ;
  assign n7406 = \a[9]  & \b[27]  ;
  assign n7407 = n635 & n7406 ;
  assign n7408 = \a[11]  & ~n7407 ;
  assign n7409 = ~n7405 & n7408 ;
  assign n7410 = n7404 & n7409 ;
  assign n7411 = ~n7399 & n7410 ;
  assign n7412 = ~n7397 & n7411 ;
  assign n7413 = ~n7405 & ~n7407 ;
  assign n7414 = n7404 & n7413 ;
  assign n7415 = ~n7399 & n7414 ;
  assign n7416 = ~n7397 & n7415 ;
  assign n7417 = ~\a[11]  & ~n7416 ;
  assign n7418 = ~n7412 & ~n7417 ;
  assign n7419 = ~n6869 & n7261 ;
  assign n7420 = ~n7019 & n7419 ;
  assign n7421 = n7266 & ~n7420 ;
  assign n7422 = n7046 & n7237 ;
  assign n7423 = ~n7231 & ~n7422 ;
  assign n7424 = n6810 & n7197 ;
  assign n7425 = ~n7047 & n7424 ;
  assign n7426 = n7202 & ~n7425 ;
  assign n7427 = n7051 & n7175 ;
  assign n7428 = ~n7174 & ~n7427 ;
  assign n7429 = ~n6792 & n7136 ;
  assign n7430 = ~n6795 & n7429 ;
  assign n7431 = n7141 & ~n7430 ;
  assign n7432 = ~n948 & n3402 ;
  assign n7433 = ~n908 & n3402 ;
  assign n7434 = ~n912 & n7433 ;
  assign n7435 = ~n7432 & ~n7434 ;
  assign n7436 = ~n951 & ~n7435 ;
  assign n7437 = \b[11]  & n3733 ;
  assign n7438 = n3730 & n7437 ;
  assign n7439 = \b[13]  & n3400 ;
  assign n7440 = \a[24]  & \b[12]  ;
  assign n7441 = n3391 & n7440 ;
  assign n7442 = ~\a[24]  & \b[12]  ;
  assign n7443 = n3394 & n7442 ;
  assign n7444 = ~n7441 & ~n7443 ;
  assign n7445 = ~n7439 & n7444 ;
  assign n7446 = ~n7438 & n7445 ;
  assign n7447 = ~\a[26]  & n7446 ;
  assign n7448 = ~n7436 & n7447 ;
  assign n7449 = \a[26]  & ~n7446 ;
  assign n7450 = \a[26]  & ~n951 ;
  assign n7451 = ~n7435 & n7450 ;
  assign n7452 = ~n7449 & ~n7451 ;
  assign n7453 = ~n7448 & n7452 ;
  assign n7454 = n7055 & n7131 ;
  assign n7455 = ~n7129 & ~n7454 ;
  assign n7456 = ~n685 & ~n3956 ;
  assign n7457 = ~n4246 & n7456 ;
  assign n7458 = n682 & n7457 ;
  assign n7459 = n685 & ~n3956 ;
  assign n7460 = ~n4246 & n7459 ;
  assign n7461 = ~n682 & n7460 ;
  assign n7462 = ~n7458 & ~n7461 ;
  assign n7463 = \b[8]  & n4647 ;
  assign n7464 = n4644 & n7463 ;
  assign n7465 = ~\a[26]  & \b[9]  ;
  assign n7466 = n4646 & n7465 ;
  assign n7467 = ~n7464 & ~n7466 ;
  assign n7468 = \b[10]  & n4247 ;
  assign n7469 = \a[27]  & \b[9]  ;
  assign n7470 = n4238 & n7469 ;
  assign n7471 = \a[29]  & ~n7470 ;
  assign n7472 = ~n7468 & n7471 ;
  assign n7473 = n7467 & n7472 ;
  assign n7474 = n7462 & n7473 ;
  assign n7475 = ~n7468 & ~n7470 ;
  assign n7476 = n7467 & n7475 ;
  assign n7477 = n7462 & n7476 ;
  assign n7478 = ~\a[29]  & ~n7477 ;
  assign n7479 = ~n7474 & ~n7478 ;
  assign n7480 = ~n380 & n5211 ;
  assign n7481 = ~n322 & n5211 ;
  assign n7482 = ~n326 & n7481 ;
  assign n7483 = ~n7480 & ~n7482 ;
  assign n7484 = ~n383 & ~n7483 ;
  assign n7485 = \b[5]  & n5595 ;
  assign n7486 = n5592 & n7485 ;
  assign n7487 = \b[7]  & n5209 ;
  assign n7488 = \a[29]  & \b[6]  ;
  assign n7489 = n5593 & n7488 ;
  assign n7490 = ~\a[30]  & \b[6]  ;
  assign n7491 = n5203 & n7490 ;
  assign n7492 = ~n7489 & ~n7491 ;
  assign n7493 = ~n7487 & n7492 ;
  assign n7494 = ~n7486 & n7493 ;
  assign n7495 = ~\a[32]  & n7494 ;
  assign n7496 = ~n7484 & n7495 ;
  assign n7497 = \a[32]  & ~n7494 ;
  assign n7498 = \a[32]  & ~n383 ;
  assign n7499 = ~n7483 & n7498 ;
  assign n7500 = ~n7497 & ~n7499 ;
  assign n7501 = ~n7496 & n7500 ;
  assign n7502 = ~n7101 & ~n7104 ;
  assign n7503 = n222 & n6309 ;
  assign n7504 = \b[4]  & n6307 ;
  assign n7505 = \a[32]  & \b[3]  ;
  assign n7506 = n6776 & n7505 ;
  assign n7507 = ~\a[33]  & \b[3]  ;
  assign n7508 = n6301 & n7507 ;
  assign n7509 = ~n7506 & ~n7508 ;
  assign n7510 = ~n7504 & n7509 ;
  assign n7511 = \b[2]  & n6778 ;
  assign n7512 = n6775 & n7511 ;
  assign n7513 = \a[35]  & ~n7512 ;
  assign n7514 = n7510 & n7513 ;
  assign n7515 = ~n7503 & n7514 ;
  assign n7516 = n7510 & ~n7512 ;
  assign n7517 = ~n7503 & n7516 ;
  assign n7518 = ~\a[35]  & ~n7517 ;
  assign n7519 = ~n7515 & ~n7518 ;
  assign n7520 = \a[38]  & \b[0]  ;
  assign n7521 = ~n7098 & n7520 ;
  assign n7522 = \a[36]  & \b[0]  ;
  assign n7523 = \a[35]  & ~\a[37]  ;
  assign n7524 = n7522 & n7523 ;
  assign n7525 = ~\a[36]  & \b[0]  ;
  assign n7526 = ~\a[35]  & \a[37]  ;
  assign n7527 = n7525 & n7526 ;
  assign n7528 = ~n7524 & ~n7527 ;
  assign n7529 = \a[37]  & ~\a[38]  ;
  assign n7530 = ~\a[37]  & \a[38]  ;
  assign n7531 = ~n7529 & ~n7530 ;
  assign n7532 = ~n7098 & n7531 ;
  assign n7533 = \b[1]  & n7532 ;
  assign n7534 = ~n7098 & ~n7531 ;
  assign n7535 = ~n137 & n7534 ;
  assign n7536 = ~n7533 & ~n7535 ;
  assign n7537 = n7528 & n7536 ;
  assign n7538 = n7521 & ~n7537 ;
  assign n7539 = ~n7521 & n7528 ;
  assign n7540 = n7536 & n7539 ;
  assign n7541 = ~n7538 & ~n7540 ;
  assign n7542 = n7519 & ~n7541 ;
  assign n7543 = ~n7519 & n7541 ;
  assign n7544 = ~n7542 & ~n7543 ;
  assign n7545 = ~n7502 & n7544 ;
  assign n7546 = n7502 & ~n7544 ;
  assign n7547 = ~n7545 & ~n7546 ;
  assign n7548 = ~n7501 & ~n7547 ;
  assign n7549 = n7501 & n7547 ;
  assign n7550 = ~n7548 & ~n7549 ;
  assign n7551 = n7479 & ~n7550 ;
  assign n7552 = n7455 & n7551 ;
  assign n7553 = n7479 & n7550 ;
  assign n7554 = ~n7455 & n7553 ;
  assign n7555 = ~n7552 & ~n7554 ;
  assign n7556 = ~n7479 & ~n7550 ;
  assign n7557 = ~n7455 & n7556 ;
  assign n7558 = ~n7479 & n7550 ;
  assign n7559 = n7455 & n7558 ;
  assign n7560 = ~n7557 & ~n7559 ;
  assign n7561 = n7555 & n7560 ;
  assign n7562 = ~n7453 & ~n7561 ;
  assign n7563 = ~n7431 & n7562 ;
  assign n7564 = ~n7453 & n7561 ;
  assign n7565 = n7431 & n7564 ;
  assign n7566 = ~n7563 & ~n7565 ;
  assign n7567 = n7453 & ~n7561 ;
  assign n7568 = n7431 & n7567 ;
  assign n7569 = n7453 & n7561 ;
  assign n7570 = ~n7431 & n7569 ;
  assign n7571 = ~n7568 & ~n7570 ;
  assign n7572 = n7566 & n7571 ;
  assign n7573 = ~n7428 & n7572 ;
  assign n7574 = ~n7174 & ~n7572 ;
  assign n7575 = ~n7427 & n7574 ;
  assign n7576 = ~n1512 & ~n2413 ;
  assign n7577 = ~n2619 & n7576 ;
  assign n7578 = n1509 & n7577 ;
  assign n7579 = n1512 & ~n2413 ;
  assign n7580 = ~n2619 & n7579 ;
  assign n7581 = ~n1509 & n7580 ;
  assign n7582 = ~n7578 & ~n7581 ;
  assign n7583 = \b[14]  & n2912 ;
  assign n7584 = n2909 & n7583 ;
  assign n7585 = \b[16]  & n2620 ;
  assign n7586 = \a[21]  & \b[15]  ;
  assign n7587 = n2611 & n7586 ;
  assign n7588 = ~\a[21]  & \b[15]  ;
  assign n7589 = n2614 & n7588 ;
  assign n7590 = ~n7587 & ~n7589 ;
  assign n7591 = ~n7585 & n7590 ;
  assign n7592 = ~n7584 & n7591 ;
  assign n7593 = n7582 & n7592 ;
  assign n7594 = ~\a[23]  & ~n7593 ;
  assign n7595 = \a[23]  & n7592 ;
  assign n7596 = n7582 & n7595 ;
  assign n7597 = ~n7594 & ~n7596 ;
  assign n7598 = ~n7575 & ~n7597 ;
  assign n7599 = ~n7573 & n7598 ;
  assign n7600 = ~n7572 & n7597 ;
  assign n7601 = n7428 & n7600 ;
  assign n7602 = n7572 & n7597 ;
  assign n7603 = ~n7428 & n7602 ;
  assign n7604 = ~n7601 & ~n7603 ;
  assign n7605 = ~n7599 & n7604 ;
  assign n7606 = n1965 & ~n2079 ;
  assign n7607 = ~n2077 & n7606 ;
  assign n7608 = \b[17]  & n2218 ;
  assign n7609 = n2216 & n7608 ;
  assign n7610 = ~\a[18]  & \b[18]  ;
  assign n7611 = n1957 & n7610 ;
  assign n7612 = ~n7609 & ~n7611 ;
  assign n7613 = \b[19]  & n1963 ;
  assign n7614 = \a[18]  & \b[18]  ;
  assign n7615 = n2210 & n7614 ;
  assign n7616 = \a[20]  & ~n7615 ;
  assign n7617 = ~n7613 & n7616 ;
  assign n7618 = n7612 & n7617 ;
  assign n7619 = ~n7607 & n7618 ;
  assign n7620 = ~n7613 & ~n7615 ;
  assign n7621 = n7612 & n7620 ;
  assign n7622 = ~n7607 & n7621 ;
  assign n7623 = ~\a[20]  & ~n7622 ;
  assign n7624 = ~n7619 & ~n7623 ;
  assign n7625 = ~n7605 & ~n7624 ;
  assign n7626 = n7426 & n7625 ;
  assign n7627 = n7605 & ~n7624 ;
  assign n7628 = ~n7426 & n7627 ;
  assign n7629 = ~n7626 & ~n7628 ;
  assign n7630 = ~n7605 & n7624 ;
  assign n7631 = ~n7426 & n7630 ;
  assign n7632 = n7605 & n7624 ;
  assign n7633 = n7426 & n7632 ;
  assign n7634 = ~n7631 & ~n7633 ;
  assign n7635 = n7629 & n7634 ;
  assign n7636 = ~n7423 & n7635 ;
  assign n7637 = ~n7231 & ~n7635 ;
  assign n7638 = ~n7422 & n7637 ;
  assign n7639 = n1467 & n2768 ;
  assign n7640 = ~n2765 & n7639 ;
  assign n7641 = n1467 & n6462 ;
  assign n7642 = ~n2764 & n7641 ;
  assign n7643 = \b[20]  & n1652 ;
  assign n7644 = n1649 & n7643 ;
  assign n7645 = ~\a[15]  & \b[21]  ;
  assign n7646 = n1459 & n7645 ;
  assign n7647 = ~n7644 & ~n7646 ;
  assign n7648 = \b[22]  & n1465 ;
  assign n7649 = \a[15]  & \b[21]  ;
  assign n7650 = n1456 & n7649 ;
  assign n7651 = \a[17]  & ~n7650 ;
  assign n7652 = ~n7648 & n7651 ;
  assign n7653 = n7647 & n7652 ;
  assign n7654 = ~n7642 & n7653 ;
  assign n7655 = ~n7640 & n7654 ;
  assign n7656 = ~n7648 & ~n7650 ;
  assign n7657 = n7647 & n7656 ;
  assign n7658 = ~n7642 & n7657 ;
  assign n7659 = ~n7640 & n7658 ;
  assign n7660 = ~\a[17]  & ~n7659 ;
  assign n7661 = ~n7655 & ~n7660 ;
  assign n7662 = ~n7638 & ~n7661 ;
  assign n7663 = ~n7636 & n7662 ;
  assign n7664 = ~n7635 & n7661 ;
  assign n7665 = n7423 & n7664 ;
  assign n7666 = n7635 & n7661 ;
  assign n7667 = ~n7423 & n7666 ;
  assign n7668 = ~n7665 & ~n7667 ;
  assign n7669 = ~n7663 & n7668 ;
  assign n7670 = n999 & ~n3567 ;
  assign n7671 = ~n3565 & n7670 ;
  assign n7672 = \b[23]  & n1182 ;
  assign n7673 = n1179 & n7672 ;
  assign n7674 = ~\a[11]  & \a[13]  ;
  assign n7675 = ~\a[12]  & \b[24]  ;
  assign n7676 = n7674 & n7675 ;
  assign n7677 = ~n7673 & ~n7676 ;
  assign n7678 = \b[25]  & n997 ;
  assign n7679 = \a[12]  & \b[24]  ;
  assign n7680 = n988 & n7679 ;
  assign n7681 = \a[14]  & ~n7680 ;
  assign n7682 = ~n7678 & n7681 ;
  assign n7683 = n7677 & n7682 ;
  assign n7684 = ~n7671 & n7683 ;
  assign n7685 = ~n7678 & ~n7680 ;
  assign n7686 = n7677 & n7685 ;
  assign n7687 = ~n7671 & n7686 ;
  assign n7688 = ~\a[14]  & ~n7687 ;
  assign n7689 = ~n7684 & ~n7688 ;
  assign n7690 = ~n7669 & ~n7689 ;
  assign n7691 = n7421 & n7690 ;
  assign n7692 = n7669 & ~n7689 ;
  assign n7693 = ~n7421 & n7692 ;
  assign n7694 = ~n7691 & ~n7693 ;
  assign n7695 = ~n7669 & n7689 ;
  assign n7696 = ~n7421 & n7695 ;
  assign n7697 = n7669 & n7689 ;
  assign n7698 = n7421 & n7697 ;
  assign n7699 = ~n7696 & ~n7698 ;
  assign n7700 = n7694 & n7699 ;
  assign n7701 = n7418 & ~n7700 ;
  assign n7702 = n7395 & n7701 ;
  assign n7703 = n7418 & n7700 ;
  assign n7704 = ~n7395 & n7703 ;
  assign n7705 = ~n7702 & ~n7704 ;
  assign n7706 = ~n7395 & n7700 ;
  assign n7707 = ~n7277 & ~n7700 ;
  assign n7708 = ~n7394 & n7707 ;
  assign n7709 = ~n7418 & ~n7708 ;
  assign n7710 = ~n7706 & n7709 ;
  assign n7711 = n7705 & ~n7710 ;
  assign n7712 = n7393 & n7711 ;
  assign n7713 = ~n7393 & ~n7711 ;
  assign n7714 = ~n7712 & ~n7713 ;
  assign n7715 = n7390 & ~n7714 ;
  assign n7716 = ~n7390 & n7714 ;
  assign n7717 = ~n7715 & ~n7716 ;
  assign n7718 = n252 & n6565 ;
  assign n7719 = ~n6562 & n7718 ;
  assign n7720 = ~n5850 & ~n6565 ;
  assign n7721 = n252 & n7720 ;
  assign n7722 = ~n6561 & n7721 ;
  assign n7723 = \b[32]  & n303 ;
  assign n7724 = n300 & n7723 ;
  assign n7725 = ~\a[3]  & \b[33]  ;
  assign n7726 = n244 & n7725 ;
  assign n7727 = ~n7724 & ~n7726 ;
  assign n7728 = \b[34]  & n250 ;
  assign n7729 = \a[3]  & \b[33]  ;
  assign n7730 = n241 & n7729 ;
  assign n7731 = \a[5]  & ~n7730 ;
  assign n7732 = ~n7728 & n7731 ;
  assign n7733 = n7727 & n7732 ;
  assign n7734 = ~n7722 & n7733 ;
  assign n7735 = ~n7719 & n7734 ;
  assign n7736 = ~n7728 & ~n7730 ;
  assign n7737 = n7727 & n7736 ;
  assign n7738 = ~n7722 & n7737 ;
  assign n7739 = ~n7719 & n7738 ;
  assign n7740 = ~\a[5]  & ~n7739 ;
  assign n7741 = ~n7735 & ~n7740 ;
  assign n7742 = ~n7717 & ~n7741 ;
  assign n7743 = ~n7373 & n7742 ;
  assign n7744 = n7717 & ~n7741 ;
  assign n7745 = n7373 & n7744 ;
  assign n7746 = ~n7743 & ~n7745 ;
  assign n7747 = ~n7717 & n7741 ;
  assign n7748 = n7373 & n7747 ;
  assign n7749 = n7717 & n7741 ;
  assign n7750 = ~n7373 & n7749 ;
  assign n7751 = ~n7748 & ~n7750 ;
  assign n7752 = n7746 & n7751 ;
  assign n7753 = ~n6605 & n7337 ;
  assign n7754 = ~n7333 & n7753 ;
  assign n7755 = ~n7336 & ~n7754 ;
  assign n7756 = ~\b[36]  & ~\b[37]  ;
  assign n7757 = \b[36]  & \b[37]  ;
  assign n7758 = ~n7756 & ~n7757 ;
  assign n7759 = ~n7755 & n7758 ;
  assign n7760 = ~n7336 & ~n7758 ;
  assign n7761 = ~n7754 & n7760 ;
  assign n7762 = n134 & ~n7761 ;
  assign n7763 = ~n7759 & n7762 ;
  assign n7764 = \a[0]  & \b[37]  ;
  assign n7765 = n133 & n7764 ;
  assign n7766 = \b[36]  & n141 ;
  assign n7767 = ~\a[1]  & \b[35]  ;
  assign n7768 = n1521 & n7767 ;
  assign n7769 = ~n7766 & ~n7768 ;
  assign n7770 = ~n7765 & n7769 ;
  assign n7771 = ~n7763 & n7770 ;
  assign n7772 = ~\a[2]  & ~n7771 ;
  assign n7773 = \a[2]  & n7770 ;
  assign n7774 = ~n7763 & n7773 ;
  assign n7775 = ~n7772 & ~n7774 ;
  assign n7776 = ~n7752 & n7775 ;
  assign n7777 = ~n7371 & n7776 ;
  assign n7778 = n7752 & n7775 ;
  assign n7779 = n7371 & n7778 ;
  assign n7780 = ~n7777 & ~n7779 ;
  assign n7781 = ~n7752 & ~n7775 ;
  assign n7782 = n7371 & n7781 ;
  assign n7783 = n7752 & ~n7775 ;
  assign n7784 = ~n7371 & n7783 ;
  assign n7785 = ~n7782 & ~n7784 ;
  assign n7786 = n7780 & n7785 ;
  assign n7787 = ~n7368 & n7786 ;
  assign n7788 = ~n7358 & ~n7786 ;
  assign n7789 = ~n7365 & n7788 ;
  assign n7790 = ~n7787 & ~n7789 ;
  assign n7791 = ~n7358 & n7785 ;
  assign n7792 = ~n7365 & n7791 ;
  assign n7793 = n7780 & ~n7792 ;
  assign n7794 = n7371 & n7752 ;
  assign n7795 = n7746 & ~n7794 ;
  assign n7796 = n7316 & ~n7716 ;
  assign n7797 = ~n7372 & n7796 ;
  assign n7798 = ~n7715 & ~n7797 ;
  assign n7799 = n252 & ~n6610 ;
  assign n7800 = ~n6608 & n7799 ;
  assign n7801 = \b[35]  & n250 ;
  assign n7802 = \a[3]  & \b[34]  ;
  assign n7803 = n241 & n7802 ;
  assign n7804 = ~n7801 & ~n7803 ;
  assign n7805 = \b[33]  & n303 ;
  assign n7806 = n300 & n7805 ;
  assign n7807 = ~\a[3]  & \b[34]  ;
  assign n7808 = n244 & n7807 ;
  assign n7809 = ~n7806 & ~n7808 ;
  assign n7810 = n7804 & n7809 ;
  assign n7811 = ~n7800 & n7810 ;
  assign n7812 = ~\a[5]  & ~n7811 ;
  assign n7813 = \a[5]  & n7810 ;
  assign n7814 = ~n7800 & n7813 ;
  assign n7815 = ~n7812 & ~n7814 ;
  assign n7816 = ~n7710 & ~n7712 ;
  assign n7817 = n430 & n5810 ;
  assign n7818 = ~n5807 & n7817 ;
  assign n7819 = n430 & ~n5810 ;
  assign n7820 = ~n5457 & n7819 ;
  assign n7821 = ~n5806 & n7820 ;
  assign n7822 = \b[30]  & n486 ;
  assign n7823 = n483 & n7822 ;
  assign n7824 = ~\a[6]  & \b[31]  ;
  assign n7825 = n422 & n7824 ;
  assign n7826 = ~n7823 & ~n7825 ;
  assign n7827 = \b[32]  & n428 ;
  assign n7828 = \a[6]  & \b[31]  ;
  assign n7829 = n419 & n7828 ;
  assign n7830 = \a[8]  & ~n7829 ;
  assign n7831 = ~n7827 & n7830 ;
  assign n7832 = n7826 & n7831 ;
  assign n7833 = ~n7821 & n7832 ;
  assign n7834 = ~n7818 & n7833 ;
  assign n7835 = ~n7827 & ~n7829 ;
  assign n7836 = n7826 & n7835 ;
  assign n7837 = ~n7821 & n7836 ;
  assign n7838 = ~n7818 & n7837 ;
  assign n7839 = ~\a[8]  & ~n7838 ;
  assign n7840 = ~n7834 & ~n7839 ;
  assign n7841 = ~n7277 & n7694 ;
  assign n7842 = ~n7394 & n7841 ;
  assign n7843 = n7699 & ~n7842 ;
  assign n7844 = n646 & ~n4502 ;
  assign n7845 = ~n4500 & n7844 ;
  assign n7846 = \b[29]  & n644 ;
  assign n7847 = \a[9]  & \b[28]  ;
  assign n7848 = n635 & n7847 ;
  assign n7849 = ~n7846 & ~n7848 ;
  assign n7850 = \b[27]  & n796 ;
  assign n7851 = n793 & n7850 ;
  assign n7852 = ~\a[9]  & \b[28]  ;
  assign n7853 = n638 & n7852 ;
  assign n7854 = ~n7851 & ~n7853 ;
  assign n7855 = n7849 & n7854 ;
  assign n7856 = ~n7845 & n7855 ;
  assign n7857 = ~\a[11]  & ~n7856 ;
  assign n7858 = \a[11]  & n7855 ;
  assign n7859 = ~n7845 & n7858 ;
  assign n7860 = ~n7857 & ~n7859 ;
  assign n7861 = n7421 & n7669 ;
  assign n7862 = ~n7663 & ~n7861 ;
  assign n7863 = n999 & ~n4141 ;
  assign n7864 = ~n4518 & n7863 ;
  assign n7865 = \b[24]  & n1182 ;
  assign n7866 = n1179 & n7865 ;
  assign n7867 = ~\a[12]  & \b[25]  ;
  assign n7868 = n7674 & n7867 ;
  assign n7869 = ~n7866 & ~n7868 ;
  assign n7870 = \b[26]  & n997 ;
  assign n7871 = \a[12]  & \b[25]  ;
  assign n7872 = n988 & n7871 ;
  assign n7873 = \a[14]  & ~n7872 ;
  assign n7874 = ~n7870 & n7873 ;
  assign n7875 = n7869 & n7874 ;
  assign n7876 = ~n7864 & n7875 ;
  assign n7877 = ~n7870 & ~n7872 ;
  assign n7878 = n7869 & n7877 ;
  assign n7879 = ~n7864 & n7878 ;
  assign n7880 = ~\a[14]  & ~n7879 ;
  assign n7881 = ~n7876 & ~n7880 ;
  assign n7882 = ~n7231 & n7629 ;
  assign n7883 = ~n7422 & n7882 ;
  assign n7884 = n7634 & ~n7883 ;
  assign n7885 = n7426 & n7605 ;
  assign n7886 = ~n7599 & ~n7885 ;
  assign n7887 = ~n7174 & n7571 ;
  assign n7888 = ~n7427 & n7887 ;
  assign n7889 = n7566 & ~n7888 ;
  assign n7890 = n7431 & n7561 ;
  assign n7891 = n7560 & ~n7890 ;
  assign n7892 = n1087 & n3402 ;
  assign n7893 = ~n1084 & n7892 ;
  assign n7894 = n1552 & n3402 ;
  assign n7895 = ~n1083 & n7894 ;
  assign n7896 = \b[12]  & n3733 ;
  assign n7897 = n3730 & n7896 ;
  assign n7898 = \b[14]  & n3400 ;
  assign n7899 = \a[24]  & \b[13]  ;
  assign n7900 = n3391 & n7899 ;
  assign n7901 = ~\a[24]  & \b[13]  ;
  assign n7902 = n3394 & n7901 ;
  assign n7903 = ~n7900 & ~n7902 ;
  assign n7904 = ~n7898 & n7903 ;
  assign n7905 = ~n7897 & n7904 ;
  assign n7906 = ~n7895 & n7905 ;
  assign n7907 = ~n7893 & n7906 ;
  assign n7908 = ~\a[26]  & ~n7907 ;
  assign n7909 = \a[26]  & n7905 ;
  assign n7910 = ~n7895 & n7909 ;
  assign n7911 = ~n7893 & n7910 ;
  assign n7912 = ~n7908 & ~n7911 ;
  assign n7913 = ~n728 & n4249 ;
  assign n7914 = ~n726 & n7913 ;
  assign n7915 = \b[9]  & n4647 ;
  assign n7916 = n4644 & n7915 ;
  assign n7917 = ~\a[26]  & \b[10]  ;
  assign n7918 = n4646 & n7917 ;
  assign n7919 = ~n7916 & ~n7918 ;
  assign n7920 = \b[11]  & n4247 ;
  assign n7921 = \a[27]  & \b[10]  ;
  assign n7922 = n4238 & n7921 ;
  assign n7923 = \a[29]  & ~n7922 ;
  assign n7924 = ~n7920 & n7923 ;
  assign n7925 = n7919 & n7924 ;
  assign n7926 = ~n7914 & n7925 ;
  assign n7927 = ~n7920 & ~n7922 ;
  assign n7928 = n7919 & n7927 ;
  assign n7929 = ~n7914 & n7928 ;
  assign n7930 = ~\a[29]  & ~n7929 ;
  assign n7931 = ~n7926 & ~n7930 ;
  assign n7932 = ~n7129 & ~n7549 ;
  assign n7933 = ~n7454 & n7932 ;
  assign n7934 = ~n7548 & ~n7933 ;
  assign n7935 = ~n7543 & ~n7545 ;
  assign n7936 = ~n270 & n6309 ;
  assign n7937 = ~n218 & n6309 ;
  assign n7938 = ~n220 & n7937 ;
  assign n7939 = ~n7936 & ~n7938 ;
  assign n7940 = ~n273 & ~n7939 ;
  assign n7941 = \b[3]  & n6778 ;
  assign n7942 = n6775 & n7941 ;
  assign n7943 = \b[5]  & n6307 ;
  assign n7944 = \a[32]  & \b[4]  ;
  assign n7945 = n6776 & n7944 ;
  assign n7946 = ~\a[33]  & \b[4]  ;
  assign n7947 = n6301 & n7946 ;
  assign n7948 = ~n7945 & ~n7947 ;
  assign n7949 = ~n7943 & n7948 ;
  assign n7950 = ~n7942 & n7949 ;
  assign n7951 = ~\a[35]  & n7950 ;
  assign n7952 = ~n7940 & n7951 ;
  assign n7953 = \a[35]  & ~n7950 ;
  assign n7954 = \a[35]  & ~n273 ;
  assign n7955 = ~n7939 & n7954 ;
  assign n7956 = ~n7953 & ~n7955 ;
  assign n7957 = ~n7952 & n7956 ;
  assign n7958 = \a[38]  & ~n7099 ;
  assign n7959 = n7528 & n7958 ;
  assign n7960 = n7536 & n7959 ;
  assign n7961 = \a[38]  & ~n7960 ;
  assign n7962 = \b[2]  & n7532 ;
  assign n7963 = ~\a[36]  & \b[1]  ;
  assign n7964 = n7526 & n7963 ;
  assign n7965 = \a[36]  & \b[1]  ;
  assign n7966 = n7523 & n7965 ;
  assign n7967 = ~n7964 & ~n7966 ;
  assign n7968 = ~n7962 & n7967 ;
  assign n7969 = n157 & n7534 ;
  assign n7970 = n7098 & ~n7531 ;
  assign n7971 = \a[36]  & ~\a[37]  ;
  assign n7972 = ~\a[36]  & \a[37]  ;
  assign n7973 = ~n7971 & ~n7972 ;
  assign n7974 = \b[0]  & n7973 ;
  assign n7975 = n7970 & n7974 ;
  assign n7976 = ~n7969 & ~n7975 ;
  assign n7977 = n7968 & n7976 ;
  assign n7978 = ~n7961 & ~n7977 ;
  assign n7979 = n7961 & n7977 ;
  assign n7980 = ~n7978 & ~n7979 ;
  assign n7981 = n7957 & ~n7980 ;
  assign n7982 = ~n7957 & n7980 ;
  assign n7983 = ~n7981 & ~n7982 ;
  assign n7984 = ~n7935 & n7983 ;
  assign n7985 = ~n505 & ~n4909 ;
  assign n7986 = ~n5208 & n7985 ;
  assign n7987 = n502 & n7986 ;
  assign n7988 = n505 & ~n4909 ;
  assign n7989 = ~n5208 & n7988 ;
  assign n7990 = ~n502 & n7989 ;
  assign n7991 = ~n7987 & ~n7990 ;
  assign n7992 = \b[6]  & n5595 ;
  assign n7993 = n5592 & n7992 ;
  assign n7994 = \b[8]  & n5209 ;
  assign n7995 = \a[29]  & \b[7]  ;
  assign n7996 = n5593 & n7995 ;
  assign n7997 = ~\a[30]  & \b[7]  ;
  assign n7998 = n5203 & n7997 ;
  assign n7999 = ~n7996 & ~n7998 ;
  assign n8000 = ~n7994 & n7999 ;
  assign n8001 = ~n7993 & n8000 ;
  assign n8002 = n7991 & n8001 ;
  assign n8003 = ~\a[32]  & ~n8002 ;
  assign n8004 = \a[32]  & n8001 ;
  assign n8005 = n7991 & n8004 ;
  assign n8006 = ~n8003 & ~n8005 ;
  assign n8007 = ~n7543 & ~n7983 ;
  assign n8008 = ~n7545 & n8007 ;
  assign n8009 = ~n8006 & ~n8008 ;
  assign n8010 = ~n7984 & n8009 ;
  assign n8011 = ~n7984 & ~n8008 ;
  assign n8012 = n8006 & ~n8011 ;
  assign n8013 = ~n8010 & ~n8012 ;
  assign n8014 = n7934 & n8013 ;
  assign n8015 = ~n7934 & ~n8013 ;
  assign n8016 = ~n8014 & ~n8015 ;
  assign n8017 = ~n7931 & n8016 ;
  assign n8018 = n7931 & ~n8016 ;
  assign n8019 = ~n8017 & ~n8018 ;
  assign n8020 = n7912 & ~n8019 ;
  assign n8021 = n7891 & n8020 ;
  assign n8022 = n7912 & n8019 ;
  assign n8023 = ~n7891 & n8022 ;
  assign n8024 = ~n8021 & ~n8023 ;
  assign n8025 = ~n7912 & ~n8019 ;
  assign n8026 = ~n7891 & n8025 ;
  assign n8027 = ~n7912 & n8019 ;
  assign n8028 = n7891 & n8027 ;
  assign n8029 = ~n8026 & ~n8028 ;
  assign n8030 = n8024 & n8029 ;
  assign n8031 = ~n1694 & n2622 ;
  assign n8032 = ~n1692 & n8031 ;
  assign n8033 = \b[15]  & n2912 ;
  assign n8034 = n2909 & n8033 ;
  assign n8035 = \b[17]  & n2620 ;
  assign n8036 = \a[21]  & \b[16]  ;
  assign n8037 = n2611 & n8036 ;
  assign n8038 = ~\a[21]  & \b[16]  ;
  assign n8039 = n2614 & n8038 ;
  assign n8040 = ~n8037 & ~n8039 ;
  assign n8041 = ~n8035 & n8040 ;
  assign n8042 = ~n8034 & n8041 ;
  assign n8043 = ~\a[23]  & n8042 ;
  assign n8044 = ~n8032 & n8043 ;
  assign n8045 = ~n8032 & n8042 ;
  assign n8046 = \a[23]  & ~n8045 ;
  assign n8047 = ~n8044 & ~n8046 ;
  assign n8048 = ~n8030 & n8047 ;
  assign n8049 = n7889 & n8048 ;
  assign n8050 = n8030 & n8047 ;
  assign n8051 = ~n7889 & n8050 ;
  assign n8052 = ~n8049 & ~n8051 ;
  assign n8053 = ~n8030 & ~n8047 ;
  assign n8054 = ~n7889 & n8053 ;
  assign n8055 = n8030 & ~n8047 ;
  assign n8056 = n7889 & n8055 ;
  assign n8057 = ~n8054 & ~n8056 ;
  assign n8058 = n8052 & n8057 ;
  assign n8059 = ~n7886 & n8058 ;
  assign n8060 = ~n7599 & ~n8058 ;
  assign n8061 = ~n7885 & n8060 ;
  assign n8062 = n1965 & n2293 ;
  assign n8063 = ~n2290 & n8062 ;
  assign n8064 = n1965 & n5705 ;
  assign n8065 = ~n2289 & n8064 ;
  assign n8066 = \b[18]  & n2218 ;
  assign n8067 = n2216 & n8066 ;
  assign n8068 = ~\a[18]  & \b[19]  ;
  assign n8069 = n1957 & n8068 ;
  assign n8070 = ~n8067 & ~n8069 ;
  assign n8071 = \b[20]  & n1963 ;
  assign n8072 = \a[18]  & \b[19]  ;
  assign n8073 = n2210 & n8072 ;
  assign n8074 = \a[20]  & ~n8073 ;
  assign n8075 = ~n8071 & n8074 ;
  assign n8076 = n8070 & n8075 ;
  assign n8077 = ~n8065 & n8076 ;
  assign n8078 = ~n8063 & n8077 ;
  assign n8079 = ~n8071 & ~n8073 ;
  assign n8080 = n8070 & n8079 ;
  assign n8081 = ~n8065 & n8080 ;
  assign n8082 = ~n8063 & n8081 ;
  assign n8083 = ~\a[20]  & ~n8082 ;
  assign n8084 = ~n8078 & ~n8083 ;
  assign n8085 = ~n8061 & ~n8084 ;
  assign n8086 = ~n8059 & n8085 ;
  assign n8087 = ~n8058 & n8084 ;
  assign n8088 = n7886 & n8087 ;
  assign n8089 = n8058 & n8084 ;
  assign n8090 = ~n7886 & n8089 ;
  assign n8091 = ~n8088 & ~n8090 ;
  assign n8092 = ~n8086 & n8091 ;
  assign n8093 = n1467 & ~n3022 ;
  assign n8094 = ~n3020 & n8093 ;
  assign n8095 = \b[21]  & n1652 ;
  assign n8096 = n1649 & n8095 ;
  assign n8097 = ~\a[15]  & \b[22]  ;
  assign n8098 = n1459 & n8097 ;
  assign n8099 = ~n8096 & ~n8098 ;
  assign n8100 = \b[23]  & n1465 ;
  assign n8101 = \a[15]  & \b[22]  ;
  assign n8102 = n1456 & n8101 ;
  assign n8103 = \a[17]  & ~n8102 ;
  assign n8104 = ~n8100 & n8103 ;
  assign n8105 = n8099 & n8104 ;
  assign n8106 = ~n8094 & n8105 ;
  assign n8107 = ~n8100 & ~n8102 ;
  assign n8108 = n8099 & n8107 ;
  assign n8109 = ~n8094 & n8108 ;
  assign n8110 = ~\a[17]  & ~n8109 ;
  assign n8111 = ~n8106 & ~n8110 ;
  assign n8112 = ~n8092 & ~n8111 ;
  assign n8113 = n7884 & n8112 ;
  assign n8114 = n8092 & ~n8111 ;
  assign n8115 = ~n7884 & n8114 ;
  assign n8116 = ~n8113 & ~n8115 ;
  assign n8117 = ~n8092 & n8111 ;
  assign n8118 = ~n7884 & n8117 ;
  assign n8119 = n8092 & n8111 ;
  assign n8120 = n7884 & n8119 ;
  assign n8121 = ~n8118 & ~n8120 ;
  assign n8122 = n8116 & n8121 ;
  assign n8123 = n7881 & ~n8122 ;
  assign n8124 = n7862 & n8123 ;
  assign n8125 = n7881 & n8122 ;
  assign n8126 = ~n7862 & n8125 ;
  assign n8127 = ~n8124 & ~n8126 ;
  assign n8128 = ~n7862 & n8122 ;
  assign n8129 = ~n7663 & ~n8122 ;
  assign n8130 = ~n7861 & n8129 ;
  assign n8131 = ~n7881 & ~n8130 ;
  assign n8132 = ~n8128 & n8131 ;
  assign n8133 = n8127 & ~n8132 ;
  assign n8134 = n7860 & ~n8133 ;
  assign n8135 = ~n7843 & n8134 ;
  assign n8136 = n7860 & n8133 ;
  assign n8137 = n7843 & n8136 ;
  assign n8138 = ~n8135 & ~n8137 ;
  assign n8139 = ~n7860 & ~n8133 ;
  assign n8140 = n7843 & n8139 ;
  assign n8141 = ~n7860 & n8133 ;
  assign n8142 = ~n7843 & n8141 ;
  assign n8143 = ~n8140 & ~n8142 ;
  assign n8144 = n8138 & n8143 ;
  assign n8145 = n7840 & ~n8144 ;
  assign n8146 = n7816 & n8145 ;
  assign n8147 = n7840 & n8144 ;
  assign n8148 = ~n7816 & n8147 ;
  assign n8149 = ~n8146 & ~n8148 ;
  assign n8150 = ~n7840 & ~n8144 ;
  assign n8151 = ~n7816 & n8150 ;
  assign n8152 = ~n7840 & n8144 ;
  assign n8153 = n7816 & n8152 ;
  assign n8154 = ~n8151 & ~n8153 ;
  assign n8155 = n8149 & n8154 ;
  assign n8156 = n7815 & ~n8155 ;
  assign n8157 = ~n7798 & n8156 ;
  assign n8158 = n7815 & n8155 ;
  assign n8159 = n7798 & n8158 ;
  assign n8160 = ~n8157 & ~n8159 ;
  assign n8161 = ~n7815 & ~n8155 ;
  assign n8162 = n7798 & n8161 ;
  assign n8163 = ~n7815 & n8155 ;
  assign n8164 = ~n7798 & n8163 ;
  assign n8165 = ~n8162 & ~n8164 ;
  assign n8166 = n8160 & n8165 ;
  assign n8167 = ~n7795 & n8166 ;
  assign n8168 = n7746 & ~n8166 ;
  assign n8169 = ~n7794 & n8168 ;
  assign n8170 = ~n7336 & ~n7757 ;
  assign n8171 = ~n7754 & n8170 ;
  assign n8172 = ~n7756 & ~n8171 ;
  assign n8173 = ~\b[37]  & ~\b[38]  ;
  assign n8174 = \b[37]  & \b[38]  ;
  assign n8175 = ~n8173 & ~n8174 ;
  assign n8176 = n134 & n8175 ;
  assign n8177 = ~n8172 & n8176 ;
  assign n8178 = n134 & ~n8175 ;
  assign n8179 = ~n7756 & n8178 ;
  assign n8180 = ~n8171 & n8179 ;
  assign n8181 = \a[0]  & \b[38]  ;
  assign n8182 = n133 & n8181 ;
  assign n8183 = \b[37]  & n141 ;
  assign n8184 = ~\a[1]  & \b[36]  ;
  assign n8185 = n1521 & n8184 ;
  assign n8186 = ~n8183 & ~n8185 ;
  assign n8187 = ~n8182 & n8186 ;
  assign n8188 = \a[2]  & n8187 ;
  assign n8189 = ~n8180 & n8188 ;
  assign n8190 = ~n8177 & n8189 ;
  assign n8191 = ~n8180 & n8187 ;
  assign n8192 = ~n8177 & n8191 ;
  assign n8193 = ~\a[2]  & ~n8192 ;
  assign n8194 = ~n8190 & ~n8193 ;
  assign n8195 = ~n8169 & ~n8194 ;
  assign n8196 = ~n8167 & n8195 ;
  assign n8197 = ~n8166 & n8194 ;
  assign n8198 = n7795 & n8197 ;
  assign n8199 = n8166 & n8194 ;
  assign n8200 = ~n7795 & n8199 ;
  assign n8201 = ~n8198 & ~n8200 ;
  assign n8202 = ~n8196 & n8201 ;
  assign n8203 = n7793 & n8202 ;
  assign n8204 = ~n7793 & ~n8202 ;
  assign n8205 = ~n8203 & ~n8204 ;
  assign n8206 = ~n8196 & ~n8203 ;
  assign n8207 = n7746 & n8165 ;
  assign n8208 = ~n7794 & n8207 ;
  assign n8209 = n8160 & ~n8208 ;
  assign n8210 = n7798 & n8155 ;
  assign n8211 = n8154 & ~n8210 ;
  assign n8212 = ~n7334 & ~n7337 ;
  assign n8213 = n252 & ~n7754 ;
  assign n8214 = ~n8212 & n8213 ;
  assign n8215 = \b[34]  & n303 ;
  assign n8216 = n300 & n8215 ;
  assign n8217 = ~\a[3]  & \b[35]  ;
  assign n8218 = n244 & n8217 ;
  assign n8219 = ~n8216 & ~n8218 ;
  assign n8220 = \b[36]  & n250 ;
  assign n8221 = \a[3]  & \b[35]  ;
  assign n8222 = n241 & n8221 ;
  assign n8223 = \a[5]  & ~n8222 ;
  assign n8224 = ~n8220 & n8223 ;
  assign n8225 = n8219 & n8224 ;
  assign n8226 = ~n8214 & n8225 ;
  assign n8227 = ~n8220 & ~n8222 ;
  assign n8228 = n8219 & n8227 ;
  assign n8229 = ~n8214 & n8228 ;
  assign n8230 = ~\a[5]  & ~n8229 ;
  assign n8231 = ~n8226 & ~n8230 ;
  assign n8232 = ~n7710 & n8143 ;
  assign n8233 = ~n7712 & n8232 ;
  assign n8234 = n8138 & ~n8233 ;
  assign n8235 = n7843 & n8133 ;
  assign n8236 = ~n8132 & ~n8235 ;
  assign n8237 = ~n7663 & n8116 ;
  assign n8238 = ~n7861 & n8237 ;
  assign n8239 = n8121 & ~n8238 ;
  assign n8240 = n7884 & n8092 ;
  assign n8241 = ~n8086 & ~n8240 ;
  assign n8242 = ~n7599 & n8052 ;
  assign n8243 = ~n7885 & n8242 ;
  assign n8244 = n8057 & ~n8243 ;
  assign n8245 = n7889 & n8030 ;
  assign n8246 = n8029 & ~n8245 ;
  assign n8247 = n7560 & ~n8017 ;
  assign n8248 = ~n7890 & n8247 ;
  assign n8249 = ~n8018 & ~n8248 ;
  assign n8250 = ~n8010 & ~n8014 ;
  assign n8251 = ~n7543 & ~n7981 ;
  assign n8252 = ~n7545 & n8251 ;
  assign n8253 = ~n7982 & ~n8252 ;
  assign n8254 = n177 & n7534 ;
  assign n8255 = \b[3]  & n7532 ;
  assign n8256 = \a[35]  & \b[2]  ;
  assign n8257 = n7971 & n8256 ;
  assign n8258 = ~\a[36]  & \b[2]  ;
  assign n8259 = n7526 & n8258 ;
  assign n8260 = ~n8257 & ~n8259 ;
  assign n8261 = ~n8255 & n8260 ;
  assign n8262 = ~n8254 & n8261 ;
  assign n8263 = \b[1]  & n7973 ;
  assign n8264 = n7970 & n8263 ;
  assign n8265 = ~\a[38]  & ~n8264 ;
  assign n8266 = n8262 & n8265 ;
  assign n8267 = n8262 & ~n8264 ;
  assign n8268 = \a[38]  & ~n8267 ;
  assign n8269 = ~n8266 & ~n8268 ;
  assign n8270 = \a[38]  & ~\a[39]  ;
  assign n8271 = ~\a[38]  & \a[39]  ;
  assign n8272 = ~n8270 & ~n8271 ;
  assign n8273 = \b[0]  & ~n8272 ;
  assign n8274 = n7960 & n7977 ;
  assign n8275 = n8273 & n8274 ;
  assign n8276 = ~n8273 & ~n8274 ;
  assign n8277 = ~n8275 & ~n8276 ;
  assign n8278 = n8269 & n8277 ;
  assign n8279 = ~n8269 & ~n8277 ;
  assign n8280 = ~n8278 & ~n8279 ;
  assign n8281 = ~n323 & ~n5952 ;
  assign n8282 = ~n6306 & n8281 ;
  assign n8283 = n320 & n8282 ;
  assign n8284 = n323 & ~n5952 ;
  assign n8285 = ~n6306 & n8284 ;
  assign n8286 = ~n320 & n8285 ;
  assign n8287 = ~n8283 & ~n8286 ;
  assign n8288 = \b[4]  & n6778 ;
  assign n8289 = n6775 & n8288 ;
  assign n8290 = \b[6]  & n6307 ;
  assign n8291 = \a[32]  & \b[5]  ;
  assign n8292 = n6776 & n8291 ;
  assign n8293 = ~\a[33]  & \b[5]  ;
  assign n8294 = n6301 & n8293 ;
  assign n8295 = ~n8292 & ~n8294 ;
  assign n8296 = ~n8290 & n8295 ;
  assign n8297 = ~n8289 & n8296 ;
  assign n8298 = n8287 & n8297 ;
  assign n8299 = ~\a[35]  & ~n8298 ;
  assign n8300 = \a[35]  & n8297 ;
  assign n8301 = n8287 & n8300 ;
  assign n8302 = ~n8299 & ~n8301 ;
  assign n8303 = n8280 & ~n8302 ;
  assign n8304 = ~n8280 & n8302 ;
  assign n8305 = ~n8303 & ~n8304 ;
  assign n8306 = ~n586 & n5211 ;
  assign n8307 = ~n504 & n5211 ;
  assign n8308 = ~n508 & n8307 ;
  assign n8309 = ~n8306 & ~n8308 ;
  assign n8310 = ~n589 & ~n8309 ;
  assign n8311 = \b[7]  & n5595 ;
  assign n8312 = n5592 & n8311 ;
  assign n8313 = \b[9]  & n5209 ;
  assign n8314 = \a[29]  & \b[8]  ;
  assign n8315 = n5593 & n8314 ;
  assign n8316 = ~\a[30]  & \b[8]  ;
  assign n8317 = n5203 & n8316 ;
  assign n8318 = ~n8315 & ~n8317 ;
  assign n8319 = ~n8313 & n8318 ;
  assign n8320 = ~n8312 & n8319 ;
  assign n8321 = ~\a[32]  & n8320 ;
  assign n8322 = ~n8310 & n8321 ;
  assign n8323 = \a[32]  & ~n8320 ;
  assign n8324 = \a[32]  & ~n589 ;
  assign n8325 = ~n8309 & n8324 ;
  assign n8326 = ~n8323 & ~n8325 ;
  assign n8327 = ~n8322 & n8326 ;
  assign n8328 = ~n8305 & n8327 ;
  assign n8329 = n8253 & n8328 ;
  assign n8330 = n8305 & n8327 ;
  assign n8331 = ~n8253 & n8330 ;
  assign n8332 = ~n8329 & ~n8331 ;
  assign n8333 = ~n8305 & ~n8327 ;
  assign n8334 = ~n8253 & n8333 ;
  assign n8335 = n8305 & ~n8327 ;
  assign n8336 = n8253 & n8335 ;
  assign n8337 = ~n8334 & ~n8336 ;
  assign n8338 = n8332 & n8337 ;
  assign n8339 = ~n909 & ~n3956 ;
  assign n8340 = ~n4246 & n8339 ;
  assign n8341 = n906 & n8340 ;
  assign n8342 = n909 & ~n3956 ;
  assign n8343 = ~n4246 & n8342 ;
  assign n8344 = ~n906 & n8343 ;
  assign n8345 = ~n8341 & ~n8344 ;
  assign n8346 = \b[10]  & n4647 ;
  assign n8347 = n4644 & n8346 ;
  assign n8348 = ~\a[26]  & \b[11]  ;
  assign n8349 = n4646 & n8348 ;
  assign n8350 = ~n8347 & ~n8349 ;
  assign n8351 = \b[12]  & n4247 ;
  assign n8352 = \a[27]  & \b[11]  ;
  assign n8353 = n4238 & n8352 ;
  assign n8354 = \a[29]  & ~n8353 ;
  assign n8355 = ~n8351 & n8354 ;
  assign n8356 = n8350 & n8355 ;
  assign n8357 = n8345 & n8356 ;
  assign n8358 = ~n8351 & ~n8353 ;
  assign n8359 = n8350 & n8358 ;
  assign n8360 = n8345 & n8359 ;
  assign n8361 = ~\a[29]  & ~n8360 ;
  assign n8362 = ~n8357 & ~n8361 ;
  assign n8363 = ~n8338 & n8362 ;
  assign n8364 = n8250 & n8363 ;
  assign n8365 = n8338 & n8362 ;
  assign n8366 = ~n8250 & n8365 ;
  assign n8367 = ~n8364 & ~n8366 ;
  assign n8368 = ~n8250 & n8338 ;
  assign n8369 = ~n8010 & ~n8338 ;
  assign n8370 = ~n8014 & n8369 ;
  assign n8371 = ~n8362 & ~n8370 ;
  assign n8372 = ~n8368 & n8371 ;
  assign n8373 = n8367 & ~n8372 ;
  assign n8374 = ~n1233 & n3402 ;
  assign n8375 = ~n1231 & n8374 ;
  assign n8376 = \b[13]  & n3733 ;
  assign n8377 = n3730 & n8376 ;
  assign n8378 = \b[15]  & n3400 ;
  assign n8379 = \a[24]  & \b[14]  ;
  assign n8380 = n3391 & n8379 ;
  assign n8381 = ~\a[24]  & \b[14]  ;
  assign n8382 = n3394 & n8381 ;
  assign n8383 = ~n8380 & ~n8382 ;
  assign n8384 = ~n8378 & n8383 ;
  assign n8385 = ~n8377 & n8384 ;
  assign n8386 = ~\a[26]  & n8385 ;
  assign n8387 = ~n8375 & n8386 ;
  assign n8388 = ~n8375 & n8385 ;
  assign n8389 = \a[26]  & ~n8388 ;
  assign n8390 = ~n8387 & ~n8389 ;
  assign n8391 = n8373 & n8390 ;
  assign n8392 = ~n8249 & n8391 ;
  assign n8393 = ~n8373 & n8390 ;
  assign n8394 = n8249 & n8393 ;
  assign n8395 = ~n8392 & ~n8394 ;
  assign n8396 = ~n8373 & ~n8390 ;
  assign n8397 = ~n8249 & n8396 ;
  assign n8398 = n8373 & ~n8390 ;
  assign n8399 = n8249 & n8398 ;
  assign n8400 = ~n8397 & ~n8399 ;
  assign n8401 = n8395 & n8400 ;
  assign n8402 = ~n8246 & n8401 ;
  assign n8403 = n1875 & n2622 ;
  assign n8404 = ~n1872 & n8403 ;
  assign n8405 = n2622 & n5000 ;
  assign n8406 = ~n1871 & n8405 ;
  assign n8407 = \b[16]  & n2912 ;
  assign n8408 = n2909 & n8407 ;
  assign n8409 = ~\a[21]  & \b[17]  ;
  assign n8410 = n2614 & n8409 ;
  assign n8411 = ~n8408 & ~n8410 ;
  assign n8412 = \b[18]  & n2620 ;
  assign n8413 = \a[21]  & \b[17]  ;
  assign n8414 = n2611 & n8413 ;
  assign n8415 = \a[23]  & ~n8414 ;
  assign n8416 = ~n8412 & n8415 ;
  assign n8417 = n8411 & n8416 ;
  assign n8418 = ~n8406 & n8417 ;
  assign n8419 = ~n8404 & n8418 ;
  assign n8420 = ~n8412 & ~n8414 ;
  assign n8421 = n8411 & n8420 ;
  assign n8422 = ~n8406 & n8421 ;
  assign n8423 = ~n8404 & n8422 ;
  assign n8424 = ~\a[23]  & ~n8423 ;
  assign n8425 = ~n8419 & ~n8424 ;
  assign n8426 = n8029 & ~n8401 ;
  assign n8427 = ~n8245 & n8426 ;
  assign n8428 = ~n8425 & ~n8427 ;
  assign n8429 = ~n8402 & n8428 ;
  assign n8430 = ~n8401 & n8425 ;
  assign n8431 = n8246 & n8430 ;
  assign n8432 = n8401 & n8425 ;
  assign n8433 = ~n8246 & n8432 ;
  assign n8434 = ~n8431 & ~n8433 ;
  assign n8435 = ~n8429 & n8434 ;
  assign n8436 = n1965 & ~n2523 ;
  assign n8437 = ~n2521 & n8436 ;
  assign n8438 = \b[19]  & n2218 ;
  assign n8439 = n2216 & n8438 ;
  assign n8440 = ~\a[18]  & \b[20]  ;
  assign n8441 = n1957 & n8440 ;
  assign n8442 = ~n8439 & ~n8441 ;
  assign n8443 = \b[21]  & n1963 ;
  assign n8444 = \a[18]  & \b[20]  ;
  assign n8445 = n2210 & n8444 ;
  assign n8446 = \a[20]  & ~n8445 ;
  assign n8447 = ~n8443 & n8446 ;
  assign n8448 = n8442 & n8447 ;
  assign n8449 = ~n8437 & n8448 ;
  assign n8450 = ~n8443 & ~n8445 ;
  assign n8451 = n8442 & n8450 ;
  assign n8452 = ~n8437 & n8451 ;
  assign n8453 = ~\a[20]  & ~n8452 ;
  assign n8454 = ~n8449 & ~n8453 ;
  assign n8455 = ~n8435 & ~n8454 ;
  assign n8456 = n8244 & n8455 ;
  assign n8457 = n8435 & ~n8454 ;
  assign n8458 = ~n8244 & n8457 ;
  assign n8459 = ~n8456 & ~n8458 ;
  assign n8460 = ~n8435 & n8454 ;
  assign n8461 = ~n8244 & n8460 ;
  assign n8462 = n8435 & n8454 ;
  assign n8463 = n8244 & n8462 ;
  assign n8464 = ~n8461 & ~n8463 ;
  assign n8465 = n8459 & n8464 ;
  assign n8466 = n1467 & n3283 ;
  assign n8467 = ~n3280 & n8466 ;
  assign n8468 = n1467 & n4107 ;
  assign n8469 = ~n3279 & n8468 ;
  assign n8470 = \b[22]  & n1652 ;
  assign n8471 = n1649 & n8470 ;
  assign n8472 = ~\a[15]  & \b[23]  ;
  assign n8473 = n1459 & n8472 ;
  assign n8474 = ~n8471 & ~n8473 ;
  assign n8475 = \b[24]  & n1465 ;
  assign n8476 = \a[15]  & \b[23]  ;
  assign n8477 = n1456 & n8476 ;
  assign n8478 = \a[17]  & ~n8477 ;
  assign n8479 = ~n8475 & n8478 ;
  assign n8480 = n8474 & n8479 ;
  assign n8481 = ~n8469 & n8480 ;
  assign n8482 = ~n8467 & n8481 ;
  assign n8483 = ~n8475 & ~n8477 ;
  assign n8484 = n8474 & n8483 ;
  assign n8485 = ~n8469 & n8484 ;
  assign n8486 = ~n8467 & n8485 ;
  assign n8487 = ~\a[17]  & ~n8486 ;
  assign n8488 = ~n8482 & ~n8487 ;
  assign n8489 = ~n8465 & n8488 ;
  assign n8490 = n8241 & n8489 ;
  assign n8491 = n8465 & n8488 ;
  assign n8492 = ~n8241 & n8491 ;
  assign n8493 = ~n8490 & ~n8492 ;
  assign n8494 = ~n8241 & n8465 ;
  assign n8495 = ~n8086 & ~n8465 ;
  assign n8496 = ~n8240 & n8495 ;
  assign n8497 = ~n8488 & ~n8496 ;
  assign n8498 = ~n8494 & n8497 ;
  assign n8499 = n8493 & ~n8498 ;
  assign n8500 = n999 & ~n4148 ;
  assign n8501 = ~n4146 & n8500 ;
  assign n8502 = \b[25]  & n1182 ;
  assign n8503 = n1179 & n8502 ;
  assign n8504 = ~\a[12]  & \b[26]  ;
  assign n8505 = n7674 & n8504 ;
  assign n8506 = ~n8503 & ~n8505 ;
  assign n8507 = \b[27]  & n997 ;
  assign n8508 = \a[12]  & \b[26]  ;
  assign n8509 = n988 & n8508 ;
  assign n8510 = \a[14]  & ~n8509 ;
  assign n8511 = ~n8507 & n8510 ;
  assign n8512 = n8506 & n8511 ;
  assign n8513 = ~n8501 & n8512 ;
  assign n8514 = ~n8507 & ~n8509 ;
  assign n8515 = n8506 & n8514 ;
  assign n8516 = ~n8501 & n8515 ;
  assign n8517 = ~\a[14]  & ~n8516 ;
  assign n8518 = ~n8513 & ~n8517 ;
  assign n8519 = ~n8499 & ~n8518 ;
  assign n8520 = n8239 & n8519 ;
  assign n8521 = n8499 & ~n8518 ;
  assign n8522 = ~n8239 & n8521 ;
  assign n8523 = ~n8520 & ~n8522 ;
  assign n8524 = ~n8499 & n8518 ;
  assign n8525 = ~n8239 & n8524 ;
  assign n8526 = n8499 & n8518 ;
  assign n8527 = n8239 & n8526 ;
  assign n8528 = ~n8525 & ~n8527 ;
  assign n8529 = n8523 & n8528 ;
  assign n8530 = ~n8236 & n8529 ;
  assign n8531 = n646 & ~n5455 ;
  assign n8532 = ~n6160 & n8531 ;
  assign n8533 = \b[28]  & n796 ;
  assign n8534 = n793 & n8533 ;
  assign n8535 = ~\a[9]  & \b[29]  ;
  assign n8536 = n638 & n8535 ;
  assign n8537 = ~n8534 & ~n8536 ;
  assign n8538 = \b[30]  & n644 ;
  assign n8539 = \a[9]  & \b[29]  ;
  assign n8540 = n635 & n8539 ;
  assign n8541 = \a[11]  & ~n8540 ;
  assign n8542 = ~n8538 & n8541 ;
  assign n8543 = n8537 & n8542 ;
  assign n8544 = ~n8532 & n8543 ;
  assign n8545 = ~n8538 & ~n8540 ;
  assign n8546 = n8537 & n8545 ;
  assign n8547 = ~n8532 & n8546 ;
  assign n8548 = ~\a[11]  & ~n8547 ;
  assign n8549 = ~n8544 & ~n8548 ;
  assign n8550 = ~n8132 & ~n8529 ;
  assign n8551 = ~n8235 & n8550 ;
  assign n8552 = ~n8549 & ~n8551 ;
  assign n8553 = ~n8530 & n8552 ;
  assign n8554 = ~n8529 & n8549 ;
  assign n8555 = n8236 & n8554 ;
  assign n8556 = n8529 & n8549 ;
  assign n8557 = ~n8236 & n8556 ;
  assign n8558 = ~n8555 & ~n8557 ;
  assign n8559 = ~n8553 & n8558 ;
  assign n8560 = n8234 & n8559 ;
  assign n8561 = ~n8234 & ~n8559 ;
  assign n8562 = ~n8560 & ~n8561 ;
  assign n8563 = n430 & ~n5855 ;
  assign n8564 = ~n5853 & n8563 ;
  assign n8565 = \b[33]  & n428 ;
  assign n8566 = \a[6]  & \b[32]  ;
  assign n8567 = n419 & n8566 ;
  assign n8568 = ~n8565 & ~n8567 ;
  assign n8569 = \b[31]  & n486 ;
  assign n8570 = n483 & n8569 ;
  assign n8571 = ~\a[6]  & \b[32]  ;
  assign n8572 = n422 & n8571 ;
  assign n8573 = ~n8570 & ~n8572 ;
  assign n8574 = n8568 & n8573 ;
  assign n8575 = ~n8564 & n8574 ;
  assign n8576 = ~\a[8]  & ~n8575 ;
  assign n8577 = \a[8]  & n8574 ;
  assign n8578 = ~n8564 & n8577 ;
  assign n8579 = ~n8576 & ~n8578 ;
  assign n8580 = n8562 & ~n8579 ;
  assign n8581 = ~n8562 & n8579 ;
  assign n8582 = ~n8580 & ~n8581 ;
  assign n8583 = n8231 & ~n8582 ;
  assign n8584 = n8211 & n8583 ;
  assign n8585 = n8231 & n8582 ;
  assign n8586 = ~n8211 & n8585 ;
  assign n8587 = ~n8584 & ~n8586 ;
  assign n8588 = ~n8231 & ~n8582 ;
  assign n8589 = ~n8211 & n8588 ;
  assign n8590 = ~n8231 & n8582 ;
  assign n8591 = n8211 & n8590 ;
  assign n8592 = ~n8589 & ~n8591 ;
  assign n8593 = n8587 & n8592 ;
  assign n8594 = ~n7756 & n8175 ;
  assign n8595 = ~n8171 & n8594 ;
  assign n8596 = ~n8174 & ~n8595 ;
  assign n8597 = ~\b[38]  & ~\b[39]  ;
  assign n8598 = \b[38]  & \b[39]  ;
  assign n8599 = ~n8597 & ~n8598 ;
  assign n8600 = ~n8596 & n8599 ;
  assign n8601 = ~n8174 & ~n8599 ;
  assign n8602 = ~n8595 & n8601 ;
  assign n8603 = n134 & ~n8602 ;
  assign n8604 = ~n8600 & n8603 ;
  assign n8605 = \a[0]  & \b[39]  ;
  assign n8606 = n133 & n8605 ;
  assign n8607 = \b[38]  & n141 ;
  assign n8608 = ~\a[1]  & \b[37]  ;
  assign n8609 = n1521 & n8608 ;
  assign n8610 = ~n8607 & ~n8609 ;
  assign n8611 = ~n8606 & n8610 ;
  assign n8612 = ~n8604 & n8611 ;
  assign n8613 = ~\a[2]  & ~n8612 ;
  assign n8614 = \a[2]  & n8611 ;
  assign n8615 = ~n8604 & n8614 ;
  assign n8616 = ~n8613 & ~n8615 ;
  assign n8617 = ~n8593 & ~n8616 ;
  assign n8618 = n8209 & n8617 ;
  assign n8619 = n8593 & ~n8616 ;
  assign n8620 = ~n8209 & n8619 ;
  assign n8621 = ~n8618 & ~n8620 ;
  assign n8622 = ~n8593 & n8616 ;
  assign n8623 = ~n8209 & n8622 ;
  assign n8624 = n8593 & n8616 ;
  assign n8625 = n8209 & n8624 ;
  assign n8626 = ~n8623 & ~n8625 ;
  assign n8627 = n8621 & n8626 ;
  assign n8628 = ~n8206 & n8627 ;
  assign n8629 = ~n8196 & ~n8627 ;
  assign n8630 = ~n8203 & n8629 ;
  assign n8631 = ~n8628 & ~n8630 ;
  assign n8632 = ~n8196 & n8621 ;
  assign n8633 = ~n8203 & n8632 ;
  assign n8634 = n8626 & ~n8633 ;
  assign n8635 = n8209 & n8593 ;
  assign n8636 = n8592 & ~n8635 ;
  assign n8637 = n8154 & ~n8580 ;
  assign n8638 = ~n8210 & n8637 ;
  assign n8639 = ~n8581 & ~n8638 ;
  assign n8640 = ~n8553 & ~n8560 ;
  assign n8641 = n430 & n6565 ;
  assign n8642 = ~n6562 & n8641 ;
  assign n8643 = n430 & n7720 ;
  assign n8644 = ~n6561 & n8643 ;
  assign n8645 = \b[32]  & n486 ;
  assign n8646 = n483 & n8645 ;
  assign n8647 = ~\a[6]  & \b[33]  ;
  assign n8648 = n422 & n8647 ;
  assign n8649 = ~n8646 & ~n8648 ;
  assign n8650 = \b[34]  & n428 ;
  assign n8651 = \a[6]  & \b[33]  ;
  assign n8652 = n419 & n8651 ;
  assign n8653 = \a[8]  & ~n8652 ;
  assign n8654 = ~n8650 & n8653 ;
  assign n8655 = n8649 & n8654 ;
  assign n8656 = ~n8644 & n8655 ;
  assign n8657 = ~n8642 & n8656 ;
  assign n8658 = ~n8650 & ~n8652 ;
  assign n8659 = n8649 & n8658 ;
  assign n8660 = ~n8644 & n8659 ;
  assign n8661 = ~n8642 & n8660 ;
  assign n8662 = ~\a[8]  & ~n8661 ;
  assign n8663 = ~n8657 & ~n8662 ;
  assign n8664 = ~n8132 & n8523 ;
  assign n8665 = ~n8235 & n8664 ;
  assign n8666 = n8528 & ~n8665 ;
  assign n8667 = n646 & ~n5462 ;
  assign n8668 = ~n5460 & n8667 ;
  assign n8669 = \b[31]  & n644 ;
  assign n8670 = \a[9]  & \b[30]  ;
  assign n8671 = n635 & n8670 ;
  assign n8672 = ~n8669 & ~n8671 ;
  assign n8673 = \b[29]  & n796 ;
  assign n8674 = n793 & n8673 ;
  assign n8675 = ~\a[9]  & \b[30]  ;
  assign n8676 = n638 & n8675 ;
  assign n8677 = ~n8674 & ~n8676 ;
  assign n8678 = n8672 & n8677 ;
  assign n8679 = ~n8668 & n8678 ;
  assign n8680 = ~\a[11]  & ~n8679 ;
  assign n8681 = \a[11]  & n8678 ;
  assign n8682 = ~n8668 & n8681 ;
  assign n8683 = ~n8680 & ~n8682 ;
  assign n8684 = n8239 & n8499 ;
  assign n8685 = ~n8498 & ~n8684 ;
  assign n8686 = ~n8086 & n8459 ;
  assign n8687 = ~n8240 & n8686 ;
  assign n8688 = n8464 & ~n8687 ;
  assign n8689 = n8244 & n8435 ;
  assign n8690 = ~n8429 & ~n8689 ;
  assign n8691 = n8029 & n8395 ;
  assign n8692 = n8400 & ~n8691 ;
  assign n8693 = n8030 & n8400 ;
  assign n8694 = n7889 & n8693 ;
  assign n8695 = ~n8692 & ~n8694 ;
  assign n8696 = n8249 & n8373 ;
  assign n8697 = ~n8372 & ~n8696 ;
  assign n8698 = ~n8010 & n8332 ;
  assign n8699 = ~n8014 & n8698 ;
  assign n8700 = n8337 & ~n8699 ;
  assign n8701 = ~n948 & n4249 ;
  assign n8702 = ~n908 & n4249 ;
  assign n8703 = ~n912 & n8702 ;
  assign n8704 = ~n8701 & ~n8703 ;
  assign n8705 = ~n951 & ~n8704 ;
  assign n8706 = \b[11]  & n4647 ;
  assign n8707 = n4644 & n8706 ;
  assign n8708 = ~\a[26]  & \b[12]  ;
  assign n8709 = n4646 & n8708 ;
  assign n8710 = ~n8707 & ~n8709 ;
  assign n8711 = \b[13]  & n4247 ;
  assign n8712 = \a[27]  & \b[12]  ;
  assign n8713 = n4238 & n8712 ;
  assign n8714 = \a[29]  & ~n8713 ;
  assign n8715 = ~n8711 & n8714 ;
  assign n8716 = n8710 & n8715 ;
  assign n8717 = ~n8705 & n8716 ;
  assign n8718 = ~n8711 & ~n8713 ;
  assign n8719 = n8710 & n8718 ;
  assign n8720 = ~\a[29]  & ~n8719 ;
  assign n8721 = ~\a[29]  & ~n951 ;
  assign n8722 = ~n8704 & n8721 ;
  assign n8723 = ~n8720 & ~n8722 ;
  assign n8724 = ~n8717 & n8723 ;
  assign n8725 = n8253 & n8305 ;
  assign n8726 = ~n8303 & ~n8725 ;
  assign n8727 = ~n8275 & ~n8278 ;
  assign n8728 = n222 & n7534 ;
  assign n8729 = \b[4]  & n7532 ;
  assign n8730 = \a[35]  & \b[3]  ;
  assign n8731 = n7971 & n8730 ;
  assign n8732 = ~\a[36]  & \b[3]  ;
  assign n8733 = n7526 & n8732 ;
  assign n8734 = ~n8731 & ~n8733 ;
  assign n8735 = ~n8729 & n8734 ;
  assign n8736 = \b[2]  & n7973 ;
  assign n8737 = n7970 & n8736 ;
  assign n8738 = \a[38]  & ~n8737 ;
  assign n8739 = n8735 & n8738 ;
  assign n8740 = ~n8728 & n8739 ;
  assign n8741 = n8735 & ~n8737 ;
  assign n8742 = ~n8728 & n8741 ;
  assign n8743 = ~\a[38]  & ~n8742 ;
  assign n8744 = ~n8740 & ~n8743 ;
  assign n8745 = \a[41]  & \b[0]  ;
  assign n8746 = ~n8272 & n8745 ;
  assign n8747 = \a[39]  & \b[0]  ;
  assign n8748 = \a[38]  & ~\a[40]  ;
  assign n8749 = n8747 & n8748 ;
  assign n8750 = ~\a[39]  & \b[0]  ;
  assign n8751 = ~\a[38]  & \a[40]  ;
  assign n8752 = n8750 & n8751 ;
  assign n8753 = ~n8749 & ~n8752 ;
  assign n8754 = \a[40]  & ~\a[41]  ;
  assign n8755 = ~\a[40]  & \a[41]  ;
  assign n8756 = ~n8754 & ~n8755 ;
  assign n8757 = ~n8272 & n8756 ;
  assign n8758 = \b[1]  & n8757 ;
  assign n8759 = ~n8272 & ~n8756 ;
  assign n8760 = ~n137 & n8759 ;
  assign n8761 = ~n8758 & ~n8760 ;
  assign n8762 = n8753 & n8761 ;
  assign n8763 = n8746 & ~n8762 ;
  assign n8764 = ~n8746 & n8753 ;
  assign n8765 = n8761 & n8764 ;
  assign n8766 = ~n8763 & ~n8765 ;
  assign n8767 = n8744 & ~n8766 ;
  assign n8768 = ~n8744 & n8766 ;
  assign n8769 = ~n8767 & ~n8768 ;
  assign n8770 = ~n8727 & n8769 ;
  assign n8771 = n8727 & ~n8769 ;
  assign n8772 = ~n8770 & ~n8771 ;
  assign n8773 = ~n380 & n6309 ;
  assign n8774 = ~n322 & n6309 ;
  assign n8775 = ~n326 & n8774 ;
  assign n8776 = ~n8773 & ~n8775 ;
  assign n8777 = ~n383 & ~n8776 ;
  assign n8778 = \b[5]  & n6778 ;
  assign n8779 = n6775 & n8778 ;
  assign n8780 = \b[7]  & n6307 ;
  assign n8781 = \a[32]  & \b[6]  ;
  assign n8782 = n6776 & n8781 ;
  assign n8783 = ~\a[33]  & \b[6]  ;
  assign n8784 = n6301 & n8783 ;
  assign n8785 = ~n8782 & ~n8784 ;
  assign n8786 = ~n8780 & n8785 ;
  assign n8787 = ~n8779 & n8786 ;
  assign n8788 = ~\a[35]  & n8787 ;
  assign n8789 = ~n8777 & n8788 ;
  assign n8790 = \a[35]  & ~n8787 ;
  assign n8791 = \a[35]  & ~n383 ;
  assign n8792 = ~n8776 & n8791 ;
  assign n8793 = ~n8790 & ~n8792 ;
  assign n8794 = ~n8789 & n8793 ;
  assign n8795 = n8772 & n8794 ;
  assign n8796 = ~n8772 & ~n8794 ;
  assign n8797 = ~n8795 & ~n8796 ;
  assign n8798 = ~n685 & ~n4909 ;
  assign n8799 = ~n5208 & n8798 ;
  assign n8800 = n682 & n8799 ;
  assign n8801 = n685 & ~n4909 ;
  assign n8802 = ~n5208 & n8801 ;
  assign n8803 = ~n682 & n8802 ;
  assign n8804 = ~n8800 & ~n8803 ;
  assign n8805 = \b[8]  & n5595 ;
  assign n8806 = n5592 & n8805 ;
  assign n8807 = \b[10]  & n5209 ;
  assign n8808 = \a[29]  & \b[9]  ;
  assign n8809 = n5593 & n8808 ;
  assign n8810 = ~\a[30]  & \b[9]  ;
  assign n8811 = n5203 & n8810 ;
  assign n8812 = ~n8809 & ~n8811 ;
  assign n8813 = ~n8807 & n8812 ;
  assign n8814 = ~n8806 & n8813 ;
  assign n8815 = n8804 & n8814 ;
  assign n8816 = ~\a[32]  & ~n8815 ;
  assign n8817 = \a[32]  & n8814 ;
  assign n8818 = n8804 & n8817 ;
  assign n8819 = ~n8816 & ~n8818 ;
  assign n8820 = ~n8797 & ~n8819 ;
  assign n8821 = ~n8726 & n8820 ;
  assign n8822 = n8797 & ~n8819 ;
  assign n8823 = n8726 & n8822 ;
  assign n8824 = ~n8821 & ~n8823 ;
  assign n8825 = ~n8797 & n8819 ;
  assign n8826 = n8726 & n8825 ;
  assign n8827 = n8797 & n8819 ;
  assign n8828 = ~n8726 & n8827 ;
  assign n8829 = ~n8826 & ~n8828 ;
  assign n8830 = n8824 & n8829 ;
  assign n8831 = n8724 & ~n8830 ;
  assign n8832 = ~n8700 & n8831 ;
  assign n8833 = n8724 & n8830 ;
  assign n8834 = n8700 & n8833 ;
  assign n8835 = ~n8832 & ~n8834 ;
  assign n8836 = ~n8724 & ~n8830 ;
  assign n8837 = n8700 & n8836 ;
  assign n8838 = ~n8724 & n8830 ;
  assign n8839 = ~n8700 & n8838 ;
  assign n8840 = ~n8837 & ~n8839 ;
  assign n8841 = n8835 & n8840 ;
  assign n8842 = ~n8697 & n8841 ;
  assign n8843 = ~n8372 & ~n8841 ;
  assign n8844 = ~n8696 & n8843 ;
  assign n8845 = ~n1512 & ~n3154 ;
  assign n8846 = ~n3399 & n8845 ;
  assign n8847 = n1509 & n8846 ;
  assign n8848 = n1512 & ~n3154 ;
  assign n8849 = ~n3399 & n8848 ;
  assign n8850 = ~n1509 & n8849 ;
  assign n8851 = ~n8847 & ~n8850 ;
  assign n8852 = \b[14]  & n3733 ;
  assign n8853 = n3730 & n8852 ;
  assign n8854 = \b[16]  & n3400 ;
  assign n8855 = \a[24]  & \b[15]  ;
  assign n8856 = n3391 & n8855 ;
  assign n8857 = ~\a[23]  & \b[15]  ;
  assign n8858 = n3732 & n8857 ;
  assign n8859 = ~n8856 & ~n8858 ;
  assign n8860 = ~n8854 & n8859 ;
  assign n8861 = ~n8853 & n8860 ;
  assign n8862 = n8851 & n8861 ;
  assign n8863 = ~\a[26]  & ~n8862 ;
  assign n8864 = \a[26]  & n8861 ;
  assign n8865 = n8851 & n8864 ;
  assign n8866 = ~n8863 & ~n8865 ;
  assign n8867 = ~n8844 & ~n8866 ;
  assign n8868 = ~n8842 & n8867 ;
  assign n8869 = ~n8841 & n8866 ;
  assign n8870 = n8697 & n8869 ;
  assign n8871 = n8841 & n8866 ;
  assign n8872 = ~n8697 & n8871 ;
  assign n8873 = ~n8870 & ~n8872 ;
  assign n8874 = ~n8868 & n8873 ;
  assign n8875 = n8695 & ~n8874 ;
  assign n8876 = ~n8695 & n8874 ;
  assign n8877 = ~n8875 & ~n8876 ;
  assign n8878 = ~n2079 & n2622 ;
  assign n8879 = ~n2077 & n8878 ;
  assign n8880 = \b[17]  & n2912 ;
  assign n8881 = n2909 & n8880 ;
  assign n8882 = \b[19]  & n2620 ;
  assign n8883 = \a[20]  & \b[18]  ;
  assign n8884 = n2910 & n8883 ;
  assign n8885 = ~\a[21]  & \b[18]  ;
  assign n8886 = n2614 & n8885 ;
  assign n8887 = ~n8884 & ~n8886 ;
  assign n8888 = ~n8882 & n8887 ;
  assign n8889 = ~n8881 & n8888 ;
  assign n8890 = ~n8879 & n8889 ;
  assign n8891 = ~\a[23]  & ~n8890 ;
  assign n8892 = \a[23]  & n8889 ;
  assign n8893 = ~n8879 & n8892 ;
  assign n8894 = ~n8891 & ~n8893 ;
  assign n8895 = n8877 & ~n8894 ;
  assign n8896 = ~n8877 & n8894 ;
  assign n8897 = ~n8895 & ~n8896 ;
  assign n8898 = ~n8690 & n8897 ;
  assign n8899 = ~n8429 & ~n8897 ;
  assign n8900 = ~n8689 & n8899 ;
  assign n8901 = n1965 & ~n2771 ;
  assign n8902 = ~n2769 & n8901 ;
  assign n8903 = \b[20]  & n2218 ;
  assign n8904 = n2216 & n8903 ;
  assign n8905 = \b[22]  & n1963 ;
  assign n8906 = \a[17]  & \b[21]  ;
  assign n8907 = n1954 & n8906 ;
  assign n8908 = ~\a[18]  & \b[21]  ;
  assign n8909 = n1957 & n8908 ;
  assign n8910 = ~n8907 & ~n8909 ;
  assign n8911 = ~n8905 & n8910 ;
  assign n8912 = ~n8904 & n8911 ;
  assign n8913 = ~n8902 & n8912 ;
  assign n8914 = ~\a[20]  & ~n8913 ;
  assign n8915 = \a[20]  & n8912 ;
  assign n8916 = ~n8902 & n8915 ;
  assign n8917 = ~n8914 & ~n8916 ;
  assign n8918 = ~n8900 & ~n8917 ;
  assign n8919 = ~n8898 & n8918 ;
  assign n8920 = ~n8897 & n8917 ;
  assign n8921 = n8690 & n8920 ;
  assign n8922 = n8897 & n8917 ;
  assign n8923 = ~n8690 & n8922 ;
  assign n8924 = ~n8921 & ~n8923 ;
  assign n8925 = ~n8919 & n8924 ;
  assign n8926 = n1467 & ~n3567 ;
  assign n8927 = ~n3565 & n8926 ;
  assign n8928 = \b[25]  & n1465 ;
  assign n8929 = \a[15]  & \b[24]  ;
  assign n8930 = n1456 & n8929 ;
  assign n8931 = ~n8928 & ~n8930 ;
  assign n8932 = \b[23]  & n1652 ;
  assign n8933 = n1649 & n8932 ;
  assign n8934 = ~\a[14]  & \b[24]  ;
  assign n8935 = n1651 & n8934 ;
  assign n8936 = ~n8933 & ~n8935 ;
  assign n8937 = n8931 & n8936 ;
  assign n8938 = ~n8927 & n8937 ;
  assign n8939 = ~\a[17]  & ~n8938 ;
  assign n8940 = \a[17]  & n8937 ;
  assign n8941 = ~n8927 & n8940 ;
  assign n8942 = ~n8939 & ~n8941 ;
  assign n8943 = ~n8925 & ~n8942 ;
  assign n8944 = n8688 & n8943 ;
  assign n8945 = n8925 & ~n8942 ;
  assign n8946 = ~n8688 & n8945 ;
  assign n8947 = ~n8944 & ~n8946 ;
  assign n8948 = ~n8925 & n8942 ;
  assign n8949 = ~n8688 & n8948 ;
  assign n8950 = n8925 & n8942 ;
  assign n8951 = n8688 & n8950 ;
  assign n8952 = ~n8949 & ~n8951 ;
  assign n8953 = n8947 & n8952 ;
  assign n8954 = ~n8685 & n8953 ;
  assign n8955 = n999 & n4456 ;
  assign n8956 = ~n4453 & n8955 ;
  assign n8957 = n999 & n5421 ;
  assign n8958 = ~n4452 & n8957 ;
  assign n8959 = \b[26]  & n1182 ;
  assign n8960 = n1179 & n8959 ;
  assign n8961 = ~\a[12]  & \b[27]  ;
  assign n8962 = n7674 & n8961 ;
  assign n8963 = ~n8960 & ~n8962 ;
  assign n8964 = \b[28]  & n997 ;
  assign n8965 = \a[12]  & \b[27]  ;
  assign n8966 = n988 & n8965 ;
  assign n8967 = \a[14]  & ~n8966 ;
  assign n8968 = ~n8964 & n8967 ;
  assign n8969 = n8963 & n8968 ;
  assign n8970 = ~n8958 & n8969 ;
  assign n8971 = ~n8956 & n8970 ;
  assign n8972 = ~n8964 & ~n8966 ;
  assign n8973 = n8963 & n8972 ;
  assign n8974 = ~n8958 & n8973 ;
  assign n8975 = ~n8956 & n8974 ;
  assign n8976 = ~\a[14]  & ~n8975 ;
  assign n8977 = ~n8971 & ~n8976 ;
  assign n8978 = ~n8498 & ~n8953 ;
  assign n8979 = ~n8684 & n8978 ;
  assign n8980 = ~n8977 & ~n8979 ;
  assign n8981 = ~n8954 & n8980 ;
  assign n8982 = ~n8953 & n8977 ;
  assign n8983 = n8685 & n8982 ;
  assign n8984 = n8953 & n8977 ;
  assign n8985 = ~n8685 & n8984 ;
  assign n8986 = ~n8983 & ~n8985 ;
  assign n8987 = ~n8981 & n8986 ;
  assign n8988 = n8683 & ~n8987 ;
  assign n8989 = ~n8666 & n8988 ;
  assign n8990 = n8683 & n8987 ;
  assign n8991 = n8666 & n8990 ;
  assign n8992 = ~n8989 & ~n8991 ;
  assign n8993 = ~n8683 & ~n8987 ;
  assign n8994 = n8666 & n8993 ;
  assign n8995 = ~n8683 & n8987 ;
  assign n8996 = ~n8666 & n8995 ;
  assign n8997 = ~n8994 & ~n8996 ;
  assign n8998 = n8992 & n8997 ;
  assign n8999 = n8663 & ~n8998 ;
  assign n9000 = n8640 & n8999 ;
  assign n9001 = n8663 & n8998 ;
  assign n9002 = ~n8640 & n9001 ;
  assign n9003 = ~n9000 & ~n9002 ;
  assign n9004 = ~n8663 & ~n8998 ;
  assign n9005 = ~n8640 & n9004 ;
  assign n9006 = ~n8663 & n8998 ;
  assign n9007 = n8640 & n9006 ;
  assign n9008 = ~n9005 & ~n9007 ;
  assign n9009 = n9003 & n9008 ;
  assign n9010 = n252 & ~n7761 ;
  assign n9011 = ~n7759 & n9010 ;
  assign n9012 = \b[35]  & n303 ;
  assign n9013 = n300 & n9012 ;
  assign n9014 = \b[37]  & n250 ;
  assign n9015 = \a[2]  & \b[36]  ;
  assign n9016 = n301 & n9015 ;
  assign n9017 = ~\a[3]  & \b[36]  ;
  assign n9018 = n244 & n9017 ;
  assign n9019 = ~n9016 & ~n9018 ;
  assign n9020 = ~n9014 & n9019 ;
  assign n9021 = ~n9013 & n9020 ;
  assign n9022 = ~n9011 & n9021 ;
  assign n9023 = ~\a[5]  & ~n9022 ;
  assign n9024 = \a[5]  & n9021 ;
  assign n9025 = ~n9011 & n9024 ;
  assign n9026 = ~n9023 & ~n9025 ;
  assign n9027 = ~n9009 & ~n9026 ;
  assign n9028 = n8639 & n9027 ;
  assign n9029 = n9009 & ~n9026 ;
  assign n9030 = ~n8639 & n9029 ;
  assign n9031 = ~n9028 & ~n9030 ;
  assign n9032 = ~n9009 & n9026 ;
  assign n9033 = ~n8639 & n9032 ;
  assign n9034 = n9009 & n9026 ;
  assign n9035 = n8639 & n9034 ;
  assign n9036 = ~n9033 & ~n9035 ;
  assign n9037 = n9031 & n9036 ;
  assign n9038 = ~n8636 & n9037 ;
  assign n9039 = ~n8174 & ~n8598 ;
  assign n9040 = ~n8595 & n9039 ;
  assign n9041 = ~n8597 & ~n9040 ;
  assign n9042 = ~\b[39]  & ~\b[40]  ;
  assign n9043 = \b[39]  & \b[40]  ;
  assign n9044 = ~n9042 & ~n9043 ;
  assign n9045 = n134 & n9044 ;
  assign n9046 = ~n9041 & n9045 ;
  assign n9047 = n134 & ~n9044 ;
  assign n9048 = ~n8597 & n9047 ;
  assign n9049 = ~n9040 & n9048 ;
  assign n9050 = \a[0]  & \b[40]  ;
  assign n9051 = n133 & n9050 ;
  assign n9052 = \b[39]  & n141 ;
  assign n9053 = ~\a[1]  & \b[38]  ;
  assign n9054 = n1521 & n9053 ;
  assign n9055 = ~n9052 & ~n9054 ;
  assign n9056 = ~n9051 & n9055 ;
  assign n9057 = \a[2]  & n9056 ;
  assign n9058 = ~n9049 & n9057 ;
  assign n9059 = ~n9046 & n9058 ;
  assign n9060 = ~n9049 & n9056 ;
  assign n9061 = ~n9046 & n9060 ;
  assign n9062 = ~\a[2]  & ~n9061 ;
  assign n9063 = ~n9059 & ~n9062 ;
  assign n9064 = n8592 & ~n9037 ;
  assign n9065 = ~n8635 & n9064 ;
  assign n9066 = ~n9063 & ~n9065 ;
  assign n9067 = ~n9038 & n9066 ;
  assign n9068 = ~n9037 & n9063 ;
  assign n9069 = n8636 & n9068 ;
  assign n9070 = n9037 & n9063 ;
  assign n9071 = ~n8636 & n9070 ;
  assign n9072 = ~n9069 & ~n9071 ;
  assign n9073 = ~n9067 & n9072 ;
  assign n9074 = n8634 & n9073 ;
  assign n9075 = ~n8634 & ~n9073 ;
  assign n9076 = ~n9074 & ~n9075 ;
  assign n9077 = ~n9067 & ~n9074 ;
  assign n9078 = n8592 & n9031 ;
  assign n9079 = ~n8635 & n9078 ;
  assign n9080 = n9036 & ~n9079 ;
  assign n9081 = n8639 & n9009 ;
  assign n9082 = n9008 & ~n9081 ;
  assign n9083 = ~n8172 & ~n8175 ;
  assign n9084 = n252 & ~n8595 ;
  assign n9085 = ~n9083 & n9084 ;
  assign n9086 = \b[36]  & n303 ;
  assign n9087 = n300 & n9086 ;
  assign n9088 = \b[38]  & n250 ;
  assign n9089 = \a[2]  & \b[37]  ;
  assign n9090 = n301 & n9089 ;
  assign n9091 = ~\a[3]  & \b[37]  ;
  assign n9092 = n244 & n9091 ;
  assign n9093 = ~n9090 & ~n9092 ;
  assign n9094 = ~n9088 & n9093 ;
  assign n9095 = ~n9087 & n9094 ;
  assign n9096 = ~n9085 & n9095 ;
  assign n9097 = ~\a[5]  & ~n9096 ;
  assign n9098 = \a[5]  & n9095 ;
  assign n9099 = ~n9085 & n9098 ;
  assign n9100 = ~n9097 & ~n9099 ;
  assign n9101 = ~n8553 & n8997 ;
  assign n9102 = ~n8560 & n9101 ;
  assign n9103 = n8992 & ~n9102 ;
  assign n9104 = n8666 & n8987 ;
  assign n9105 = ~n8981 & ~n9104 ;
  assign n9106 = n646 & n5810 ;
  assign n9107 = ~n5807 & n9106 ;
  assign n9108 = n646 & ~n5810 ;
  assign n9109 = ~n5457 & n9108 ;
  assign n9110 = ~n5806 & n9109 ;
  assign n9111 = \b[30]  & n796 ;
  assign n9112 = n793 & n9111 ;
  assign n9113 = \b[32]  & n644 ;
  assign n9114 = \a[8]  & \b[31]  ;
  assign n9115 = n794 & n9114 ;
  assign n9116 = ~\a[9]  & \b[31]  ;
  assign n9117 = n638 & n9116 ;
  assign n9118 = ~n9115 & ~n9117 ;
  assign n9119 = ~n9113 & n9118 ;
  assign n9120 = ~n9112 & n9119 ;
  assign n9121 = ~n9110 & n9120 ;
  assign n9122 = ~n9107 & n9121 ;
  assign n9123 = ~\a[11]  & ~n9122 ;
  assign n9124 = \a[11]  & n9120 ;
  assign n9125 = ~n9110 & n9124 ;
  assign n9126 = ~n9107 & n9125 ;
  assign n9127 = ~n9123 & ~n9126 ;
  assign n9128 = ~n8498 & n8947 ;
  assign n9129 = ~n8684 & n9128 ;
  assign n9130 = n8952 & ~n9129 ;
  assign n9131 = n999 & ~n4502 ;
  assign n9132 = ~n4500 & n9131 ;
  assign n9133 = \b[27]  & n1182 ;
  assign n9134 = n1179 & n9133 ;
  assign n9135 = \b[29]  & n997 ;
  assign n9136 = \a[11]  & \b[28]  ;
  assign n9137 = n1180 & n9136 ;
  assign n9138 = ~\a[12]  & \b[28]  ;
  assign n9139 = n7674 & n9138 ;
  assign n9140 = ~n9137 & ~n9139 ;
  assign n9141 = ~n9135 & n9140 ;
  assign n9142 = ~n9134 & n9141 ;
  assign n9143 = ~n9132 & n9142 ;
  assign n9144 = ~\a[14]  & ~n9143 ;
  assign n9145 = \a[14]  & n9142 ;
  assign n9146 = ~n9132 & n9145 ;
  assign n9147 = ~n9144 & ~n9146 ;
  assign n9148 = n8688 & n8925 ;
  assign n9149 = ~n8919 & ~n9148 ;
  assign n9150 = n1467 & ~n4141 ;
  assign n9151 = ~n4518 & n9150 ;
  assign n9152 = \b[24]  & n1652 ;
  assign n9153 = n1649 & n9152 ;
  assign n9154 = ~\a[14]  & \b[25]  ;
  assign n9155 = n1651 & n9154 ;
  assign n9156 = ~n9153 & ~n9155 ;
  assign n9157 = \b[26]  & n1465 ;
  assign n9158 = \a[15]  & \b[25]  ;
  assign n9159 = n1456 & n9158 ;
  assign n9160 = \a[17]  & ~n9159 ;
  assign n9161 = ~n9157 & n9160 ;
  assign n9162 = n9156 & n9161 ;
  assign n9163 = ~n9151 & n9162 ;
  assign n9164 = ~n9157 & ~n9159 ;
  assign n9165 = n9156 & n9164 ;
  assign n9166 = ~n9151 & n9165 ;
  assign n9167 = ~\a[17]  & ~n9166 ;
  assign n9168 = ~n9163 & ~n9167 ;
  assign n9169 = ~n8429 & ~n8895 ;
  assign n9170 = ~n8689 & n9169 ;
  assign n9171 = ~n8896 & ~n9170 ;
  assign n9172 = ~n8868 & ~n8876 ;
  assign n9173 = ~n8372 & n8840 ;
  assign n9174 = ~n8696 & n9173 ;
  assign n9175 = n8835 & ~n9174 ;
  assign n9176 = ~n1694 & n3402 ;
  assign n9177 = ~n1692 & n9176 ;
  assign n9178 = \b[15]  & n3733 ;
  assign n9179 = n3730 & n9178 ;
  assign n9180 = ~\a[24]  & \b[16]  ;
  assign n9181 = n3394 & n9180 ;
  assign n9182 = ~n9179 & ~n9181 ;
  assign n9183 = \b[17]  & n3400 ;
  assign n9184 = \a[24]  & \b[16]  ;
  assign n9185 = n3391 & n9184 ;
  assign n9186 = \a[26]  & ~n9185 ;
  assign n9187 = ~n9183 & n9186 ;
  assign n9188 = n9182 & n9187 ;
  assign n9189 = ~n9177 & n9188 ;
  assign n9190 = ~n9183 & ~n9185 ;
  assign n9191 = n9182 & n9190 ;
  assign n9192 = ~n9177 & n9191 ;
  assign n9193 = ~\a[26]  & ~n9192 ;
  assign n9194 = ~n9189 & ~n9193 ;
  assign n9195 = n8700 & n8830 ;
  assign n9196 = n8824 & ~n9195 ;
  assign n9197 = n1087 & n4249 ;
  assign n9198 = ~n1084 & n9197 ;
  assign n9199 = ~n1087 & n4249 ;
  assign n9200 = ~n946 & n9199 ;
  assign n9201 = ~n1083 & n9200 ;
  assign n9202 = \b[12]  & n4647 ;
  assign n9203 = n4644 & n9202 ;
  assign n9204 = ~\a[27]  & \b[13]  ;
  assign n9205 = n4241 & n9204 ;
  assign n9206 = ~n9203 & ~n9205 ;
  assign n9207 = \b[14]  & n4247 ;
  assign n9208 = \a[27]  & \b[13]  ;
  assign n9209 = n4238 & n9208 ;
  assign n9210 = \a[29]  & ~n9209 ;
  assign n9211 = ~n9207 & n9210 ;
  assign n9212 = n9206 & n9211 ;
  assign n9213 = ~n9201 & n9212 ;
  assign n9214 = ~n9198 & n9213 ;
  assign n9215 = ~n9207 & ~n9209 ;
  assign n9216 = n9206 & n9215 ;
  assign n9217 = ~n9201 & n9216 ;
  assign n9218 = ~n9198 & n9217 ;
  assign n9219 = ~\a[29]  & ~n9218 ;
  assign n9220 = ~n9214 & ~n9219 ;
  assign n9221 = ~n725 & n5211 ;
  assign n9222 = ~n684 & n5211 ;
  assign n9223 = ~n721 & n9222 ;
  assign n9224 = ~n9221 & ~n9223 ;
  assign n9225 = ~n728 & ~n9224 ;
  assign n9226 = \b[9]  & n5595 ;
  assign n9227 = n5592 & n9226 ;
  assign n9228 = \b[11]  & n5209 ;
  assign n9229 = \a[30]  & \b[10]  ;
  assign n9230 = n5200 & n9229 ;
  assign n9231 = ~\a[30]  & \b[10]  ;
  assign n9232 = n5203 & n9231 ;
  assign n9233 = ~n9230 & ~n9232 ;
  assign n9234 = ~n9228 & n9233 ;
  assign n9235 = ~n9227 & n9234 ;
  assign n9236 = ~\a[32]  & n9235 ;
  assign n9237 = ~n9225 & n9236 ;
  assign n9238 = \a[32]  & ~n9235 ;
  assign n9239 = \a[32]  & ~n728 ;
  assign n9240 = ~n9224 & n9239 ;
  assign n9241 = ~n9238 & ~n9240 ;
  assign n9242 = ~n9237 & n9241 ;
  assign n9243 = ~n8303 & ~n8795 ;
  assign n9244 = ~n8725 & n9243 ;
  assign n9245 = ~n8796 & ~n9244 ;
  assign n9246 = ~n505 & ~n5952 ;
  assign n9247 = ~n6306 & n9246 ;
  assign n9248 = n502 & n9247 ;
  assign n9249 = n505 & ~n5952 ;
  assign n9250 = ~n6306 & n9249 ;
  assign n9251 = ~n502 & n9250 ;
  assign n9252 = ~n9248 & ~n9251 ;
  assign n9253 = \b[6]  & n6778 ;
  assign n9254 = n6775 & n9253 ;
  assign n9255 = \b[8]  & n6307 ;
  assign n9256 = \a[32]  & \b[7]  ;
  assign n9257 = n6776 & n9256 ;
  assign n9258 = ~\a[33]  & \b[7]  ;
  assign n9259 = n6301 & n9258 ;
  assign n9260 = ~n9257 & ~n9259 ;
  assign n9261 = ~n9255 & n9260 ;
  assign n9262 = ~n9254 & n9261 ;
  assign n9263 = n9252 & n9262 ;
  assign n9264 = ~\a[35]  & ~n9263 ;
  assign n9265 = \a[35]  & n9262 ;
  assign n9266 = n9252 & n9265 ;
  assign n9267 = ~n9264 & ~n9266 ;
  assign n9268 = ~n8768 & ~n8770 ;
  assign n9269 = ~n273 & n7534 ;
  assign n9270 = ~n271 & n9269 ;
  assign n9271 = \b[3]  & n7973 ;
  assign n9272 = n7970 & n9271 ;
  assign n9273 = \b[5]  & n7532 ;
  assign n9274 = \a[35]  & \b[4]  ;
  assign n9275 = n7971 & n9274 ;
  assign n9276 = ~\a[36]  & \b[4]  ;
  assign n9277 = n7526 & n9276 ;
  assign n9278 = ~n9275 & ~n9277 ;
  assign n9279 = ~n9273 & n9278 ;
  assign n9280 = ~n9272 & n9279 ;
  assign n9281 = ~\a[38]  & n9280 ;
  assign n9282 = ~n9270 & n9281 ;
  assign n9283 = ~n9270 & n9280 ;
  assign n9284 = \a[38]  & ~n9283 ;
  assign n9285 = ~n9282 & ~n9284 ;
  assign n9286 = \a[41]  & ~n8273 ;
  assign n9287 = n8753 & n9286 ;
  assign n9288 = n8761 & n9287 ;
  assign n9289 = \a[41]  & ~n9288 ;
  assign n9290 = \b[2]  & n8757 ;
  assign n9291 = ~\a[39]  & \b[1]  ;
  assign n9292 = n8751 & n9291 ;
  assign n9293 = \a[39]  & \b[1]  ;
  assign n9294 = n8748 & n9293 ;
  assign n9295 = ~n9292 & ~n9294 ;
  assign n9296 = ~n9290 & n9295 ;
  assign n9297 = n157 & n8759 ;
  assign n9298 = n8272 & ~n8756 ;
  assign n9299 = \a[39]  & ~\a[40]  ;
  assign n9300 = ~\a[39]  & \a[40]  ;
  assign n9301 = ~n9299 & ~n9300 ;
  assign n9302 = \b[0]  & n9301 ;
  assign n9303 = n9298 & n9302 ;
  assign n9304 = ~n9297 & ~n9303 ;
  assign n9305 = n9296 & n9304 ;
  assign n9306 = ~n9289 & ~n9305 ;
  assign n9307 = n9289 & n9305 ;
  assign n9308 = ~n9306 & ~n9307 ;
  assign n9309 = n9285 & ~n9308 ;
  assign n9310 = ~n9285 & n9308 ;
  assign n9311 = ~n9309 & ~n9310 ;
  assign n9312 = ~n9268 & n9311 ;
  assign n9313 = n9268 & ~n9311 ;
  assign n9314 = ~n9312 & ~n9313 ;
  assign n9315 = ~n9267 & n9314 ;
  assign n9316 = n9267 & ~n9314 ;
  assign n9317 = ~n9315 & ~n9316 ;
  assign n9318 = n9245 & n9317 ;
  assign n9319 = ~n9245 & ~n9317 ;
  assign n9320 = ~n9318 & ~n9319 ;
  assign n9321 = ~n9242 & ~n9320 ;
  assign n9322 = n9242 & n9320 ;
  assign n9323 = ~n9321 & ~n9322 ;
  assign n9324 = n9220 & ~n9323 ;
  assign n9325 = n9196 & n9324 ;
  assign n9326 = n9220 & n9323 ;
  assign n9327 = ~n9196 & n9326 ;
  assign n9328 = ~n9325 & ~n9327 ;
  assign n9329 = ~n9220 & ~n9323 ;
  assign n9330 = ~n9196 & n9329 ;
  assign n9331 = ~n9220 & n9323 ;
  assign n9332 = n9196 & n9331 ;
  assign n9333 = ~n9330 & ~n9332 ;
  assign n9334 = n9328 & n9333 ;
  assign n9335 = n9194 & ~n9334 ;
  assign n9336 = ~n9175 & n9335 ;
  assign n9337 = n9194 & n9334 ;
  assign n9338 = n9175 & n9337 ;
  assign n9339 = ~n9336 & ~n9338 ;
  assign n9340 = ~n9194 & ~n9334 ;
  assign n9341 = n9175 & n9340 ;
  assign n9342 = ~n9194 & n9334 ;
  assign n9343 = ~n9175 & n9342 ;
  assign n9344 = ~n9341 & ~n9343 ;
  assign n9345 = n9339 & n9344 ;
  assign n9346 = n2293 & n2622 ;
  assign n9347 = ~n2290 & n9346 ;
  assign n9348 = n2622 & n5705 ;
  assign n9349 = ~n2289 & n9348 ;
  assign n9350 = \b[20]  & n2620 ;
  assign n9351 = \a[20]  & \b[19]  ;
  assign n9352 = n2910 & n9351 ;
  assign n9353 = ~\a[21]  & \b[19]  ;
  assign n9354 = n2614 & n9353 ;
  assign n9355 = ~n9352 & ~n9354 ;
  assign n9356 = ~n9350 & n9355 ;
  assign n9357 = \b[18]  & n2912 ;
  assign n9358 = n2909 & n9357 ;
  assign n9359 = \a[23]  & ~n9358 ;
  assign n9360 = n9356 & n9359 ;
  assign n9361 = ~n9349 & n9360 ;
  assign n9362 = ~n9347 & n9361 ;
  assign n9363 = n9356 & ~n9358 ;
  assign n9364 = ~n9349 & n9363 ;
  assign n9365 = ~n9347 & n9364 ;
  assign n9366 = ~\a[23]  & ~n9365 ;
  assign n9367 = ~n9362 & ~n9366 ;
  assign n9368 = ~n9345 & ~n9367 ;
  assign n9369 = ~n9172 & n9368 ;
  assign n9370 = n9345 & ~n9367 ;
  assign n9371 = n9172 & n9370 ;
  assign n9372 = ~n9369 & ~n9371 ;
  assign n9373 = ~n9345 & n9367 ;
  assign n9374 = n9172 & n9373 ;
  assign n9375 = n9345 & n9367 ;
  assign n9376 = ~n9172 & n9375 ;
  assign n9377 = ~n9374 & ~n9376 ;
  assign n9378 = n9372 & n9377 ;
  assign n9379 = ~n9171 & ~n9378 ;
  assign n9380 = ~n8896 & n9378 ;
  assign n9381 = ~n9170 & n9380 ;
  assign n9382 = n1965 & ~n3022 ;
  assign n9383 = ~n3020 & n9382 ;
  assign n9384 = \b[23]  & n1963 ;
  assign n9385 = \a[18]  & \b[22]  ;
  assign n9386 = n2210 & n9385 ;
  assign n9387 = ~n9384 & ~n9386 ;
  assign n9388 = \b[21]  & n2218 ;
  assign n9389 = n2216 & n9388 ;
  assign n9390 = ~\a[18]  & \b[22]  ;
  assign n9391 = n1957 & n9390 ;
  assign n9392 = ~n9389 & ~n9391 ;
  assign n9393 = n9387 & n9392 ;
  assign n9394 = ~n9383 & n9393 ;
  assign n9395 = ~\a[20]  & ~n9394 ;
  assign n9396 = \a[20]  & n9393 ;
  assign n9397 = ~n9383 & n9396 ;
  assign n9398 = ~n9395 & ~n9397 ;
  assign n9399 = ~n9381 & ~n9398 ;
  assign n9400 = ~n9379 & n9399 ;
  assign n9401 = ~n9378 & n9398 ;
  assign n9402 = ~n9171 & n9401 ;
  assign n9403 = n9378 & n9398 ;
  assign n9404 = n9171 & n9403 ;
  assign n9405 = ~n9402 & ~n9404 ;
  assign n9406 = ~n9400 & n9405 ;
  assign n9407 = n9168 & ~n9406 ;
  assign n9408 = n9149 & n9407 ;
  assign n9409 = n9168 & n9406 ;
  assign n9410 = ~n9149 & n9409 ;
  assign n9411 = ~n9408 & ~n9410 ;
  assign n9412 = ~n9149 & n9406 ;
  assign n9413 = ~n8919 & ~n9406 ;
  assign n9414 = ~n9148 & n9413 ;
  assign n9415 = ~n9168 & ~n9414 ;
  assign n9416 = ~n9412 & n9415 ;
  assign n9417 = n9411 & ~n9416 ;
  assign n9418 = n9147 & ~n9417 ;
  assign n9419 = ~n9130 & n9418 ;
  assign n9420 = n9147 & n9417 ;
  assign n9421 = n9130 & n9420 ;
  assign n9422 = ~n9419 & ~n9421 ;
  assign n9423 = ~n9147 & ~n9417 ;
  assign n9424 = n9130 & n9423 ;
  assign n9425 = ~n9147 & n9417 ;
  assign n9426 = ~n9130 & n9425 ;
  assign n9427 = ~n9424 & ~n9426 ;
  assign n9428 = n9422 & n9427 ;
  assign n9429 = n9127 & ~n9428 ;
  assign n9430 = n9105 & n9429 ;
  assign n9431 = n9127 & n9428 ;
  assign n9432 = ~n9105 & n9431 ;
  assign n9433 = ~n9430 & ~n9432 ;
  assign n9434 = ~n9105 & n9428 ;
  assign n9435 = ~n8981 & ~n9428 ;
  assign n9436 = ~n9104 & n9435 ;
  assign n9437 = ~n9127 & ~n9436 ;
  assign n9438 = ~n9434 & n9437 ;
  assign n9439 = n9433 & ~n9438 ;
  assign n9440 = n9103 & n9439 ;
  assign n9441 = ~n9103 & ~n9439 ;
  assign n9442 = ~n9440 & ~n9441 ;
  assign n9443 = n430 & ~n6610 ;
  assign n9444 = ~n6608 & n9443 ;
  assign n9445 = \b[33]  & n486 ;
  assign n9446 = n483 & n9445 ;
  assign n9447 = \b[35]  & n428 ;
  assign n9448 = \a[5]  & \b[34]  ;
  assign n9449 = n484 & n9448 ;
  assign n9450 = ~\a[6]  & \b[34]  ;
  assign n9451 = n422 & n9450 ;
  assign n9452 = ~n9449 & ~n9451 ;
  assign n9453 = ~n9447 & n9452 ;
  assign n9454 = ~n9446 & n9453 ;
  assign n9455 = ~n9444 & n9454 ;
  assign n9456 = ~\a[8]  & ~n9455 ;
  assign n9457 = \a[8]  & n9454 ;
  assign n9458 = ~n9444 & n9457 ;
  assign n9459 = ~n9456 & ~n9458 ;
  assign n9460 = n9442 & ~n9459 ;
  assign n9461 = ~n9442 & n9459 ;
  assign n9462 = ~n9460 & ~n9461 ;
  assign n9463 = ~n9100 & ~n9462 ;
  assign n9464 = ~n9082 & n9463 ;
  assign n9465 = ~n9100 & n9462 ;
  assign n9466 = n9082 & n9465 ;
  assign n9467 = ~n9464 & ~n9466 ;
  assign n9468 = n9100 & ~n9462 ;
  assign n9469 = n9082 & n9468 ;
  assign n9470 = n9100 & n9462 ;
  assign n9471 = ~n9082 & n9470 ;
  assign n9472 = ~n9469 & ~n9471 ;
  assign n9473 = n9467 & n9472 ;
  assign n9474 = ~n8597 & n9044 ;
  assign n9475 = ~n9040 & n9474 ;
  assign n9476 = ~n9043 & ~n9475 ;
  assign n9477 = ~\b[40]  & ~\b[41]  ;
  assign n9478 = \b[40]  & \b[41]  ;
  assign n9479 = ~n9477 & ~n9478 ;
  assign n9480 = ~n9476 & n9479 ;
  assign n9481 = ~n9043 & ~n9479 ;
  assign n9482 = ~n9475 & n9481 ;
  assign n9483 = n134 & ~n9482 ;
  assign n9484 = ~n9480 & n9483 ;
  assign n9485 = \a[0]  & \b[41]  ;
  assign n9486 = n133 & n9485 ;
  assign n9487 = \b[40]  & n141 ;
  assign n9488 = ~\a[1]  & \b[39]  ;
  assign n9489 = n1521 & n9488 ;
  assign n9490 = ~n9487 & ~n9489 ;
  assign n9491 = ~n9486 & n9490 ;
  assign n9492 = ~n9484 & n9491 ;
  assign n9493 = ~\a[2]  & ~n9492 ;
  assign n9494 = \a[2]  & n9491 ;
  assign n9495 = ~n9484 & n9494 ;
  assign n9496 = ~n9493 & ~n9495 ;
  assign n9497 = ~n9473 & n9496 ;
  assign n9498 = ~n9080 & n9497 ;
  assign n9499 = n9473 & n9496 ;
  assign n9500 = n9080 & n9499 ;
  assign n9501 = ~n9498 & ~n9500 ;
  assign n9502 = ~n9473 & ~n9496 ;
  assign n9503 = n9080 & n9502 ;
  assign n9504 = n9473 & ~n9496 ;
  assign n9505 = ~n9080 & n9504 ;
  assign n9506 = ~n9503 & ~n9505 ;
  assign n9507 = n9501 & n9506 ;
  assign n9508 = ~n9077 & n9507 ;
  assign n9509 = ~n9067 & ~n9507 ;
  assign n9510 = ~n9074 & n9509 ;
  assign n9511 = ~n9508 & ~n9510 ;
  assign n9512 = ~n9067 & n9506 ;
  assign n9513 = ~n9074 & n9512 ;
  assign n9514 = n9501 & ~n9513 ;
  assign n9515 = n9080 & n9473 ;
  assign n9516 = n9467 & ~n9515 ;
  assign n9517 = n9008 & ~n9460 ;
  assign n9518 = ~n9081 & n9517 ;
  assign n9519 = ~n9461 & ~n9518 ;
  assign n9520 = n252 & ~n8602 ;
  assign n9521 = ~n8600 & n9520 ;
  assign n9522 = \b[39]  & n250 ;
  assign n9523 = \a[3]  & \b[38]  ;
  assign n9524 = n241 & n9523 ;
  assign n9525 = ~n9522 & ~n9524 ;
  assign n9526 = \b[37]  & n303 ;
  assign n9527 = n300 & n9526 ;
  assign n9528 = ~\a[3]  & \b[38]  ;
  assign n9529 = n244 & n9528 ;
  assign n9530 = ~n9527 & ~n9529 ;
  assign n9531 = n9525 & n9530 ;
  assign n9532 = ~n9521 & n9531 ;
  assign n9533 = ~\a[5]  & ~n9532 ;
  assign n9534 = \a[5]  & n9531 ;
  assign n9535 = ~n9521 & n9534 ;
  assign n9536 = ~n9533 & ~n9535 ;
  assign n9537 = ~n9438 & ~n9440 ;
  assign n9538 = n430 & n7337 ;
  assign n9539 = ~n7334 & n9538 ;
  assign n9540 = n430 & ~n7337 ;
  assign n9541 = ~n6605 & n9540 ;
  assign n9542 = ~n7333 & n9541 ;
  assign n9543 = \b[34]  & n486 ;
  assign n9544 = n483 & n9543 ;
  assign n9545 = ~\a[5]  & \b[35]  ;
  assign n9546 = n485 & n9545 ;
  assign n9547 = ~n9544 & ~n9546 ;
  assign n9548 = \b[36]  & n428 ;
  assign n9549 = \a[6]  & \b[35]  ;
  assign n9550 = n419 & n9549 ;
  assign n9551 = \a[8]  & ~n9550 ;
  assign n9552 = ~n9548 & n9551 ;
  assign n9553 = n9547 & n9552 ;
  assign n9554 = ~n9542 & n9553 ;
  assign n9555 = ~n9539 & n9554 ;
  assign n9556 = ~n9548 & ~n9550 ;
  assign n9557 = n9547 & n9556 ;
  assign n9558 = ~n9542 & n9557 ;
  assign n9559 = ~n9539 & n9558 ;
  assign n9560 = ~\a[8]  & ~n9559 ;
  assign n9561 = ~n9555 & ~n9560 ;
  assign n9562 = ~n8981 & n9427 ;
  assign n9563 = n9422 & ~n9562 ;
  assign n9564 = n8987 & n9422 ;
  assign n9565 = n8666 & n9564 ;
  assign n9566 = ~n9563 & ~n9565 ;
  assign n9567 = n9130 & n9417 ;
  assign n9568 = ~n9416 & ~n9567 ;
  assign n9569 = ~n8919 & ~n9400 ;
  assign n9570 = ~n9148 & n9569 ;
  assign n9571 = n9405 & ~n9570 ;
  assign n9572 = n9372 & ~n9381 ;
  assign n9573 = ~n8868 & n9344 ;
  assign n9574 = ~n8876 & n9573 ;
  assign n9575 = n9339 & ~n9574 ;
  assign n9576 = n9175 & n9334 ;
  assign n9577 = n9333 & ~n9576 ;
  assign n9578 = n8824 & ~n9322 ;
  assign n9579 = ~n9195 & n9578 ;
  assign n9580 = ~n9321 & ~n9579 ;
  assign n9581 = ~n1233 & n4249 ;
  assign n9582 = ~n1231 & n9581 ;
  assign n9583 = \b[13]  & n4647 ;
  assign n9584 = n4644 & n9583 ;
  assign n9585 = ~\a[27]  & \b[14]  ;
  assign n9586 = n4241 & n9585 ;
  assign n9587 = ~n9584 & ~n9586 ;
  assign n9588 = \b[15]  & n4247 ;
  assign n9589 = \a[27]  & \b[14]  ;
  assign n9590 = n4238 & n9589 ;
  assign n9591 = \a[29]  & ~n9590 ;
  assign n9592 = ~n9588 & n9591 ;
  assign n9593 = n9587 & n9592 ;
  assign n9594 = ~n9582 & n9593 ;
  assign n9595 = ~n9588 & ~n9590 ;
  assign n9596 = n9587 & n9595 ;
  assign n9597 = ~n9582 & n9596 ;
  assign n9598 = ~\a[29]  & ~n9597 ;
  assign n9599 = ~n9594 & ~n9598 ;
  assign n9600 = ~n9315 & ~n9318 ;
  assign n9601 = ~n909 & ~n4909 ;
  assign n9602 = ~n5208 & n9601 ;
  assign n9603 = n906 & n9602 ;
  assign n9604 = n909 & ~n4909 ;
  assign n9605 = ~n5208 & n9604 ;
  assign n9606 = ~n906 & n9605 ;
  assign n9607 = ~n9603 & ~n9606 ;
  assign n9608 = \b[10]  & n5595 ;
  assign n9609 = n5592 & n9608 ;
  assign n9610 = ~\a[30]  & \b[11]  ;
  assign n9611 = n5203 & n9610 ;
  assign n9612 = ~n9609 & ~n9611 ;
  assign n9613 = \b[12]  & n5209 ;
  assign n9614 = \a[30]  & \b[11]  ;
  assign n9615 = n5200 & n9614 ;
  assign n9616 = \a[32]  & ~n9615 ;
  assign n9617 = ~n9613 & n9616 ;
  assign n9618 = n9612 & n9617 ;
  assign n9619 = n9607 & n9618 ;
  assign n9620 = ~n9613 & ~n9615 ;
  assign n9621 = n9612 & n9620 ;
  assign n9622 = n9607 & n9621 ;
  assign n9623 = ~\a[32]  & ~n9622 ;
  assign n9624 = ~n9619 & ~n9623 ;
  assign n9625 = ~n8768 & ~n9309 ;
  assign n9626 = ~n8770 & n9625 ;
  assign n9627 = ~n9310 & ~n9626 ;
  assign n9628 = n177 & n8759 ;
  assign n9629 = \b[3]  & n8757 ;
  assign n9630 = \a[38]  & \b[2]  ;
  assign n9631 = n9299 & n9630 ;
  assign n9632 = ~\a[39]  & \b[2]  ;
  assign n9633 = n8751 & n9632 ;
  assign n9634 = ~n9631 & ~n9633 ;
  assign n9635 = ~n9629 & n9634 ;
  assign n9636 = ~n9628 & n9635 ;
  assign n9637 = \b[1]  & n9301 ;
  assign n9638 = n9298 & n9637 ;
  assign n9639 = ~\a[41]  & ~n9638 ;
  assign n9640 = n9636 & n9639 ;
  assign n9641 = n9636 & ~n9638 ;
  assign n9642 = \a[41]  & ~n9641 ;
  assign n9643 = ~n9640 & ~n9642 ;
  assign n9644 = \a[41]  & ~\a[42]  ;
  assign n9645 = ~\a[41]  & \a[42]  ;
  assign n9646 = ~n9644 & ~n9645 ;
  assign n9647 = \b[0]  & ~n9646 ;
  assign n9648 = n9288 & n9305 ;
  assign n9649 = n9647 & n9648 ;
  assign n9650 = ~n9647 & ~n9648 ;
  assign n9651 = ~n9649 & ~n9650 ;
  assign n9652 = n9643 & n9651 ;
  assign n9653 = ~n9643 & ~n9651 ;
  assign n9654 = ~n9652 & ~n9653 ;
  assign n9655 = ~n323 & ~n7098 ;
  assign n9656 = ~n7531 & n9655 ;
  assign n9657 = n320 & n9656 ;
  assign n9658 = n323 & ~n7098 ;
  assign n9659 = ~n7531 & n9658 ;
  assign n9660 = ~n320 & n9659 ;
  assign n9661 = ~n9657 & ~n9660 ;
  assign n9662 = \b[4]  & n7973 ;
  assign n9663 = n7970 & n9662 ;
  assign n9664 = \b[6]  & n7532 ;
  assign n9665 = \a[35]  & \b[5]  ;
  assign n9666 = n7971 & n9665 ;
  assign n9667 = ~\a[36]  & \b[5]  ;
  assign n9668 = n7526 & n9667 ;
  assign n9669 = ~n9666 & ~n9668 ;
  assign n9670 = ~n9664 & n9669 ;
  assign n9671 = ~n9663 & n9670 ;
  assign n9672 = n9661 & n9671 ;
  assign n9673 = ~\a[38]  & ~n9672 ;
  assign n9674 = \a[38]  & n9671 ;
  assign n9675 = n9661 & n9674 ;
  assign n9676 = ~n9673 & ~n9675 ;
  assign n9677 = n9654 & ~n9676 ;
  assign n9678 = ~n9654 & n9676 ;
  assign n9679 = ~n9677 & ~n9678 ;
  assign n9680 = ~n9627 & ~n9679 ;
  assign n9681 = n9627 & n9679 ;
  assign n9682 = ~n9680 & ~n9681 ;
  assign n9683 = ~n589 & n6309 ;
  assign n9684 = ~n587 & n9683 ;
  assign n9685 = \b[7]  & n6778 ;
  assign n9686 = n6775 & n9685 ;
  assign n9687 = \b[9]  & n6307 ;
  assign n9688 = \a[33]  & \b[8]  ;
  assign n9689 = n6298 & n9688 ;
  assign n9690 = ~\a[33]  & \b[8]  ;
  assign n9691 = n6301 & n9690 ;
  assign n9692 = ~n9689 & ~n9691 ;
  assign n9693 = ~n9687 & n9692 ;
  assign n9694 = ~n9686 & n9693 ;
  assign n9695 = ~\a[35]  & n9694 ;
  assign n9696 = ~n9684 & n9695 ;
  assign n9697 = ~n9684 & n9694 ;
  assign n9698 = \a[35]  & ~n9697 ;
  assign n9699 = ~n9696 & ~n9698 ;
  assign n9700 = ~n9682 & ~n9699 ;
  assign n9701 = n9682 & n9699 ;
  assign n9702 = ~n9700 & ~n9701 ;
  assign n9703 = ~n9624 & ~n9702 ;
  assign n9704 = ~n9600 & n9703 ;
  assign n9705 = ~n9624 & n9702 ;
  assign n9706 = n9600 & n9705 ;
  assign n9707 = ~n9704 & ~n9706 ;
  assign n9708 = n9624 & ~n9702 ;
  assign n9709 = n9600 & n9708 ;
  assign n9710 = n9624 & n9702 ;
  assign n9711 = ~n9600 & n9710 ;
  assign n9712 = ~n9709 & ~n9711 ;
  assign n9713 = n9707 & n9712 ;
  assign n9714 = ~n9599 & ~n9713 ;
  assign n9715 = n9580 & n9714 ;
  assign n9716 = ~n9599 & n9713 ;
  assign n9717 = ~n9580 & n9716 ;
  assign n9718 = ~n9715 & ~n9717 ;
  assign n9719 = n9599 & ~n9713 ;
  assign n9720 = ~n9580 & n9719 ;
  assign n9721 = n9599 & n9713 ;
  assign n9722 = n9580 & n9721 ;
  assign n9723 = ~n9720 & ~n9722 ;
  assign n9724 = n9718 & n9723 ;
  assign n9725 = ~n9577 & n9724 ;
  assign n9726 = n1875 & n3402 ;
  assign n9727 = ~n1872 & n9726 ;
  assign n9728 = n3402 & n5000 ;
  assign n9729 = ~n1871 & n9728 ;
  assign n9730 = \b[16]  & n3733 ;
  assign n9731 = n3730 & n9730 ;
  assign n9732 = ~\a[24]  & \b[17]  ;
  assign n9733 = n3394 & n9732 ;
  assign n9734 = ~n9731 & ~n9733 ;
  assign n9735 = \b[18]  & n3400 ;
  assign n9736 = \a[24]  & \b[17]  ;
  assign n9737 = n3391 & n9736 ;
  assign n9738 = \a[26]  & ~n9737 ;
  assign n9739 = ~n9735 & n9738 ;
  assign n9740 = n9734 & n9739 ;
  assign n9741 = ~n9729 & n9740 ;
  assign n9742 = ~n9727 & n9741 ;
  assign n9743 = ~n9735 & ~n9737 ;
  assign n9744 = n9734 & n9743 ;
  assign n9745 = ~n9729 & n9744 ;
  assign n9746 = ~n9727 & n9745 ;
  assign n9747 = ~\a[26]  & ~n9746 ;
  assign n9748 = ~n9742 & ~n9747 ;
  assign n9749 = n9333 & ~n9724 ;
  assign n9750 = ~n9576 & n9749 ;
  assign n9751 = ~n9748 & ~n9750 ;
  assign n9752 = ~n9725 & n9751 ;
  assign n9753 = ~n9724 & n9748 ;
  assign n9754 = n9577 & n9753 ;
  assign n9755 = n9724 & n9748 ;
  assign n9756 = ~n9577 & n9755 ;
  assign n9757 = ~n9754 & ~n9756 ;
  assign n9758 = ~n9752 & n9757 ;
  assign n9759 = n9575 & n9758 ;
  assign n9760 = ~n9575 & ~n9758 ;
  assign n9761 = ~n9759 & ~n9760 ;
  assign n9762 = ~n2523 & n2622 ;
  assign n9763 = ~n2521 & n9762 ;
  assign n9764 = \b[19]  & n2912 ;
  assign n9765 = n2909 & n9764 ;
  assign n9766 = \b[21]  & n2620 ;
  assign n9767 = \a[20]  & \b[20]  ;
  assign n9768 = n2910 & n9767 ;
  assign n9769 = ~\a[21]  & \b[20]  ;
  assign n9770 = n2614 & n9769 ;
  assign n9771 = ~n9768 & ~n9770 ;
  assign n9772 = ~n9766 & n9771 ;
  assign n9773 = ~n9765 & n9772 ;
  assign n9774 = ~n9763 & n9773 ;
  assign n9775 = ~\a[23]  & ~n9774 ;
  assign n9776 = \a[23]  & n9773 ;
  assign n9777 = ~n9763 & n9776 ;
  assign n9778 = ~n9775 & ~n9777 ;
  assign n9779 = n9761 & ~n9778 ;
  assign n9780 = ~n9761 & n9778 ;
  assign n9781 = ~n9779 & ~n9780 ;
  assign n9782 = n1965 & n3283 ;
  assign n9783 = ~n3280 & n9782 ;
  assign n9784 = n1965 & n4107 ;
  assign n9785 = ~n3279 & n9784 ;
  assign n9786 = \b[22]  & n2218 ;
  assign n9787 = n2216 & n9786 ;
  assign n9788 = ~\a[18]  & \b[23]  ;
  assign n9789 = n1957 & n9788 ;
  assign n9790 = ~n9787 & ~n9789 ;
  assign n9791 = \b[24]  & n1963 ;
  assign n9792 = \a[18]  & \b[23]  ;
  assign n9793 = n2210 & n9792 ;
  assign n9794 = \a[20]  & ~n9793 ;
  assign n9795 = ~n9791 & n9794 ;
  assign n9796 = n9790 & n9795 ;
  assign n9797 = ~n9785 & n9796 ;
  assign n9798 = ~n9783 & n9797 ;
  assign n9799 = ~n9791 & ~n9793 ;
  assign n9800 = n9790 & n9799 ;
  assign n9801 = ~n9785 & n9800 ;
  assign n9802 = ~n9783 & n9801 ;
  assign n9803 = ~\a[20]  & ~n9802 ;
  assign n9804 = ~n9798 & ~n9803 ;
  assign n9805 = ~n9781 & n9804 ;
  assign n9806 = n9572 & n9805 ;
  assign n9807 = n9781 & n9804 ;
  assign n9808 = ~n9572 & n9807 ;
  assign n9809 = ~n9806 & ~n9808 ;
  assign n9810 = ~n9781 & ~n9804 ;
  assign n9811 = ~n9572 & n9810 ;
  assign n9812 = n9781 & ~n9804 ;
  assign n9813 = n9572 & n9812 ;
  assign n9814 = ~n9811 & ~n9813 ;
  assign n9815 = n9809 & n9814 ;
  assign n9816 = ~n9571 & ~n9815 ;
  assign n9817 = n9405 & n9815 ;
  assign n9818 = ~n9570 & n9817 ;
  assign n9819 = n1467 & ~n4148 ;
  assign n9820 = ~n4146 & n9819 ;
  assign n9821 = \b[25]  & n1652 ;
  assign n9822 = n1649 & n9821 ;
  assign n9823 = ~\a[15]  & \b[26]  ;
  assign n9824 = n1459 & n9823 ;
  assign n9825 = ~n9822 & ~n9824 ;
  assign n9826 = \b[27]  & n1465 ;
  assign n9827 = \a[15]  & \b[26]  ;
  assign n9828 = n1456 & n9827 ;
  assign n9829 = \a[17]  & ~n9828 ;
  assign n9830 = ~n9826 & n9829 ;
  assign n9831 = n9825 & n9830 ;
  assign n9832 = ~n9820 & n9831 ;
  assign n9833 = ~n9826 & ~n9828 ;
  assign n9834 = n9825 & n9833 ;
  assign n9835 = ~n9820 & n9834 ;
  assign n9836 = ~\a[17]  & ~n9835 ;
  assign n9837 = ~n9832 & ~n9836 ;
  assign n9838 = ~n9818 & ~n9837 ;
  assign n9839 = ~n9816 & n9838 ;
  assign n9840 = ~n9815 & n9837 ;
  assign n9841 = ~n9571 & n9840 ;
  assign n9842 = n9815 & n9837 ;
  assign n9843 = n9571 & n9842 ;
  assign n9844 = ~n9841 & ~n9843 ;
  assign n9845 = ~n9839 & n9844 ;
  assign n9846 = ~n9568 & n9845 ;
  assign n9847 = n999 & n5105 ;
  assign n9848 = ~n5102 & n9847 ;
  assign n9849 = n999 & ~n5105 ;
  assign n9850 = ~n4497 & n9849 ;
  assign n9851 = ~n5101 & n9850 ;
  assign n9852 = \b[28]  & n1182 ;
  assign n9853 = n1179 & n9852 ;
  assign n9854 = \b[30]  & n997 ;
  assign n9855 = \a[11]  & \b[29]  ;
  assign n9856 = n1180 & n9855 ;
  assign n9857 = ~\a[12]  & \b[29]  ;
  assign n9858 = n7674 & n9857 ;
  assign n9859 = ~n9856 & ~n9858 ;
  assign n9860 = ~n9854 & n9859 ;
  assign n9861 = ~n9853 & n9860 ;
  assign n9862 = ~n9851 & n9861 ;
  assign n9863 = ~n9848 & n9862 ;
  assign n9864 = ~\a[14]  & ~n9863 ;
  assign n9865 = \a[14]  & n9861 ;
  assign n9866 = ~n9851 & n9865 ;
  assign n9867 = ~n9848 & n9866 ;
  assign n9868 = ~n9864 & ~n9867 ;
  assign n9869 = ~n9416 & ~n9845 ;
  assign n9870 = ~n9567 & n9869 ;
  assign n9871 = ~n9868 & ~n9870 ;
  assign n9872 = ~n9846 & n9871 ;
  assign n9873 = ~n9845 & n9868 ;
  assign n9874 = n9568 & n9873 ;
  assign n9875 = n9845 & n9868 ;
  assign n9876 = ~n9568 & n9875 ;
  assign n9877 = ~n9874 & ~n9876 ;
  assign n9878 = ~n9872 & n9877 ;
  assign n9879 = ~n9566 & n9878 ;
  assign n9880 = n9566 & ~n9878 ;
  assign n9881 = ~n9879 & ~n9880 ;
  assign n9882 = n646 & ~n5855 ;
  assign n9883 = ~n5853 & n9882 ;
  assign n9884 = \b[31]  & n796 ;
  assign n9885 = n793 & n9884 ;
  assign n9886 = \b[33]  & n644 ;
  assign n9887 = \a[8]  & \b[32]  ;
  assign n9888 = n794 & n9887 ;
  assign n9889 = ~\a[9]  & \b[32]  ;
  assign n9890 = n638 & n9889 ;
  assign n9891 = ~n9888 & ~n9890 ;
  assign n9892 = ~n9886 & n9891 ;
  assign n9893 = ~n9885 & n9892 ;
  assign n9894 = ~n9883 & n9893 ;
  assign n9895 = ~\a[11]  & ~n9894 ;
  assign n9896 = \a[11]  & n9893 ;
  assign n9897 = ~n9883 & n9896 ;
  assign n9898 = ~n9895 & ~n9897 ;
  assign n9899 = n9881 & ~n9898 ;
  assign n9900 = ~n9881 & n9898 ;
  assign n9901 = ~n9899 & ~n9900 ;
  assign n9902 = n9561 & ~n9901 ;
  assign n9903 = n9537 & n9902 ;
  assign n9904 = n9561 & n9901 ;
  assign n9905 = ~n9537 & n9904 ;
  assign n9906 = ~n9903 & ~n9905 ;
  assign n9907 = ~n9561 & ~n9901 ;
  assign n9908 = ~n9537 & n9907 ;
  assign n9909 = ~n9561 & n9901 ;
  assign n9910 = n9537 & n9909 ;
  assign n9911 = ~n9908 & ~n9910 ;
  assign n9912 = n9906 & n9911 ;
  assign n9913 = ~n9536 & ~n9912 ;
  assign n9914 = n9519 & n9913 ;
  assign n9915 = ~n9536 & n9912 ;
  assign n9916 = ~n9519 & n9915 ;
  assign n9917 = ~n9914 & ~n9916 ;
  assign n9918 = n9536 & ~n9912 ;
  assign n9919 = ~n9519 & n9918 ;
  assign n9920 = n9536 & n9912 ;
  assign n9921 = n9519 & n9920 ;
  assign n9922 = ~n9919 & ~n9921 ;
  assign n9923 = n9917 & n9922 ;
  assign n9924 = ~n9516 & n9923 ;
  assign n9925 = ~n9043 & ~n9478 ;
  assign n9926 = ~n9475 & n9925 ;
  assign n9927 = ~n9477 & ~n9926 ;
  assign n9928 = ~\b[41]  & ~\b[42]  ;
  assign n9929 = \b[41]  & \b[42]  ;
  assign n9930 = ~n9928 & ~n9929 ;
  assign n9931 = n134 & n9930 ;
  assign n9932 = ~n9927 & n9931 ;
  assign n9933 = n134 & ~n9930 ;
  assign n9934 = ~n9477 & n9933 ;
  assign n9935 = ~n9926 & n9934 ;
  assign n9936 = \a[0]  & \b[42]  ;
  assign n9937 = n133 & n9936 ;
  assign n9938 = \b[41]  & n141 ;
  assign n9939 = ~\a[1]  & \b[40]  ;
  assign n9940 = n1521 & n9939 ;
  assign n9941 = ~n9938 & ~n9940 ;
  assign n9942 = ~n9937 & n9941 ;
  assign n9943 = \a[2]  & n9942 ;
  assign n9944 = ~n9935 & n9943 ;
  assign n9945 = ~n9932 & n9944 ;
  assign n9946 = ~n9935 & n9942 ;
  assign n9947 = ~n9932 & n9946 ;
  assign n9948 = ~\a[2]  & ~n9947 ;
  assign n9949 = ~n9945 & ~n9948 ;
  assign n9950 = n9467 & ~n9923 ;
  assign n9951 = ~n9515 & n9950 ;
  assign n9952 = ~n9949 & ~n9951 ;
  assign n9953 = ~n9924 & n9952 ;
  assign n9954 = ~n9923 & n9949 ;
  assign n9955 = n9516 & n9954 ;
  assign n9956 = n9923 & n9949 ;
  assign n9957 = ~n9516 & n9956 ;
  assign n9958 = ~n9955 & ~n9957 ;
  assign n9959 = ~n9953 & n9958 ;
  assign n9960 = n9514 & n9959 ;
  assign n9961 = ~n9514 & ~n9959 ;
  assign n9962 = ~n9960 & ~n9961 ;
  assign n9963 = ~n9953 & ~n9960 ;
  assign n9964 = n9467 & n9917 ;
  assign n9965 = ~n9515 & n9964 ;
  assign n9966 = n9922 & ~n9965 ;
  assign n9967 = n9519 & n9912 ;
  assign n9968 = n9911 & ~n9967 ;
  assign n9969 = n252 & n9044 ;
  assign n9970 = ~n9041 & n9969 ;
  assign n9971 = n252 & ~n9044 ;
  assign n9972 = ~n8597 & n9971 ;
  assign n9973 = ~n9040 & n9972 ;
  assign n9974 = \b[38]  & n303 ;
  assign n9975 = n300 & n9974 ;
  assign n9976 = ~\a[3]  & \b[39]  ;
  assign n9977 = n244 & n9976 ;
  assign n9978 = ~n9975 & ~n9977 ;
  assign n9979 = \b[40]  & n250 ;
  assign n9980 = \a[3]  & \b[39]  ;
  assign n9981 = n241 & n9980 ;
  assign n9982 = \a[5]  & ~n9981 ;
  assign n9983 = ~n9979 & n9982 ;
  assign n9984 = n9978 & n9983 ;
  assign n9985 = ~n9973 & n9984 ;
  assign n9986 = ~n9970 & n9985 ;
  assign n9987 = ~n9979 & ~n9981 ;
  assign n9988 = n9978 & n9987 ;
  assign n9989 = ~n9973 & n9988 ;
  assign n9990 = ~n9970 & n9989 ;
  assign n9991 = ~\a[5]  & ~n9990 ;
  assign n9992 = ~n9986 & ~n9991 ;
  assign n9993 = ~n9438 & ~n9899 ;
  assign n9994 = ~n9440 & n9993 ;
  assign n9995 = ~n9900 & ~n9994 ;
  assign n9996 = ~n9872 & ~n9879 ;
  assign n9997 = ~n9416 & ~n9839 ;
  assign n9998 = ~n9567 & n9997 ;
  assign n9999 = n9844 & ~n9998 ;
  assign n10000 = n999 & ~n5462 ;
  assign n10001 = ~n5460 & n10000 ;
  assign n10002 = \b[29]  & n1182 ;
  assign n10003 = n1179 & n10002 ;
  assign n10004 = \b[31]  & n997 ;
  assign n10005 = \a[11]  & \b[30]  ;
  assign n10006 = n1180 & n10005 ;
  assign n10007 = ~\a[12]  & \b[30]  ;
  assign n10008 = n7674 & n10007 ;
  assign n10009 = ~n10006 & ~n10008 ;
  assign n10010 = ~n10004 & n10009 ;
  assign n10011 = ~n10003 & n10010 ;
  assign n10012 = ~n10001 & n10011 ;
  assign n10013 = ~\a[14]  & ~n10012 ;
  assign n10014 = \a[14]  & n10011 ;
  assign n10015 = ~n10001 & n10014 ;
  assign n10016 = ~n10013 & ~n10015 ;
  assign n10017 = n9814 & ~n9818 ;
  assign n10018 = n9372 & ~n9779 ;
  assign n10019 = ~n9381 & n10018 ;
  assign n10020 = ~n9780 & ~n10019 ;
  assign n10021 = ~n9752 & ~n9759 ;
  assign n10022 = n9333 & n9718 ;
  assign n10023 = ~n9576 & n10022 ;
  assign n10024 = n9723 & ~n10023 ;
  assign n10025 = n9580 & n9713 ;
  assign n10026 = n9707 & ~n10025 ;
  assign n10027 = ~n9315 & ~n9701 ;
  assign n10028 = ~n9318 & n10027 ;
  assign n10029 = ~n9700 & ~n10028 ;
  assign n10030 = ~n951 & n5211 ;
  assign n10031 = ~n949 & n10030 ;
  assign n10032 = \b[11]  & n5595 ;
  assign n10033 = n5592 & n10032 ;
  assign n10034 = ~\a[30]  & \b[12]  ;
  assign n10035 = n5203 & n10034 ;
  assign n10036 = ~n10033 & ~n10035 ;
  assign n10037 = \b[13]  & n5209 ;
  assign n10038 = \a[30]  & \b[12]  ;
  assign n10039 = n5200 & n10038 ;
  assign n10040 = \a[32]  & ~n10039 ;
  assign n10041 = ~n10037 & n10040 ;
  assign n10042 = n10036 & n10041 ;
  assign n10043 = ~n10031 & n10042 ;
  assign n10044 = ~n10037 & ~n10039 ;
  assign n10045 = n10036 & n10044 ;
  assign n10046 = ~n10031 & n10045 ;
  assign n10047 = ~\a[32]  & ~n10046 ;
  assign n10048 = ~n10043 & ~n10047 ;
  assign n10049 = ~n9677 & ~n9681 ;
  assign n10050 = ~n9649 & ~n9652 ;
  assign n10051 = n222 & n8759 ;
  assign n10052 = \b[4]  & n8757 ;
  assign n10053 = \a[38]  & \b[3]  ;
  assign n10054 = n9299 & n10053 ;
  assign n10055 = ~\a[39]  & \b[3]  ;
  assign n10056 = n8751 & n10055 ;
  assign n10057 = ~n10054 & ~n10056 ;
  assign n10058 = ~n10052 & n10057 ;
  assign n10059 = \b[2]  & n9301 ;
  assign n10060 = n9298 & n10059 ;
  assign n10061 = \a[41]  & ~n10060 ;
  assign n10062 = n10058 & n10061 ;
  assign n10063 = ~n10051 & n10062 ;
  assign n10064 = n10058 & ~n10060 ;
  assign n10065 = ~n10051 & n10064 ;
  assign n10066 = ~\a[41]  & ~n10065 ;
  assign n10067 = ~n10063 & ~n10066 ;
  assign n10068 = \a[44]  & \b[0]  ;
  assign n10069 = ~n9646 & n10068 ;
  assign n10070 = \a[42]  & \b[0]  ;
  assign n10071 = \a[41]  & ~\a[43]  ;
  assign n10072 = n10070 & n10071 ;
  assign n10073 = ~\a[42]  & \b[0]  ;
  assign n10074 = ~\a[41]  & \a[43]  ;
  assign n10075 = n10073 & n10074 ;
  assign n10076 = ~n10072 & ~n10075 ;
  assign n10077 = \a[43]  & ~\a[44]  ;
  assign n10078 = ~\a[43]  & \a[44]  ;
  assign n10079 = ~n10077 & ~n10078 ;
  assign n10080 = ~n9646 & n10079 ;
  assign n10081 = \b[1]  & n10080 ;
  assign n10082 = ~n9646 & ~n10079 ;
  assign n10083 = ~n137 & n10082 ;
  assign n10084 = ~n10081 & ~n10083 ;
  assign n10085 = n10076 & n10084 ;
  assign n10086 = n10069 & ~n10085 ;
  assign n10087 = ~n10069 & n10076 ;
  assign n10088 = n10084 & n10087 ;
  assign n10089 = ~n10086 & ~n10088 ;
  assign n10090 = n10067 & ~n10089 ;
  assign n10091 = ~n10067 & n10089 ;
  assign n10092 = ~n10090 & ~n10091 ;
  assign n10093 = ~n10050 & n10092 ;
  assign n10094 = n10050 & ~n10092 ;
  assign n10095 = ~n10093 & ~n10094 ;
  assign n10096 = ~n383 & n7534 ;
  assign n10097 = ~n381 & n10096 ;
  assign n10098 = \b[5]  & n7973 ;
  assign n10099 = n7970 & n10098 ;
  assign n10100 = \b[7]  & n7532 ;
  assign n10101 = \a[35]  & \b[6]  ;
  assign n10102 = n7971 & n10101 ;
  assign n10103 = ~\a[36]  & \b[6]  ;
  assign n10104 = n7526 & n10103 ;
  assign n10105 = ~n10102 & ~n10104 ;
  assign n10106 = ~n10100 & n10105 ;
  assign n10107 = ~n10099 & n10106 ;
  assign n10108 = ~\a[38]  & n10107 ;
  assign n10109 = ~n10097 & n10108 ;
  assign n10110 = ~n10097 & n10107 ;
  assign n10111 = \a[38]  & ~n10110 ;
  assign n10112 = ~n10109 & ~n10111 ;
  assign n10113 = n10095 & n10112 ;
  assign n10114 = ~n10095 & ~n10112 ;
  assign n10115 = ~n10113 & ~n10114 ;
  assign n10116 = ~n685 & ~n5952 ;
  assign n10117 = ~n6306 & n10116 ;
  assign n10118 = n682 & n10117 ;
  assign n10119 = n685 & ~n5952 ;
  assign n10120 = ~n6306 & n10119 ;
  assign n10121 = ~n682 & n10120 ;
  assign n10122 = ~n10118 & ~n10121 ;
  assign n10123 = \b[8]  & n6778 ;
  assign n10124 = n6775 & n10123 ;
  assign n10125 = \b[10]  & n6307 ;
  assign n10126 = \a[33]  & \b[9]  ;
  assign n10127 = n6298 & n10126 ;
  assign n10128 = ~\a[33]  & \b[9]  ;
  assign n10129 = n6301 & n10128 ;
  assign n10130 = ~n10127 & ~n10129 ;
  assign n10131 = ~n10125 & n10130 ;
  assign n10132 = ~n10124 & n10131 ;
  assign n10133 = n10122 & n10132 ;
  assign n10134 = ~\a[35]  & ~n10133 ;
  assign n10135 = \a[35]  & n10132 ;
  assign n10136 = n10122 & n10135 ;
  assign n10137 = ~n10134 & ~n10136 ;
  assign n10138 = ~n10115 & ~n10137 ;
  assign n10139 = ~n10049 & n10138 ;
  assign n10140 = n10115 & ~n10137 ;
  assign n10141 = n10049 & n10140 ;
  assign n10142 = ~n10139 & ~n10141 ;
  assign n10143 = ~n10115 & n10137 ;
  assign n10144 = n10049 & n10143 ;
  assign n10145 = n10115 & n10137 ;
  assign n10146 = ~n10049 & n10145 ;
  assign n10147 = ~n10144 & ~n10146 ;
  assign n10148 = n10142 & n10147 ;
  assign n10149 = n10048 & ~n10148 ;
  assign n10150 = ~n10029 & n10149 ;
  assign n10151 = n10048 & n10148 ;
  assign n10152 = n10029 & n10151 ;
  assign n10153 = ~n10150 & ~n10152 ;
  assign n10154 = ~n10048 & ~n10148 ;
  assign n10155 = n10029 & n10154 ;
  assign n10156 = ~n10048 & n10148 ;
  assign n10157 = ~n10029 & n10156 ;
  assign n10158 = ~n10155 & ~n10157 ;
  assign n10159 = n10153 & n10158 ;
  assign n10160 = ~n10026 & n10159 ;
  assign n10161 = n9707 & ~n10159 ;
  assign n10162 = ~n10025 & n10161 ;
  assign n10163 = n1512 & n4249 ;
  assign n10164 = ~n1509 & n10163 ;
  assign n10165 = ~n1228 & ~n1512 ;
  assign n10166 = n4249 & n10165 ;
  assign n10167 = ~n1508 & n10166 ;
  assign n10168 = \b[14]  & n4647 ;
  assign n10169 = n4644 & n10168 ;
  assign n10170 = ~\a[27]  & \b[15]  ;
  assign n10171 = n4241 & n10170 ;
  assign n10172 = ~n10169 & ~n10171 ;
  assign n10173 = \b[16]  & n4247 ;
  assign n10174 = \a[27]  & \b[15]  ;
  assign n10175 = n4238 & n10174 ;
  assign n10176 = \a[29]  & ~n10175 ;
  assign n10177 = ~n10173 & n10176 ;
  assign n10178 = n10172 & n10177 ;
  assign n10179 = ~n10167 & n10178 ;
  assign n10180 = ~n10164 & n10179 ;
  assign n10181 = ~n10173 & ~n10175 ;
  assign n10182 = n10172 & n10181 ;
  assign n10183 = ~n10167 & n10182 ;
  assign n10184 = ~n10164 & n10183 ;
  assign n10185 = ~\a[29]  & ~n10184 ;
  assign n10186 = ~n10180 & ~n10185 ;
  assign n10187 = ~n10162 & ~n10186 ;
  assign n10188 = ~n10160 & n10187 ;
  assign n10189 = ~n10159 & n10186 ;
  assign n10190 = n10026 & n10189 ;
  assign n10191 = n10159 & n10186 ;
  assign n10192 = ~n10026 & n10191 ;
  assign n10193 = ~n10190 & ~n10192 ;
  assign n10194 = ~n10188 & n10193 ;
  assign n10195 = ~n2079 & n3402 ;
  assign n10196 = ~n2077 & n10195 ;
  assign n10197 = \b[17]  & n3733 ;
  assign n10198 = n3730 & n10197 ;
  assign n10199 = ~\a[24]  & \b[18]  ;
  assign n10200 = n3394 & n10199 ;
  assign n10201 = ~n10198 & ~n10200 ;
  assign n10202 = \b[19]  & n3400 ;
  assign n10203 = \a[24]  & \b[18]  ;
  assign n10204 = n3391 & n10203 ;
  assign n10205 = \a[26]  & ~n10204 ;
  assign n10206 = ~n10202 & n10205 ;
  assign n10207 = n10201 & n10206 ;
  assign n10208 = ~n10196 & n10207 ;
  assign n10209 = ~n10202 & ~n10204 ;
  assign n10210 = n10201 & n10209 ;
  assign n10211 = ~n10196 & n10210 ;
  assign n10212 = ~\a[26]  & ~n10211 ;
  assign n10213 = ~n10208 & ~n10212 ;
  assign n10214 = ~n10194 & ~n10213 ;
  assign n10215 = n10024 & n10214 ;
  assign n10216 = n10194 & ~n10213 ;
  assign n10217 = ~n10024 & n10216 ;
  assign n10218 = ~n10215 & ~n10217 ;
  assign n10219 = ~n10194 & n10213 ;
  assign n10220 = ~n10024 & n10219 ;
  assign n10221 = n10194 & n10213 ;
  assign n10222 = n10024 & n10221 ;
  assign n10223 = ~n10220 & ~n10222 ;
  assign n10224 = n10218 & n10223 ;
  assign n10225 = n2622 & ~n2771 ;
  assign n10226 = ~n2769 & n10225 ;
  assign n10227 = \b[20]  & n2912 ;
  assign n10228 = n2909 & n10227 ;
  assign n10229 = \b[22]  & n2620 ;
  assign n10230 = \a[20]  & \b[21]  ;
  assign n10231 = n2910 & n10230 ;
  assign n10232 = ~\a[21]  & \b[21]  ;
  assign n10233 = n2614 & n10232 ;
  assign n10234 = ~n10231 & ~n10233 ;
  assign n10235 = ~n10229 & n10234 ;
  assign n10236 = ~n10228 & n10235 ;
  assign n10237 = ~n10226 & n10236 ;
  assign n10238 = ~\a[23]  & ~n10237 ;
  assign n10239 = \a[23]  & n10236 ;
  assign n10240 = ~n10226 & n10239 ;
  assign n10241 = ~n10238 & ~n10240 ;
  assign n10242 = ~n10224 & ~n10241 ;
  assign n10243 = ~n10021 & n10242 ;
  assign n10244 = n10224 & ~n10241 ;
  assign n10245 = n10021 & n10244 ;
  assign n10246 = ~n10243 & ~n10245 ;
  assign n10247 = ~n10224 & n10241 ;
  assign n10248 = n10021 & n10247 ;
  assign n10249 = n10224 & n10241 ;
  assign n10250 = ~n10021 & n10249 ;
  assign n10251 = ~n10248 & ~n10250 ;
  assign n10252 = n10246 & n10251 ;
  assign n10253 = n1965 & ~n3567 ;
  assign n10254 = ~n3565 & n10253 ;
  assign n10255 = \b[25]  & n1963 ;
  assign n10256 = \a[18]  & \b[24]  ;
  assign n10257 = n2210 & n10256 ;
  assign n10258 = ~n10255 & ~n10257 ;
  assign n10259 = \b[23]  & n2218 ;
  assign n10260 = n2216 & n10259 ;
  assign n10261 = ~\a[18]  & \b[24]  ;
  assign n10262 = n1957 & n10261 ;
  assign n10263 = ~n10260 & ~n10262 ;
  assign n10264 = n10258 & n10263 ;
  assign n10265 = ~n10254 & n10264 ;
  assign n10266 = ~\a[20]  & ~n10265 ;
  assign n10267 = \a[20]  & n10264 ;
  assign n10268 = ~n10254 & n10267 ;
  assign n10269 = ~n10266 & ~n10268 ;
  assign n10270 = ~n10252 & ~n10269 ;
  assign n10271 = n10020 & n10270 ;
  assign n10272 = n10252 & ~n10269 ;
  assign n10273 = ~n10020 & n10272 ;
  assign n10274 = ~n10271 & ~n10273 ;
  assign n10275 = ~n10252 & n10269 ;
  assign n10276 = ~n10020 & n10275 ;
  assign n10277 = n10252 & n10269 ;
  assign n10278 = n10020 & n10277 ;
  assign n10279 = ~n10276 & ~n10278 ;
  assign n10280 = n10274 & n10279 ;
  assign n10281 = ~n10017 & n10280 ;
  assign n10282 = n1467 & n4456 ;
  assign n10283 = ~n4453 & n10282 ;
  assign n10284 = n1467 & ~n4456 ;
  assign n10285 = ~n4143 & n10284 ;
  assign n10286 = ~n4452 & n10285 ;
  assign n10287 = \b[26]  & n1652 ;
  assign n10288 = n1649 & n10287 ;
  assign n10289 = ~\a[15]  & \b[27]  ;
  assign n10290 = n1459 & n10289 ;
  assign n10291 = ~n10288 & ~n10290 ;
  assign n10292 = \b[28]  & n1465 ;
  assign n10293 = \a[15]  & \b[27]  ;
  assign n10294 = n1456 & n10293 ;
  assign n10295 = \a[17]  & ~n10294 ;
  assign n10296 = ~n10292 & n10295 ;
  assign n10297 = n10291 & n10296 ;
  assign n10298 = ~n10286 & n10297 ;
  assign n10299 = ~n10283 & n10298 ;
  assign n10300 = ~n10292 & ~n10294 ;
  assign n10301 = n10291 & n10300 ;
  assign n10302 = ~n10286 & n10301 ;
  assign n10303 = ~n10283 & n10302 ;
  assign n10304 = ~\a[17]  & ~n10303 ;
  assign n10305 = ~n10299 & ~n10304 ;
  assign n10306 = n9814 & ~n10280 ;
  assign n10307 = ~n9818 & n10306 ;
  assign n10308 = ~n10305 & ~n10307 ;
  assign n10309 = ~n10281 & n10308 ;
  assign n10310 = ~n10280 & n10305 ;
  assign n10311 = n10017 & n10310 ;
  assign n10312 = n10280 & n10305 ;
  assign n10313 = ~n10017 & n10312 ;
  assign n10314 = ~n10311 & ~n10313 ;
  assign n10315 = ~n10309 & n10314 ;
  assign n10316 = n10016 & ~n10315 ;
  assign n10317 = ~n9999 & n10316 ;
  assign n10318 = n10016 & n10315 ;
  assign n10319 = n9999 & n10318 ;
  assign n10320 = ~n10317 & ~n10319 ;
  assign n10321 = ~n9999 & ~n10315 ;
  assign n10322 = n9844 & n10315 ;
  assign n10323 = ~n9998 & n10322 ;
  assign n10324 = ~n10016 & ~n10323 ;
  assign n10325 = ~n10321 & n10324 ;
  assign n10326 = n10320 & ~n10325 ;
  assign n10327 = ~n551 & ~n5850 ;
  assign n10328 = ~n6565 & n10327 ;
  assign n10329 = ~n6561 & n10328 ;
  assign n10330 = ~n643 & n10329 ;
  assign n10331 = n646 & n6565 ;
  assign n10332 = ~n6562 & n10331 ;
  assign n10333 = ~n10330 & ~n10332 ;
  assign n10334 = \b[32]  & n796 ;
  assign n10335 = n793 & n10334 ;
  assign n10336 = ~\a[9]  & \b[33]  ;
  assign n10337 = n638 & n10336 ;
  assign n10338 = ~n10335 & ~n10337 ;
  assign n10339 = \b[34]  & n644 ;
  assign n10340 = \a[9]  & \b[33]  ;
  assign n10341 = n635 & n10340 ;
  assign n10342 = \a[11]  & ~n10341 ;
  assign n10343 = ~n10339 & n10342 ;
  assign n10344 = n10338 & n10343 ;
  assign n10345 = n10333 & n10344 ;
  assign n10346 = ~n10339 & ~n10341 ;
  assign n10347 = n10338 & n10346 ;
  assign n10348 = n10333 & n10347 ;
  assign n10349 = ~\a[11]  & ~n10348 ;
  assign n10350 = ~n10345 & ~n10349 ;
  assign n10351 = ~n10326 & ~n10350 ;
  assign n10352 = ~n9996 & n10351 ;
  assign n10353 = n10326 & ~n10350 ;
  assign n10354 = n9996 & n10353 ;
  assign n10355 = ~n10352 & ~n10354 ;
  assign n10356 = ~n10326 & n10350 ;
  assign n10357 = n9996 & n10356 ;
  assign n10358 = n10326 & n10350 ;
  assign n10359 = ~n9996 & n10358 ;
  assign n10360 = ~n10357 & ~n10359 ;
  assign n10361 = n10355 & n10360 ;
  assign n10362 = n430 & ~n7761 ;
  assign n10363 = ~n7759 & n10362 ;
  assign n10364 = \b[35]  & n486 ;
  assign n10365 = n483 & n10364 ;
  assign n10366 = \b[37]  & n428 ;
  assign n10367 = \a[6]  & \b[36]  ;
  assign n10368 = n419 & n10367 ;
  assign n10369 = ~\a[6]  & \b[36]  ;
  assign n10370 = n422 & n10369 ;
  assign n10371 = ~n10368 & ~n10370 ;
  assign n10372 = ~n10366 & n10371 ;
  assign n10373 = ~n10365 & n10372 ;
  assign n10374 = ~n10363 & n10373 ;
  assign n10375 = ~\a[8]  & ~n10374 ;
  assign n10376 = \a[8]  & n10373 ;
  assign n10377 = ~n10363 & n10376 ;
  assign n10378 = ~n10375 & ~n10377 ;
  assign n10379 = ~n10361 & ~n10378 ;
  assign n10380 = n9995 & n10379 ;
  assign n10381 = n10361 & ~n10378 ;
  assign n10382 = ~n9995 & n10381 ;
  assign n10383 = ~n10380 & ~n10382 ;
  assign n10384 = ~n10361 & n10378 ;
  assign n10385 = ~n9995 & n10384 ;
  assign n10386 = n10361 & n10378 ;
  assign n10387 = n9995 & n10386 ;
  assign n10388 = ~n10385 & ~n10387 ;
  assign n10389 = n10383 & n10388 ;
  assign n10390 = n9992 & ~n10389 ;
  assign n10391 = n9968 & n10390 ;
  assign n10392 = n9992 & n10389 ;
  assign n10393 = ~n9968 & n10392 ;
  assign n10394 = ~n10391 & ~n10393 ;
  assign n10395 = ~n9968 & n10389 ;
  assign n10396 = n9911 & ~n10389 ;
  assign n10397 = ~n9967 & n10396 ;
  assign n10398 = ~n9992 & ~n10397 ;
  assign n10399 = ~n10395 & n10398 ;
  assign n10400 = n10394 & ~n10399 ;
  assign n10401 = ~n9477 & n9930 ;
  assign n10402 = ~n9926 & n10401 ;
  assign n10403 = ~n9929 & ~n10402 ;
  assign n10404 = ~\b[42]  & ~\b[43]  ;
  assign n10405 = \b[42]  & \b[43]  ;
  assign n10406 = ~n10404 & ~n10405 ;
  assign n10407 = ~n10403 & n10406 ;
  assign n10408 = ~n9929 & ~n10406 ;
  assign n10409 = ~n10402 & n10408 ;
  assign n10410 = n134 & ~n10409 ;
  assign n10411 = ~n10407 & n10410 ;
  assign n10412 = \a[0]  & \b[43]  ;
  assign n10413 = n133 & n10412 ;
  assign n10414 = \b[42]  & n141 ;
  assign n10415 = ~\a[1]  & \b[41]  ;
  assign n10416 = ~\a[0]  & \a[2]  ;
  assign n10417 = n10415 & n10416 ;
  assign n10418 = ~n10414 & ~n10417 ;
  assign n10419 = ~n10413 & n10418 ;
  assign n10420 = ~n10411 & n10419 ;
  assign n10421 = ~\a[2]  & ~n10420 ;
  assign n10422 = \a[2]  & n10419 ;
  assign n10423 = ~n10411 & n10422 ;
  assign n10424 = ~n10421 & ~n10423 ;
  assign n10425 = ~n10400 & ~n10424 ;
  assign n10426 = n9966 & n10425 ;
  assign n10427 = n10400 & ~n10424 ;
  assign n10428 = ~n9966 & n10427 ;
  assign n10429 = ~n10426 & ~n10428 ;
  assign n10430 = ~n10400 & n10424 ;
  assign n10431 = ~n9966 & n10430 ;
  assign n10432 = n10400 & n10424 ;
  assign n10433 = n9966 & n10432 ;
  assign n10434 = ~n10431 & ~n10433 ;
  assign n10435 = n10429 & n10434 ;
  assign n10436 = ~n9963 & n10435 ;
  assign n10437 = ~n9953 & ~n10435 ;
  assign n10438 = ~n9960 & n10437 ;
  assign n10439 = ~n10436 & ~n10438 ;
  assign n10440 = ~n9953 & n10429 ;
  assign n10441 = n10434 & ~n10440 ;
  assign n10442 = n9959 & n10434 ;
  assign n10443 = n9514 & n10442 ;
  assign n10444 = ~n10441 & ~n10443 ;
  assign n10445 = n9966 & n10400 ;
  assign n10446 = ~n10399 & ~n10445 ;
  assign n10447 = n252 & ~n9482 ;
  assign n10448 = ~n9480 & n10447 ;
  assign n10449 = \b[41]  & n250 ;
  assign n10450 = \a[3]  & \b[40]  ;
  assign n10451 = n241 & n10450 ;
  assign n10452 = ~n10449 & ~n10451 ;
  assign n10453 = \b[39]  & n303 ;
  assign n10454 = n300 & n10453 ;
  assign n10455 = ~\a[3]  & \b[40]  ;
  assign n10456 = n244 & n10455 ;
  assign n10457 = ~n10454 & ~n10456 ;
  assign n10458 = n10452 & n10457 ;
  assign n10459 = ~n10448 & n10458 ;
  assign n10460 = ~\a[5]  & ~n10459 ;
  assign n10461 = \a[5]  & n10458 ;
  assign n10462 = ~n10448 & n10461 ;
  assign n10463 = ~n10460 & ~n10462 ;
  assign n10464 = n9911 & n10383 ;
  assign n10465 = n10388 & ~n10464 ;
  assign n10466 = n9912 & n10388 ;
  assign n10467 = n9519 & n10466 ;
  assign n10468 = ~n10465 & ~n10467 ;
  assign n10469 = n9995 & n10361 ;
  assign n10470 = n10355 & ~n10469 ;
  assign n10471 = ~n9872 & ~n10325 ;
  assign n10472 = ~n9879 & n10471 ;
  assign n10473 = n10320 & ~n10472 ;
  assign n10474 = ~n10309 & ~n10323 ;
  assign n10475 = n999 & n5810 ;
  assign n10476 = ~n5807 & n10475 ;
  assign n10477 = n999 & ~n5810 ;
  assign n10478 = ~n5457 & n10477 ;
  assign n10479 = ~n5806 & n10478 ;
  assign n10480 = \b[30]  & n1182 ;
  assign n10481 = n1179 & n10480 ;
  assign n10482 = \b[32]  & n997 ;
  assign n10483 = \a[11]  & \b[31]  ;
  assign n10484 = n1180 & n10483 ;
  assign n10485 = ~\a[12]  & \b[31]  ;
  assign n10486 = n7674 & n10485 ;
  assign n10487 = ~n10484 & ~n10486 ;
  assign n10488 = ~n10482 & n10487 ;
  assign n10489 = ~n10481 & n10488 ;
  assign n10490 = ~n10479 & n10489 ;
  assign n10491 = ~n10476 & n10490 ;
  assign n10492 = ~\a[14]  & ~n10491 ;
  assign n10493 = \a[14]  & n10489 ;
  assign n10494 = ~n10479 & n10493 ;
  assign n10495 = ~n10476 & n10494 ;
  assign n10496 = ~n10492 & ~n10495 ;
  assign n10497 = n9814 & n10274 ;
  assign n10498 = ~n9818 & n10497 ;
  assign n10499 = n10279 & ~n10498 ;
  assign n10500 = n1467 & ~n4502 ;
  assign n10501 = ~n4500 & n10500 ;
  assign n10502 = \b[29]  & n1465 ;
  assign n10503 = \a[15]  & \b[28]  ;
  assign n10504 = n1456 & n10503 ;
  assign n10505 = ~n10502 & ~n10504 ;
  assign n10506 = \b[27]  & n1652 ;
  assign n10507 = n1649 & n10506 ;
  assign n10508 = ~\a[15]  & \b[28]  ;
  assign n10509 = n1459 & n10508 ;
  assign n10510 = ~n10507 & ~n10509 ;
  assign n10511 = n10505 & n10510 ;
  assign n10512 = ~n10501 & n10511 ;
  assign n10513 = ~\a[17]  & ~n10512 ;
  assign n10514 = \a[17]  & n10511 ;
  assign n10515 = ~n10501 & n10514 ;
  assign n10516 = ~n10513 & ~n10515 ;
  assign n10517 = n10020 & n10252 ;
  assign n10518 = n10246 & ~n10517 ;
  assign n10519 = n1965 & n3604 ;
  assign n10520 = ~n3601 & n10519 ;
  assign n10521 = n1965 & ~n3604 ;
  assign n10522 = ~n3562 & n10521 ;
  assign n10523 = ~n3600 & n10522 ;
  assign n10524 = \b[24]  & n2218 ;
  assign n10525 = n2216 & n10524 ;
  assign n10526 = ~\a[18]  & \b[25]  ;
  assign n10527 = n1957 & n10526 ;
  assign n10528 = ~n10525 & ~n10527 ;
  assign n10529 = \b[26]  & n1963 ;
  assign n10530 = \a[18]  & \b[25]  ;
  assign n10531 = n2210 & n10530 ;
  assign n10532 = \a[20]  & ~n10531 ;
  assign n10533 = ~n10529 & n10532 ;
  assign n10534 = n10528 & n10533 ;
  assign n10535 = ~n10523 & n10534 ;
  assign n10536 = ~n10520 & n10535 ;
  assign n10537 = ~n10529 & ~n10531 ;
  assign n10538 = n10528 & n10537 ;
  assign n10539 = ~n10523 & n10538 ;
  assign n10540 = ~n10520 & n10539 ;
  assign n10541 = ~\a[20]  & ~n10540 ;
  assign n10542 = ~n10536 & ~n10541 ;
  assign n10543 = ~n9752 & n10218 ;
  assign n10544 = ~n9759 & n10543 ;
  assign n10545 = n10223 & ~n10544 ;
  assign n10546 = n10024 & n10194 ;
  assign n10547 = ~n10188 & ~n10546 ;
  assign n10548 = n9707 & n10158 ;
  assign n10549 = ~n10025 & n10548 ;
  assign n10550 = n10153 & ~n10549 ;
  assign n10551 = ~n1691 & n4249 ;
  assign n10552 = ~n1511 & n4249 ;
  assign n10553 = ~n1515 & n10552 ;
  assign n10554 = ~n10551 & ~n10553 ;
  assign n10555 = ~n1694 & ~n10554 ;
  assign n10556 = \b[15]  & n4647 ;
  assign n10557 = n4644 & n10556 ;
  assign n10558 = ~\a[27]  & \b[16]  ;
  assign n10559 = n4241 & n10558 ;
  assign n10560 = ~n10557 & ~n10559 ;
  assign n10561 = \b[17]  & n4247 ;
  assign n10562 = \a[27]  & \b[16]  ;
  assign n10563 = n4238 & n10562 ;
  assign n10564 = \a[29]  & ~n10563 ;
  assign n10565 = ~n10561 & n10564 ;
  assign n10566 = n10560 & n10565 ;
  assign n10567 = ~n10555 & n10566 ;
  assign n10568 = ~n10561 & ~n10563 ;
  assign n10569 = n10560 & n10568 ;
  assign n10570 = ~\a[29]  & ~n10569 ;
  assign n10571 = ~\a[29]  & ~n1694 ;
  assign n10572 = ~n10554 & n10571 ;
  assign n10573 = ~n10570 & ~n10572 ;
  assign n10574 = ~n10567 & n10573 ;
  assign n10575 = n10029 & n10148 ;
  assign n10576 = n10142 & ~n10575 ;
  assign n10577 = n1087 & n5211 ;
  assign n10578 = ~n1084 & n10577 ;
  assign n10579 = ~n1087 & n5211 ;
  assign n10580 = ~n946 & n10579 ;
  assign n10581 = ~n1083 & n10580 ;
  assign n10582 = \b[12]  & n5595 ;
  assign n10583 = n5592 & n10582 ;
  assign n10584 = ~\a[30]  & \b[13]  ;
  assign n10585 = n5203 & n10584 ;
  assign n10586 = ~n10583 & ~n10585 ;
  assign n10587 = \b[14]  & n5209 ;
  assign n10588 = \a[30]  & \b[13]  ;
  assign n10589 = n5200 & n10588 ;
  assign n10590 = \a[32]  & ~n10589 ;
  assign n10591 = ~n10587 & n10590 ;
  assign n10592 = n10586 & n10591 ;
  assign n10593 = ~n10581 & n10592 ;
  assign n10594 = ~n10578 & n10593 ;
  assign n10595 = ~n10587 & ~n10589 ;
  assign n10596 = n10586 & n10595 ;
  assign n10597 = ~n10581 & n10596 ;
  assign n10598 = ~n10578 & n10597 ;
  assign n10599 = ~\a[32]  & ~n10598 ;
  assign n10600 = ~n10594 & ~n10599 ;
  assign n10601 = ~n725 & n6309 ;
  assign n10602 = ~n684 & n6309 ;
  assign n10603 = ~n721 & n10602 ;
  assign n10604 = ~n10601 & ~n10603 ;
  assign n10605 = ~n728 & ~n10604 ;
  assign n10606 = \b[9]  & n6778 ;
  assign n10607 = n6775 & n10606 ;
  assign n10608 = \b[11]  & n6307 ;
  assign n10609 = \a[33]  & \b[10]  ;
  assign n10610 = n6298 & n10609 ;
  assign n10611 = ~\a[33]  & \b[10]  ;
  assign n10612 = n6301 & n10611 ;
  assign n10613 = ~n10610 & ~n10612 ;
  assign n10614 = ~n10608 & n10613 ;
  assign n10615 = ~n10607 & n10614 ;
  assign n10616 = ~\a[35]  & n10615 ;
  assign n10617 = ~n10605 & n10616 ;
  assign n10618 = \a[35]  & ~n10615 ;
  assign n10619 = \a[35]  & ~n728 ;
  assign n10620 = ~n10604 & n10619 ;
  assign n10621 = ~n10618 & ~n10620 ;
  assign n10622 = ~n10617 & n10621 ;
  assign n10623 = ~n9677 & ~n10113 ;
  assign n10624 = ~n9681 & n10623 ;
  assign n10625 = ~n10114 & ~n10624 ;
  assign n10626 = ~n505 & ~n7098 ;
  assign n10627 = ~n7531 & n10626 ;
  assign n10628 = n502 & n10627 ;
  assign n10629 = n505 & ~n7098 ;
  assign n10630 = ~n7531 & n10629 ;
  assign n10631 = ~n502 & n10630 ;
  assign n10632 = ~n10628 & ~n10631 ;
  assign n10633 = \b[6]  & n7973 ;
  assign n10634 = n7970 & n10633 ;
  assign n10635 = \b[8]  & n7532 ;
  assign n10636 = \a[35]  & \b[7]  ;
  assign n10637 = n7971 & n10636 ;
  assign n10638 = ~\a[36]  & \b[7]  ;
  assign n10639 = n7526 & n10638 ;
  assign n10640 = ~n10637 & ~n10639 ;
  assign n10641 = ~n10635 & n10640 ;
  assign n10642 = ~n10634 & n10641 ;
  assign n10643 = n10632 & n10642 ;
  assign n10644 = ~\a[38]  & ~n10643 ;
  assign n10645 = \a[38]  & n10642 ;
  assign n10646 = n10632 & n10645 ;
  assign n10647 = ~n10644 & ~n10646 ;
  assign n10648 = ~n10091 & ~n10093 ;
  assign n10649 = ~n273 & n8759 ;
  assign n10650 = ~n271 & n10649 ;
  assign n10651 = \b[3]  & n9301 ;
  assign n10652 = n9298 & n10651 ;
  assign n10653 = \b[5]  & n8757 ;
  assign n10654 = \a[38]  & \b[4]  ;
  assign n10655 = n9299 & n10654 ;
  assign n10656 = ~\a[39]  & \b[4]  ;
  assign n10657 = n8751 & n10656 ;
  assign n10658 = ~n10655 & ~n10657 ;
  assign n10659 = ~n10653 & n10658 ;
  assign n10660 = ~n10652 & n10659 ;
  assign n10661 = ~n10650 & n10660 ;
  assign n10662 = ~\a[41]  & ~n10661 ;
  assign n10663 = \a[41]  & n10660 ;
  assign n10664 = ~n10650 & n10663 ;
  assign n10665 = ~n10662 & ~n10664 ;
  assign n10666 = \a[44]  & ~n9647 ;
  assign n10667 = n10076 & n10666 ;
  assign n10668 = n10084 & n10667 ;
  assign n10669 = \a[44]  & ~n10668 ;
  assign n10670 = \b[2]  & n10080 ;
  assign n10671 = ~\a[42]  & \b[1]  ;
  assign n10672 = n10074 & n10671 ;
  assign n10673 = \a[42]  & \b[1]  ;
  assign n10674 = n10071 & n10673 ;
  assign n10675 = ~n10672 & ~n10674 ;
  assign n10676 = ~n10670 & n10675 ;
  assign n10677 = n157 & n10082 ;
  assign n10678 = n9646 & ~n10079 ;
  assign n10679 = \a[42]  & ~\a[43]  ;
  assign n10680 = ~\a[42]  & \a[43]  ;
  assign n10681 = ~n10679 & ~n10680 ;
  assign n10682 = \b[0]  & n10681 ;
  assign n10683 = n10678 & n10682 ;
  assign n10684 = ~n10677 & ~n10683 ;
  assign n10685 = n10676 & n10684 ;
  assign n10686 = ~n10669 & ~n10685 ;
  assign n10687 = n10669 & n10685 ;
  assign n10688 = ~n10686 & ~n10687 ;
  assign n10689 = ~n10665 & ~n10688 ;
  assign n10690 = n10665 & n10688 ;
  assign n10691 = ~n10689 & ~n10690 ;
  assign n10692 = ~n10648 & n10691 ;
  assign n10693 = n10648 & ~n10691 ;
  assign n10694 = ~n10692 & ~n10693 ;
  assign n10695 = ~n10647 & n10694 ;
  assign n10696 = n10647 & ~n10694 ;
  assign n10697 = ~n10695 & ~n10696 ;
  assign n10698 = n10625 & n10697 ;
  assign n10699 = ~n10625 & ~n10697 ;
  assign n10700 = ~n10698 & ~n10699 ;
  assign n10701 = ~n10622 & ~n10700 ;
  assign n10702 = n10622 & n10700 ;
  assign n10703 = ~n10701 & ~n10702 ;
  assign n10704 = n10600 & ~n10703 ;
  assign n10705 = n10576 & n10704 ;
  assign n10706 = n10600 & n10703 ;
  assign n10707 = ~n10576 & n10706 ;
  assign n10708 = ~n10705 & ~n10707 ;
  assign n10709 = ~n10600 & ~n10703 ;
  assign n10710 = ~n10576 & n10709 ;
  assign n10711 = ~n10600 & n10703 ;
  assign n10712 = n10576 & n10711 ;
  assign n10713 = ~n10710 & ~n10712 ;
  assign n10714 = n10708 & n10713 ;
  assign n10715 = n10574 & ~n10714 ;
  assign n10716 = ~n10550 & n10715 ;
  assign n10717 = n10574 & n10714 ;
  assign n10718 = n10550 & n10717 ;
  assign n10719 = ~n10716 & ~n10718 ;
  assign n10720 = ~n10574 & ~n10714 ;
  assign n10721 = n10550 & n10720 ;
  assign n10722 = ~n10574 & n10714 ;
  assign n10723 = ~n10550 & n10722 ;
  assign n10724 = ~n10721 & ~n10723 ;
  assign n10725 = n10719 & n10724 ;
  assign n10726 = ~n10547 & n10725 ;
  assign n10727 = ~n10188 & ~n10725 ;
  assign n10728 = ~n10546 & n10727 ;
  assign n10729 = n2293 & n3402 ;
  assign n10730 = ~n2290 & n10729 ;
  assign n10731 = n3402 & n5705 ;
  assign n10732 = ~n2289 & n10731 ;
  assign n10733 = \b[18]  & n3733 ;
  assign n10734 = n3730 & n10733 ;
  assign n10735 = ~\a[24]  & \b[19]  ;
  assign n10736 = n3394 & n10735 ;
  assign n10737 = ~n10734 & ~n10736 ;
  assign n10738 = \b[20]  & n3400 ;
  assign n10739 = \a[24]  & \b[19]  ;
  assign n10740 = n3391 & n10739 ;
  assign n10741 = \a[26]  & ~n10740 ;
  assign n10742 = ~n10738 & n10741 ;
  assign n10743 = n10737 & n10742 ;
  assign n10744 = ~n10732 & n10743 ;
  assign n10745 = ~n10730 & n10744 ;
  assign n10746 = ~n10738 & ~n10740 ;
  assign n10747 = n10737 & n10746 ;
  assign n10748 = ~n10732 & n10747 ;
  assign n10749 = ~n10730 & n10748 ;
  assign n10750 = ~\a[26]  & ~n10749 ;
  assign n10751 = ~n10745 & ~n10750 ;
  assign n10752 = ~n10728 & ~n10751 ;
  assign n10753 = ~n10726 & n10752 ;
  assign n10754 = ~n10725 & n10751 ;
  assign n10755 = n10547 & n10754 ;
  assign n10756 = n10725 & n10751 ;
  assign n10757 = ~n10547 & n10756 ;
  assign n10758 = ~n10755 & ~n10757 ;
  assign n10759 = ~n10753 & n10758 ;
  assign n10760 = ~n10545 & ~n10759 ;
  assign n10761 = n10545 & n10759 ;
  assign n10762 = ~n10760 & ~n10761 ;
  assign n10763 = n2622 & ~n3022 ;
  assign n10764 = ~n3020 & n10763 ;
  assign n10765 = \b[21]  & n2912 ;
  assign n10766 = n2909 & n10765 ;
  assign n10767 = \b[23]  & n2620 ;
  assign n10768 = \a[20]  & \b[22]  ;
  assign n10769 = n2910 & n10768 ;
  assign n10770 = ~\a[21]  & \b[22]  ;
  assign n10771 = n2614 & n10770 ;
  assign n10772 = ~n10769 & ~n10771 ;
  assign n10773 = ~n10767 & n10772 ;
  assign n10774 = ~n10766 & n10773 ;
  assign n10775 = ~\a[23]  & n10774 ;
  assign n10776 = ~n10764 & n10775 ;
  assign n10777 = ~n10764 & n10774 ;
  assign n10778 = \a[23]  & ~n10777 ;
  assign n10779 = ~n10776 & ~n10778 ;
  assign n10780 = n10762 & n10779 ;
  assign n10781 = ~n10762 & ~n10779 ;
  assign n10782 = ~n10780 & ~n10781 ;
  assign n10783 = n10542 & ~n10782 ;
  assign n10784 = n10518 & n10783 ;
  assign n10785 = n10542 & n10782 ;
  assign n10786 = ~n10518 & n10785 ;
  assign n10787 = ~n10784 & ~n10786 ;
  assign n10788 = ~n10542 & ~n10782 ;
  assign n10789 = ~n10518 & n10788 ;
  assign n10790 = ~n10542 & n10782 ;
  assign n10791 = n10518 & n10790 ;
  assign n10792 = ~n10789 & ~n10791 ;
  assign n10793 = n10787 & n10792 ;
  assign n10794 = n10516 & ~n10793 ;
  assign n10795 = ~n10499 & n10794 ;
  assign n10796 = n10516 & n10793 ;
  assign n10797 = n10499 & n10796 ;
  assign n10798 = ~n10795 & ~n10797 ;
  assign n10799 = ~n10516 & ~n10793 ;
  assign n10800 = n10499 & n10799 ;
  assign n10801 = ~n10516 & n10793 ;
  assign n10802 = ~n10499 & n10801 ;
  assign n10803 = ~n10800 & ~n10802 ;
  assign n10804 = n10798 & n10803 ;
  assign n10805 = n10496 & ~n10804 ;
  assign n10806 = n10474 & n10805 ;
  assign n10807 = n10496 & n10804 ;
  assign n10808 = ~n10474 & n10807 ;
  assign n10809 = ~n10806 & ~n10808 ;
  assign n10810 = ~n10474 & n10804 ;
  assign n10811 = ~n10309 & ~n10804 ;
  assign n10812 = ~n10323 & n10811 ;
  assign n10813 = ~n10496 & ~n10812 ;
  assign n10814 = ~n10810 & n10813 ;
  assign n10815 = n10809 & ~n10814 ;
  assign n10816 = n646 & ~n6610 ;
  assign n10817 = ~n6608 & n10816 ;
  assign n10818 = \b[35]  & n644 ;
  assign n10819 = \a[9]  & \b[34]  ;
  assign n10820 = n635 & n10819 ;
  assign n10821 = ~n10818 & ~n10820 ;
  assign n10822 = \b[33]  & n796 ;
  assign n10823 = n793 & n10822 ;
  assign n10824 = ~\a[9]  & \b[34]  ;
  assign n10825 = n638 & n10824 ;
  assign n10826 = ~n10823 & ~n10825 ;
  assign n10827 = n10821 & n10826 ;
  assign n10828 = ~n10817 & n10827 ;
  assign n10829 = ~\a[11]  & ~n10828 ;
  assign n10830 = \a[11]  & n10827 ;
  assign n10831 = ~n10817 & n10830 ;
  assign n10832 = ~n10829 & ~n10831 ;
  assign n10833 = ~n10815 & ~n10832 ;
  assign n10834 = n10473 & n10833 ;
  assign n10835 = n10815 & ~n10832 ;
  assign n10836 = ~n10473 & n10835 ;
  assign n10837 = ~n10834 & ~n10836 ;
  assign n10838 = ~n10815 & n10832 ;
  assign n10839 = ~n10473 & n10838 ;
  assign n10840 = n10815 & n10832 ;
  assign n10841 = n10473 & n10840 ;
  assign n10842 = ~n10839 & ~n10841 ;
  assign n10843 = n10837 & n10842 ;
  assign n10844 = ~n10470 & n10843 ;
  assign n10845 = n10355 & ~n10843 ;
  assign n10846 = ~n10469 & n10845 ;
  assign n10847 = n430 & n8175 ;
  assign n10848 = ~n8172 & n10847 ;
  assign n10849 = n430 & ~n8175 ;
  assign n10850 = ~n7756 & n10849 ;
  assign n10851 = ~n8171 & n10850 ;
  assign n10852 = \b[36]  & n486 ;
  assign n10853 = n483 & n10852 ;
  assign n10854 = \b[38]  & n428 ;
  assign n10855 = \a[6]  & \b[37]  ;
  assign n10856 = n419 & n10855 ;
  assign n10857 = ~\a[6]  & \b[37]  ;
  assign n10858 = n422 & n10857 ;
  assign n10859 = ~n10856 & ~n10858 ;
  assign n10860 = ~n10854 & n10859 ;
  assign n10861 = ~n10853 & n10860 ;
  assign n10862 = ~n10851 & n10861 ;
  assign n10863 = ~n10848 & n10862 ;
  assign n10864 = ~\a[8]  & ~n10863 ;
  assign n10865 = \a[8]  & n10861 ;
  assign n10866 = ~n10851 & n10865 ;
  assign n10867 = ~n10848 & n10866 ;
  assign n10868 = ~n10864 & ~n10867 ;
  assign n10869 = ~n10846 & ~n10868 ;
  assign n10870 = ~n10844 & n10869 ;
  assign n10871 = ~n10843 & n10868 ;
  assign n10872 = n10470 & n10871 ;
  assign n10873 = n10843 & n10868 ;
  assign n10874 = ~n10470 & n10873 ;
  assign n10875 = ~n10872 & ~n10874 ;
  assign n10876 = ~n10870 & n10875 ;
  assign n10877 = ~n10468 & n10876 ;
  assign n10878 = n10468 & ~n10876 ;
  assign n10879 = ~n10877 & ~n10878 ;
  assign n10880 = ~n10463 & n10879 ;
  assign n10881 = n10463 & ~n10879 ;
  assign n10882 = ~n10880 & ~n10881 ;
  assign n10883 = ~n10446 & n10882 ;
  assign n10884 = ~n9929 & ~n10405 ;
  assign n10885 = ~n10402 & n10884 ;
  assign n10886 = ~n10404 & ~n10885 ;
  assign n10887 = ~\b[43]  & ~\b[44]  ;
  assign n10888 = \b[43]  & \b[44]  ;
  assign n10889 = ~n10887 & ~n10888 ;
  assign n10890 = ~n10886 & ~n10889 ;
  assign n10891 = ~n10404 & n10889 ;
  assign n10892 = ~n10885 & n10891 ;
  assign n10893 = n134 & ~n10892 ;
  assign n10894 = ~n10890 & n10893 ;
  assign n10895 = \a[0]  & \b[44]  ;
  assign n10896 = n133 & n10895 ;
  assign n10897 = \b[43]  & n141 ;
  assign n10898 = ~\a[1]  & \b[42]  ;
  assign n10899 = n10416 & n10898 ;
  assign n10900 = ~n10897 & ~n10899 ;
  assign n10901 = ~n10896 & n10900 ;
  assign n10902 = \a[2]  & n10901 ;
  assign n10903 = ~n10894 & n10902 ;
  assign n10904 = ~n10894 & n10901 ;
  assign n10905 = ~\a[2]  & ~n10904 ;
  assign n10906 = ~n10903 & ~n10905 ;
  assign n10907 = ~n10399 & ~n10882 ;
  assign n10908 = ~n10445 & n10907 ;
  assign n10909 = ~n10906 & ~n10908 ;
  assign n10910 = ~n10883 & n10909 ;
  assign n10911 = ~n10882 & n10906 ;
  assign n10912 = n10446 & n10911 ;
  assign n10913 = n10882 & n10906 ;
  assign n10914 = ~n10446 & n10913 ;
  assign n10915 = ~n10912 & ~n10914 ;
  assign n10916 = ~n10910 & n10915 ;
  assign n10917 = ~n10444 & n10916 ;
  assign n10918 = n10444 & ~n10916 ;
  assign n10919 = ~n10917 & ~n10918 ;
  assign n10920 = ~n10910 & ~n10917 ;
  assign n10921 = ~n10399 & ~n10880 ;
  assign n10922 = ~n10445 & n10921 ;
  assign n10923 = ~n10881 & ~n10922 ;
  assign n10924 = ~n10870 & ~n10877 ;
  assign n10925 = n10355 & n10837 ;
  assign n10926 = ~n10469 & n10925 ;
  assign n10927 = n10842 & ~n10926 ;
  assign n10928 = n10473 & n10815 ;
  assign n10929 = ~n10814 & ~n10928 ;
  assign n10930 = ~n10309 & n10803 ;
  assign n10931 = ~n10323 & n10930 ;
  assign n10932 = n10798 & ~n10931 ;
  assign n10933 = n10499 & n10793 ;
  assign n10934 = n10792 & ~n10933 ;
  assign n10935 = n10246 & ~n10780 ;
  assign n10936 = ~n10517 & n10935 ;
  assign n10937 = ~n10781 & ~n10936 ;
  assign n10938 = ~n10753 & ~n10761 ;
  assign n10939 = ~n10188 & n10724 ;
  assign n10940 = ~n10546 & n10939 ;
  assign n10941 = n10719 & ~n10940 ;
  assign n10942 = n10550 & n10714 ;
  assign n10943 = n10713 & ~n10942 ;
  assign n10944 = n10142 & ~n10702 ;
  assign n10945 = ~n10575 & n10944 ;
  assign n10946 = ~n10701 & ~n10945 ;
  assign n10947 = ~n1233 & n5211 ;
  assign n10948 = ~n1231 & n10947 ;
  assign n10949 = \b[13]  & n5595 ;
  assign n10950 = n5592 & n10949 ;
  assign n10951 = ~\a[30]  & \b[14]  ;
  assign n10952 = n5203 & n10951 ;
  assign n10953 = ~n10950 & ~n10952 ;
  assign n10954 = \b[15]  & n5209 ;
  assign n10955 = \a[30]  & \b[14]  ;
  assign n10956 = n5200 & n10955 ;
  assign n10957 = \a[32]  & ~n10956 ;
  assign n10958 = ~n10954 & n10957 ;
  assign n10959 = n10953 & n10958 ;
  assign n10960 = ~n10948 & n10959 ;
  assign n10961 = ~n10954 & ~n10956 ;
  assign n10962 = n10953 & n10961 ;
  assign n10963 = ~n10948 & n10962 ;
  assign n10964 = ~\a[32]  & ~n10963 ;
  assign n10965 = ~n10960 & ~n10964 ;
  assign n10966 = ~n10695 & ~n10698 ;
  assign n10967 = ~n10091 & ~n10689 ;
  assign n10968 = ~n10093 & n10967 ;
  assign n10969 = ~n10690 & ~n10968 ;
  assign n10970 = n177 & n10082 ;
  assign n10971 = \b[3]  & n10080 ;
  assign n10972 = \a[41]  & \b[2]  ;
  assign n10973 = n10679 & n10972 ;
  assign n10974 = ~\a[42]  & \b[2]  ;
  assign n10975 = n10074 & n10974 ;
  assign n10976 = ~n10973 & ~n10975 ;
  assign n10977 = ~n10971 & n10976 ;
  assign n10978 = ~n10970 & n10977 ;
  assign n10979 = \b[1]  & n10681 ;
  assign n10980 = n10678 & n10979 ;
  assign n10981 = ~\a[44]  & ~n10980 ;
  assign n10982 = n10978 & n10981 ;
  assign n10983 = n10978 & ~n10980 ;
  assign n10984 = \a[44]  & ~n10983 ;
  assign n10985 = ~n10982 & ~n10984 ;
  assign n10986 = \a[44]  & ~\a[45]  ;
  assign n10987 = ~\a[44]  & \a[45]  ;
  assign n10988 = ~n10986 & ~n10987 ;
  assign n10989 = \b[0]  & ~n10988 ;
  assign n10990 = n10668 & n10685 ;
  assign n10991 = n10989 & n10990 ;
  assign n10992 = ~n10989 & ~n10990 ;
  assign n10993 = ~n10991 & ~n10992 ;
  assign n10994 = n10985 & n10993 ;
  assign n10995 = ~n10985 & ~n10993 ;
  assign n10996 = ~n10994 & ~n10995 ;
  assign n10997 = ~n323 & ~n8272 ;
  assign n10998 = ~n8756 & n10997 ;
  assign n10999 = n320 & n10998 ;
  assign n11000 = n323 & ~n8272 ;
  assign n11001 = ~n8756 & n11000 ;
  assign n11002 = ~n320 & n11001 ;
  assign n11003 = ~n10999 & ~n11002 ;
  assign n11004 = \b[4]  & n9301 ;
  assign n11005 = n9298 & n11004 ;
  assign n11006 = ~\a[39]  & \b[5]  ;
  assign n11007 = n8751 & n11006 ;
  assign n11008 = ~n11005 & ~n11007 ;
  assign n11009 = \b[6]  & n8757 ;
  assign n11010 = \a[39]  & \b[5]  ;
  assign n11011 = n8748 & n11010 ;
  assign n11012 = \a[41]  & ~n11011 ;
  assign n11013 = ~n11009 & n11012 ;
  assign n11014 = n11008 & n11013 ;
  assign n11015 = n11003 & n11014 ;
  assign n11016 = ~n11009 & ~n11011 ;
  assign n11017 = n11008 & n11016 ;
  assign n11018 = n11003 & n11017 ;
  assign n11019 = ~\a[41]  & ~n11018 ;
  assign n11020 = ~n11015 & ~n11019 ;
  assign n11021 = n10996 & ~n11020 ;
  assign n11022 = ~n10996 & n11020 ;
  assign n11023 = ~n11021 & ~n11022 ;
  assign n11024 = ~n586 & n7534 ;
  assign n11025 = ~n504 & n7534 ;
  assign n11026 = ~n508 & n11025 ;
  assign n11027 = ~n11024 & ~n11026 ;
  assign n11028 = ~n589 & ~n11027 ;
  assign n11029 = \b[7]  & n7973 ;
  assign n11030 = n7970 & n11029 ;
  assign n11031 = \b[9]  & n7532 ;
  assign n11032 = \a[36]  & \b[8]  ;
  assign n11033 = n7523 & n11032 ;
  assign n11034 = ~\a[36]  & \b[8]  ;
  assign n11035 = n7526 & n11034 ;
  assign n11036 = ~n11033 & ~n11035 ;
  assign n11037 = ~n11031 & n11036 ;
  assign n11038 = ~n11030 & n11037 ;
  assign n11039 = ~\a[38]  & n11038 ;
  assign n11040 = ~n11028 & n11039 ;
  assign n11041 = \a[38]  & ~n11038 ;
  assign n11042 = \a[38]  & ~n589 ;
  assign n11043 = ~n11027 & n11042 ;
  assign n11044 = ~n11041 & ~n11043 ;
  assign n11045 = ~n11040 & n11044 ;
  assign n11046 = ~n11023 & ~n11045 ;
  assign n11047 = ~n10969 & n11046 ;
  assign n11048 = n11023 & ~n11045 ;
  assign n11049 = n10969 & n11048 ;
  assign n11050 = ~n11047 & ~n11049 ;
  assign n11051 = ~n11023 & n11045 ;
  assign n11052 = n10969 & n11051 ;
  assign n11053 = n11023 & n11045 ;
  assign n11054 = ~n10969 & n11053 ;
  assign n11055 = ~n11052 & ~n11054 ;
  assign n11056 = n11050 & n11055 ;
  assign n11057 = ~n10966 & n11056 ;
  assign n11058 = ~n909 & ~n5952 ;
  assign n11059 = ~n6306 & n11058 ;
  assign n11060 = n906 & n11059 ;
  assign n11061 = n909 & ~n5952 ;
  assign n11062 = ~n6306 & n11061 ;
  assign n11063 = ~n906 & n11062 ;
  assign n11064 = ~n11060 & ~n11063 ;
  assign n11065 = \b[10]  & n6778 ;
  assign n11066 = n6775 & n11065 ;
  assign n11067 = \b[12]  & n6307 ;
  assign n11068 = \a[33]  & \b[11]  ;
  assign n11069 = n6298 & n11068 ;
  assign n11070 = ~\a[33]  & \b[11]  ;
  assign n11071 = n6301 & n11070 ;
  assign n11072 = ~n11069 & ~n11071 ;
  assign n11073 = ~n11067 & n11072 ;
  assign n11074 = ~n11066 & n11073 ;
  assign n11075 = n11064 & n11074 ;
  assign n11076 = ~\a[35]  & ~n11075 ;
  assign n11077 = \a[35]  & n11074 ;
  assign n11078 = n11064 & n11077 ;
  assign n11079 = ~n11076 & ~n11078 ;
  assign n11080 = ~n10695 & ~n11056 ;
  assign n11081 = ~n10698 & n11080 ;
  assign n11082 = ~n11079 & ~n11081 ;
  assign n11083 = ~n11057 & n11082 ;
  assign n11084 = ~n11056 & n11079 ;
  assign n11085 = n10966 & n11084 ;
  assign n11086 = n11056 & n11079 ;
  assign n11087 = ~n10966 & n11086 ;
  assign n11088 = ~n11085 & ~n11087 ;
  assign n11089 = ~n11083 & n11088 ;
  assign n11090 = ~n10965 & ~n11089 ;
  assign n11091 = n10946 & n11090 ;
  assign n11092 = ~n10965 & n11089 ;
  assign n11093 = ~n10946 & n11092 ;
  assign n11094 = ~n11091 & ~n11093 ;
  assign n11095 = n10965 & ~n11089 ;
  assign n11096 = ~n10946 & n11095 ;
  assign n11097 = n10965 & n11089 ;
  assign n11098 = n10946 & n11097 ;
  assign n11099 = ~n11096 & ~n11098 ;
  assign n11100 = n11094 & n11099 ;
  assign n11101 = ~n10943 & n11100 ;
  assign n11102 = n1875 & n4249 ;
  assign n11103 = ~n1872 & n11102 ;
  assign n11104 = n4249 & n5000 ;
  assign n11105 = ~n1871 & n11104 ;
  assign n11106 = \b[16]  & n4647 ;
  assign n11107 = n4644 & n11106 ;
  assign n11108 = ~\a[27]  & \b[17]  ;
  assign n11109 = n4241 & n11108 ;
  assign n11110 = ~n11107 & ~n11109 ;
  assign n11111 = \b[18]  & n4247 ;
  assign n11112 = \a[27]  & \b[17]  ;
  assign n11113 = n4238 & n11112 ;
  assign n11114 = \a[29]  & ~n11113 ;
  assign n11115 = ~n11111 & n11114 ;
  assign n11116 = n11110 & n11115 ;
  assign n11117 = ~n11105 & n11116 ;
  assign n11118 = ~n11103 & n11117 ;
  assign n11119 = ~n11111 & ~n11113 ;
  assign n11120 = n11110 & n11119 ;
  assign n11121 = ~n11105 & n11120 ;
  assign n11122 = ~n11103 & n11121 ;
  assign n11123 = ~\a[29]  & ~n11122 ;
  assign n11124 = ~n11118 & ~n11123 ;
  assign n11125 = n10713 & ~n11100 ;
  assign n11126 = ~n10942 & n11125 ;
  assign n11127 = ~n11124 & ~n11126 ;
  assign n11128 = ~n11101 & n11127 ;
  assign n11129 = ~n11100 & n11124 ;
  assign n11130 = n10943 & n11129 ;
  assign n11131 = n11100 & n11124 ;
  assign n11132 = ~n10943 & n11131 ;
  assign n11133 = ~n11130 & ~n11132 ;
  assign n11134 = ~n11128 & n11133 ;
  assign n11135 = ~n2520 & n3402 ;
  assign n11136 = ~n2292 & n3402 ;
  assign n11137 = ~n2516 & n11136 ;
  assign n11138 = ~n11135 & ~n11137 ;
  assign n11139 = ~n2523 & ~n11138 ;
  assign n11140 = \b[19]  & n3733 ;
  assign n11141 = n3730 & n11140 ;
  assign n11142 = ~\a[24]  & \b[20]  ;
  assign n11143 = n3394 & n11142 ;
  assign n11144 = ~n11141 & ~n11143 ;
  assign n11145 = \b[21]  & n3400 ;
  assign n11146 = \a[24]  & \b[20]  ;
  assign n11147 = n3391 & n11146 ;
  assign n11148 = \a[26]  & ~n11147 ;
  assign n11149 = ~n11145 & n11148 ;
  assign n11150 = n11144 & n11149 ;
  assign n11151 = ~n11139 & n11150 ;
  assign n11152 = ~n11145 & ~n11147 ;
  assign n11153 = n11144 & n11152 ;
  assign n11154 = ~\a[26]  & ~n11153 ;
  assign n11155 = ~\a[26]  & ~n2523 ;
  assign n11156 = ~n11138 & n11155 ;
  assign n11157 = ~n11154 & ~n11156 ;
  assign n11158 = ~n11151 & n11157 ;
  assign n11159 = ~n11134 & ~n11158 ;
  assign n11160 = n10941 & n11159 ;
  assign n11161 = n11134 & ~n11158 ;
  assign n11162 = ~n10941 & n11161 ;
  assign n11163 = ~n11160 & ~n11162 ;
  assign n11164 = ~n11134 & n11158 ;
  assign n11165 = ~n10941 & n11164 ;
  assign n11166 = n11134 & n11158 ;
  assign n11167 = n10941 & n11166 ;
  assign n11168 = ~n11165 & ~n11167 ;
  assign n11169 = n11163 & n11168 ;
  assign n11170 = ~n3280 & ~n3283 ;
  assign n11171 = n2622 & ~n3560 ;
  assign n11172 = ~n11170 & n11171 ;
  assign n11173 = \b[22]  & n2912 ;
  assign n11174 = n2909 & n11173 ;
  assign n11175 = \b[24]  & n2620 ;
  assign n11176 = \a[21]  & \b[23]  ;
  assign n11177 = n2611 & n11176 ;
  assign n11178 = ~\a[21]  & \b[23]  ;
  assign n11179 = n2614 & n11178 ;
  assign n11180 = ~n11177 & ~n11179 ;
  assign n11181 = ~n11175 & n11180 ;
  assign n11182 = ~n11174 & n11181 ;
  assign n11183 = ~n11172 & n11182 ;
  assign n11184 = ~\a[23]  & ~n11183 ;
  assign n11185 = \a[23]  & n11182 ;
  assign n11186 = ~n11172 & n11185 ;
  assign n11187 = ~n11184 & ~n11186 ;
  assign n11188 = ~n11169 & n11187 ;
  assign n11189 = n10938 & n11188 ;
  assign n11190 = n11169 & n11187 ;
  assign n11191 = ~n10938 & n11190 ;
  assign n11192 = ~n11189 & ~n11191 ;
  assign n11193 = ~n11169 & ~n11187 ;
  assign n11194 = ~n10938 & n11193 ;
  assign n11195 = n11169 & ~n11187 ;
  assign n11196 = n10938 & n11195 ;
  assign n11197 = ~n11194 & ~n11196 ;
  assign n11198 = n11192 & n11197 ;
  assign n11199 = ~n1805 & ~n1962 ;
  assign n11200 = ~n4148 & n11199 ;
  assign n11201 = ~n4146 & n11200 ;
  assign n11202 = \b[25]  & n2218 ;
  assign n11203 = n2216 & n11202 ;
  assign n11204 = ~\a[18]  & \b[26]  ;
  assign n11205 = n1957 & n11204 ;
  assign n11206 = ~n11203 & ~n11205 ;
  assign n11207 = \b[27]  & n1963 ;
  assign n11208 = \a[18]  & \b[26]  ;
  assign n11209 = n2210 & n11208 ;
  assign n11210 = \a[20]  & ~n11209 ;
  assign n11211 = ~n11207 & n11210 ;
  assign n11212 = n11206 & n11211 ;
  assign n11213 = ~n11201 & n11212 ;
  assign n11214 = ~n11207 & ~n11209 ;
  assign n11215 = n11206 & n11214 ;
  assign n11216 = ~n11201 & n11215 ;
  assign n11217 = ~\a[20]  & ~n11216 ;
  assign n11218 = ~n11213 & ~n11217 ;
  assign n11219 = ~n11198 & ~n11218 ;
  assign n11220 = n10937 & n11219 ;
  assign n11221 = n11198 & ~n11218 ;
  assign n11222 = ~n10937 & n11221 ;
  assign n11223 = ~n11220 & ~n11222 ;
  assign n11224 = ~n11198 & n11218 ;
  assign n11225 = ~n10937 & n11224 ;
  assign n11226 = n11198 & n11218 ;
  assign n11227 = n10937 & n11226 ;
  assign n11228 = ~n11225 & ~n11227 ;
  assign n11229 = n11223 & n11228 ;
  assign n11230 = ~n10934 & n11229 ;
  assign n11231 = n1467 & n5105 ;
  assign n11232 = ~n5102 & n11231 ;
  assign n11233 = n1467 & ~n5105 ;
  assign n11234 = ~n4497 & n11233 ;
  assign n11235 = ~n5101 & n11234 ;
  assign n11236 = \b[28]  & n1652 ;
  assign n11237 = n1649 & n11236 ;
  assign n11238 = ~\a[15]  & \b[29]  ;
  assign n11239 = n1459 & n11238 ;
  assign n11240 = ~n11237 & ~n11239 ;
  assign n11241 = \b[30]  & n1465 ;
  assign n11242 = \a[15]  & \b[29]  ;
  assign n11243 = n1456 & n11242 ;
  assign n11244 = \a[17]  & ~n11243 ;
  assign n11245 = ~n11241 & n11244 ;
  assign n11246 = n11240 & n11245 ;
  assign n11247 = ~n11235 & n11246 ;
  assign n11248 = ~n11232 & n11247 ;
  assign n11249 = ~n11241 & ~n11243 ;
  assign n11250 = n11240 & n11249 ;
  assign n11251 = ~n11235 & n11250 ;
  assign n11252 = ~n11232 & n11251 ;
  assign n11253 = ~\a[17]  & ~n11252 ;
  assign n11254 = ~n11248 & ~n11253 ;
  assign n11255 = n10792 & ~n11229 ;
  assign n11256 = ~n10933 & n11255 ;
  assign n11257 = ~n11254 & ~n11256 ;
  assign n11258 = ~n11230 & n11257 ;
  assign n11259 = ~n11229 & n11254 ;
  assign n11260 = n10934 & n11259 ;
  assign n11261 = n11229 & n11254 ;
  assign n11262 = ~n10934 & n11261 ;
  assign n11263 = ~n11260 & ~n11262 ;
  assign n11264 = ~n11258 & n11263 ;
  assign n11265 = n999 & ~n5855 ;
  assign n11266 = ~n5853 & n11265 ;
  assign n11267 = \b[31]  & n1182 ;
  assign n11268 = n1179 & n11267 ;
  assign n11269 = \b[33]  & n997 ;
  assign n11270 = \a[11]  & \b[32]  ;
  assign n11271 = n1180 & n11270 ;
  assign n11272 = ~\a[12]  & \b[32]  ;
  assign n11273 = n7674 & n11272 ;
  assign n11274 = ~n11271 & ~n11273 ;
  assign n11275 = ~n11269 & n11274 ;
  assign n11276 = ~n11268 & n11275 ;
  assign n11277 = ~n11266 & n11276 ;
  assign n11278 = ~\a[14]  & ~n11277 ;
  assign n11279 = \a[14]  & n11276 ;
  assign n11280 = ~n11266 & n11279 ;
  assign n11281 = ~n11278 & ~n11280 ;
  assign n11282 = ~n11264 & ~n11281 ;
  assign n11283 = n10932 & n11282 ;
  assign n11284 = n11264 & ~n11281 ;
  assign n11285 = ~n10932 & n11284 ;
  assign n11286 = ~n11283 & ~n11285 ;
  assign n11287 = ~n11264 & n11281 ;
  assign n11288 = ~n10932 & n11287 ;
  assign n11289 = n11264 & n11281 ;
  assign n11290 = n10932 & n11289 ;
  assign n11291 = ~n11288 & ~n11290 ;
  assign n11292 = n11286 & n11291 ;
  assign n11293 = ~n10929 & n11292 ;
  assign n11294 = n646 & n7337 ;
  assign n11295 = ~n7334 & n11294 ;
  assign n11296 = n646 & ~n7337 ;
  assign n11297 = ~n6605 & n11296 ;
  assign n11298 = ~n7333 & n11297 ;
  assign n11299 = \b[34]  & n796 ;
  assign n11300 = n793 & n11299 ;
  assign n11301 = ~\a[9]  & \b[35]  ;
  assign n11302 = n638 & n11301 ;
  assign n11303 = ~n11300 & ~n11302 ;
  assign n11304 = \b[36]  & n644 ;
  assign n11305 = \a[9]  & \b[35]  ;
  assign n11306 = n635 & n11305 ;
  assign n11307 = \a[11]  & ~n11306 ;
  assign n11308 = ~n11304 & n11307 ;
  assign n11309 = n11303 & n11308 ;
  assign n11310 = ~n11298 & n11309 ;
  assign n11311 = ~n11295 & n11310 ;
  assign n11312 = ~n11304 & ~n11306 ;
  assign n11313 = n11303 & n11312 ;
  assign n11314 = ~n11298 & n11313 ;
  assign n11315 = ~n11295 & n11314 ;
  assign n11316 = ~\a[11]  & ~n11315 ;
  assign n11317 = ~n11311 & ~n11316 ;
  assign n11318 = ~n10814 & ~n11292 ;
  assign n11319 = ~n10928 & n11318 ;
  assign n11320 = ~n11317 & ~n11319 ;
  assign n11321 = ~n11293 & n11320 ;
  assign n11322 = ~n11292 & n11317 ;
  assign n11323 = n10929 & n11322 ;
  assign n11324 = n11292 & n11317 ;
  assign n11325 = ~n10929 & n11324 ;
  assign n11326 = ~n11323 & ~n11325 ;
  assign n11327 = ~n11321 & n11326 ;
  assign n11328 = n430 & ~n8602 ;
  assign n11329 = ~n8600 & n11328 ;
  assign n11330 = \b[37]  & n486 ;
  assign n11331 = n483 & n11330 ;
  assign n11332 = \b[39]  & n428 ;
  assign n11333 = \a[6]  & \b[38]  ;
  assign n11334 = n419 & n11333 ;
  assign n11335 = ~\a[6]  & \b[38]  ;
  assign n11336 = n422 & n11335 ;
  assign n11337 = ~n11334 & ~n11336 ;
  assign n11338 = ~n11332 & n11337 ;
  assign n11339 = ~n11331 & n11338 ;
  assign n11340 = ~n11329 & n11339 ;
  assign n11341 = ~\a[8]  & ~n11340 ;
  assign n11342 = \a[8]  & n11339 ;
  assign n11343 = ~n11329 & n11342 ;
  assign n11344 = ~n11341 & ~n11343 ;
  assign n11345 = ~n11327 & ~n11344 ;
  assign n11346 = n10927 & n11345 ;
  assign n11347 = n11327 & ~n11344 ;
  assign n11348 = ~n10927 & n11347 ;
  assign n11349 = ~n11346 & ~n11348 ;
  assign n11350 = ~n11327 & n11344 ;
  assign n11351 = ~n10927 & n11350 ;
  assign n11352 = n11327 & n11344 ;
  assign n11353 = n10927 & n11352 ;
  assign n11354 = ~n11351 & ~n11353 ;
  assign n11355 = n11349 & n11354 ;
  assign n11356 = n252 & n9930 ;
  assign n11357 = ~n9927 & n11356 ;
  assign n11358 = ~n9477 & ~n9930 ;
  assign n11359 = n252 & n11358 ;
  assign n11360 = ~n9926 & n11359 ;
  assign n11361 = \b[40]  & n303 ;
  assign n11362 = n300 & n11361 ;
  assign n11363 = ~\a[3]  & \b[41]  ;
  assign n11364 = n244 & n11363 ;
  assign n11365 = ~n11362 & ~n11364 ;
  assign n11366 = \b[42]  & n250 ;
  assign n11367 = \a[3]  & \b[41]  ;
  assign n11368 = n241 & n11367 ;
  assign n11369 = \a[5]  & ~n11368 ;
  assign n11370 = ~n11366 & n11369 ;
  assign n11371 = n11365 & n11370 ;
  assign n11372 = ~n11360 & n11371 ;
  assign n11373 = ~n11357 & n11372 ;
  assign n11374 = ~n11366 & ~n11368 ;
  assign n11375 = n11365 & n11374 ;
  assign n11376 = ~n11360 & n11375 ;
  assign n11377 = ~n11357 & n11376 ;
  assign n11378 = ~\a[5]  & ~n11377 ;
  assign n11379 = ~n11373 & ~n11378 ;
  assign n11380 = ~n11355 & ~n11379 ;
  assign n11381 = ~n10924 & n11380 ;
  assign n11382 = n11355 & ~n11379 ;
  assign n11383 = n10924 & n11382 ;
  assign n11384 = ~n11381 & ~n11383 ;
  assign n11385 = ~n11355 & n11379 ;
  assign n11386 = n10924 & n11385 ;
  assign n11387 = n11355 & n11379 ;
  assign n11388 = ~n10924 & n11387 ;
  assign n11389 = ~n11386 & ~n11388 ;
  assign n11390 = n11384 & n11389 ;
  assign n11391 = ~n10888 & ~n10892 ;
  assign n11392 = ~\b[44]  & ~\b[45]  ;
  assign n11393 = \b[44]  & \b[45]  ;
  assign n11394 = ~n11392 & ~n11393 ;
  assign n11395 = ~n11391 & n11394 ;
  assign n11396 = ~n10888 & ~n11394 ;
  assign n11397 = ~n10892 & n11396 ;
  assign n11398 = n134 & ~n11397 ;
  assign n11399 = ~n11395 & n11398 ;
  assign n11400 = \a[0]  & \b[45]  ;
  assign n11401 = n133 & n11400 ;
  assign n11402 = \b[44]  & n141 ;
  assign n11403 = ~\a[1]  & \b[43]  ;
  assign n11404 = n10416 & n11403 ;
  assign n11405 = ~n11402 & ~n11404 ;
  assign n11406 = ~n11401 & n11405 ;
  assign n11407 = ~n11399 & n11406 ;
  assign n11408 = ~\a[2]  & ~n11407 ;
  assign n11409 = \a[2]  & n11406 ;
  assign n11410 = ~n11399 & n11409 ;
  assign n11411 = ~n11408 & ~n11410 ;
  assign n11412 = ~n11390 & n11411 ;
  assign n11413 = ~n10923 & n11412 ;
  assign n11414 = n11390 & n11411 ;
  assign n11415 = n10923 & n11414 ;
  assign n11416 = ~n11413 & ~n11415 ;
  assign n11417 = ~n10923 & ~n11390 ;
  assign n11418 = ~n10881 & n11390 ;
  assign n11419 = ~n10922 & n11418 ;
  assign n11420 = ~n11411 & ~n11419 ;
  assign n11421 = ~n11417 & n11420 ;
  assign n11422 = n11416 & ~n11421 ;
  assign n11423 = ~n10920 & n11422 ;
  assign n11424 = n10920 & ~n11422 ;
  assign n11425 = ~n11423 & ~n11424 ;
  assign n11426 = ~n10910 & ~n11421 ;
  assign n11427 = ~n10917 & n11426 ;
  assign n11428 = n11416 & ~n11427 ;
  assign n11429 = n11384 & ~n11419 ;
  assign n11430 = n252 & ~n10409 ;
  assign n11431 = ~n10407 & n11430 ;
  assign n11432 = \b[43]  & n250 ;
  assign n11433 = \a[3]  & \b[42]  ;
  assign n11434 = n241 & n11433 ;
  assign n11435 = ~n11432 & ~n11434 ;
  assign n11436 = \b[41]  & n303 ;
  assign n11437 = n300 & n11436 ;
  assign n11438 = ~\a[3]  & \b[42]  ;
  assign n11439 = n244 & n11438 ;
  assign n11440 = ~n11437 & ~n11439 ;
  assign n11441 = n11435 & n11440 ;
  assign n11442 = ~n11431 & n11441 ;
  assign n11443 = ~\a[5]  & ~n11442 ;
  assign n11444 = \a[5]  & n11441 ;
  assign n11445 = ~n11431 & n11444 ;
  assign n11446 = ~n11443 & ~n11445 ;
  assign n11447 = ~n10870 & n11349 ;
  assign n11448 = ~n10877 & n11447 ;
  assign n11449 = n11354 & ~n11448 ;
  assign n11450 = n10927 & n11327 ;
  assign n11451 = ~n11321 & ~n11450 ;
  assign n11452 = ~n10814 & n11286 ;
  assign n11453 = ~n10928 & n11452 ;
  assign n11454 = n11291 & ~n11453 ;
  assign n11455 = n10932 & n11264 ;
  assign n11456 = ~n11258 & ~n11455 ;
  assign n11457 = n10792 & n11223 ;
  assign n11458 = ~n10933 & n11457 ;
  assign n11459 = n11228 & ~n11458 ;
  assign n11460 = n1467 & ~n5462 ;
  assign n11461 = ~n5460 & n11460 ;
  assign n11462 = \b[31]  & n1465 ;
  assign n11463 = \a[15]  & \b[30]  ;
  assign n11464 = n1456 & n11463 ;
  assign n11465 = ~n11462 & ~n11464 ;
  assign n11466 = \b[29]  & n1652 ;
  assign n11467 = n1649 & n11466 ;
  assign n11468 = ~\a[15]  & \b[30]  ;
  assign n11469 = n1459 & n11468 ;
  assign n11470 = ~n11467 & ~n11469 ;
  assign n11471 = n11465 & n11470 ;
  assign n11472 = ~n11461 & n11471 ;
  assign n11473 = ~\a[17]  & ~n11472 ;
  assign n11474 = \a[17]  & n11471 ;
  assign n11475 = ~n11461 & n11474 ;
  assign n11476 = ~n11473 & ~n11475 ;
  assign n11477 = n10937 & n11198 ;
  assign n11478 = n11197 & ~n11477 ;
  assign n11479 = n1965 & n4456 ;
  assign n11480 = ~n4453 & n11479 ;
  assign n11481 = n1965 & ~n4456 ;
  assign n11482 = ~n4143 & n11481 ;
  assign n11483 = ~n4452 & n11482 ;
  assign n11484 = \b[26]  & n2218 ;
  assign n11485 = n2216 & n11484 ;
  assign n11486 = ~\a[18]  & \b[27]  ;
  assign n11487 = n1957 & n11486 ;
  assign n11488 = ~n11485 & ~n11487 ;
  assign n11489 = \b[28]  & n1963 ;
  assign n11490 = \a[18]  & \b[27]  ;
  assign n11491 = n2210 & n11490 ;
  assign n11492 = \a[20]  & ~n11491 ;
  assign n11493 = ~n11489 & n11492 ;
  assign n11494 = n11488 & n11493 ;
  assign n11495 = ~n11483 & n11494 ;
  assign n11496 = ~n11480 & n11495 ;
  assign n11497 = ~n11489 & ~n11491 ;
  assign n11498 = n11488 & n11497 ;
  assign n11499 = ~n11483 & n11498 ;
  assign n11500 = ~n11480 & n11499 ;
  assign n11501 = ~\a[20]  & ~n11500 ;
  assign n11502 = ~n11496 & ~n11501 ;
  assign n11503 = ~n10753 & n11163 ;
  assign n11504 = ~n10761 & n11503 ;
  assign n11505 = n11168 & ~n11504 ;
  assign n11506 = n10941 & n11134 ;
  assign n11507 = ~n11128 & ~n11506 ;
  assign n11508 = n10713 & n11094 ;
  assign n11509 = ~n10942 & n11508 ;
  assign n11510 = n11099 & ~n11509 ;
  assign n11511 = n10946 & n11089 ;
  assign n11512 = ~n11083 & ~n11511 ;
  assign n11513 = ~n10695 & n11055 ;
  assign n11514 = ~n10698 & n11513 ;
  assign n11515 = n11050 & ~n11514 ;
  assign n11516 = ~n948 & n6309 ;
  assign n11517 = ~n908 & n6309 ;
  assign n11518 = ~n912 & n11517 ;
  assign n11519 = ~n11516 & ~n11518 ;
  assign n11520 = ~n951 & ~n11519 ;
  assign n11521 = \b[11]  & n6778 ;
  assign n11522 = n6775 & n11521 ;
  assign n11523 = \b[13]  & n6307 ;
  assign n11524 = \a[33]  & \b[12]  ;
  assign n11525 = n6298 & n11524 ;
  assign n11526 = ~\a[33]  & \b[12]  ;
  assign n11527 = n6301 & n11526 ;
  assign n11528 = ~n11525 & ~n11527 ;
  assign n11529 = ~n11523 & n11528 ;
  assign n11530 = ~n11522 & n11529 ;
  assign n11531 = ~\a[35]  & n11530 ;
  assign n11532 = ~n11520 & n11531 ;
  assign n11533 = \a[35]  & ~n11530 ;
  assign n11534 = \a[35]  & ~n951 ;
  assign n11535 = ~n11519 & n11534 ;
  assign n11536 = ~n11533 & ~n11535 ;
  assign n11537 = ~n11532 & n11536 ;
  assign n11538 = n10969 & n11023 ;
  assign n11539 = ~n11021 & ~n11538 ;
  assign n11540 = ~n10991 & ~n10994 ;
  assign n11541 = n222 & n10082 ;
  assign n11542 = \b[4]  & n10080 ;
  assign n11543 = \a[41]  & \b[3]  ;
  assign n11544 = n10679 & n11543 ;
  assign n11545 = ~\a[42]  & \b[3]  ;
  assign n11546 = n10074 & n11545 ;
  assign n11547 = ~n11544 & ~n11546 ;
  assign n11548 = ~n11542 & n11547 ;
  assign n11549 = \b[2]  & n10681 ;
  assign n11550 = n10678 & n11549 ;
  assign n11551 = \a[44]  & ~n11550 ;
  assign n11552 = n11548 & n11551 ;
  assign n11553 = ~n11541 & n11552 ;
  assign n11554 = n11548 & ~n11550 ;
  assign n11555 = ~n11541 & n11554 ;
  assign n11556 = ~\a[44]  & ~n11555 ;
  assign n11557 = ~n11553 & ~n11556 ;
  assign n11558 = \a[47]  & \b[0]  ;
  assign n11559 = ~n10988 & n11558 ;
  assign n11560 = \a[45]  & \b[0]  ;
  assign n11561 = \a[44]  & ~\a[46]  ;
  assign n11562 = n11560 & n11561 ;
  assign n11563 = ~\a[45]  & \b[0]  ;
  assign n11564 = ~\a[44]  & \a[46]  ;
  assign n11565 = n11563 & n11564 ;
  assign n11566 = ~n11562 & ~n11565 ;
  assign n11567 = \a[46]  & ~\a[47]  ;
  assign n11568 = ~\a[46]  & \a[47]  ;
  assign n11569 = ~n11567 & ~n11568 ;
  assign n11570 = ~n10988 & n11569 ;
  assign n11571 = \b[1]  & n11570 ;
  assign n11572 = ~n10988 & ~n11569 ;
  assign n11573 = ~n137 & n11572 ;
  assign n11574 = ~n11571 & ~n11573 ;
  assign n11575 = n11566 & n11574 ;
  assign n11576 = ~n11559 & ~n11575 ;
  assign n11577 = n11559 & n11566 ;
  assign n11578 = n11574 & n11577 ;
  assign n11579 = ~n11576 & ~n11578 ;
  assign n11580 = n11557 & n11579 ;
  assign n11581 = ~n11557 & ~n11579 ;
  assign n11582 = ~n11580 & ~n11581 ;
  assign n11583 = ~n11540 & n11582 ;
  assign n11584 = n11540 & ~n11582 ;
  assign n11585 = ~n11583 & ~n11584 ;
  assign n11586 = ~n383 & n8759 ;
  assign n11587 = ~n381 & n11586 ;
  assign n11588 = \b[5]  & n9301 ;
  assign n11589 = n9298 & n11588 ;
  assign n11590 = ~\a[39]  & \b[6]  ;
  assign n11591 = n8751 & n11590 ;
  assign n11592 = ~n11589 & ~n11591 ;
  assign n11593 = \b[7]  & n8757 ;
  assign n11594 = \a[39]  & \b[6]  ;
  assign n11595 = n8748 & n11594 ;
  assign n11596 = \a[41]  & ~n11595 ;
  assign n11597 = ~n11593 & n11596 ;
  assign n11598 = n11592 & n11597 ;
  assign n11599 = ~n11587 & n11598 ;
  assign n11600 = ~n11593 & ~n11595 ;
  assign n11601 = n11592 & n11600 ;
  assign n11602 = ~n11587 & n11601 ;
  assign n11603 = ~\a[41]  & ~n11602 ;
  assign n11604 = ~n11599 & ~n11603 ;
  assign n11605 = n11585 & ~n11604 ;
  assign n11606 = ~n11585 & n11604 ;
  assign n11607 = ~n11605 & ~n11606 ;
  assign n11608 = n685 & n7534 ;
  assign n11609 = ~n682 & n11608 ;
  assign n11610 = ~n584 & ~n685 ;
  assign n11611 = n7534 & n11610 ;
  assign n11612 = ~n681 & n11611 ;
  assign n11613 = \b[8]  & n7973 ;
  assign n11614 = n7970 & n11613 ;
  assign n11615 = \b[10]  & n7532 ;
  assign n11616 = \a[36]  & \b[9]  ;
  assign n11617 = n7523 & n11616 ;
  assign n11618 = ~\a[36]  & \b[9]  ;
  assign n11619 = n7526 & n11618 ;
  assign n11620 = ~n11617 & ~n11619 ;
  assign n11621 = ~n11615 & n11620 ;
  assign n11622 = ~n11614 & n11621 ;
  assign n11623 = ~n11612 & n11622 ;
  assign n11624 = ~n11609 & n11623 ;
  assign n11625 = ~\a[38]  & ~n11624 ;
  assign n11626 = \a[38]  & n11622 ;
  assign n11627 = ~n11612 & n11626 ;
  assign n11628 = ~n11609 & n11627 ;
  assign n11629 = ~n11625 & ~n11628 ;
  assign n11630 = ~n11607 & ~n11629 ;
  assign n11631 = ~n11539 & n11630 ;
  assign n11632 = n11607 & ~n11629 ;
  assign n11633 = n11539 & n11632 ;
  assign n11634 = ~n11631 & ~n11633 ;
  assign n11635 = ~n11607 & n11629 ;
  assign n11636 = n11539 & n11635 ;
  assign n11637 = n11607 & n11629 ;
  assign n11638 = ~n11539 & n11637 ;
  assign n11639 = ~n11636 & ~n11638 ;
  assign n11640 = n11634 & n11639 ;
  assign n11641 = ~n11537 & ~n11640 ;
  assign n11642 = ~n11515 & n11641 ;
  assign n11643 = ~n11537 & n11640 ;
  assign n11644 = n11515 & n11643 ;
  assign n11645 = ~n11642 & ~n11644 ;
  assign n11646 = n11537 & ~n11640 ;
  assign n11647 = n11515 & n11646 ;
  assign n11648 = n11537 & n11640 ;
  assign n11649 = ~n11515 & n11648 ;
  assign n11650 = ~n11647 & ~n11649 ;
  assign n11651 = n11645 & n11650 ;
  assign n11652 = ~n11512 & n11651 ;
  assign n11653 = ~n11083 & ~n11651 ;
  assign n11654 = ~n11511 & n11653 ;
  assign n11655 = n1512 & n5211 ;
  assign n11656 = ~n1509 & n11655 ;
  assign n11657 = n5211 & n10165 ;
  assign n11658 = ~n1508 & n11657 ;
  assign n11659 = \b[14]  & n5595 ;
  assign n11660 = n5592 & n11659 ;
  assign n11661 = ~\a[30]  & \b[15]  ;
  assign n11662 = n5203 & n11661 ;
  assign n11663 = ~n11660 & ~n11662 ;
  assign n11664 = \b[16]  & n5209 ;
  assign n11665 = \a[30]  & \b[15]  ;
  assign n11666 = n5200 & n11665 ;
  assign n11667 = \a[32]  & ~n11666 ;
  assign n11668 = ~n11664 & n11667 ;
  assign n11669 = n11663 & n11668 ;
  assign n11670 = ~n11658 & n11669 ;
  assign n11671 = ~n11656 & n11670 ;
  assign n11672 = ~n11664 & ~n11666 ;
  assign n11673 = n11663 & n11672 ;
  assign n11674 = ~n11658 & n11673 ;
  assign n11675 = ~n11656 & n11674 ;
  assign n11676 = ~\a[32]  & ~n11675 ;
  assign n11677 = ~n11671 & ~n11676 ;
  assign n11678 = ~n11654 & ~n11677 ;
  assign n11679 = ~n11652 & n11678 ;
  assign n11680 = ~n11651 & n11677 ;
  assign n11681 = n11512 & n11680 ;
  assign n11682 = n11651 & n11677 ;
  assign n11683 = ~n11512 & n11682 ;
  assign n11684 = ~n11681 & ~n11683 ;
  assign n11685 = ~n11679 & n11684 ;
  assign n11686 = ~n2076 & n4249 ;
  assign n11687 = ~n1874 & n4249 ;
  assign n11688 = ~n1878 & n11687 ;
  assign n11689 = ~n11686 & ~n11688 ;
  assign n11690 = ~n2079 & ~n11689 ;
  assign n11691 = \b[17]  & n4647 ;
  assign n11692 = n4644 & n11691 ;
  assign n11693 = ~\a[27]  & \b[18]  ;
  assign n11694 = n4241 & n11693 ;
  assign n11695 = ~n11692 & ~n11694 ;
  assign n11696 = \b[19]  & n4247 ;
  assign n11697 = \a[27]  & \b[18]  ;
  assign n11698 = n4238 & n11697 ;
  assign n11699 = \a[29]  & ~n11698 ;
  assign n11700 = ~n11696 & n11699 ;
  assign n11701 = n11695 & n11700 ;
  assign n11702 = ~n11690 & n11701 ;
  assign n11703 = ~n11696 & ~n11698 ;
  assign n11704 = n11695 & n11703 ;
  assign n11705 = ~\a[29]  & ~n11704 ;
  assign n11706 = ~\a[29]  & ~n2079 ;
  assign n11707 = ~n11689 & n11706 ;
  assign n11708 = ~n11705 & ~n11707 ;
  assign n11709 = ~n11702 & n11708 ;
  assign n11710 = ~n11685 & ~n11709 ;
  assign n11711 = n11510 & n11710 ;
  assign n11712 = n11685 & ~n11709 ;
  assign n11713 = ~n11510 & n11712 ;
  assign n11714 = ~n11711 & ~n11713 ;
  assign n11715 = ~n11685 & n11709 ;
  assign n11716 = ~n11510 & n11715 ;
  assign n11717 = n11685 & n11709 ;
  assign n11718 = n11510 & n11717 ;
  assign n11719 = ~n11716 & ~n11718 ;
  assign n11720 = n11714 & n11719 ;
  assign n11721 = ~n11507 & n11720 ;
  assign n11722 = ~n11128 & ~n11720 ;
  assign n11723 = ~n11506 & n11722 ;
  assign n11724 = ~n2768 & ~n3154 ;
  assign n11725 = ~n3399 & n11724 ;
  assign n11726 = n2765 & n11725 ;
  assign n11727 = n2768 & ~n3154 ;
  assign n11728 = ~n3399 & n11727 ;
  assign n11729 = ~n2765 & n11728 ;
  assign n11730 = ~n11726 & ~n11729 ;
  assign n11731 = \b[20]  & n3733 ;
  assign n11732 = n3730 & n11731 ;
  assign n11733 = ~\a[24]  & \b[21]  ;
  assign n11734 = n3394 & n11733 ;
  assign n11735 = ~n11732 & ~n11734 ;
  assign n11736 = \b[22]  & n3400 ;
  assign n11737 = \a[24]  & \b[21]  ;
  assign n11738 = n3391 & n11737 ;
  assign n11739 = \a[26]  & ~n11738 ;
  assign n11740 = ~n11736 & n11739 ;
  assign n11741 = n11735 & n11740 ;
  assign n11742 = n11730 & n11741 ;
  assign n11743 = ~n11736 & ~n11738 ;
  assign n11744 = n11735 & n11743 ;
  assign n11745 = n11730 & n11744 ;
  assign n11746 = ~\a[26]  & ~n11745 ;
  assign n11747 = ~n11742 & ~n11746 ;
  assign n11748 = ~n11723 & ~n11747 ;
  assign n11749 = ~n11721 & n11748 ;
  assign n11750 = ~n11720 & n11747 ;
  assign n11751 = n11507 & n11750 ;
  assign n11752 = n11720 & n11747 ;
  assign n11753 = ~n11507 & n11752 ;
  assign n11754 = ~n11751 & ~n11753 ;
  assign n11755 = ~n11749 & n11754 ;
  assign n11756 = ~n11505 & ~n11755 ;
  assign n11757 = n11505 & n11755 ;
  assign n11758 = ~n11756 & ~n11757 ;
  assign n11759 = n2622 & ~n3567 ;
  assign n11760 = ~n3565 & n11759 ;
  assign n11761 = \b[23]  & n2912 ;
  assign n11762 = n2909 & n11761 ;
  assign n11763 = \b[25]  & n2620 ;
  assign n11764 = \a[21]  & \b[24]  ;
  assign n11765 = n2611 & n11764 ;
  assign n11766 = ~\a[21]  & \b[24]  ;
  assign n11767 = n2614 & n11766 ;
  assign n11768 = ~n11765 & ~n11767 ;
  assign n11769 = ~n11763 & n11768 ;
  assign n11770 = ~n11762 & n11769 ;
  assign n11771 = ~\a[23]  & n11770 ;
  assign n11772 = ~n11760 & n11771 ;
  assign n11773 = ~n11760 & n11770 ;
  assign n11774 = \a[23]  & ~n11773 ;
  assign n11775 = ~n11772 & ~n11774 ;
  assign n11776 = n11758 & n11775 ;
  assign n11777 = ~n11758 & ~n11775 ;
  assign n11778 = ~n11776 & ~n11777 ;
  assign n11779 = ~n11502 & ~n11778 ;
  assign n11780 = ~n11478 & n11779 ;
  assign n11781 = ~n11502 & n11778 ;
  assign n11782 = n11478 & n11781 ;
  assign n11783 = ~n11780 & ~n11782 ;
  assign n11784 = n11502 & ~n11778 ;
  assign n11785 = n11478 & n11784 ;
  assign n11786 = n11502 & n11778 ;
  assign n11787 = ~n11478 & n11786 ;
  assign n11788 = ~n11785 & ~n11787 ;
  assign n11789 = n11783 & n11788 ;
  assign n11790 = n11476 & ~n11789 ;
  assign n11791 = ~n11459 & n11790 ;
  assign n11792 = n11476 & n11789 ;
  assign n11793 = n11459 & n11792 ;
  assign n11794 = ~n11791 & ~n11793 ;
  assign n11795 = ~n11476 & ~n11789 ;
  assign n11796 = n11459 & n11795 ;
  assign n11797 = ~n11476 & n11789 ;
  assign n11798 = ~n11459 & n11797 ;
  assign n11799 = ~n11796 & ~n11798 ;
  assign n11800 = n11794 & n11799 ;
  assign n11801 = ~n11456 & n11800 ;
  assign n11802 = ~n11258 & ~n11800 ;
  assign n11803 = ~n11455 & n11802 ;
  assign n11804 = ~n847 & ~n5850 ;
  assign n11805 = ~n6565 & n11804 ;
  assign n11806 = ~n6561 & n11805 ;
  assign n11807 = ~n996 & n11806 ;
  assign n11808 = n999 & n6565 ;
  assign n11809 = ~n6562 & n11808 ;
  assign n11810 = ~n11807 & ~n11809 ;
  assign n11811 = \b[32]  & n1182 ;
  assign n11812 = n1179 & n11811 ;
  assign n11813 = \b[34]  & n997 ;
  assign n11814 = \a[11]  & \b[33]  ;
  assign n11815 = n1180 & n11814 ;
  assign n11816 = ~\a[12]  & \b[33]  ;
  assign n11817 = n7674 & n11816 ;
  assign n11818 = ~n11815 & ~n11817 ;
  assign n11819 = ~n11813 & n11818 ;
  assign n11820 = ~n11812 & n11819 ;
  assign n11821 = n11810 & n11820 ;
  assign n11822 = ~\a[14]  & ~n11821 ;
  assign n11823 = \a[14]  & n11820 ;
  assign n11824 = n11810 & n11823 ;
  assign n11825 = ~n11822 & ~n11824 ;
  assign n11826 = ~n11803 & ~n11825 ;
  assign n11827 = ~n11801 & n11826 ;
  assign n11828 = ~n11800 & n11825 ;
  assign n11829 = n11456 & n11828 ;
  assign n11830 = n11800 & n11825 ;
  assign n11831 = ~n11456 & n11830 ;
  assign n11832 = ~n11829 & ~n11831 ;
  assign n11833 = ~n11827 & n11832 ;
  assign n11834 = n646 & ~n7761 ;
  assign n11835 = ~n7759 & n11834 ;
  assign n11836 = \b[37]  & n644 ;
  assign n11837 = \a[9]  & \b[36]  ;
  assign n11838 = n635 & n11837 ;
  assign n11839 = ~n11836 & ~n11838 ;
  assign n11840 = \b[35]  & n796 ;
  assign n11841 = n793 & n11840 ;
  assign n11842 = ~\a[9]  & \b[36]  ;
  assign n11843 = n638 & n11842 ;
  assign n11844 = ~n11841 & ~n11843 ;
  assign n11845 = n11839 & n11844 ;
  assign n11846 = ~n11835 & n11845 ;
  assign n11847 = ~\a[11]  & ~n11846 ;
  assign n11848 = \a[11]  & n11845 ;
  assign n11849 = ~n11835 & n11848 ;
  assign n11850 = ~n11847 & ~n11849 ;
  assign n11851 = ~n11833 & ~n11850 ;
  assign n11852 = n11454 & n11851 ;
  assign n11853 = n11833 & ~n11850 ;
  assign n11854 = ~n11454 & n11853 ;
  assign n11855 = ~n11852 & ~n11854 ;
  assign n11856 = ~n11833 & n11850 ;
  assign n11857 = ~n11454 & n11856 ;
  assign n11858 = n11833 & n11850 ;
  assign n11859 = n11454 & n11858 ;
  assign n11860 = ~n11857 & ~n11859 ;
  assign n11861 = n11855 & n11860 ;
  assign n11862 = ~n11451 & n11861 ;
  assign n11863 = ~n11321 & ~n11861 ;
  assign n11864 = ~n11450 & n11863 ;
  assign n11865 = n430 & n9044 ;
  assign n11866 = ~n9041 & n11865 ;
  assign n11867 = n430 & ~n9044 ;
  assign n11868 = ~n8597 & n11867 ;
  assign n11869 = ~n9040 & n11868 ;
  assign n11870 = \b[38]  & n486 ;
  assign n11871 = n483 & n11870 ;
  assign n11872 = \b[40]  & n428 ;
  assign n11873 = \a[6]  & \b[39]  ;
  assign n11874 = n419 & n11873 ;
  assign n11875 = ~\a[6]  & \b[39]  ;
  assign n11876 = n422 & n11875 ;
  assign n11877 = ~n11874 & ~n11876 ;
  assign n11878 = ~n11872 & n11877 ;
  assign n11879 = ~n11871 & n11878 ;
  assign n11880 = ~n11869 & n11879 ;
  assign n11881 = ~n11866 & n11880 ;
  assign n11882 = ~\a[8]  & ~n11881 ;
  assign n11883 = \a[8]  & n11879 ;
  assign n11884 = ~n11869 & n11883 ;
  assign n11885 = ~n11866 & n11884 ;
  assign n11886 = ~n11882 & ~n11885 ;
  assign n11887 = ~n11864 & ~n11886 ;
  assign n11888 = ~n11862 & n11887 ;
  assign n11889 = ~n11861 & n11886 ;
  assign n11890 = n11451 & n11889 ;
  assign n11891 = n11861 & n11886 ;
  assign n11892 = ~n11451 & n11891 ;
  assign n11893 = ~n11890 & ~n11892 ;
  assign n11894 = ~n11888 & n11893 ;
  assign n11895 = n11449 & n11894 ;
  assign n11896 = ~n11449 & ~n11894 ;
  assign n11897 = ~n11895 & ~n11896 ;
  assign n11898 = ~n11446 & n11897 ;
  assign n11899 = n11446 & ~n11897 ;
  assign n11900 = ~n11898 & ~n11899 ;
  assign n11901 = ~n10888 & ~n11393 ;
  assign n11902 = ~n10892 & n11901 ;
  assign n11903 = ~n11392 & ~n11902 ;
  assign n11904 = ~\b[45]  & ~\b[46]  ;
  assign n11905 = \b[45]  & \b[46]  ;
  assign n11906 = ~n11904 & ~n11905 ;
  assign n11907 = n134 & n11906 ;
  assign n11908 = ~n11903 & n11907 ;
  assign n11909 = n134 & ~n11906 ;
  assign n11910 = ~n11392 & n11909 ;
  assign n11911 = ~n11902 & n11910 ;
  assign n11912 = \a[0]  & \b[46]  ;
  assign n11913 = n133 & n11912 ;
  assign n11914 = \b[45]  & n141 ;
  assign n11915 = ~\a[1]  & \b[44]  ;
  assign n11916 = n10416 & n11915 ;
  assign n11917 = ~n11914 & ~n11916 ;
  assign n11918 = ~n11913 & n11917 ;
  assign n11919 = \a[2]  & n11918 ;
  assign n11920 = ~n11911 & n11919 ;
  assign n11921 = ~n11908 & n11920 ;
  assign n11922 = ~n11911 & n11918 ;
  assign n11923 = ~n11908 & n11922 ;
  assign n11924 = ~\a[2]  & ~n11923 ;
  assign n11925 = ~n11921 & ~n11924 ;
  assign n11926 = ~n11900 & ~n11925 ;
  assign n11927 = ~n11429 & n11926 ;
  assign n11928 = n11900 & ~n11925 ;
  assign n11929 = n11429 & n11928 ;
  assign n11930 = ~n11927 & ~n11929 ;
  assign n11931 = ~n11900 & n11925 ;
  assign n11932 = n11429 & n11931 ;
  assign n11933 = n11900 & n11925 ;
  assign n11934 = ~n11429 & n11933 ;
  assign n11935 = ~n11932 & ~n11934 ;
  assign n11936 = n11930 & n11935 ;
  assign n11937 = n11428 & n11936 ;
  assign n11938 = ~n11428 & ~n11936 ;
  assign n11939 = ~n11937 & ~n11938 ;
  assign n11940 = n11930 & ~n11937 ;
  assign n11941 = n11384 & ~n11898 ;
  assign n11942 = ~n11419 & n11941 ;
  assign n11943 = ~n11899 & ~n11942 ;
  assign n11944 = ~n11888 & ~n11895 ;
  assign n11945 = n252 & ~n10892 ;
  assign n11946 = ~n10890 & n11945 ;
  assign n11947 = \b[42]  & n303 ;
  assign n11948 = n300 & n11947 ;
  assign n11949 = ~\a[3]  & \b[43]  ;
  assign n11950 = n244 & n11949 ;
  assign n11951 = ~n11948 & ~n11950 ;
  assign n11952 = \b[44]  & n250 ;
  assign n11953 = \a[3]  & \b[43]  ;
  assign n11954 = n241 & n11953 ;
  assign n11955 = \a[5]  & ~n11954 ;
  assign n11956 = ~n11952 & n11955 ;
  assign n11957 = n11951 & n11956 ;
  assign n11958 = ~n11946 & n11957 ;
  assign n11959 = ~n11952 & ~n11954 ;
  assign n11960 = n11951 & n11959 ;
  assign n11961 = ~n11946 & n11960 ;
  assign n11962 = ~\a[5]  & ~n11961 ;
  assign n11963 = ~n11958 & ~n11962 ;
  assign n11964 = ~n11321 & n11855 ;
  assign n11965 = ~n11450 & n11964 ;
  assign n11966 = n11860 & ~n11965 ;
  assign n11967 = n11454 & n11833 ;
  assign n11968 = ~n11827 & ~n11967 ;
  assign n11969 = ~n11258 & n11799 ;
  assign n11970 = ~n11455 & n11969 ;
  assign n11971 = n11794 & ~n11970 ;
  assign n11972 = n11459 & n11789 ;
  assign n11973 = n11783 & ~n11972 ;
  assign n11974 = n1467 & n5810 ;
  assign n11975 = ~n5807 & n11974 ;
  assign n11976 = n1467 & ~n5810 ;
  assign n11977 = ~n5457 & n11976 ;
  assign n11978 = ~n5806 & n11977 ;
  assign n11979 = \b[30]  & n1652 ;
  assign n11980 = n1649 & n11979 ;
  assign n11981 = ~\a[15]  & \b[31]  ;
  assign n11982 = n1459 & n11981 ;
  assign n11983 = ~n11980 & ~n11982 ;
  assign n11984 = \b[32]  & n1465 ;
  assign n11985 = \a[15]  & \b[31]  ;
  assign n11986 = n1456 & n11985 ;
  assign n11987 = \a[17]  & ~n11986 ;
  assign n11988 = ~n11984 & n11987 ;
  assign n11989 = n11983 & n11988 ;
  assign n11990 = ~n11978 & n11989 ;
  assign n11991 = ~n11975 & n11990 ;
  assign n11992 = ~n11984 & ~n11986 ;
  assign n11993 = n11983 & n11992 ;
  assign n11994 = ~n11978 & n11993 ;
  assign n11995 = ~n11975 & n11994 ;
  assign n11996 = ~\a[17]  & ~n11995 ;
  assign n11997 = ~n11991 & ~n11996 ;
  assign n11998 = n11197 & ~n11776 ;
  assign n11999 = ~n11477 & n11998 ;
  assign n12000 = ~n11777 & ~n11999 ;
  assign n12001 = n1965 & ~n4502 ;
  assign n12002 = ~n4500 & n12001 ;
  assign n12003 = \b[29]  & n1963 ;
  assign n12004 = \a[18]  & \b[28]  ;
  assign n12005 = n2210 & n12004 ;
  assign n12006 = ~n12003 & ~n12005 ;
  assign n12007 = \b[27]  & n2218 ;
  assign n12008 = n2216 & n12007 ;
  assign n12009 = ~\a[18]  & \b[28]  ;
  assign n12010 = n1957 & n12009 ;
  assign n12011 = ~n12008 & ~n12010 ;
  assign n12012 = n12006 & n12011 ;
  assign n12013 = ~n12002 & n12012 ;
  assign n12014 = ~\a[20]  & ~n12013 ;
  assign n12015 = \a[20]  & n12012 ;
  assign n12016 = ~n12002 & n12015 ;
  assign n12017 = ~n12014 & ~n12016 ;
  assign n12018 = ~n11749 & ~n11757 ;
  assign n12019 = n2622 & n3604 ;
  assign n12020 = ~n3601 & n12019 ;
  assign n12021 = ~n3562 & ~n3604 ;
  assign n12022 = n2622 & n12021 ;
  assign n12023 = ~n3600 & n12022 ;
  assign n12024 = \b[24]  & n2912 ;
  assign n12025 = n2909 & n12024 ;
  assign n12026 = ~\a[21]  & \b[25]  ;
  assign n12027 = n2614 & n12026 ;
  assign n12028 = ~n12025 & ~n12027 ;
  assign n12029 = \b[26]  & n2620 ;
  assign n12030 = \a[21]  & \b[25]  ;
  assign n12031 = n2611 & n12030 ;
  assign n12032 = \a[23]  & ~n12031 ;
  assign n12033 = ~n12029 & n12032 ;
  assign n12034 = n12028 & n12033 ;
  assign n12035 = ~n12023 & n12034 ;
  assign n12036 = ~n12020 & n12035 ;
  assign n12037 = ~n12029 & ~n12031 ;
  assign n12038 = n12028 & n12037 ;
  assign n12039 = ~n12023 & n12038 ;
  assign n12040 = ~n12020 & n12039 ;
  assign n12041 = ~\a[23]  & ~n12040 ;
  assign n12042 = ~n12036 & ~n12041 ;
  assign n12043 = ~n11128 & n11714 ;
  assign n12044 = ~n11506 & n12043 ;
  assign n12045 = n11719 & ~n12044 ;
  assign n12046 = n11510 & n11685 ;
  assign n12047 = ~n11679 & ~n12046 ;
  assign n12048 = ~n11083 & n11650 ;
  assign n12049 = ~n11511 & n12048 ;
  assign n12050 = n11645 & ~n12049 ;
  assign n12051 = ~n1691 & n5211 ;
  assign n12052 = ~n1511 & n5211 ;
  assign n12053 = ~n1515 & n12052 ;
  assign n12054 = ~n12051 & ~n12053 ;
  assign n12055 = ~n1694 & ~n12054 ;
  assign n12056 = \b[15]  & n5595 ;
  assign n12057 = n5592 & n12056 ;
  assign n12058 = ~\a[30]  & \b[16]  ;
  assign n12059 = n5203 & n12058 ;
  assign n12060 = ~n12057 & ~n12059 ;
  assign n12061 = \b[17]  & n5209 ;
  assign n12062 = \a[30]  & \b[16]  ;
  assign n12063 = n5200 & n12062 ;
  assign n12064 = \a[32]  & ~n12063 ;
  assign n12065 = ~n12061 & n12064 ;
  assign n12066 = n12060 & n12065 ;
  assign n12067 = ~n12055 & n12066 ;
  assign n12068 = ~n12061 & ~n12063 ;
  assign n12069 = n12060 & n12068 ;
  assign n12070 = ~\a[32]  & ~n12069 ;
  assign n12071 = ~\a[32]  & ~n1694 ;
  assign n12072 = ~n12054 & n12071 ;
  assign n12073 = ~n12070 & ~n12072 ;
  assign n12074 = ~n12067 & n12073 ;
  assign n12075 = n11515 & n11640 ;
  assign n12076 = n11634 & ~n12075 ;
  assign n12077 = ~n725 & n7534 ;
  assign n12078 = ~n684 & n7534 ;
  assign n12079 = ~n721 & n12078 ;
  assign n12080 = ~n12077 & ~n12079 ;
  assign n12081 = ~n728 & ~n12080 ;
  assign n12082 = \b[9]  & n7973 ;
  assign n12083 = n7970 & n12082 ;
  assign n12084 = \b[11]  & n7532 ;
  assign n12085 = \a[36]  & \b[10]  ;
  assign n12086 = n7523 & n12085 ;
  assign n12087 = ~\a[36]  & \b[10]  ;
  assign n12088 = n7526 & n12087 ;
  assign n12089 = ~n12086 & ~n12088 ;
  assign n12090 = ~n12084 & n12089 ;
  assign n12091 = ~n12083 & n12090 ;
  assign n12092 = ~\a[38]  & n12091 ;
  assign n12093 = ~n12081 & n12092 ;
  assign n12094 = \a[38]  & ~n12091 ;
  assign n12095 = \a[38]  & ~n728 ;
  assign n12096 = ~n12080 & n12095 ;
  assign n12097 = ~n12094 & ~n12096 ;
  assign n12098 = ~n12093 & n12097 ;
  assign n12099 = ~n11021 & ~n11605 ;
  assign n12100 = ~n11538 & n12099 ;
  assign n12101 = ~n11606 & ~n12100 ;
  assign n12102 = ~n505 & ~n8272 ;
  assign n12103 = ~n8756 & n12102 ;
  assign n12104 = n502 & n12103 ;
  assign n12105 = n505 & ~n8272 ;
  assign n12106 = ~n8756 & n12105 ;
  assign n12107 = ~n502 & n12106 ;
  assign n12108 = ~n12104 & ~n12107 ;
  assign n12109 = \b[6]  & n9301 ;
  assign n12110 = n9298 & n12109 ;
  assign n12111 = ~\a[39]  & \b[7]  ;
  assign n12112 = n8751 & n12111 ;
  assign n12113 = ~n12110 & ~n12112 ;
  assign n12114 = \b[8]  & n8757 ;
  assign n12115 = \a[39]  & \b[7]  ;
  assign n12116 = n8748 & n12115 ;
  assign n12117 = \a[41]  & ~n12116 ;
  assign n12118 = ~n12114 & n12117 ;
  assign n12119 = n12113 & n12118 ;
  assign n12120 = n12108 & n12119 ;
  assign n12121 = ~n12114 & ~n12116 ;
  assign n12122 = n12113 & n12121 ;
  assign n12123 = n12108 & n12122 ;
  assign n12124 = ~\a[41]  & ~n12123 ;
  assign n12125 = ~n12120 & ~n12124 ;
  assign n12126 = ~n11581 & ~n11583 ;
  assign n12127 = ~n273 & n10082 ;
  assign n12128 = ~n271 & n12127 ;
  assign n12129 = \b[3]  & n10681 ;
  assign n12130 = n10678 & n12129 ;
  assign n12131 = \b[5]  & n10080 ;
  assign n12132 = \a[41]  & \b[4]  ;
  assign n12133 = n10679 & n12132 ;
  assign n12134 = ~\a[42]  & \b[4]  ;
  assign n12135 = n10074 & n12134 ;
  assign n12136 = ~n12133 & ~n12135 ;
  assign n12137 = ~n12131 & n12136 ;
  assign n12138 = ~n12130 & n12137 ;
  assign n12139 = ~n12128 & n12138 ;
  assign n12140 = ~\a[44]  & ~n12139 ;
  assign n12141 = \a[44]  & n12138 ;
  assign n12142 = ~n12128 & n12141 ;
  assign n12143 = ~n12140 & ~n12142 ;
  assign n12144 = \a[47]  & ~n10989 ;
  assign n12145 = n11566 & n12144 ;
  assign n12146 = n11574 & n12145 ;
  assign n12147 = \a[47]  & ~n12146 ;
  assign n12148 = \b[2]  & n11570 ;
  assign n12149 = ~\a[45]  & \b[1]  ;
  assign n12150 = n11564 & n12149 ;
  assign n12151 = \a[45]  & \b[1]  ;
  assign n12152 = n11561 & n12151 ;
  assign n12153 = ~n12150 & ~n12152 ;
  assign n12154 = ~n12148 & n12153 ;
  assign n12155 = n157 & n11572 ;
  assign n12156 = n10988 & ~n11569 ;
  assign n12157 = \a[45]  & ~\a[46]  ;
  assign n12158 = ~\a[45]  & \a[46]  ;
  assign n12159 = ~n12157 & ~n12158 ;
  assign n12160 = \b[0]  & n12159 ;
  assign n12161 = n12156 & n12160 ;
  assign n12162 = ~n12155 & ~n12161 ;
  assign n12163 = n12154 & n12162 ;
  assign n12164 = ~n12147 & ~n12163 ;
  assign n12165 = n12147 & n12163 ;
  assign n12166 = ~n12164 & ~n12165 ;
  assign n12167 = ~n12143 & ~n12166 ;
  assign n12168 = n12143 & n12166 ;
  assign n12169 = ~n12167 & ~n12168 ;
  assign n12170 = ~n12126 & n12169 ;
  assign n12171 = n12126 & ~n12169 ;
  assign n12172 = ~n12170 & ~n12171 ;
  assign n12173 = ~n12125 & n12172 ;
  assign n12174 = n12125 & ~n12172 ;
  assign n12175 = ~n12173 & ~n12174 ;
  assign n12176 = n12101 & n12175 ;
  assign n12177 = ~n12101 & ~n12175 ;
  assign n12178 = ~n12176 & ~n12177 ;
  assign n12179 = ~n12098 & ~n12178 ;
  assign n12180 = n12098 & n12178 ;
  assign n12181 = ~n12179 & ~n12180 ;
  assign n12182 = n1087 & n6309 ;
  assign n12183 = ~n1084 & n12182 ;
  assign n12184 = n1552 & n6309 ;
  assign n12185 = ~n1083 & n12184 ;
  assign n12186 = \b[12]  & n6778 ;
  assign n12187 = n6775 & n12186 ;
  assign n12188 = \b[14]  & n6307 ;
  assign n12189 = \a[33]  & \b[13]  ;
  assign n12190 = n6298 & n12189 ;
  assign n12191 = ~\a[33]  & \b[13]  ;
  assign n12192 = n6301 & n12191 ;
  assign n12193 = ~n12190 & ~n12192 ;
  assign n12194 = ~n12188 & n12193 ;
  assign n12195 = ~n12187 & n12194 ;
  assign n12196 = ~n12185 & n12195 ;
  assign n12197 = ~n12183 & n12196 ;
  assign n12198 = ~\a[35]  & ~n12197 ;
  assign n12199 = \a[35]  & n12195 ;
  assign n12200 = ~n12185 & n12199 ;
  assign n12201 = ~n12183 & n12200 ;
  assign n12202 = ~n12198 & ~n12201 ;
  assign n12203 = ~n12181 & ~n12202 ;
  assign n12204 = ~n12076 & n12203 ;
  assign n12205 = n12181 & ~n12202 ;
  assign n12206 = n12076 & n12205 ;
  assign n12207 = ~n12204 & ~n12206 ;
  assign n12208 = ~n12181 & n12202 ;
  assign n12209 = n12076 & n12208 ;
  assign n12210 = n12181 & n12202 ;
  assign n12211 = ~n12076 & n12210 ;
  assign n12212 = ~n12209 & ~n12211 ;
  assign n12213 = n12207 & n12212 ;
  assign n12214 = ~n12074 & ~n12213 ;
  assign n12215 = n12050 & n12214 ;
  assign n12216 = ~n12074 & n12213 ;
  assign n12217 = ~n12050 & n12216 ;
  assign n12218 = ~n12215 & ~n12217 ;
  assign n12219 = n12074 & ~n12213 ;
  assign n12220 = ~n12050 & n12219 ;
  assign n12221 = n12074 & n12213 ;
  assign n12222 = n12050 & n12221 ;
  assign n12223 = ~n12220 & ~n12222 ;
  assign n12224 = n12218 & n12223 ;
  assign n12225 = ~n12047 & n12224 ;
  assign n12226 = n2293 & n4249 ;
  assign n12227 = ~n2290 & n12226 ;
  assign n12228 = ~n2293 & n4249 ;
  assign n12229 = ~n2074 & n12228 ;
  assign n12230 = ~n2289 & n12229 ;
  assign n12231 = \b[18]  & n4647 ;
  assign n12232 = n4644 & n12231 ;
  assign n12233 = ~\a[27]  & \b[19]  ;
  assign n12234 = n4241 & n12233 ;
  assign n12235 = ~n12232 & ~n12234 ;
  assign n12236 = \b[20]  & n4247 ;
  assign n12237 = \a[27]  & \b[19]  ;
  assign n12238 = n4238 & n12237 ;
  assign n12239 = \a[29]  & ~n12238 ;
  assign n12240 = ~n12236 & n12239 ;
  assign n12241 = n12235 & n12240 ;
  assign n12242 = ~n12230 & n12241 ;
  assign n12243 = ~n12227 & n12242 ;
  assign n12244 = ~n12236 & ~n12238 ;
  assign n12245 = n12235 & n12244 ;
  assign n12246 = ~n12230 & n12245 ;
  assign n12247 = ~n12227 & n12246 ;
  assign n12248 = ~\a[29]  & ~n12247 ;
  assign n12249 = ~n12243 & ~n12248 ;
  assign n12250 = ~n11679 & ~n12224 ;
  assign n12251 = ~n12046 & n12250 ;
  assign n12252 = ~n12249 & ~n12251 ;
  assign n12253 = ~n12225 & n12252 ;
  assign n12254 = ~n12224 & n12249 ;
  assign n12255 = n12047 & n12254 ;
  assign n12256 = n12224 & n12249 ;
  assign n12257 = ~n12047 & n12256 ;
  assign n12258 = ~n12255 & ~n12257 ;
  assign n12259 = ~n12253 & n12258 ;
  assign n12260 = ~n3019 & n3402 ;
  assign n12261 = ~n2767 & n3402 ;
  assign n12262 = ~n2771 & n12261 ;
  assign n12263 = ~n12260 & ~n12262 ;
  assign n12264 = ~n3022 & ~n12263 ;
  assign n12265 = \b[21]  & n3733 ;
  assign n12266 = n3730 & n12265 ;
  assign n12267 = ~\a[24]  & \b[22]  ;
  assign n12268 = n3394 & n12267 ;
  assign n12269 = ~n12266 & ~n12268 ;
  assign n12270 = \b[23]  & n3400 ;
  assign n12271 = \a[24]  & \b[22]  ;
  assign n12272 = n3391 & n12271 ;
  assign n12273 = \a[26]  & ~n12272 ;
  assign n12274 = ~n12270 & n12273 ;
  assign n12275 = n12269 & n12274 ;
  assign n12276 = ~n12264 & n12275 ;
  assign n12277 = ~n12270 & ~n12272 ;
  assign n12278 = n12269 & n12277 ;
  assign n12279 = ~\a[26]  & ~n12278 ;
  assign n12280 = ~\a[26]  & ~n3022 ;
  assign n12281 = ~n12263 & n12280 ;
  assign n12282 = ~n12279 & ~n12281 ;
  assign n12283 = ~n12276 & n12282 ;
  assign n12284 = ~n12259 & ~n12283 ;
  assign n12285 = n12045 & n12284 ;
  assign n12286 = n12259 & ~n12283 ;
  assign n12287 = ~n12045 & n12286 ;
  assign n12288 = ~n12285 & ~n12287 ;
  assign n12289 = ~n12259 & n12283 ;
  assign n12290 = ~n12045 & n12289 ;
  assign n12291 = n12259 & n12283 ;
  assign n12292 = n12045 & n12291 ;
  assign n12293 = ~n12290 & ~n12292 ;
  assign n12294 = n12288 & n12293 ;
  assign n12295 = n12042 & ~n12294 ;
  assign n12296 = n12018 & n12295 ;
  assign n12297 = n12042 & n12294 ;
  assign n12298 = ~n12018 & n12297 ;
  assign n12299 = ~n12296 & ~n12298 ;
  assign n12300 = ~n12042 & ~n12294 ;
  assign n12301 = ~n12018 & n12300 ;
  assign n12302 = ~n12042 & n12294 ;
  assign n12303 = n12018 & n12302 ;
  assign n12304 = ~n12301 & ~n12303 ;
  assign n12305 = n12299 & n12304 ;
  assign n12306 = n12017 & ~n12305 ;
  assign n12307 = ~n12000 & n12306 ;
  assign n12308 = n12017 & n12305 ;
  assign n12309 = n12000 & n12308 ;
  assign n12310 = ~n12307 & ~n12309 ;
  assign n12311 = ~n12017 & ~n12305 ;
  assign n12312 = n12000 & n12311 ;
  assign n12313 = ~n12017 & n12305 ;
  assign n12314 = ~n12000 & n12313 ;
  assign n12315 = ~n12312 & ~n12314 ;
  assign n12316 = n12310 & n12315 ;
  assign n12317 = n11997 & ~n12316 ;
  assign n12318 = n11973 & n12317 ;
  assign n12319 = n11997 & n12316 ;
  assign n12320 = ~n11973 & n12319 ;
  assign n12321 = ~n12318 & ~n12320 ;
  assign n12322 = ~n11973 & n12316 ;
  assign n12323 = n11783 & ~n12316 ;
  assign n12324 = ~n11972 & n12323 ;
  assign n12325 = ~n11997 & ~n12324 ;
  assign n12326 = ~n12322 & n12325 ;
  assign n12327 = n12321 & ~n12326 ;
  assign n12328 = n999 & ~n6610 ;
  assign n12329 = ~n6608 & n12328 ;
  assign n12330 = \b[33]  & n1182 ;
  assign n12331 = n1179 & n12330 ;
  assign n12332 = \b[35]  & n997 ;
  assign n12333 = \a[11]  & \b[34]  ;
  assign n12334 = n1180 & n12333 ;
  assign n12335 = ~\a[12]  & \b[34]  ;
  assign n12336 = n7674 & n12335 ;
  assign n12337 = ~n12334 & ~n12336 ;
  assign n12338 = ~n12332 & n12337 ;
  assign n12339 = ~n12331 & n12338 ;
  assign n12340 = ~n12329 & n12339 ;
  assign n12341 = ~\a[14]  & ~n12340 ;
  assign n12342 = \a[14]  & n12339 ;
  assign n12343 = ~n12329 & n12342 ;
  assign n12344 = ~n12341 & ~n12343 ;
  assign n12345 = ~n12327 & ~n12344 ;
  assign n12346 = n11971 & n12345 ;
  assign n12347 = n12327 & ~n12344 ;
  assign n12348 = ~n11971 & n12347 ;
  assign n12349 = ~n12346 & ~n12348 ;
  assign n12350 = ~n12327 & n12344 ;
  assign n12351 = ~n11971 & n12350 ;
  assign n12352 = n12327 & n12344 ;
  assign n12353 = n11971 & n12352 ;
  assign n12354 = ~n12351 & ~n12353 ;
  assign n12355 = n12349 & n12354 ;
  assign n12356 = ~n11968 & n12355 ;
  assign n12357 = ~n11827 & ~n12355 ;
  assign n12358 = ~n11967 & n12357 ;
  assign n12359 = n646 & n8175 ;
  assign n12360 = ~n8172 & n12359 ;
  assign n12361 = n646 & ~n8175 ;
  assign n12362 = ~n7756 & n12361 ;
  assign n12363 = ~n8171 & n12362 ;
  assign n12364 = \b[36]  & n796 ;
  assign n12365 = n793 & n12364 ;
  assign n12366 = ~\a[9]  & \b[37]  ;
  assign n12367 = n638 & n12366 ;
  assign n12368 = ~n12365 & ~n12367 ;
  assign n12369 = \b[38]  & n644 ;
  assign n12370 = \a[9]  & \b[37]  ;
  assign n12371 = n635 & n12370 ;
  assign n12372 = \a[11]  & ~n12371 ;
  assign n12373 = ~n12369 & n12372 ;
  assign n12374 = n12368 & n12373 ;
  assign n12375 = ~n12363 & n12374 ;
  assign n12376 = ~n12360 & n12375 ;
  assign n12377 = ~n12369 & ~n12371 ;
  assign n12378 = n12368 & n12377 ;
  assign n12379 = ~n12363 & n12378 ;
  assign n12380 = ~n12360 & n12379 ;
  assign n12381 = ~\a[11]  & ~n12380 ;
  assign n12382 = ~n12376 & ~n12381 ;
  assign n12383 = ~n12358 & ~n12382 ;
  assign n12384 = ~n12356 & n12383 ;
  assign n12385 = ~n12355 & n12382 ;
  assign n12386 = n11968 & n12385 ;
  assign n12387 = n12355 & n12382 ;
  assign n12388 = ~n11968 & n12387 ;
  assign n12389 = ~n12386 & ~n12388 ;
  assign n12390 = ~n12384 & n12389 ;
  assign n12391 = n430 & ~n9482 ;
  assign n12392 = ~n9480 & n12391 ;
  assign n12393 = \b[39]  & n486 ;
  assign n12394 = n483 & n12393 ;
  assign n12395 = \b[41]  & n428 ;
  assign n12396 = \a[6]  & \b[40]  ;
  assign n12397 = n419 & n12396 ;
  assign n12398 = ~\a[6]  & \b[40]  ;
  assign n12399 = n422 & n12398 ;
  assign n12400 = ~n12397 & ~n12399 ;
  assign n12401 = ~n12395 & n12400 ;
  assign n12402 = ~n12394 & n12401 ;
  assign n12403 = ~n12392 & n12402 ;
  assign n12404 = ~\a[8]  & ~n12403 ;
  assign n12405 = \a[8]  & n12402 ;
  assign n12406 = ~n12392 & n12405 ;
  assign n12407 = ~n12404 & ~n12406 ;
  assign n12408 = ~n12390 & ~n12407 ;
  assign n12409 = n11966 & n12408 ;
  assign n12410 = n12390 & ~n12407 ;
  assign n12411 = ~n11966 & n12410 ;
  assign n12412 = ~n12409 & ~n12411 ;
  assign n12413 = ~n12390 & n12407 ;
  assign n12414 = ~n11966 & n12413 ;
  assign n12415 = n12390 & n12407 ;
  assign n12416 = n11966 & n12415 ;
  assign n12417 = ~n12414 & ~n12416 ;
  assign n12418 = n12412 & n12417 ;
  assign n12419 = n11963 & ~n12418 ;
  assign n12420 = n11944 & n12419 ;
  assign n12421 = n11963 & n12418 ;
  assign n12422 = ~n11944 & n12421 ;
  assign n12423 = ~n12420 & ~n12422 ;
  assign n12424 = ~n11963 & ~n12418 ;
  assign n12425 = ~n11944 & n12424 ;
  assign n12426 = ~n11963 & n12418 ;
  assign n12427 = n11944 & n12426 ;
  assign n12428 = ~n12425 & ~n12427 ;
  assign n12429 = n12423 & n12428 ;
  assign n12430 = ~n11392 & n11906 ;
  assign n12431 = ~n11902 & n12430 ;
  assign n12432 = ~n11905 & ~n12431 ;
  assign n12433 = ~\b[46]  & ~\b[47]  ;
  assign n12434 = \b[46]  & \b[47]  ;
  assign n12435 = ~n12433 & ~n12434 ;
  assign n12436 = ~n12432 & n12435 ;
  assign n12437 = ~n11905 & ~n12435 ;
  assign n12438 = ~n12431 & n12437 ;
  assign n12439 = n134 & ~n12438 ;
  assign n12440 = ~n12436 & n12439 ;
  assign n12441 = \a[0]  & \b[47]  ;
  assign n12442 = n133 & n12441 ;
  assign n12443 = \b[46]  & n141 ;
  assign n12444 = ~\a[1]  & \b[45]  ;
  assign n12445 = n10416 & n12444 ;
  assign n12446 = ~n12443 & ~n12445 ;
  assign n12447 = ~n12442 & n12446 ;
  assign n12448 = ~n12440 & n12447 ;
  assign n12449 = ~\a[2]  & ~n12448 ;
  assign n12450 = \a[2]  & n12447 ;
  assign n12451 = ~n12440 & n12450 ;
  assign n12452 = ~n12449 & ~n12451 ;
  assign n12453 = ~n12429 & ~n12452 ;
  assign n12454 = n11943 & n12453 ;
  assign n12455 = n12429 & ~n12452 ;
  assign n12456 = ~n11943 & n12455 ;
  assign n12457 = ~n12454 & ~n12456 ;
  assign n12458 = ~n12429 & n12452 ;
  assign n12459 = ~n11943 & n12458 ;
  assign n12460 = n12429 & n12452 ;
  assign n12461 = n11943 & n12460 ;
  assign n12462 = ~n12459 & ~n12461 ;
  assign n12463 = n12457 & n12462 ;
  assign n12464 = ~n11940 & n12463 ;
  assign n12465 = n11930 & ~n12463 ;
  assign n12466 = ~n11937 & n12465 ;
  assign n12467 = ~n12464 & ~n12466 ;
  assign n12468 = n11930 & n12457 ;
  assign n12469 = ~n11937 & n12468 ;
  assign n12470 = n12462 & ~n12469 ;
  assign n12471 = n11943 & n12429 ;
  assign n12472 = n12428 & ~n12471 ;
  assign n12473 = ~n11905 & ~n12434 ;
  assign n12474 = ~n12431 & n12473 ;
  assign n12475 = ~n12433 & ~n12474 ;
  assign n12476 = ~\b[47]  & ~\b[48]  ;
  assign n12477 = \b[47]  & \b[48]  ;
  assign n12478 = ~n12476 & ~n12477 ;
  assign n12479 = n134 & n12478 ;
  assign n12480 = ~n12475 & n12479 ;
  assign n12481 = n134 & ~n12478 ;
  assign n12482 = ~n12433 & n12481 ;
  assign n12483 = ~n12474 & n12482 ;
  assign n12484 = \a[0]  & \b[48]  ;
  assign n12485 = n133 & n12484 ;
  assign n12486 = \b[47]  & n141 ;
  assign n12487 = ~\a[1]  & \b[46]  ;
  assign n12488 = n10416 & n12487 ;
  assign n12489 = ~n12486 & ~n12488 ;
  assign n12490 = ~n12485 & n12489 ;
  assign n12491 = \a[2]  & n12490 ;
  assign n12492 = ~n12483 & n12491 ;
  assign n12493 = ~n12480 & n12492 ;
  assign n12494 = ~n12483 & n12490 ;
  assign n12495 = ~n12480 & n12494 ;
  assign n12496 = ~\a[2]  & ~n12495 ;
  assign n12497 = ~n12493 & ~n12496 ;
  assign n12498 = n252 & ~n11397 ;
  assign n12499 = ~n11395 & n12498 ;
  assign n12500 = \b[45]  & n250 ;
  assign n12501 = \a[3]  & \b[44]  ;
  assign n12502 = n241 & n12501 ;
  assign n12503 = ~n12500 & ~n12502 ;
  assign n12504 = \b[43]  & n303 ;
  assign n12505 = n300 & n12504 ;
  assign n12506 = ~\a[3]  & \b[44]  ;
  assign n12507 = n244 & n12506 ;
  assign n12508 = ~n12505 & ~n12507 ;
  assign n12509 = n12503 & n12508 ;
  assign n12510 = ~n12499 & n12509 ;
  assign n12511 = ~\a[5]  & ~n12510 ;
  assign n12512 = \a[5]  & n12509 ;
  assign n12513 = ~n12499 & n12512 ;
  assign n12514 = ~n12511 & ~n12513 ;
  assign n12515 = ~n11888 & n12412 ;
  assign n12516 = ~n11895 & n12515 ;
  assign n12517 = n12417 & ~n12516 ;
  assign n12518 = n11966 & n12390 ;
  assign n12519 = ~n12384 & ~n12518 ;
  assign n12520 = ~n11827 & n12349 ;
  assign n12521 = ~n11967 & n12520 ;
  assign n12522 = n12354 & ~n12521 ;
  assign n12523 = n11971 & n12327 ;
  assign n12524 = ~n12326 & ~n12523 ;
  assign n12525 = n11783 & n12315 ;
  assign n12526 = ~n11972 & n12525 ;
  assign n12527 = n12310 & ~n12526 ;
  assign n12528 = n12000 & n12305 ;
  assign n12529 = n12304 & ~n12528 ;
  assign n12530 = n1965 & n5105 ;
  assign n12531 = ~n5102 & n12530 ;
  assign n12532 = n1965 & ~n5105 ;
  assign n12533 = ~n4497 & n12532 ;
  assign n12534 = ~n5101 & n12533 ;
  assign n12535 = \b[28]  & n2218 ;
  assign n12536 = n2216 & n12535 ;
  assign n12537 = ~\a[18]  & \b[29]  ;
  assign n12538 = n1957 & n12537 ;
  assign n12539 = ~n12536 & ~n12538 ;
  assign n12540 = \b[30]  & n1963 ;
  assign n12541 = \a[18]  & \b[29]  ;
  assign n12542 = n2210 & n12541 ;
  assign n12543 = \a[20]  & ~n12542 ;
  assign n12544 = ~n12540 & n12543 ;
  assign n12545 = n12539 & n12544 ;
  assign n12546 = ~n12534 & n12545 ;
  assign n12547 = ~n12531 & n12546 ;
  assign n12548 = ~n12540 & ~n12542 ;
  assign n12549 = n12539 & n12548 ;
  assign n12550 = ~n12534 & n12549 ;
  assign n12551 = ~n12531 & n12550 ;
  assign n12552 = ~\a[20]  & ~n12551 ;
  assign n12553 = ~n12547 & ~n12552 ;
  assign n12554 = ~n11749 & n12288 ;
  assign n12555 = ~n11757 & n12554 ;
  assign n12556 = n12293 & ~n12555 ;
  assign n12557 = n12045 & n12259 ;
  assign n12558 = ~n12253 & ~n12557 ;
  assign n12559 = ~n11679 & n12218 ;
  assign n12560 = ~n12046 & n12559 ;
  assign n12561 = n12223 & ~n12560 ;
  assign n12562 = n12050 & n12213 ;
  assign n12563 = n12207 & ~n12562 ;
  assign n12564 = n11634 & ~n12180 ;
  assign n12565 = ~n12075 & n12564 ;
  assign n12566 = ~n12179 & ~n12565 ;
  assign n12567 = ~n1233 & n6309 ;
  assign n12568 = ~n1231 & n12567 ;
  assign n12569 = \b[13]  & n6778 ;
  assign n12570 = n6775 & n12569 ;
  assign n12571 = \b[15]  & n6307 ;
  assign n12572 = \a[33]  & \b[14]  ;
  assign n12573 = n6298 & n12572 ;
  assign n12574 = ~\a[33]  & \b[14]  ;
  assign n12575 = n6301 & n12574 ;
  assign n12576 = ~n12573 & ~n12575 ;
  assign n12577 = ~n12571 & n12576 ;
  assign n12578 = ~n12570 & n12577 ;
  assign n12579 = ~\a[35]  & n12578 ;
  assign n12580 = ~n12568 & n12579 ;
  assign n12581 = ~n12568 & n12578 ;
  assign n12582 = \a[35]  & ~n12581 ;
  assign n12583 = ~n12580 & ~n12582 ;
  assign n12584 = ~n12173 & ~n12176 ;
  assign n12585 = ~n11581 & ~n12167 ;
  assign n12586 = ~n11583 & n12585 ;
  assign n12587 = ~n12168 & ~n12586 ;
  assign n12588 = n177 & n11572 ;
  assign n12589 = \b[3]  & n11570 ;
  assign n12590 = \a[45]  & \b[2]  ;
  assign n12591 = n11561 & n12590 ;
  assign n12592 = ~\a[44]  & \b[2]  ;
  assign n12593 = n12158 & n12592 ;
  assign n12594 = ~n12591 & ~n12593 ;
  assign n12595 = ~n12589 & n12594 ;
  assign n12596 = ~n12588 & n12595 ;
  assign n12597 = \b[1]  & n12159 ;
  assign n12598 = n12156 & n12597 ;
  assign n12599 = ~\a[47]  & ~n12598 ;
  assign n12600 = n12596 & n12599 ;
  assign n12601 = n12596 & ~n12598 ;
  assign n12602 = \a[47]  & ~n12601 ;
  assign n12603 = ~n12600 & ~n12602 ;
  assign n12604 = \a[47]  & ~\a[48]  ;
  assign n12605 = ~\a[47]  & \a[48]  ;
  assign n12606 = ~n12604 & ~n12605 ;
  assign n12607 = \b[0]  & ~n12606 ;
  assign n12608 = n12146 & n12163 ;
  assign n12609 = n12607 & n12608 ;
  assign n12610 = ~n12607 & ~n12608 ;
  assign n12611 = ~n12609 & ~n12610 ;
  assign n12612 = n12603 & n12611 ;
  assign n12613 = ~n12603 & ~n12611 ;
  assign n12614 = ~n12612 & ~n12613 ;
  assign n12615 = ~n323 & ~n9646 ;
  assign n12616 = ~n10079 & n12615 ;
  assign n12617 = n320 & n12616 ;
  assign n12618 = n323 & ~n9646 ;
  assign n12619 = ~n10079 & n12618 ;
  assign n12620 = ~n320 & n12619 ;
  assign n12621 = ~n12617 & ~n12620 ;
  assign n12622 = \b[4]  & n10681 ;
  assign n12623 = n10678 & n12622 ;
  assign n12624 = \b[6]  & n10080 ;
  assign n12625 = \a[41]  & \b[5]  ;
  assign n12626 = n10679 & n12625 ;
  assign n12627 = ~\a[42]  & \b[5]  ;
  assign n12628 = n10074 & n12627 ;
  assign n12629 = ~n12626 & ~n12628 ;
  assign n12630 = ~n12624 & n12629 ;
  assign n12631 = ~n12623 & n12630 ;
  assign n12632 = n12621 & n12631 ;
  assign n12633 = ~\a[44]  & ~n12632 ;
  assign n12634 = \a[44]  & n12631 ;
  assign n12635 = n12621 & n12634 ;
  assign n12636 = ~n12633 & ~n12635 ;
  assign n12637 = n12614 & ~n12636 ;
  assign n12638 = ~n12614 & n12636 ;
  assign n12639 = ~n12637 & ~n12638 ;
  assign n12640 = ~n586 & n8759 ;
  assign n12641 = ~n504 & n8759 ;
  assign n12642 = ~n508 & n12641 ;
  assign n12643 = ~n12640 & ~n12642 ;
  assign n12644 = ~n589 & ~n12643 ;
  assign n12645 = \b[7]  & n9301 ;
  assign n12646 = n9298 & n12645 ;
  assign n12647 = ~\a[39]  & \b[8]  ;
  assign n12648 = n8751 & n12647 ;
  assign n12649 = ~n12646 & ~n12648 ;
  assign n12650 = \b[9]  & n8757 ;
  assign n12651 = \a[39]  & \b[8]  ;
  assign n12652 = n8748 & n12651 ;
  assign n12653 = \a[41]  & ~n12652 ;
  assign n12654 = ~n12650 & n12653 ;
  assign n12655 = n12649 & n12654 ;
  assign n12656 = ~n12644 & n12655 ;
  assign n12657 = ~n12650 & ~n12652 ;
  assign n12658 = n12649 & n12657 ;
  assign n12659 = ~\a[41]  & ~n12658 ;
  assign n12660 = ~\a[41]  & ~n589 ;
  assign n12661 = ~n12643 & n12660 ;
  assign n12662 = ~n12659 & ~n12661 ;
  assign n12663 = ~n12656 & n12662 ;
  assign n12664 = ~n12639 & n12663 ;
  assign n12665 = ~n12587 & n12664 ;
  assign n12666 = n12639 & n12663 ;
  assign n12667 = n12587 & n12666 ;
  assign n12668 = ~n12665 & ~n12667 ;
  assign n12669 = ~n12639 & ~n12663 ;
  assign n12670 = n12587 & n12669 ;
  assign n12671 = n12639 & ~n12663 ;
  assign n12672 = ~n12587 & n12671 ;
  assign n12673 = ~n12670 & ~n12672 ;
  assign n12674 = n12668 & n12673 ;
  assign n12675 = ~n12584 & n12674 ;
  assign n12676 = ~n909 & ~n7098 ;
  assign n12677 = ~n7531 & n12676 ;
  assign n12678 = n906 & n12677 ;
  assign n12679 = n909 & ~n7098 ;
  assign n12680 = ~n7531 & n12679 ;
  assign n12681 = ~n906 & n12680 ;
  assign n12682 = ~n12678 & ~n12681 ;
  assign n12683 = \b[10]  & n7973 ;
  assign n12684 = n7970 & n12683 ;
  assign n12685 = \b[12]  & n7532 ;
  assign n12686 = \a[36]  & \b[11]  ;
  assign n12687 = n7523 & n12686 ;
  assign n12688 = ~\a[36]  & \b[11]  ;
  assign n12689 = n7526 & n12688 ;
  assign n12690 = ~n12687 & ~n12689 ;
  assign n12691 = ~n12685 & n12690 ;
  assign n12692 = ~n12684 & n12691 ;
  assign n12693 = n12682 & n12692 ;
  assign n12694 = ~\a[38]  & ~n12693 ;
  assign n12695 = \a[38]  & n12692 ;
  assign n12696 = n12682 & n12695 ;
  assign n12697 = ~n12694 & ~n12696 ;
  assign n12698 = ~n12173 & ~n12674 ;
  assign n12699 = ~n12176 & n12698 ;
  assign n12700 = ~n12697 & ~n12699 ;
  assign n12701 = ~n12675 & n12700 ;
  assign n12702 = ~n12674 & n12697 ;
  assign n12703 = n12584 & n12702 ;
  assign n12704 = n12674 & n12697 ;
  assign n12705 = ~n12584 & n12704 ;
  assign n12706 = ~n12703 & ~n12705 ;
  assign n12707 = ~n12701 & n12706 ;
  assign n12708 = n12583 & ~n12707 ;
  assign n12709 = n12566 & n12708 ;
  assign n12710 = n12583 & n12707 ;
  assign n12711 = ~n12566 & n12710 ;
  assign n12712 = ~n12709 & ~n12711 ;
  assign n12713 = ~n12583 & ~n12707 ;
  assign n12714 = ~n12566 & n12713 ;
  assign n12715 = ~n12583 & n12707 ;
  assign n12716 = n12566 & n12715 ;
  assign n12717 = ~n12714 & ~n12716 ;
  assign n12718 = n12712 & n12717 ;
  assign n12719 = ~n12563 & n12718 ;
  assign n12720 = n12207 & ~n12718 ;
  assign n12721 = ~n12562 & n12720 ;
  assign n12722 = n1875 & n5211 ;
  assign n12723 = ~n1872 & n12722 ;
  assign n12724 = n5000 & n5211 ;
  assign n12725 = ~n1871 & n12724 ;
  assign n12726 = \b[16]  & n5595 ;
  assign n12727 = n5592 & n12726 ;
  assign n12728 = ~\a[30]  & \b[17]  ;
  assign n12729 = n5203 & n12728 ;
  assign n12730 = ~n12727 & ~n12729 ;
  assign n12731 = \b[18]  & n5209 ;
  assign n12732 = \a[30]  & \b[17]  ;
  assign n12733 = n5200 & n12732 ;
  assign n12734 = \a[32]  & ~n12733 ;
  assign n12735 = ~n12731 & n12734 ;
  assign n12736 = n12730 & n12735 ;
  assign n12737 = ~n12725 & n12736 ;
  assign n12738 = ~n12723 & n12737 ;
  assign n12739 = ~n12731 & ~n12733 ;
  assign n12740 = n12730 & n12739 ;
  assign n12741 = ~n12725 & n12740 ;
  assign n12742 = ~n12723 & n12741 ;
  assign n12743 = ~\a[32]  & ~n12742 ;
  assign n12744 = ~n12738 & ~n12743 ;
  assign n12745 = ~n12721 & ~n12744 ;
  assign n12746 = ~n12719 & n12745 ;
  assign n12747 = ~n12718 & n12744 ;
  assign n12748 = n12563 & n12747 ;
  assign n12749 = n12718 & n12744 ;
  assign n12750 = ~n12563 & n12749 ;
  assign n12751 = ~n12748 & ~n12750 ;
  assign n12752 = ~n12746 & n12751 ;
  assign n12753 = ~n2523 & n4249 ;
  assign n12754 = ~n2521 & n12753 ;
  assign n12755 = \b[21]  & n4247 ;
  assign n12756 = \a[27]  & \b[20]  ;
  assign n12757 = n4238 & n12756 ;
  assign n12758 = ~n12755 & ~n12757 ;
  assign n12759 = \b[19]  & n4647 ;
  assign n12760 = n4644 & n12759 ;
  assign n12761 = ~\a[27]  & \b[20]  ;
  assign n12762 = n4241 & n12761 ;
  assign n12763 = ~n12760 & ~n12762 ;
  assign n12764 = n12758 & n12763 ;
  assign n12765 = ~n12754 & n12764 ;
  assign n12766 = ~\a[29]  & ~n12765 ;
  assign n12767 = \a[29]  & n12764 ;
  assign n12768 = ~n12754 & n12767 ;
  assign n12769 = ~n12766 & ~n12768 ;
  assign n12770 = ~n12752 & ~n12769 ;
  assign n12771 = n12561 & n12770 ;
  assign n12772 = n12752 & ~n12769 ;
  assign n12773 = ~n12561 & n12772 ;
  assign n12774 = ~n12771 & ~n12773 ;
  assign n12775 = ~n12752 & n12769 ;
  assign n12776 = ~n12561 & n12775 ;
  assign n12777 = n12752 & n12769 ;
  assign n12778 = n12561 & n12777 ;
  assign n12779 = ~n12776 & ~n12778 ;
  assign n12780 = n12774 & n12779 ;
  assign n12781 = ~n3154 & ~n3283 ;
  assign n12782 = ~n3399 & n12781 ;
  assign n12783 = n3280 & n12782 ;
  assign n12784 = ~n3154 & n3283 ;
  assign n12785 = ~n3399 & n12784 ;
  assign n12786 = ~n3280 & n12785 ;
  assign n12787 = ~n12783 & ~n12786 ;
  assign n12788 = \b[22]  & n3733 ;
  assign n12789 = n3730 & n12788 ;
  assign n12790 = ~\a[24]  & \b[23]  ;
  assign n12791 = n3394 & n12790 ;
  assign n12792 = ~n12789 & ~n12791 ;
  assign n12793 = \b[24]  & n3400 ;
  assign n12794 = \a[24]  & \b[23]  ;
  assign n12795 = n3391 & n12794 ;
  assign n12796 = \a[26]  & ~n12795 ;
  assign n12797 = ~n12793 & n12796 ;
  assign n12798 = n12792 & n12797 ;
  assign n12799 = n12787 & n12798 ;
  assign n12800 = ~n12793 & ~n12795 ;
  assign n12801 = n12792 & n12800 ;
  assign n12802 = n12787 & n12801 ;
  assign n12803 = ~\a[26]  & ~n12802 ;
  assign n12804 = ~n12799 & ~n12803 ;
  assign n12805 = ~n12780 & n12804 ;
  assign n12806 = n12558 & n12805 ;
  assign n12807 = n12780 & n12804 ;
  assign n12808 = ~n12558 & n12807 ;
  assign n12809 = ~n12806 & ~n12808 ;
  assign n12810 = ~n12558 & n12780 ;
  assign n12811 = ~n12253 & ~n12780 ;
  assign n12812 = ~n12557 & n12811 ;
  assign n12813 = ~n12804 & ~n12812 ;
  assign n12814 = ~n12810 & n12813 ;
  assign n12815 = n12809 & ~n12814 ;
  assign n12816 = n12556 & n12815 ;
  assign n12817 = ~n12556 & ~n12815 ;
  assign n12818 = ~n12816 & ~n12817 ;
  assign n12819 = ~n2413 & ~n2619 ;
  assign n12820 = ~n4148 & n12819 ;
  assign n12821 = ~n4146 & n12820 ;
  assign n12822 = \b[25]  & n2912 ;
  assign n12823 = n2909 & n12822 ;
  assign n12824 = ~\a[21]  & \b[26]  ;
  assign n12825 = n2614 & n12824 ;
  assign n12826 = ~n12823 & ~n12825 ;
  assign n12827 = \b[27]  & n2620 ;
  assign n12828 = \a[21]  & \b[26]  ;
  assign n12829 = n2611 & n12828 ;
  assign n12830 = \a[23]  & ~n12829 ;
  assign n12831 = ~n12827 & n12830 ;
  assign n12832 = n12826 & n12831 ;
  assign n12833 = ~n12821 & n12832 ;
  assign n12834 = ~n12827 & ~n12829 ;
  assign n12835 = n12826 & n12834 ;
  assign n12836 = ~n12821 & n12835 ;
  assign n12837 = ~\a[23]  & ~n12836 ;
  assign n12838 = ~n12833 & ~n12837 ;
  assign n12839 = n12818 & ~n12838 ;
  assign n12840 = ~n12818 & n12838 ;
  assign n12841 = ~n12839 & ~n12840 ;
  assign n12842 = ~n12553 & ~n12841 ;
  assign n12843 = ~n12529 & n12842 ;
  assign n12844 = ~n12553 & n12841 ;
  assign n12845 = n12529 & n12844 ;
  assign n12846 = ~n12843 & ~n12845 ;
  assign n12847 = n12553 & ~n12841 ;
  assign n12848 = n12529 & n12847 ;
  assign n12849 = n12553 & n12841 ;
  assign n12850 = ~n12529 & n12849 ;
  assign n12851 = ~n12848 & ~n12850 ;
  assign n12852 = n12846 & n12851 ;
  assign n12853 = n1467 & ~n5855 ;
  assign n12854 = ~n5853 & n12853 ;
  assign n12855 = \b[33]  & n1465 ;
  assign n12856 = \a[15]  & \b[32]  ;
  assign n12857 = n1456 & n12856 ;
  assign n12858 = ~n12855 & ~n12857 ;
  assign n12859 = \b[31]  & n1652 ;
  assign n12860 = n1649 & n12859 ;
  assign n12861 = ~\a[15]  & \b[32]  ;
  assign n12862 = n1459 & n12861 ;
  assign n12863 = ~n12860 & ~n12862 ;
  assign n12864 = n12858 & n12863 ;
  assign n12865 = ~n12854 & n12864 ;
  assign n12866 = ~\a[17]  & ~n12865 ;
  assign n12867 = \a[17]  & n12864 ;
  assign n12868 = ~n12854 & n12867 ;
  assign n12869 = ~n12866 & ~n12868 ;
  assign n12870 = ~n12852 & ~n12869 ;
  assign n12871 = n12527 & n12870 ;
  assign n12872 = n12852 & ~n12869 ;
  assign n12873 = ~n12527 & n12872 ;
  assign n12874 = ~n12871 & ~n12873 ;
  assign n12875 = ~n12852 & n12869 ;
  assign n12876 = ~n12527 & n12875 ;
  assign n12877 = n12852 & n12869 ;
  assign n12878 = n12527 & n12877 ;
  assign n12879 = ~n12876 & ~n12878 ;
  assign n12880 = n12874 & n12879 ;
  assign n12881 = ~n12524 & n12880 ;
  assign n12882 = n999 & n7337 ;
  assign n12883 = ~n7334 & n12882 ;
  assign n12884 = n999 & ~n7337 ;
  assign n12885 = ~n6605 & n12884 ;
  assign n12886 = ~n7333 & n12885 ;
  assign n12887 = \b[34]  & n1182 ;
  assign n12888 = n1179 & n12887 ;
  assign n12889 = \b[36]  & n997 ;
  assign n12890 = \a[11]  & \b[35]  ;
  assign n12891 = n1180 & n12890 ;
  assign n12892 = ~\a[12]  & \b[35]  ;
  assign n12893 = n7674 & n12892 ;
  assign n12894 = ~n12891 & ~n12893 ;
  assign n12895 = ~n12889 & n12894 ;
  assign n12896 = ~n12888 & n12895 ;
  assign n12897 = ~n12886 & n12896 ;
  assign n12898 = ~n12883 & n12897 ;
  assign n12899 = ~\a[14]  & ~n12898 ;
  assign n12900 = \a[14]  & n12896 ;
  assign n12901 = ~n12886 & n12900 ;
  assign n12902 = ~n12883 & n12901 ;
  assign n12903 = ~n12899 & ~n12902 ;
  assign n12904 = ~n12326 & ~n12880 ;
  assign n12905 = ~n12523 & n12904 ;
  assign n12906 = ~n12903 & ~n12905 ;
  assign n12907 = ~n12881 & n12906 ;
  assign n12908 = ~n12880 & n12903 ;
  assign n12909 = n12524 & n12908 ;
  assign n12910 = n12880 & n12903 ;
  assign n12911 = ~n12524 & n12910 ;
  assign n12912 = ~n12909 & ~n12911 ;
  assign n12913 = ~n12907 & n12912 ;
  assign n12914 = n646 & ~n8602 ;
  assign n12915 = ~n8600 & n12914 ;
  assign n12916 = \b[39]  & n644 ;
  assign n12917 = \a[9]  & \b[38]  ;
  assign n12918 = n635 & n12917 ;
  assign n12919 = ~n12916 & ~n12918 ;
  assign n12920 = \b[37]  & n796 ;
  assign n12921 = n793 & n12920 ;
  assign n12922 = ~\a[9]  & \b[38]  ;
  assign n12923 = n638 & n12922 ;
  assign n12924 = ~n12921 & ~n12923 ;
  assign n12925 = n12919 & n12924 ;
  assign n12926 = ~n12915 & n12925 ;
  assign n12927 = ~\a[11]  & ~n12926 ;
  assign n12928 = \a[11]  & n12925 ;
  assign n12929 = ~n12915 & n12928 ;
  assign n12930 = ~n12927 & ~n12929 ;
  assign n12931 = ~n12913 & ~n12930 ;
  assign n12932 = n12522 & n12931 ;
  assign n12933 = n12913 & ~n12930 ;
  assign n12934 = ~n12522 & n12933 ;
  assign n12935 = ~n12932 & ~n12934 ;
  assign n12936 = ~n12913 & n12930 ;
  assign n12937 = ~n12522 & n12936 ;
  assign n12938 = n12913 & n12930 ;
  assign n12939 = n12522 & n12938 ;
  assign n12940 = ~n12937 & ~n12939 ;
  assign n12941 = n12935 & n12940 ;
  assign n12942 = ~n12519 & n12941 ;
  assign n12943 = ~n12384 & ~n12941 ;
  assign n12944 = ~n12518 & n12943 ;
  assign n12945 = n430 & n9930 ;
  assign n12946 = ~n9927 & n12945 ;
  assign n12947 = n430 & ~n9930 ;
  assign n12948 = ~n9477 & n12947 ;
  assign n12949 = ~n9926 & n12948 ;
  assign n12950 = \b[40]  & n486 ;
  assign n12951 = n483 & n12950 ;
  assign n12952 = \b[42]  & n428 ;
  assign n12953 = \a[6]  & \b[41]  ;
  assign n12954 = n419 & n12953 ;
  assign n12955 = ~\a[6]  & \b[41]  ;
  assign n12956 = n422 & n12955 ;
  assign n12957 = ~n12954 & ~n12956 ;
  assign n12958 = ~n12952 & n12957 ;
  assign n12959 = ~n12951 & n12958 ;
  assign n12960 = ~n12949 & n12959 ;
  assign n12961 = ~n12946 & n12960 ;
  assign n12962 = ~\a[8]  & ~n12961 ;
  assign n12963 = \a[8]  & n12959 ;
  assign n12964 = ~n12949 & n12963 ;
  assign n12965 = ~n12946 & n12964 ;
  assign n12966 = ~n12962 & ~n12965 ;
  assign n12967 = ~n12944 & ~n12966 ;
  assign n12968 = ~n12942 & n12967 ;
  assign n12969 = ~n12941 & n12966 ;
  assign n12970 = n12519 & n12969 ;
  assign n12971 = n12941 & n12966 ;
  assign n12972 = ~n12519 & n12971 ;
  assign n12973 = ~n12970 & ~n12972 ;
  assign n12974 = ~n12968 & n12973 ;
  assign n12975 = n12517 & n12974 ;
  assign n12976 = ~n12517 & ~n12974 ;
  assign n12977 = ~n12975 & ~n12976 ;
  assign n12978 = ~n12514 & n12977 ;
  assign n12979 = n12514 & ~n12977 ;
  assign n12980 = ~n12978 & ~n12979 ;
  assign n12981 = n12497 & ~n12980 ;
  assign n12982 = n12472 & n12981 ;
  assign n12983 = n12497 & n12980 ;
  assign n12984 = ~n12472 & n12983 ;
  assign n12985 = ~n12982 & ~n12984 ;
  assign n12986 = ~n12497 & ~n12980 ;
  assign n12987 = ~n12472 & n12986 ;
  assign n12988 = ~n12497 & n12980 ;
  assign n12989 = n12472 & n12988 ;
  assign n12990 = ~n12987 & ~n12989 ;
  assign n12991 = n12985 & n12990 ;
  assign n12992 = n12470 & n12991 ;
  assign n12993 = ~n12470 & ~n12991 ;
  assign n12994 = ~n12992 & ~n12993 ;
  assign n12995 = n12990 & ~n12992 ;
  assign n12996 = n12428 & ~n12978 ;
  assign n12997 = ~n12471 & n12996 ;
  assign n12998 = ~n12979 & ~n12997 ;
  assign n12999 = ~n12968 & ~n12975 ;
  assign n13000 = ~n12384 & n12935 ;
  assign n13001 = ~n12518 & n13000 ;
  assign n13002 = n12940 & ~n13001 ;
  assign n13003 = n12522 & n12913 ;
  assign n13004 = ~n12907 & ~n13003 ;
  assign n13005 = ~n12326 & n12874 ;
  assign n13006 = ~n12523 & n13005 ;
  assign n13007 = n12879 & ~n13006 ;
  assign n13008 = n12527 & n12852 ;
  assign n13009 = n12846 & ~n13008 ;
  assign n13010 = n12304 & ~n12839 ;
  assign n13011 = ~n12528 & n13010 ;
  assign n13012 = ~n12840 & ~n13011 ;
  assign n13013 = n1965 & ~n5462 ;
  assign n13014 = ~n5460 & n13013 ;
  assign n13015 = \b[31]  & n1963 ;
  assign n13016 = \a[18]  & \b[30]  ;
  assign n13017 = n2210 & n13016 ;
  assign n13018 = ~n13015 & ~n13017 ;
  assign n13019 = \b[29]  & n2218 ;
  assign n13020 = n2216 & n13019 ;
  assign n13021 = ~\a[18]  & \b[30]  ;
  assign n13022 = n1957 & n13021 ;
  assign n13023 = ~n13020 & ~n13022 ;
  assign n13024 = n13018 & n13023 ;
  assign n13025 = ~n13014 & n13024 ;
  assign n13026 = ~\a[20]  & ~n13025 ;
  assign n13027 = \a[20]  & n13024 ;
  assign n13028 = ~n13014 & n13027 ;
  assign n13029 = ~n13026 & ~n13028 ;
  assign n13030 = ~n12814 & ~n12816 ;
  assign n13031 = n2622 & n4456 ;
  assign n13032 = ~n4453 & n13031 ;
  assign n13033 = n2622 & ~n4456 ;
  assign n13034 = ~n4143 & n13033 ;
  assign n13035 = ~n4452 & n13034 ;
  assign n13036 = \b[26]  & n2912 ;
  assign n13037 = n2909 & n13036 ;
  assign n13038 = ~\a[21]  & \b[27]  ;
  assign n13039 = n2614 & n13038 ;
  assign n13040 = ~n13037 & ~n13039 ;
  assign n13041 = \b[28]  & n2620 ;
  assign n13042 = \a[21]  & \b[27]  ;
  assign n13043 = n2611 & n13042 ;
  assign n13044 = \a[23]  & ~n13043 ;
  assign n13045 = ~n13041 & n13044 ;
  assign n13046 = n13040 & n13045 ;
  assign n13047 = ~n13035 & n13046 ;
  assign n13048 = ~n13032 & n13047 ;
  assign n13049 = ~n13041 & ~n13043 ;
  assign n13050 = n13040 & n13049 ;
  assign n13051 = ~n13035 & n13050 ;
  assign n13052 = ~n13032 & n13051 ;
  assign n13053 = ~\a[23]  & ~n13052 ;
  assign n13054 = ~n13048 & ~n13053 ;
  assign n13055 = ~n12253 & n12774 ;
  assign n13056 = ~n12557 & n13055 ;
  assign n13057 = n12779 & ~n13056 ;
  assign n13058 = n12561 & n12752 ;
  assign n13059 = ~n12746 & ~n13058 ;
  assign n13060 = n12207 & n12712 ;
  assign n13061 = n12717 & ~n13060 ;
  assign n13062 = n12213 & n12717 ;
  assign n13063 = n12050 & n13062 ;
  assign n13064 = ~n13061 & ~n13063 ;
  assign n13065 = n12566 & n12707 ;
  assign n13066 = ~n12701 & ~n13065 ;
  assign n13067 = ~n12173 & n12673 ;
  assign n13068 = ~n12176 & n13067 ;
  assign n13069 = n12668 & ~n13068 ;
  assign n13070 = ~n948 & n7534 ;
  assign n13071 = ~n908 & n7534 ;
  assign n13072 = ~n912 & n13071 ;
  assign n13073 = ~n13070 & ~n13072 ;
  assign n13074 = ~n951 & ~n13073 ;
  assign n13075 = \b[11]  & n7973 ;
  assign n13076 = n7970 & n13075 ;
  assign n13077 = \b[13]  & n7532 ;
  assign n13078 = \a[36]  & \b[12]  ;
  assign n13079 = n7523 & n13078 ;
  assign n13080 = ~\a[36]  & \b[12]  ;
  assign n13081 = n7526 & n13080 ;
  assign n13082 = ~n13079 & ~n13081 ;
  assign n13083 = ~n13077 & n13082 ;
  assign n13084 = ~n13076 & n13083 ;
  assign n13085 = ~\a[38]  & n13084 ;
  assign n13086 = ~n13074 & n13085 ;
  assign n13087 = \a[38]  & ~n13084 ;
  assign n13088 = \a[38]  & ~n951 ;
  assign n13089 = ~n13073 & n13088 ;
  assign n13090 = ~n13087 & ~n13089 ;
  assign n13091 = ~n13086 & n13090 ;
  assign n13092 = n12587 & n12639 ;
  assign n13093 = ~n12637 & ~n13092 ;
  assign n13094 = ~n12609 & ~n12612 ;
  assign n13095 = n222 & n11572 ;
  assign n13096 = \b[4]  & n11570 ;
  assign n13097 = ~\a[45]  & \b[3]  ;
  assign n13098 = n11564 & n13097 ;
  assign n13099 = \a[45]  & \b[3]  ;
  assign n13100 = n11561 & n13099 ;
  assign n13101 = ~n13098 & ~n13100 ;
  assign n13102 = ~n13096 & n13101 ;
  assign n13103 = \b[2]  & n12159 ;
  assign n13104 = n12156 & n13103 ;
  assign n13105 = \a[47]  & ~n13104 ;
  assign n13106 = n13102 & n13105 ;
  assign n13107 = ~n13095 & n13106 ;
  assign n13108 = n13102 & ~n13104 ;
  assign n13109 = ~n13095 & n13108 ;
  assign n13110 = ~\a[47]  & ~n13109 ;
  assign n13111 = ~n13107 & ~n13110 ;
  assign n13112 = \a[50]  & \b[0]  ;
  assign n13113 = ~n12606 & n13112 ;
  assign n13114 = \a[48]  & ~\a[49]  ;
  assign n13115 = n11558 & n13114 ;
  assign n13116 = ~\a[48]  & \b[0]  ;
  assign n13117 = ~\a[47]  & \a[49]  ;
  assign n13118 = n13116 & n13117 ;
  assign n13119 = ~n13115 & ~n13118 ;
  assign n13120 = \a[49]  & ~\a[50]  ;
  assign n13121 = ~\a[49]  & \a[50]  ;
  assign n13122 = ~n13120 & ~n13121 ;
  assign n13123 = ~n12606 & n13122 ;
  assign n13124 = \b[1]  & n13123 ;
  assign n13125 = ~n12606 & ~n13122 ;
  assign n13126 = ~n137 & n13125 ;
  assign n13127 = ~n13124 & ~n13126 ;
  assign n13128 = n13119 & n13127 ;
  assign n13129 = ~n13113 & ~n13128 ;
  assign n13130 = n13113 & n13119 ;
  assign n13131 = n13127 & n13130 ;
  assign n13132 = ~n13129 & ~n13131 ;
  assign n13133 = n13111 & n13132 ;
  assign n13134 = ~n13111 & ~n13132 ;
  assign n13135 = ~n13133 & ~n13134 ;
  assign n13136 = ~n13094 & n13135 ;
  assign n13137 = n13094 & ~n13135 ;
  assign n13138 = ~n13136 & ~n13137 ;
  assign n13139 = ~n383 & n10082 ;
  assign n13140 = ~n381 & n13139 ;
  assign n13141 = \b[5]  & n10681 ;
  assign n13142 = n10678 & n13141 ;
  assign n13143 = \b[7]  & n10080 ;
  assign n13144 = \a[41]  & \b[6]  ;
  assign n13145 = n10679 & n13144 ;
  assign n13146 = ~\a[42]  & \b[6]  ;
  assign n13147 = n10074 & n13146 ;
  assign n13148 = ~n13145 & ~n13147 ;
  assign n13149 = ~n13143 & n13148 ;
  assign n13150 = ~n13142 & n13149 ;
  assign n13151 = ~\a[44]  & n13150 ;
  assign n13152 = ~n13140 & n13151 ;
  assign n13153 = ~n13140 & n13150 ;
  assign n13154 = \a[44]  & ~n13153 ;
  assign n13155 = ~n13152 & ~n13154 ;
  assign n13156 = n13138 & n13155 ;
  assign n13157 = ~n13138 & ~n13155 ;
  assign n13158 = ~n13156 & ~n13157 ;
  assign n13159 = n685 & n8759 ;
  assign n13160 = ~n682 & n13159 ;
  assign n13161 = ~n685 & n8759 ;
  assign n13162 = ~n584 & n13161 ;
  assign n13163 = ~n681 & n13162 ;
  assign n13164 = \b[8]  & n9301 ;
  assign n13165 = n9298 & n13164 ;
  assign n13166 = ~\a[39]  & \b[9]  ;
  assign n13167 = n8751 & n13166 ;
  assign n13168 = ~n13165 & ~n13167 ;
  assign n13169 = \b[10]  & n8757 ;
  assign n13170 = \a[39]  & \b[9]  ;
  assign n13171 = n8748 & n13170 ;
  assign n13172 = \a[41]  & ~n13171 ;
  assign n13173 = ~n13169 & n13172 ;
  assign n13174 = n13168 & n13173 ;
  assign n13175 = ~n13163 & n13174 ;
  assign n13176 = ~n13160 & n13175 ;
  assign n13177 = ~n13169 & ~n13171 ;
  assign n13178 = n13168 & n13177 ;
  assign n13179 = ~n13163 & n13178 ;
  assign n13180 = ~n13160 & n13179 ;
  assign n13181 = ~\a[41]  & ~n13180 ;
  assign n13182 = ~n13176 & ~n13181 ;
  assign n13183 = ~n13158 & ~n13182 ;
  assign n13184 = ~n13093 & n13183 ;
  assign n13185 = n13158 & ~n13182 ;
  assign n13186 = n13093 & n13185 ;
  assign n13187 = ~n13184 & ~n13186 ;
  assign n13188 = ~n13158 & n13182 ;
  assign n13189 = n13093 & n13188 ;
  assign n13190 = n13158 & n13182 ;
  assign n13191 = ~n13093 & n13190 ;
  assign n13192 = ~n13189 & ~n13191 ;
  assign n13193 = n13187 & n13192 ;
  assign n13194 = ~n13091 & ~n13193 ;
  assign n13195 = ~n13069 & n13194 ;
  assign n13196 = ~n13091 & n13193 ;
  assign n13197 = n13069 & n13196 ;
  assign n13198 = ~n13195 & ~n13197 ;
  assign n13199 = n13091 & ~n13193 ;
  assign n13200 = n13069 & n13199 ;
  assign n13201 = n13091 & n13193 ;
  assign n13202 = ~n13069 & n13201 ;
  assign n13203 = ~n13200 & ~n13202 ;
  assign n13204 = n13198 & n13203 ;
  assign n13205 = ~n13066 & n13204 ;
  assign n13206 = ~n12701 & ~n13204 ;
  assign n13207 = ~n13065 & n13206 ;
  assign n13208 = n1512 & n6309 ;
  assign n13209 = ~n1509 & n13208 ;
  assign n13210 = n6309 & n10165 ;
  assign n13211 = ~n1508 & n13210 ;
  assign n13212 = \b[14]  & n6778 ;
  assign n13213 = n6775 & n13212 ;
  assign n13214 = ~\a[33]  & \b[15]  ;
  assign n13215 = n6301 & n13214 ;
  assign n13216 = ~n13213 & ~n13215 ;
  assign n13217 = \b[16]  & n6307 ;
  assign n13218 = \a[33]  & \b[15]  ;
  assign n13219 = n6298 & n13218 ;
  assign n13220 = \a[35]  & ~n13219 ;
  assign n13221 = ~n13217 & n13220 ;
  assign n13222 = n13216 & n13221 ;
  assign n13223 = ~n13211 & n13222 ;
  assign n13224 = ~n13209 & n13223 ;
  assign n13225 = ~n13217 & ~n13219 ;
  assign n13226 = n13216 & n13225 ;
  assign n13227 = ~n13211 & n13226 ;
  assign n13228 = ~n13209 & n13227 ;
  assign n13229 = ~\a[35]  & ~n13228 ;
  assign n13230 = ~n13224 & ~n13229 ;
  assign n13231 = ~n13207 & ~n13230 ;
  assign n13232 = ~n13205 & n13231 ;
  assign n13233 = ~n13204 & n13230 ;
  assign n13234 = n13066 & n13233 ;
  assign n13235 = n13204 & n13230 ;
  assign n13236 = ~n13066 & n13235 ;
  assign n13237 = ~n13234 & ~n13236 ;
  assign n13238 = ~n13232 & n13237 ;
  assign n13239 = n13064 & ~n13238 ;
  assign n13240 = ~n13064 & n13238 ;
  assign n13241 = ~n13239 & ~n13240 ;
  assign n13242 = ~n2076 & n5211 ;
  assign n13243 = ~n1874 & n5211 ;
  assign n13244 = ~n1878 & n13243 ;
  assign n13245 = ~n13242 & ~n13244 ;
  assign n13246 = ~n2079 & ~n13245 ;
  assign n13247 = \b[17]  & n5595 ;
  assign n13248 = n5592 & n13247 ;
  assign n13249 = ~\a[30]  & \b[18]  ;
  assign n13250 = n5203 & n13249 ;
  assign n13251 = ~n13248 & ~n13250 ;
  assign n13252 = \b[19]  & n5209 ;
  assign n13253 = \a[30]  & \b[18]  ;
  assign n13254 = n5200 & n13253 ;
  assign n13255 = \a[32]  & ~n13254 ;
  assign n13256 = ~n13252 & n13255 ;
  assign n13257 = n13251 & n13256 ;
  assign n13258 = ~n13246 & n13257 ;
  assign n13259 = ~n13252 & ~n13254 ;
  assign n13260 = n13251 & n13259 ;
  assign n13261 = ~\a[32]  & ~n13260 ;
  assign n13262 = ~\a[32]  & ~n2079 ;
  assign n13263 = ~n13245 & n13262 ;
  assign n13264 = ~n13261 & ~n13263 ;
  assign n13265 = ~n13258 & n13264 ;
  assign n13266 = n13241 & ~n13265 ;
  assign n13267 = ~n13241 & n13265 ;
  assign n13268 = ~n13266 & ~n13267 ;
  assign n13269 = ~n13059 & n13268 ;
  assign n13270 = ~n12746 & ~n13268 ;
  assign n13271 = ~n13058 & n13270 ;
  assign n13272 = n2768 & n4249 ;
  assign n13273 = ~n2765 & n13272 ;
  assign n13274 = n4249 & n6462 ;
  assign n13275 = ~n2764 & n13274 ;
  assign n13276 = \b[20]  & n4647 ;
  assign n13277 = n4644 & n13276 ;
  assign n13278 = ~\a[27]  & \b[21]  ;
  assign n13279 = n4241 & n13278 ;
  assign n13280 = ~n13277 & ~n13279 ;
  assign n13281 = \b[22]  & n4247 ;
  assign n13282 = \a[27]  & \b[21]  ;
  assign n13283 = n4238 & n13282 ;
  assign n13284 = \a[29]  & ~n13283 ;
  assign n13285 = ~n13281 & n13284 ;
  assign n13286 = n13280 & n13285 ;
  assign n13287 = ~n13275 & n13286 ;
  assign n13288 = ~n13273 & n13287 ;
  assign n13289 = ~n13281 & ~n13283 ;
  assign n13290 = n13280 & n13289 ;
  assign n13291 = ~n13275 & n13290 ;
  assign n13292 = ~n13273 & n13291 ;
  assign n13293 = ~\a[29]  & ~n13292 ;
  assign n13294 = ~n13288 & ~n13293 ;
  assign n13295 = ~n13271 & ~n13294 ;
  assign n13296 = ~n13269 & n13295 ;
  assign n13297 = ~n13268 & n13294 ;
  assign n13298 = n13059 & n13297 ;
  assign n13299 = n13268 & n13294 ;
  assign n13300 = ~n13059 & n13299 ;
  assign n13301 = ~n13298 & ~n13300 ;
  assign n13302 = ~n13296 & n13301 ;
  assign n13303 = n3402 & ~n3567 ;
  assign n13304 = ~n3565 & n13303 ;
  assign n13305 = \b[23]  & n3733 ;
  assign n13306 = n3730 & n13305 ;
  assign n13307 = ~\a[24]  & \b[24]  ;
  assign n13308 = n3394 & n13307 ;
  assign n13309 = ~n13306 & ~n13308 ;
  assign n13310 = \b[25]  & n3400 ;
  assign n13311 = \a[24]  & \b[24]  ;
  assign n13312 = n3391 & n13311 ;
  assign n13313 = \a[26]  & ~n13312 ;
  assign n13314 = ~n13310 & n13313 ;
  assign n13315 = n13309 & n13314 ;
  assign n13316 = ~n13304 & n13315 ;
  assign n13317 = ~n13310 & ~n13312 ;
  assign n13318 = n13309 & n13317 ;
  assign n13319 = ~n13304 & n13318 ;
  assign n13320 = ~\a[26]  & ~n13319 ;
  assign n13321 = ~n13316 & ~n13320 ;
  assign n13322 = ~n13302 & ~n13321 ;
  assign n13323 = n13057 & n13322 ;
  assign n13324 = n13302 & ~n13321 ;
  assign n13325 = ~n13057 & n13324 ;
  assign n13326 = ~n13323 & ~n13325 ;
  assign n13327 = ~n13302 & n13321 ;
  assign n13328 = ~n13057 & n13327 ;
  assign n13329 = n13302 & n13321 ;
  assign n13330 = n13057 & n13329 ;
  assign n13331 = ~n13328 & ~n13330 ;
  assign n13332 = n13326 & n13331 ;
  assign n13333 = ~n13054 & ~n13332 ;
  assign n13334 = ~n13030 & n13333 ;
  assign n13335 = ~n13054 & n13332 ;
  assign n13336 = n13030 & n13335 ;
  assign n13337 = ~n13334 & ~n13336 ;
  assign n13338 = n13054 & ~n13332 ;
  assign n13339 = n13030 & n13338 ;
  assign n13340 = n13054 & n13332 ;
  assign n13341 = ~n13030 & n13340 ;
  assign n13342 = ~n13339 & ~n13341 ;
  assign n13343 = n13337 & n13342 ;
  assign n13344 = ~n13029 & ~n13343 ;
  assign n13345 = n13012 & n13344 ;
  assign n13346 = ~n13029 & n13343 ;
  assign n13347 = ~n13012 & n13346 ;
  assign n13348 = ~n13345 & ~n13347 ;
  assign n13349 = n13029 & ~n13343 ;
  assign n13350 = ~n13012 & n13349 ;
  assign n13351 = n13029 & n13343 ;
  assign n13352 = n13012 & n13351 ;
  assign n13353 = ~n13350 & ~n13352 ;
  assign n13354 = n13348 & n13353 ;
  assign n13355 = ~n13009 & n13354 ;
  assign n13356 = n12846 & ~n13354 ;
  assign n13357 = ~n13008 & n13356 ;
  assign n13358 = ~n1304 & ~n5850 ;
  assign n13359 = ~n6565 & n13358 ;
  assign n13360 = ~n6561 & n13359 ;
  assign n13361 = ~n1464 & n13360 ;
  assign n13362 = n1467 & n6565 ;
  assign n13363 = ~n6562 & n13362 ;
  assign n13364 = ~n13361 & ~n13363 ;
  assign n13365 = \b[32]  & n1652 ;
  assign n13366 = n1649 & n13365 ;
  assign n13367 = ~\a[15]  & \b[33]  ;
  assign n13368 = n1459 & n13367 ;
  assign n13369 = ~n13366 & ~n13368 ;
  assign n13370 = \b[34]  & n1465 ;
  assign n13371 = \a[15]  & \b[33]  ;
  assign n13372 = n1456 & n13371 ;
  assign n13373 = \a[17]  & ~n13372 ;
  assign n13374 = ~n13370 & n13373 ;
  assign n13375 = n13369 & n13374 ;
  assign n13376 = n13364 & n13375 ;
  assign n13377 = ~n13370 & ~n13372 ;
  assign n13378 = n13369 & n13377 ;
  assign n13379 = n13364 & n13378 ;
  assign n13380 = ~\a[17]  & ~n13379 ;
  assign n13381 = ~n13376 & ~n13380 ;
  assign n13382 = ~n13357 & ~n13381 ;
  assign n13383 = ~n13355 & n13382 ;
  assign n13384 = ~n13354 & n13381 ;
  assign n13385 = n13009 & n13384 ;
  assign n13386 = n13354 & n13381 ;
  assign n13387 = ~n13009 & n13386 ;
  assign n13388 = ~n13385 & ~n13387 ;
  assign n13389 = ~n13383 & n13388 ;
  assign n13390 = n999 & ~n7761 ;
  assign n13391 = ~n7759 & n13390 ;
  assign n13392 = \b[35]  & n1182 ;
  assign n13393 = n1179 & n13392 ;
  assign n13394 = \b[37]  & n997 ;
  assign n13395 = \a[11]  & \b[36]  ;
  assign n13396 = n1180 & n13395 ;
  assign n13397 = ~\a[12]  & \b[36]  ;
  assign n13398 = n7674 & n13397 ;
  assign n13399 = ~n13396 & ~n13398 ;
  assign n13400 = ~n13394 & n13399 ;
  assign n13401 = ~n13393 & n13400 ;
  assign n13402 = ~n13391 & n13401 ;
  assign n13403 = ~\a[14]  & ~n13402 ;
  assign n13404 = \a[14]  & n13401 ;
  assign n13405 = ~n13391 & n13404 ;
  assign n13406 = ~n13403 & ~n13405 ;
  assign n13407 = ~n13389 & ~n13406 ;
  assign n13408 = n13007 & n13407 ;
  assign n13409 = n13389 & ~n13406 ;
  assign n13410 = ~n13007 & n13409 ;
  assign n13411 = ~n13408 & ~n13410 ;
  assign n13412 = ~n13389 & n13406 ;
  assign n13413 = ~n13007 & n13412 ;
  assign n13414 = n13389 & n13406 ;
  assign n13415 = n13007 & n13414 ;
  assign n13416 = ~n13413 & ~n13415 ;
  assign n13417 = n13411 & n13416 ;
  assign n13418 = ~n13004 & n13417 ;
  assign n13419 = ~n12907 & ~n13417 ;
  assign n13420 = ~n13003 & n13419 ;
  assign n13421 = n646 & n9044 ;
  assign n13422 = ~n9041 & n13421 ;
  assign n13423 = n646 & ~n9044 ;
  assign n13424 = ~n8597 & n13423 ;
  assign n13425 = ~n9040 & n13424 ;
  assign n13426 = \b[38]  & n796 ;
  assign n13427 = n793 & n13426 ;
  assign n13428 = ~\a[9]  & \b[39]  ;
  assign n13429 = n638 & n13428 ;
  assign n13430 = ~n13427 & ~n13429 ;
  assign n13431 = \b[40]  & n644 ;
  assign n13432 = \a[9]  & \b[39]  ;
  assign n13433 = n635 & n13432 ;
  assign n13434 = \a[11]  & ~n13433 ;
  assign n13435 = ~n13431 & n13434 ;
  assign n13436 = n13430 & n13435 ;
  assign n13437 = ~n13425 & n13436 ;
  assign n13438 = ~n13422 & n13437 ;
  assign n13439 = ~n13431 & ~n13433 ;
  assign n13440 = n13430 & n13439 ;
  assign n13441 = ~n13425 & n13440 ;
  assign n13442 = ~n13422 & n13441 ;
  assign n13443 = ~\a[11]  & ~n13442 ;
  assign n13444 = ~n13438 & ~n13443 ;
  assign n13445 = ~n13420 & ~n13444 ;
  assign n13446 = ~n13418 & n13445 ;
  assign n13447 = ~n13417 & n13444 ;
  assign n13448 = n13004 & n13447 ;
  assign n13449 = n13417 & n13444 ;
  assign n13450 = ~n13004 & n13449 ;
  assign n13451 = ~n13448 & ~n13450 ;
  assign n13452 = ~n13446 & n13451 ;
  assign n13453 = n430 & ~n10409 ;
  assign n13454 = ~n10407 & n13453 ;
  assign n13455 = \b[41]  & n486 ;
  assign n13456 = n483 & n13455 ;
  assign n13457 = \b[43]  & n428 ;
  assign n13458 = \a[6]  & \b[42]  ;
  assign n13459 = n419 & n13458 ;
  assign n13460 = ~\a[6]  & \b[42]  ;
  assign n13461 = n422 & n13460 ;
  assign n13462 = ~n13459 & ~n13461 ;
  assign n13463 = ~n13457 & n13462 ;
  assign n13464 = ~n13456 & n13463 ;
  assign n13465 = ~n13454 & n13464 ;
  assign n13466 = ~\a[8]  & ~n13465 ;
  assign n13467 = \a[8]  & n13464 ;
  assign n13468 = ~n13454 & n13467 ;
  assign n13469 = ~n13466 & ~n13468 ;
  assign n13470 = ~n13452 & ~n13469 ;
  assign n13471 = n13002 & n13470 ;
  assign n13472 = n13452 & ~n13469 ;
  assign n13473 = ~n13002 & n13472 ;
  assign n13474 = ~n13471 & ~n13473 ;
  assign n13475 = ~n13452 & n13469 ;
  assign n13476 = ~n13002 & n13475 ;
  assign n13477 = n13452 & n13469 ;
  assign n13478 = n13002 & n13477 ;
  assign n13479 = ~n13476 & ~n13478 ;
  assign n13480 = n13474 & n13479 ;
  assign n13481 = n252 & n11906 ;
  assign n13482 = ~n11903 & n13481 ;
  assign n13483 = ~n11392 & ~n11906 ;
  assign n13484 = n252 & n13483 ;
  assign n13485 = ~n11902 & n13484 ;
  assign n13486 = \b[44]  & n303 ;
  assign n13487 = n300 & n13486 ;
  assign n13488 = ~\a[3]  & \b[45]  ;
  assign n13489 = n244 & n13488 ;
  assign n13490 = ~n13487 & ~n13489 ;
  assign n13491 = \b[46]  & n250 ;
  assign n13492 = \a[3]  & \b[45]  ;
  assign n13493 = n241 & n13492 ;
  assign n13494 = \a[5]  & ~n13493 ;
  assign n13495 = ~n13491 & n13494 ;
  assign n13496 = n13490 & n13495 ;
  assign n13497 = ~n13485 & n13496 ;
  assign n13498 = ~n13482 & n13497 ;
  assign n13499 = ~n13491 & ~n13493 ;
  assign n13500 = n13490 & n13499 ;
  assign n13501 = ~n13485 & n13500 ;
  assign n13502 = ~n13482 & n13501 ;
  assign n13503 = ~\a[5]  & ~n13502 ;
  assign n13504 = ~n13498 & ~n13503 ;
  assign n13505 = ~n13480 & ~n13504 ;
  assign n13506 = ~n12999 & n13505 ;
  assign n13507 = n13480 & ~n13504 ;
  assign n13508 = n12999 & n13507 ;
  assign n13509 = ~n13506 & ~n13508 ;
  assign n13510 = ~n13480 & n13504 ;
  assign n13511 = n12999 & n13510 ;
  assign n13512 = n13480 & n13504 ;
  assign n13513 = ~n12999 & n13512 ;
  assign n13514 = ~n13511 & ~n13513 ;
  assign n13515 = n13509 & n13514 ;
  assign n13516 = ~n12433 & n12478 ;
  assign n13517 = ~n12474 & n13516 ;
  assign n13518 = ~n12477 & ~n13517 ;
  assign n13519 = ~\b[48]  & ~\b[49]  ;
  assign n13520 = \b[48]  & \b[49]  ;
  assign n13521 = ~n13519 & ~n13520 ;
  assign n13522 = ~n13518 & n13521 ;
  assign n13523 = ~n12477 & ~n13521 ;
  assign n13524 = ~n13517 & n13523 ;
  assign n13525 = n134 & ~n13524 ;
  assign n13526 = ~n13522 & n13525 ;
  assign n13527 = \a[0]  & \b[49]  ;
  assign n13528 = n133 & n13527 ;
  assign n13529 = \b[48]  & n141 ;
  assign n13530 = ~\a[1]  & \b[47]  ;
  assign n13531 = n10416 & n13530 ;
  assign n13532 = ~n13529 & ~n13531 ;
  assign n13533 = ~n13528 & n13532 ;
  assign n13534 = ~n13526 & n13533 ;
  assign n13535 = ~\a[2]  & ~n13534 ;
  assign n13536 = \a[2]  & n13533 ;
  assign n13537 = ~n13526 & n13536 ;
  assign n13538 = ~n13535 & ~n13537 ;
  assign n13539 = ~n13515 & n13538 ;
  assign n13540 = ~n12998 & n13539 ;
  assign n13541 = n13515 & n13538 ;
  assign n13542 = n12998 & n13541 ;
  assign n13543 = ~n13540 & ~n13542 ;
  assign n13544 = ~n13515 & ~n13538 ;
  assign n13545 = n12998 & n13544 ;
  assign n13546 = n13515 & ~n13538 ;
  assign n13547 = ~n12998 & n13546 ;
  assign n13548 = ~n13545 & ~n13547 ;
  assign n13549 = n13543 & n13548 ;
  assign n13550 = ~n12995 & n13549 ;
  assign n13551 = n12990 & ~n13549 ;
  assign n13552 = ~n12992 & n13551 ;
  assign n13553 = ~n13550 & ~n13552 ;
  assign n13554 = n12990 & n13548 ;
  assign n13555 = ~n12992 & n13554 ;
  assign n13556 = n13543 & ~n13555 ;
  assign n13557 = n12998 & n13515 ;
  assign n13558 = n13509 & ~n13557 ;
  assign n13559 = n252 & ~n12438 ;
  assign n13560 = ~n12436 & n13559 ;
  assign n13561 = \b[47]  & n250 ;
  assign n13562 = \a[3]  & \b[46]  ;
  assign n13563 = n241 & n13562 ;
  assign n13564 = ~n13561 & ~n13563 ;
  assign n13565 = \b[45]  & n303 ;
  assign n13566 = n300 & n13565 ;
  assign n13567 = ~\a[3]  & \b[46]  ;
  assign n13568 = n244 & n13567 ;
  assign n13569 = ~n13566 & ~n13568 ;
  assign n13570 = n13564 & n13569 ;
  assign n13571 = ~n13560 & n13570 ;
  assign n13572 = ~\a[5]  & ~n13571 ;
  assign n13573 = \a[5]  & n13570 ;
  assign n13574 = ~n13560 & n13573 ;
  assign n13575 = ~n13572 & ~n13574 ;
  assign n13576 = ~n12968 & n13474 ;
  assign n13577 = ~n12975 & n13576 ;
  assign n13578 = n13479 & ~n13577 ;
  assign n13579 = n13002 & n13452 ;
  assign n13580 = ~n13446 & ~n13579 ;
  assign n13581 = ~n12907 & n13411 ;
  assign n13582 = ~n13003 & n13581 ;
  assign n13583 = n13416 & ~n13582 ;
  assign n13584 = n13007 & n13389 ;
  assign n13585 = ~n13383 & ~n13584 ;
  assign n13586 = n12846 & n13348 ;
  assign n13587 = n13353 & ~n13586 ;
  assign n13588 = n12852 & n13353 ;
  assign n13589 = n12527 & n13588 ;
  assign n13590 = ~n13587 & ~n13589 ;
  assign n13591 = n13012 & n13343 ;
  assign n13592 = n13337 & ~n13591 ;
  assign n13593 = n1965 & n5810 ;
  assign n13594 = ~n5807 & n13593 ;
  assign n13595 = n1965 & ~n5810 ;
  assign n13596 = ~n5457 & n13595 ;
  assign n13597 = ~n5806 & n13596 ;
  assign n13598 = \b[30]  & n2218 ;
  assign n13599 = n2216 & n13598 ;
  assign n13600 = ~\a[18]  & \b[31]  ;
  assign n13601 = n1957 & n13600 ;
  assign n13602 = ~n13599 & ~n13601 ;
  assign n13603 = \b[32]  & n1963 ;
  assign n13604 = \a[18]  & \b[31]  ;
  assign n13605 = n2210 & n13604 ;
  assign n13606 = \a[20]  & ~n13605 ;
  assign n13607 = ~n13603 & n13606 ;
  assign n13608 = n13602 & n13607 ;
  assign n13609 = ~n13597 & n13608 ;
  assign n13610 = ~n13594 & n13609 ;
  assign n13611 = ~n13603 & ~n13605 ;
  assign n13612 = n13602 & n13611 ;
  assign n13613 = ~n13597 & n13612 ;
  assign n13614 = ~n13594 & n13613 ;
  assign n13615 = ~\a[20]  & ~n13614 ;
  assign n13616 = ~n13610 & ~n13615 ;
  assign n13617 = n2622 & ~n4502 ;
  assign n13618 = ~n4500 & n13617 ;
  assign n13619 = \b[29]  & n2620 ;
  assign n13620 = \a[21]  & \b[28]  ;
  assign n13621 = n2611 & n13620 ;
  assign n13622 = ~n13619 & ~n13621 ;
  assign n13623 = \b[27]  & n2912 ;
  assign n13624 = n2909 & n13623 ;
  assign n13625 = ~\a[21]  & \b[28]  ;
  assign n13626 = n2614 & n13625 ;
  assign n13627 = ~n13624 & ~n13626 ;
  assign n13628 = n13622 & n13627 ;
  assign n13629 = ~n13618 & n13628 ;
  assign n13630 = ~\a[23]  & ~n13629 ;
  assign n13631 = \a[23]  & n13628 ;
  assign n13632 = ~n13618 & n13631 ;
  assign n13633 = ~n13630 & ~n13632 ;
  assign n13634 = ~n12814 & n13326 ;
  assign n13635 = ~n12816 & n13634 ;
  assign n13636 = n13331 & ~n13635 ;
  assign n13637 = n13057 & n13302 ;
  assign n13638 = ~n13296 & ~n13637 ;
  assign n13639 = ~n3154 & ~n3562 ;
  assign n13640 = ~n3604 & n13639 ;
  assign n13641 = ~n3600 & n13640 ;
  assign n13642 = ~n3399 & n13641 ;
  assign n13643 = n3402 & n3604 ;
  assign n13644 = ~n3601 & n13643 ;
  assign n13645 = ~n13642 & ~n13644 ;
  assign n13646 = \b[24]  & n3733 ;
  assign n13647 = n3730 & n13646 ;
  assign n13648 = ~\a[24]  & \b[25]  ;
  assign n13649 = n3394 & n13648 ;
  assign n13650 = ~n13647 & ~n13649 ;
  assign n13651 = \b[26]  & n3400 ;
  assign n13652 = \a[24]  & \b[25]  ;
  assign n13653 = n3391 & n13652 ;
  assign n13654 = \a[26]  & ~n13653 ;
  assign n13655 = ~n13651 & n13654 ;
  assign n13656 = n13650 & n13655 ;
  assign n13657 = n13645 & n13656 ;
  assign n13658 = ~n13651 & ~n13653 ;
  assign n13659 = n13650 & n13658 ;
  assign n13660 = n13645 & n13659 ;
  assign n13661 = ~\a[26]  & ~n13660 ;
  assign n13662 = ~n13657 & ~n13661 ;
  assign n13663 = ~n12746 & ~n13266 ;
  assign n13664 = ~n13058 & n13663 ;
  assign n13665 = ~n13267 & ~n13664 ;
  assign n13666 = ~n13232 & ~n13240 ;
  assign n13667 = n2293 & n5211 ;
  assign n13668 = ~n2290 & n13667 ;
  assign n13669 = n5211 & n5705 ;
  assign n13670 = ~n2289 & n13669 ;
  assign n13671 = \b[18]  & n5595 ;
  assign n13672 = n5592 & n13671 ;
  assign n13673 = ~\a[30]  & \b[19]  ;
  assign n13674 = n5203 & n13673 ;
  assign n13675 = ~n13672 & ~n13674 ;
  assign n13676 = \b[20]  & n5209 ;
  assign n13677 = \a[30]  & \b[19]  ;
  assign n13678 = n5200 & n13677 ;
  assign n13679 = \a[32]  & ~n13678 ;
  assign n13680 = ~n13676 & n13679 ;
  assign n13681 = n13675 & n13680 ;
  assign n13682 = ~n13670 & n13681 ;
  assign n13683 = ~n13668 & n13682 ;
  assign n13684 = ~n13676 & ~n13678 ;
  assign n13685 = n13675 & n13684 ;
  assign n13686 = ~n13670 & n13685 ;
  assign n13687 = ~n13668 & n13686 ;
  assign n13688 = ~\a[32]  & ~n13687 ;
  assign n13689 = ~n13683 & ~n13688 ;
  assign n13690 = ~n12701 & n13203 ;
  assign n13691 = ~n13065 & n13690 ;
  assign n13692 = n13198 & ~n13691 ;
  assign n13693 = ~n1691 & n6309 ;
  assign n13694 = ~n1511 & n6309 ;
  assign n13695 = ~n1515 & n13694 ;
  assign n13696 = ~n13693 & ~n13695 ;
  assign n13697 = ~n1694 & ~n13696 ;
  assign n13698 = \b[15]  & n6778 ;
  assign n13699 = n6775 & n13698 ;
  assign n13700 = ~\a[33]  & \b[16]  ;
  assign n13701 = n6301 & n13700 ;
  assign n13702 = ~n13699 & ~n13701 ;
  assign n13703 = \b[17]  & n6307 ;
  assign n13704 = \a[33]  & \b[16]  ;
  assign n13705 = n6298 & n13704 ;
  assign n13706 = \a[35]  & ~n13705 ;
  assign n13707 = ~n13703 & n13706 ;
  assign n13708 = n13702 & n13707 ;
  assign n13709 = ~n13697 & n13708 ;
  assign n13710 = ~n13703 & ~n13705 ;
  assign n13711 = n13702 & n13710 ;
  assign n13712 = ~\a[35]  & ~n13711 ;
  assign n13713 = ~\a[35]  & ~n1694 ;
  assign n13714 = ~n13696 & n13713 ;
  assign n13715 = ~n13712 & ~n13714 ;
  assign n13716 = ~n13709 & n13715 ;
  assign n13717 = n13069 & n13193 ;
  assign n13718 = n13187 & ~n13717 ;
  assign n13719 = ~n728 & n8759 ;
  assign n13720 = ~n726 & n13719 ;
  assign n13721 = \b[11]  & n8757 ;
  assign n13722 = \a[39]  & \b[10]  ;
  assign n13723 = n8748 & n13722 ;
  assign n13724 = ~n13721 & ~n13723 ;
  assign n13725 = \b[9]  & n9301 ;
  assign n13726 = n9298 & n13725 ;
  assign n13727 = ~\a[39]  & \b[10]  ;
  assign n13728 = n8751 & n13727 ;
  assign n13729 = ~n13726 & ~n13728 ;
  assign n13730 = n13724 & n13729 ;
  assign n13731 = ~n13720 & n13730 ;
  assign n13732 = ~\a[41]  & ~n13731 ;
  assign n13733 = \a[41]  & n13730 ;
  assign n13734 = ~n13720 & n13733 ;
  assign n13735 = ~n13732 & ~n13734 ;
  assign n13736 = ~n12637 & ~n13156 ;
  assign n13737 = ~n13092 & n13736 ;
  assign n13738 = ~n13157 & ~n13737 ;
  assign n13739 = ~n505 & ~n9646 ;
  assign n13740 = ~n10079 & n13739 ;
  assign n13741 = n502 & n13740 ;
  assign n13742 = n505 & ~n9646 ;
  assign n13743 = ~n10079 & n13742 ;
  assign n13744 = ~n502 & n13743 ;
  assign n13745 = ~n13741 & ~n13744 ;
  assign n13746 = \b[6]  & n10681 ;
  assign n13747 = n10678 & n13746 ;
  assign n13748 = \b[8]  & n10080 ;
  assign n13749 = \a[41]  & \b[7]  ;
  assign n13750 = n10679 & n13749 ;
  assign n13751 = ~\a[42]  & \b[7]  ;
  assign n13752 = n10074 & n13751 ;
  assign n13753 = ~n13750 & ~n13752 ;
  assign n13754 = ~n13748 & n13753 ;
  assign n13755 = ~n13747 & n13754 ;
  assign n13756 = n13745 & n13755 ;
  assign n13757 = ~\a[44]  & ~n13756 ;
  assign n13758 = \a[44]  & n13755 ;
  assign n13759 = n13745 & n13758 ;
  assign n13760 = ~n13757 & ~n13759 ;
  assign n13761 = ~n13134 & ~n13136 ;
  assign n13762 = ~n273 & n11572 ;
  assign n13763 = ~n271 & n13762 ;
  assign n13764 = \b[5]  & n11570 ;
  assign n13765 = \a[45]  & \b[4]  ;
  assign n13766 = n11561 & n13765 ;
  assign n13767 = ~n13764 & ~n13766 ;
  assign n13768 = \b[3]  & n12159 ;
  assign n13769 = n12156 & n13768 ;
  assign n13770 = ~\a[45]  & \b[4]  ;
  assign n13771 = n11564 & n13770 ;
  assign n13772 = ~n13769 & ~n13771 ;
  assign n13773 = n13767 & n13772 ;
  assign n13774 = ~n13763 & n13773 ;
  assign n13775 = ~\a[47]  & ~n13774 ;
  assign n13776 = \a[47]  & n13773 ;
  assign n13777 = ~n13763 & n13776 ;
  assign n13778 = ~n13775 & ~n13777 ;
  assign n13779 = \a[50]  & ~n12607 ;
  assign n13780 = n13119 & n13779 ;
  assign n13781 = n13127 & n13780 ;
  assign n13782 = \a[50]  & ~n13781 ;
  assign n13783 = \b[2]  & n13123 ;
  assign n13784 = ~\a[48]  & \b[1]  ;
  assign n13785 = n13117 & n13784 ;
  assign n13786 = \a[47]  & ~\a[49]  ;
  assign n13787 = \a[48]  & \b[1]  ;
  assign n13788 = n13786 & n13787 ;
  assign n13789 = ~n13785 & ~n13788 ;
  assign n13790 = ~n13783 & n13789 ;
  assign n13791 = n157 & n13125 ;
  assign n13792 = n12606 & ~n13122 ;
  assign n13793 = ~\a[48]  & \a[49]  ;
  assign n13794 = ~n13114 & ~n13793 ;
  assign n13795 = \b[0]  & n13794 ;
  assign n13796 = n13792 & n13795 ;
  assign n13797 = ~n13791 & ~n13796 ;
  assign n13798 = n13790 & n13797 ;
  assign n13799 = ~n13782 & ~n13798 ;
  assign n13800 = n13782 & n13798 ;
  assign n13801 = ~n13799 & ~n13800 ;
  assign n13802 = ~n13778 & ~n13801 ;
  assign n13803 = n13778 & n13801 ;
  assign n13804 = ~n13802 & ~n13803 ;
  assign n13805 = ~n13761 & n13804 ;
  assign n13806 = n13761 & ~n13804 ;
  assign n13807 = ~n13805 & ~n13806 ;
  assign n13808 = ~n13760 & n13807 ;
  assign n13809 = n13760 & ~n13807 ;
  assign n13810 = ~n13808 & ~n13809 ;
  assign n13811 = n13738 & n13810 ;
  assign n13812 = ~n13738 & ~n13810 ;
  assign n13813 = ~n13811 & ~n13812 ;
  assign n13814 = n13735 & ~n13813 ;
  assign n13815 = ~n13735 & n13813 ;
  assign n13816 = ~n13814 & ~n13815 ;
  assign n13817 = n1087 & n7534 ;
  assign n13818 = ~n1084 & n13817 ;
  assign n13819 = n1552 & n7534 ;
  assign n13820 = ~n1083 & n13819 ;
  assign n13821 = \b[12]  & n7973 ;
  assign n13822 = n7970 & n13821 ;
  assign n13823 = \b[14]  & n7532 ;
  assign n13824 = \a[36]  & \b[13]  ;
  assign n13825 = n7523 & n13824 ;
  assign n13826 = ~\a[36]  & \b[13]  ;
  assign n13827 = n7526 & n13826 ;
  assign n13828 = ~n13825 & ~n13827 ;
  assign n13829 = ~n13823 & n13828 ;
  assign n13830 = ~n13822 & n13829 ;
  assign n13831 = ~n13820 & n13830 ;
  assign n13832 = ~n13818 & n13831 ;
  assign n13833 = ~\a[38]  & ~n13832 ;
  assign n13834 = \a[38]  & n13830 ;
  assign n13835 = ~n13820 & n13834 ;
  assign n13836 = ~n13818 & n13835 ;
  assign n13837 = ~n13833 & ~n13836 ;
  assign n13838 = ~n13816 & ~n13837 ;
  assign n13839 = ~n13718 & n13838 ;
  assign n13840 = n13816 & ~n13837 ;
  assign n13841 = n13718 & n13840 ;
  assign n13842 = ~n13839 & ~n13841 ;
  assign n13843 = ~n13816 & n13837 ;
  assign n13844 = n13718 & n13843 ;
  assign n13845 = n13816 & n13837 ;
  assign n13846 = ~n13718 & n13845 ;
  assign n13847 = ~n13844 & ~n13846 ;
  assign n13848 = n13842 & n13847 ;
  assign n13849 = ~n13716 & ~n13848 ;
  assign n13850 = n13692 & n13849 ;
  assign n13851 = ~n13716 & n13848 ;
  assign n13852 = ~n13692 & n13851 ;
  assign n13853 = ~n13850 & ~n13852 ;
  assign n13854 = n13716 & ~n13848 ;
  assign n13855 = ~n13692 & n13854 ;
  assign n13856 = n13716 & n13848 ;
  assign n13857 = n13692 & n13856 ;
  assign n13858 = ~n13855 & ~n13857 ;
  assign n13859 = n13853 & n13858 ;
  assign n13860 = ~n13689 & ~n13859 ;
  assign n13861 = ~n13666 & n13860 ;
  assign n13862 = ~n13689 & n13859 ;
  assign n13863 = n13666 & n13862 ;
  assign n13864 = ~n13861 & ~n13863 ;
  assign n13865 = n13689 & ~n13859 ;
  assign n13866 = n13666 & n13865 ;
  assign n13867 = n13689 & n13859 ;
  assign n13868 = ~n13666 & n13867 ;
  assign n13869 = ~n13866 & ~n13868 ;
  assign n13870 = n13864 & n13869 ;
  assign n13871 = ~n13665 & ~n13870 ;
  assign n13872 = ~n13267 & n13870 ;
  assign n13873 = ~n13664 & n13872 ;
  assign n13874 = ~n3022 & n4249 ;
  assign n13875 = ~n3020 & n13874 ;
  assign n13876 = \b[23]  & n4247 ;
  assign n13877 = \a[27]  & \b[22]  ;
  assign n13878 = n4238 & n13877 ;
  assign n13879 = ~n13876 & ~n13878 ;
  assign n13880 = \b[21]  & n4647 ;
  assign n13881 = n4644 & n13880 ;
  assign n13882 = ~\a[27]  & \b[22]  ;
  assign n13883 = n4241 & n13882 ;
  assign n13884 = ~n13881 & ~n13883 ;
  assign n13885 = n13879 & n13884 ;
  assign n13886 = ~n13875 & n13885 ;
  assign n13887 = ~\a[29]  & ~n13886 ;
  assign n13888 = \a[29]  & n13885 ;
  assign n13889 = ~n13875 & n13888 ;
  assign n13890 = ~n13887 & ~n13889 ;
  assign n13891 = ~n13873 & ~n13890 ;
  assign n13892 = ~n13871 & n13891 ;
  assign n13893 = ~n13870 & n13890 ;
  assign n13894 = ~n13665 & n13893 ;
  assign n13895 = n13870 & n13890 ;
  assign n13896 = n13665 & n13895 ;
  assign n13897 = ~n13894 & ~n13896 ;
  assign n13898 = ~n13892 & n13897 ;
  assign n13899 = n13662 & ~n13898 ;
  assign n13900 = n13638 & n13899 ;
  assign n13901 = n13662 & n13898 ;
  assign n13902 = ~n13638 & n13901 ;
  assign n13903 = ~n13900 & ~n13902 ;
  assign n13904 = ~n13638 & n13898 ;
  assign n13905 = ~n13296 & ~n13898 ;
  assign n13906 = ~n13637 & n13905 ;
  assign n13907 = ~n13662 & ~n13906 ;
  assign n13908 = ~n13904 & n13907 ;
  assign n13909 = n13903 & ~n13908 ;
  assign n13910 = n13636 & n13909 ;
  assign n13911 = ~n13636 & ~n13909 ;
  assign n13912 = ~n13910 & ~n13911 ;
  assign n13913 = n13633 & ~n13912 ;
  assign n13914 = ~n13633 & n13912 ;
  assign n13915 = ~n13913 & ~n13914 ;
  assign n13916 = n13616 & ~n13915 ;
  assign n13917 = n13592 & n13916 ;
  assign n13918 = n13616 & n13915 ;
  assign n13919 = ~n13592 & n13918 ;
  assign n13920 = ~n13917 & ~n13919 ;
  assign n13921 = ~n13616 & ~n13915 ;
  assign n13922 = ~n13592 & n13921 ;
  assign n13923 = ~n13616 & n13915 ;
  assign n13924 = n13592 & n13923 ;
  assign n13925 = ~n13922 & ~n13924 ;
  assign n13926 = n13920 & n13925 ;
  assign n13927 = ~n13590 & n13926 ;
  assign n13928 = n13590 & ~n13926 ;
  assign n13929 = ~n13927 & ~n13928 ;
  assign n13930 = n1467 & ~n6610 ;
  assign n13931 = ~n6608 & n13930 ;
  assign n13932 = \b[35]  & n1465 ;
  assign n13933 = \a[15]  & \b[34]  ;
  assign n13934 = n1456 & n13933 ;
  assign n13935 = ~n13932 & ~n13934 ;
  assign n13936 = \b[33]  & n1652 ;
  assign n13937 = n1649 & n13936 ;
  assign n13938 = ~\a[15]  & \b[34]  ;
  assign n13939 = n1459 & n13938 ;
  assign n13940 = ~n13937 & ~n13939 ;
  assign n13941 = n13935 & n13940 ;
  assign n13942 = ~n13931 & n13941 ;
  assign n13943 = ~\a[17]  & ~n13942 ;
  assign n13944 = \a[17]  & n13941 ;
  assign n13945 = ~n13931 & n13944 ;
  assign n13946 = ~n13943 & ~n13945 ;
  assign n13947 = n13929 & ~n13946 ;
  assign n13948 = ~n13929 & n13946 ;
  assign n13949 = ~n13947 & ~n13948 ;
  assign n13950 = ~n13585 & n13949 ;
  assign n13951 = ~n13383 & ~n13949 ;
  assign n13952 = ~n13584 & n13951 ;
  assign n13953 = n999 & n8175 ;
  assign n13954 = ~n8172 & n13953 ;
  assign n13955 = n999 & ~n8175 ;
  assign n13956 = ~n7756 & n13955 ;
  assign n13957 = ~n8171 & n13956 ;
  assign n13958 = \b[36]  & n1182 ;
  assign n13959 = n1179 & n13958 ;
  assign n13960 = \b[38]  & n997 ;
  assign n13961 = \a[11]  & \b[37]  ;
  assign n13962 = n1180 & n13961 ;
  assign n13963 = ~\a[12]  & \b[37]  ;
  assign n13964 = n7674 & n13963 ;
  assign n13965 = ~n13962 & ~n13964 ;
  assign n13966 = ~n13960 & n13965 ;
  assign n13967 = ~n13959 & n13966 ;
  assign n13968 = ~n13957 & n13967 ;
  assign n13969 = ~n13954 & n13968 ;
  assign n13970 = ~\a[14]  & ~n13969 ;
  assign n13971 = \a[14]  & n13967 ;
  assign n13972 = ~n13957 & n13971 ;
  assign n13973 = ~n13954 & n13972 ;
  assign n13974 = ~n13970 & ~n13973 ;
  assign n13975 = ~n13952 & ~n13974 ;
  assign n13976 = ~n13950 & n13975 ;
  assign n13977 = ~n13949 & n13974 ;
  assign n13978 = n13585 & n13977 ;
  assign n13979 = n13949 & n13974 ;
  assign n13980 = ~n13585 & n13979 ;
  assign n13981 = ~n13978 & ~n13980 ;
  assign n13982 = ~n13976 & n13981 ;
  assign n13983 = n646 & ~n9482 ;
  assign n13984 = ~n9480 & n13983 ;
  assign n13985 = \b[41]  & n644 ;
  assign n13986 = \a[9]  & \b[40]  ;
  assign n13987 = n635 & n13986 ;
  assign n13988 = ~n13985 & ~n13987 ;
  assign n13989 = \b[39]  & n796 ;
  assign n13990 = n793 & n13989 ;
  assign n13991 = ~\a[9]  & \b[40]  ;
  assign n13992 = n638 & n13991 ;
  assign n13993 = ~n13990 & ~n13992 ;
  assign n13994 = n13988 & n13993 ;
  assign n13995 = ~n13984 & n13994 ;
  assign n13996 = ~\a[11]  & ~n13995 ;
  assign n13997 = \a[11]  & n13994 ;
  assign n13998 = ~n13984 & n13997 ;
  assign n13999 = ~n13996 & ~n13998 ;
  assign n14000 = ~n13982 & ~n13999 ;
  assign n14001 = n13583 & n14000 ;
  assign n14002 = n13982 & ~n13999 ;
  assign n14003 = ~n13583 & n14002 ;
  assign n14004 = ~n14001 & ~n14003 ;
  assign n14005 = ~n13982 & n13999 ;
  assign n14006 = ~n13583 & n14005 ;
  assign n14007 = n13982 & n13999 ;
  assign n14008 = n13583 & n14007 ;
  assign n14009 = ~n14006 & ~n14008 ;
  assign n14010 = n14004 & n14009 ;
  assign n14011 = ~n13580 & n14010 ;
  assign n14012 = ~n13446 & ~n14010 ;
  assign n14013 = ~n13579 & n14012 ;
  assign n14014 = n430 & ~n10892 ;
  assign n14015 = ~n10890 & n14014 ;
  assign n14016 = \b[42]  & n486 ;
  assign n14017 = n483 & n14016 ;
  assign n14018 = ~\a[6]  & \b[43]  ;
  assign n14019 = n422 & n14018 ;
  assign n14020 = ~n14017 & ~n14019 ;
  assign n14021 = \b[44]  & n428 ;
  assign n14022 = \a[6]  & \b[43]  ;
  assign n14023 = n419 & n14022 ;
  assign n14024 = \a[8]  & ~n14023 ;
  assign n14025 = ~n14021 & n14024 ;
  assign n14026 = n14020 & n14025 ;
  assign n14027 = ~n14015 & n14026 ;
  assign n14028 = ~n14021 & ~n14023 ;
  assign n14029 = n14020 & n14028 ;
  assign n14030 = ~n14015 & n14029 ;
  assign n14031 = ~\a[8]  & ~n14030 ;
  assign n14032 = ~n14027 & ~n14031 ;
  assign n14033 = ~n14013 & ~n14032 ;
  assign n14034 = ~n14011 & n14033 ;
  assign n14035 = ~n14010 & n14032 ;
  assign n14036 = n13580 & n14035 ;
  assign n14037 = n14010 & n14032 ;
  assign n14038 = ~n13580 & n14037 ;
  assign n14039 = ~n14036 & ~n14038 ;
  assign n14040 = ~n14034 & n14039 ;
  assign n14041 = n13578 & n14040 ;
  assign n14042 = ~n13578 & ~n14040 ;
  assign n14043 = ~n14041 & ~n14042 ;
  assign n14044 = ~n13575 & n14043 ;
  assign n14045 = n13575 & ~n14043 ;
  assign n14046 = ~n14044 & ~n14045 ;
  assign n14047 = ~n12477 & ~n13520 ;
  assign n14048 = ~n13517 & n14047 ;
  assign n14049 = ~n13519 & ~n14048 ;
  assign n14050 = ~\b[49]  & ~\b[50]  ;
  assign n14051 = \b[49]  & \b[50]  ;
  assign n14052 = ~n14050 & ~n14051 ;
  assign n14053 = n134 & n14052 ;
  assign n14054 = ~n14049 & n14053 ;
  assign n14055 = n134 & ~n14052 ;
  assign n14056 = ~n13519 & n14055 ;
  assign n14057 = ~n14048 & n14056 ;
  assign n14058 = \a[0]  & \b[50]  ;
  assign n14059 = n133 & n14058 ;
  assign n14060 = \b[49]  & n141 ;
  assign n14061 = ~\a[1]  & \b[48]  ;
  assign n14062 = n10416 & n14061 ;
  assign n14063 = ~n14060 & ~n14062 ;
  assign n14064 = ~n14059 & n14063 ;
  assign n14065 = \a[2]  & n14064 ;
  assign n14066 = ~n14057 & n14065 ;
  assign n14067 = ~n14054 & n14066 ;
  assign n14068 = ~n14057 & n14064 ;
  assign n14069 = ~n14054 & n14068 ;
  assign n14070 = ~\a[2]  & ~n14069 ;
  assign n14071 = ~n14067 & ~n14070 ;
  assign n14072 = ~n14046 & ~n14071 ;
  assign n14073 = ~n13558 & n14072 ;
  assign n14074 = n14046 & ~n14071 ;
  assign n14075 = n13558 & n14074 ;
  assign n14076 = ~n14073 & ~n14075 ;
  assign n14077 = ~n14046 & n14071 ;
  assign n14078 = n13558 & n14077 ;
  assign n14079 = n14046 & n14071 ;
  assign n14080 = ~n13558 & n14079 ;
  assign n14081 = ~n14078 & ~n14080 ;
  assign n14082 = n14076 & n14081 ;
  assign n14083 = n13556 & n14082 ;
  assign n14084 = ~n13556 & ~n14082 ;
  assign n14085 = ~n14083 & ~n14084 ;
  assign n14086 = n14076 & ~n14083 ;
  assign n14087 = n13509 & ~n14044 ;
  assign n14088 = ~n13557 & n14087 ;
  assign n14089 = ~n14045 & ~n14088 ;
  assign n14090 = ~n13519 & n14052 ;
  assign n14091 = ~n14048 & n14090 ;
  assign n14092 = ~n14051 & ~n14091 ;
  assign n14093 = ~\b[50]  & ~\b[51]  ;
  assign n14094 = \b[50]  & \b[51]  ;
  assign n14095 = ~n14093 & ~n14094 ;
  assign n14096 = ~n14092 & n14095 ;
  assign n14097 = ~n14051 & ~n14095 ;
  assign n14098 = ~n14091 & n14097 ;
  assign n14099 = n134 & ~n14098 ;
  assign n14100 = ~n14096 & n14099 ;
  assign n14101 = \a[0]  & \b[51]  ;
  assign n14102 = n133 & n14101 ;
  assign n14103 = \b[50]  & n141 ;
  assign n14104 = ~\a[1]  & \b[49]  ;
  assign n14105 = n10416 & n14104 ;
  assign n14106 = ~n14103 & ~n14105 ;
  assign n14107 = ~n14102 & n14106 ;
  assign n14108 = ~n14100 & n14107 ;
  assign n14109 = ~\a[2]  & ~n14108 ;
  assign n14110 = \a[2]  & n14107 ;
  assign n14111 = ~n14100 & n14110 ;
  assign n14112 = ~n14109 & ~n14111 ;
  assign n14113 = ~n14034 & ~n14041 ;
  assign n14114 = n252 & n12478 ;
  assign n14115 = ~n12475 & n14114 ;
  assign n14116 = n252 & ~n12478 ;
  assign n14117 = ~n12433 & n14116 ;
  assign n14118 = ~n12474 & n14117 ;
  assign n14119 = \b[46]  & n303 ;
  assign n14120 = n300 & n14119 ;
  assign n14121 = ~\a[3]  & \b[47]  ;
  assign n14122 = n244 & n14121 ;
  assign n14123 = ~n14120 & ~n14122 ;
  assign n14124 = \b[48]  & n250 ;
  assign n14125 = \a[3]  & \b[47]  ;
  assign n14126 = n241 & n14125 ;
  assign n14127 = \a[5]  & ~n14126 ;
  assign n14128 = ~n14124 & n14127 ;
  assign n14129 = n14123 & n14128 ;
  assign n14130 = ~n14118 & n14129 ;
  assign n14131 = ~n14115 & n14130 ;
  assign n14132 = ~n14124 & ~n14126 ;
  assign n14133 = n14123 & n14132 ;
  assign n14134 = ~n14118 & n14133 ;
  assign n14135 = ~n14115 & n14134 ;
  assign n14136 = ~\a[5]  & ~n14135 ;
  assign n14137 = ~n14131 & ~n14136 ;
  assign n14138 = n13583 & n13982 ;
  assign n14139 = ~n13976 & ~n14138 ;
  assign n14140 = ~n13383 & ~n13947 ;
  assign n14141 = ~n13584 & n14140 ;
  assign n14142 = ~n13948 & ~n14141 ;
  assign n14143 = n13925 & ~n13927 ;
  assign n14144 = n1467 & n7337 ;
  assign n14145 = ~n7334 & n14144 ;
  assign n14146 = n1467 & ~n7337 ;
  assign n14147 = ~n6605 & n14146 ;
  assign n14148 = ~n7333 & n14147 ;
  assign n14149 = \b[34]  & n1652 ;
  assign n14150 = n1649 & n14149 ;
  assign n14151 = ~\a[15]  & \b[35]  ;
  assign n14152 = n1459 & n14151 ;
  assign n14153 = ~n14150 & ~n14152 ;
  assign n14154 = \b[36]  & n1465 ;
  assign n14155 = \a[15]  & \b[35]  ;
  assign n14156 = n1456 & n14155 ;
  assign n14157 = \a[17]  & ~n14156 ;
  assign n14158 = ~n14154 & n14157 ;
  assign n14159 = n14153 & n14158 ;
  assign n14160 = ~n14148 & n14159 ;
  assign n14161 = ~n14145 & n14160 ;
  assign n14162 = ~n14154 & ~n14156 ;
  assign n14163 = n14153 & n14162 ;
  assign n14164 = ~n14148 & n14163 ;
  assign n14165 = ~n14145 & n14164 ;
  assign n14166 = ~\a[17]  & ~n14165 ;
  assign n14167 = ~n14161 & ~n14166 ;
  assign n14168 = n13337 & ~n13914 ;
  assign n14169 = ~n13591 & n14168 ;
  assign n14170 = ~n13913 & ~n14169 ;
  assign n14171 = ~n13908 & ~n13910 ;
  assign n14172 = n2622 & n5105 ;
  assign n14173 = ~n5102 & n14172 ;
  assign n14174 = n2622 & ~n5105 ;
  assign n14175 = ~n4497 & n14174 ;
  assign n14176 = ~n5101 & n14175 ;
  assign n14177 = \b[28]  & n2912 ;
  assign n14178 = n2909 & n14177 ;
  assign n14179 = ~\a[21]  & \b[29]  ;
  assign n14180 = n2614 & n14179 ;
  assign n14181 = ~n14178 & ~n14180 ;
  assign n14182 = \b[30]  & n2620 ;
  assign n14183 = \a[21]  & \b[29]  ;
  assign n14184 = n2611 & n14183 ;
  assign n14185 = \a[23]  & ~n14184 ;
  assign n14186 = ~n14182 & n14185 ;
  assign n14187 = n14181 & n14186 ;
  assign n14188 = ~n14176 & n14187 ;
  assign n14189 = ~n14173 & n14188 ;
  assign n14190 = ~n14182 & ~n14184 ;
  assign n14191 = n14181 & n14190 ;
  assign n14192 = ~n14176 & n14191 ;
  assign n14193 = ~n14173 & n14192 ;
  assign n14194 = ~\a[23]  & ~n14193 ;
  assign n14195 = ~n14189 & ~n14194 ;
  assign n14196 = ~n13296 & ~n13892 ;
  assign n14197 = ~n13637 & n14196 ;
  assign n14198 = n13897 & ~n14197 ;
  assign n14199 = n13864 & ~n13873 ;
  assign n14200 = ~n13232 & n13853 ;
  assign n14201 = ~n13240 & n14200 ;
  assign n14202 = n13858 & ~n14201 ;
  assign n14203 = n13692 & n13848 ;
  assign n14204 = n13842 & ~n14203 ;
  assign n14205 = n13187 & ~n13815 ;
  assign n14206 = ~n13717 & n14205 ;
  assign n14207 = ~n13814 & ~n14206 ;
  assign n14208 = ~n1230 & n7534 ;
  assign n14209 = ~n1086 & n7534 ;
  assign n14210 = ~n1226 & n14209 ;
  assign n14211 = ~n14208 & ~n14210 ;
  assign n14212 = ~n1233 & ~n14211 ;
  assign n14213 = \b[13]  & n7973 ;
  assign n14214 = n7970 & n14213 ;
  assign n14215 = \b[15]  & n7532 ;
  assign n14216 = \a[36]  & \b[14]  ;
  assign n14217 = n7523 & n14216 ;
  assign n14218 = ~\a[36]  & \b[14]  ;
  assign n14219 = n7526 & n14218 ;
  assign n14220 = ~n14217 & ~n14219 ;
  assign n14221 = ~n14215 & n14220 ;
  assign n14222 = ~n14214 & n14221 ;
  assign n14223 = ~\a[38]  & n14222 ;
  assign n14224 = ~n14212 & n14223 ;
  assign n14225 = \a[38]  & ~n14222 ;
  assign n14226 = \a[38]  & ~n1233 ;
  assign n14227 = ~n14211 & n14226 ;
  assign n14228 = ~n14225 & ~n14227 ;
  assign n14229 = ~n14224 & n14228 ;
  assign n14230 = ~n13808 & ~n13811 ;
  assign n14231 = ~n909 & ~n8272 ;
  assign n14232 = ~n8756 & n14231 ;
  assign n14233 = n906 & n14232 ;
  assign n14234 = n909 & ~n8272 ;
  assign n14235 = ~n8756 & n14234 ;
  assign n14236 = ~n906 & n14235 ;
  assign n14237 = ~n14233 & ~n14236 ;
  assign n14238 = \b[10]  & n9301 ;
  assign n14239 = n9298 & n14238 ;
  assign n14240 = ~\a[39]  & \b[11]  ;
  assign n14241 = n8751 & n14240 ;
  assign n14242 = ~n14239 & ~n14241 ;
  assign n14243 = \b[12]  & n8757 ;
  assign n14244 = \a[39]  & \b[11]  ;
  assign n14245 = n8748 & n14244 ;
  assign n14246 = \a[41]  & ~n14245 ;
  assign n14247 = ~n14243 & n14246 ;
  assign n14248 = n14242 & n14247 ;
  assign n14249 = n14237 & n14248 ;
  assign n14250 = ~n14243 & ~n14245 ;
  assign n14251 = n14242 & n14250 ;
  assign n14252 = n14237 & n14251 ;
  assign n14253 = ~\a[41]  & ~n14252 ;
  assign n14254 = ~n14249 & ~n14253 ;
  assign n14255 = ~n13134 & ~n13802 ;
  assign n14256 = ~n13136 & n14255 ;
  assign n14257 = ~n13803 & ~n14256 ;
  assign n14258 = n177 & n13125 ;
  assign n14259 = \b[3]  & n13123 ;
  assign n14260 = \a[47]  & \b[2]  ;
  assign n14261 = n13114 & n14260 ;
  assign n14262 = ~\a[48]  & \b[2]  ;
  assign n14263 = n13117 & n14262 ;
  assign n14264 = ~n14261 & ~n14263 ;
  assign n14265 = ~n14259 & n14264 ;
  assign n14266 = ~n14258 & n14265 ;
  assign n14267 = \b[1]  & n13794 ;
  assign n14268 = n13792 & n14267 ;
  assign n14269 = ~\a[50]  & ~n14268 ;
  assign n14270 = n14266 & n14269 ;
  assign n14271 = n14266 & ~n14268 ;
  assign n14272 = \a[50]  & ~n14271 ;
  assign n14273 = ~n14270 & ~n14272 ;
  assign n14274 = \a[50]  & ~\a[51]  ;
  assign n14275 = ~\a[50]  & \a[51]  ;
  assign n14276 = ~n14274 & ~n14275 ;
  assign n14277 = \b[0]  & ~n14276 ;
  assign n14278 = n13781 & n13798 ;
  assign n14279 = n14277 & n14278 ;
  assign n14280 = ~n14277 & ~n14278 ;
  assign n14281 = ~n14279 & ~n14280 ;
  assign n14282 = n14273 & n14281 ;
  assign n14283 = ~n14273 & ~n14281 ;
  assign n14284 = ~n14282 & ~n14283 ;
  assign n14285 = ~n323 & ~n10988 ;
  assign n14286 = ~n11569 & n14285 ;
  assign n14287 = n320 & n14286 ;
  assign n14288 = n323 & ~n10988 ;
  assign n14289 = ~n11569 & n14288 ;
  assign n14290 = ~n320 & n14289 ;
  assign n14291 = ~n14287 & ~n14290 ;
  assign n14292 = \b[4]  & n12159 ;
  assign n14293 = n12156 & n14292 ;
  assign n14294 = ~\a[45]  & \b[5]  ;
  assign n14295 = n11564 & n14294 ;
  assign n14296 = ~n14293 & ~n14295 ;
  assign n14297 = \b[6]  & n11570 ;
  assign n14298 = \a[45]  & \b[5]  ;
  assign n14299 = n11561 & n14298 ;
  assign n14300 = \a[47]  & ~n14299 ;
  assign n14301 = ~n14297 & n14300 ;
  assign n14302 = n14296 & n14301 ;
  assign n14303 = n14291 & n14302 ;
  assign n14304 = ~n14297 & ~n14299 ;
  assign n14305 = n14296 & n14304 ;
  assign n14306 = n14291 & n14305 ;
  assign n14307 = ~\a[47]  & ~n14306 ;
  assign n14308 = ~n14303 & ~n14307 ;
  assign n14309 = n14284 & ~n14308 ;
  assign n14310 = ~n14284 & n14308 ;
  assign n14311 = ~n14309 & ~n14310 ;
  assign n14312 = ~n14257 & ~n14311 ;
  assign n14313 = n14257 & n14311 ;
  assign n14314 = ~n14312 & ~n14313 ;
  assign n14315 = ~n589 & n10082 ;
  assign n14316 = ~n587 & n14315 ;
  assign n14317 = \b[7]  & n10681 ;
  assign n14318 = n10678 & n14317 ;
  assign n14319 = \b[9]  & n10080 ;
  assign n14320 = \a[41]  & \b[8]  ;
  assign n14321 = n10679 & n14320 ;
  assign n14322 = ~\a[42]  & \b[8]  ;
  assign n14323 = n10074 & n14322 ;
  assign n14324 = ~n14321 & ~n14323 ;
  assign n14325 = ~n14319 & n14324 ;
  assign n14326 = ~n14318 & n14325 ;
  assign n14327 = ~n14316 & n14326 ;
  assign n14328 = ~\a[44]  & ~n14327 ;
  assign n14329 = \a[44]  & n14326 ;
  assign n14330 = ~n14316 & n14329 ;
  assign n14331 = ~n14328 & ~n14330 ;
  assign n14332 = ~n14314 & n14331 ;
  assign n14333 = n14314 & ~n14331 ;
  assign n14334 = ~n14332 & ~n14333 ;
  assign n14335 = ~n14254 & ~n14334 ;
  assign n14336 = ~n14230 & n14335 ;
  assign n14337 = ~n14254 & n14334 ;
  assign n14338 = n14230 & n14337 ;
  assign n14339 = ~n14336 & ~n14338 ;
  assign n14340 = n14254 & ~n14334 ;
  assign n14341 = n14230 & n14340 ;
  assign n14342 = n14254 & n14334 ;
  assign n14343 = ~n14230 & n14342 ;
  assign n14344 = ~n14341 & ~n14343 ;
  assign n14345 = n14339 & n14344 ;
  assign n14346 = n14229 & ~n14345 ;
  assign n14347 = n14207 & n14346 ;
  assign n14348 = n14229 & n14345 ;
  assign n14349 = ~n14207 & n14348 ;
  assign n14350 = ~n14347 & ~n14349 ;
  assign n14351 = ~n14229 & ~n14345 ;
  assign n14352 = ~n14207 & n14351 ;
  assign n14353 = ~n14229 & n14345 ;
  assign n14354 = n14207 & n14353 ;
  assign n14355 = ~n14352 & ~n14354 ;
  assign n14356 = n14350 & n14355 ;
  assign n14357 = ~n14204 & n14356 ;
  assign n14358 = n1875 & n6309 ;
  assign n14359 = ~n1872 & n14358 ;
  assign n14360 = n5000 & n6309 ;
  assign n14361 = ~n1871 & n14360 ;
  assign n14362 = \b[16]  & n6778 ;
  assign n14363 = n6775 & n14362 ;
  assign n14364 = ~\a[33]  & \b[17]  ;
  assign n14365 = n6301 & n14364 ;
  assign n14366 = ~n14363 & ~n14365 ;
  assign n14367 = \b[18]  & n6307 ;
  assign n14368 = \a[33]  & \b[17]  ;
  assign n14369 = n6298 & n14368 ;
  assign n14370 = \a[35]  & ~n14369 ;
  assign n14371 = ~n14367 & n14370 ;
  assign n14372 = n14366 & n14371 ;
  assign n14373 = ~n14361 & n14372 ;
  assign n14374 = ~n14359 & n14373 ;
  assign n14375 = ~n14367 & ~n14369 ;
  assign n14376 = n14366 & n14375 ;
  assign n14377 = ~n14361 & n14376 ;
  assign n14378 = ~n14359 & n14377 ;
  assign n14379 = ~\a[35]  & ~n14378 ;
  assign n14380 = ~n14374 & ~n14379 ;
  assign n14381 = n13842 & ~n14356 ;
  assign n14382 = ~n14203 & n14381 ;
  assign n14383 = ~n14380 & ~n14382 ;
  assign n14384 = ~n14357 & n14383 ;
  assign n14385 = ~n14356 & n14380 ;
  assign n14386 = n14204 & n14385 ;
  assign n14387 = n14356 & n14380 ;
  assign n14388 = ~n14204 & n14387 ;
  assign n14389 = ~n14386 & ~n14388 ;
  assign n14390 = ~n14384 & n14389 ;
  assign n14391 = n14202 & n14390 ;
  assign n14392 = ~n14202 & ~n14390 ;
  assign n14393 = ~n14391 & ~n14392 ;
  assign n14394 = ~n2520 & n5211 ;
  assign n14395 = ~n2292 & n5211 ;
  assign n14396 = ~n2516 & n14395 ;
  assign n14397 = ~n14394 & ~n14396 ;
  assign n14398 = ~n2523 & ~n14397 ;
  assign n14399 = \b[19]  & n5595 ;
  assign n14400 = n5592 & n14399 ;
  assign n14401 = ~\a[30]  & \b[20]  ;
  assign n14402 = n5203 & n14401 ;
  assign n14403 = ~n14400 & ~n14402 ;
  assign n14404 = \b[21]  & n5209 ;
  assign n14405 = \a[30]  & \b[20]  ;
  assign n14406 = n5200 & n14405 ;
  assign n14407 = \a[32]  & ~n14406 ;
  assign n14408 = ~n14404 & n14407 ;
  assign n14409 = n14403 & n14408 ;
  assign n14410 = ~n14398 & n14409 ;
  assign n14411 = ~n14404 & ~n14406 ;
  assign n14412 = n14403 & n14411 ;
  assign n14413 = ~\a[32]  & ~n14412 ;
  assign n14414 = ~\a[32]  & ~n2523 ;
  assign n14415 = ~n14397 & n14414 ;
  assign n14416 = ~n14413 & ~n14415 ;
  assign n14417 = ~n14410 & n14416 ;
  assign n14418 = n14393 & ~n14417 ;
  assign n14419 = ~n14393 & n14417 ;
  assign n14420 = ~n14418 & ~n14419 ;
  assign n14421 = n3283 & n4249 ;
  assign n14422 = ~n3280 & n14421 ;
  assign n14423 = ~n3283 & n4249 ;
  assign n14424 = ~n3017 & n14423 ;
  assign n14425 = ~n3279 & n14424 ;
  assign n14426 = \b[22]  & n4647 ;
  assign n14427 = n4644 & n14426 ;
  assign n14428 = ~\a[27]  & \b[23]  ;
  assign n14429 = n4241 & n14428 ;
  assign n14430 = ~n14427 & ~n14429 ;
  assign n14431 = \b[24]  & n4247 ;
  assign n14432 = \a[27]  & \b[23]  ;
  assign n14433 = n4238 & n14432 ;
  assign n14434 = \a[29]  & ~n14433 ;
  assign n14435 = ~n14431 & n14434 ;
  assign n14436 = n14430 & n14435 ;
  assign n14437 = ~n14425 & n14436 ;
  assign n14438 = ~n14422 & n14437 ;
  assign n14439 = ~n14431 & ~n14433 ;
  assign n14440 = n14430 & n14439 ;
  assign n14441 = ~n14425 & n14440 ;
  assign n14442 = ~n14422 & n14441 ;
  assign n14443 = ~\a[29]  & ~n14442 ;
  assign n14444 = ~n14438 & ~n14443 ;
  assign n14445 = ~n14420 & n14444 ;
  assign n14446 = n14199 & n14445 ;
  assign n14447 = n14420 & n14444 ;
  assign n14448 = ~n14199 & n14447 ;
  assign n14449 = ~n14446 & ~n14448 ;
  assign n14450 = ~n14420 & ~n14444 ;
  assign n14451 = ~n14199 & n14450 ;
  assign n14452 = n14420 & ~n14444 ;
  assign n14453 = n14199 & n14452 ;
  assign n14454 = ~n14451 & ~n14453 ;
  assign n14455 = n14449 & n14454 ;
  assign n14456 = ~n14198 & ~n14455 ;
  assign n14457 = n13897 & n14455 ;
  assign n14458 = ~n14197 & n14457 ;
  assign n14459 = ~n3154 & ~n3399 ;
  assign n14460 = ~n4148 & n14459 ;
  assign n14461 = ~n4146 & n14460 ;
  assign n14462 = \b[25]  & n3733 ;
  assign n14463 = n3730 & n14462 ;
  assign n14464 = ~\a[24]  & \b[26]  ;
  assign n14465 = n3394 & n14464 ;
  assign n14466 = ~n14463 & ~n14465 ;
  assign n14467 = \b[27]  & n3400 ;
  assign n14468 = \a[24]  & \b[26]  ;
  assign n14469 = n3391 & n14468 ;
  assign n14470 = \a[26]  & ~n14469 ;
  assign n14471 = ~n14467 & n14470 ;
  assign n14472 = n14466 & n14471 ;
  assign n14473 = ~n14461 & n14472 ;
  assign n14474 = ~n14467 & ~n14469 ;
  assign n14475 = n14466 & n14474 ;
  assign n14476 = ~n14461 & n14475 ;
  assign n14477 = ~\a[26]  & ~n14476 ;
  assign n14478 = ~n14473 & ~n14477 ;
  assign n14479 = ~n14458 & ~n14478 ;
  assign n14480 = ~n14456 & n14479 ;
  assign n14481 = ~n14455 & n14478 ;
  assign n14482 = ~n14198 & n14481 ;
  assign n14483 = n14455 & n14478 ;
  assign n14484 = n14198 & n14483 ;
  assign n14485 = ~n14482 & ~n14484 ;
  assign n14486 = ~n14480 & n14485 ;
  assign n14487 = ~n14195 & ~n14486 ;
  assign n14488 = ~n14171 & n14487 ;
  assign n14489 = ~n14195 & n14486 ;
  assign n14490 = n14171 & n14489 ;
  assign n14491 = ~n14488 & ~n14490 ;
  assign n14492 = n14195 & ~n14486 ;
  assign n14493 = n14171 & n14492 ;
  assign n14494 = n14195 & n14486 ;
  assign n14495 = ~n14171 & n14494 ;
  assign n14496 = ~n14493 & ~n14495 ;
  assign n14497 = n14491 & n14496 ;
  assign n14498 = n1965 & ~n5855 ;
  assign n14499 = ~n5853 & n14498 ;
  assign n14500 = \b[33]  & n1963 ;
  assign n14501 = \a[18]  & \b[32]  ;
  assign n14502 = n2210 & n14501 ;
  assign n14503 = ~n14500 & ~n14502 ;
  assign n14504 = \b[31]  & n2218 ;
  assign n14505 = n2216 & n14504 ;
  assign n14506 = ~\a[18]  & \b[32]  ;
  assign n14507 = n1957 & n14506 ;
  assign n14508 = ~n14505 & ~n14507 ;
  assign n14509 = n14503 & n14508 ;
  assign n14510 = ~n14499 & n14509 ;
  assign n14511 = ~\a[20]  & ~n14510 ;
  assign n14512 = \a[20]  & n14509 ;
  assign n14513 = ~n14499 & n14512 ;
  assign n14514 = ~n14511 & ~n14513 ;
  assign n14515 = ~n14497 & ~n14514 ;
  assign n14516 = n14170 & n14515 ;
  assign n14517 = n14497 & ~n14514 ;
  assign n14518 = ~n14170 & n14517 ;
  assign n14519 = ~n14516 & ~n14518 ;
  assign n14520 = ~n14497 & n14514 ;
  assign n14521 = ~n14170 & n14520 ;
  assign n14522 = n14497 & n14514 ;
  assign n14523 = n14170 & n14522 ;
  assign n14524 = ~n14521 & ~n14523 ;
  assign n14525 = n14519 & n14524 ;
  assign n14526 = ~n14167 & ~n14525 ;
  assign n14527 = ~n14143 & n14526 ;
  assign n14528 = ~n14167 & n14525 ;
  assign n14529 = n14143 & n14528 ;
  assign n14530 = ~n14527 & ~n14529 ;
  assign n14531 = n14167 & ~n14525 ;
  assign n14532 = n14143 & n14531 ;
  assign n14533 = n14167 & n14525 ;
  assign n14534 = ~n14143 & n14533 ;
  assign n14535 = ~n14532 & ~n14534 ;
  assign n14536 = n14530 & n14535 ;
  assign n14537 = ~n14142 & ~n14536 ;
  assign n14538 = ~n13948 & n14536 ;
  assign n14539 = ~n14141 & n14538 ;
  assign n14540 = n999 & ~n8602 ;
  assign n14541 = ~n8600 & n14540 ;
  assign n14542 = \b[37]  & n1182 ;
  assign n14543 = n1179 & n14542 ;
  assign n14544 = \b[39]  & n997 ;
  assign n14545 = \a[11]  & \b[38]  ;
  assign n14546 = n1180 & n14545 ;
  assign n14547 = ~\a[12]  & \b[38]  ;
  assign n14548 = n7674 & n14547 ;
  assign n14549 = ~n14546 & ~n14548 ;
  assign n14550 = ~n14544 & n14549 ;
  assign n14551 = ~n14543 & n14550 ;
  assign n14552 = ~n14541 & n14551 ;
  assign n14553 = ~\a[14]  & ~n14552 ;
  assign n14554 = \a[14]  & n14551 ;
  assign n14555 = ~n14541 & n14554 ;
  assign n14556 = ~n14553 & ~n14555 ;
  assign n14557 = ~n14539 & ~n14556 ;
  assign n14558 = ~n14537 & n14557 ;
  assign n14559 = ~n14536 & n14556 ;
  assign n14560 = ~n14142 & n14559 ;
  assign n14561 = n14536 & n14556 ;
  assign n14562 = n14142 & n14561 ;
  assign n14563 = ~n14560 & ~n14562 ;
  assign n14564 = ~n14558 & n14563 ;
  assign n14565 = n646 & n9930 ;
  assign n14566 = ~n9927 & n14565 ;
  assign n14567 = n646 & ~n9930 ;
  assign n14568 = ~n9477 & n14567 ;
  assign n14569 = ~n9926 & n14568 ;
  assign n14570 = \b[40]  & n796 ;
  assign n14571 = n793 & n14570 ;
  assign n14572 = ~\a[9]  & \b[41]  ;
  assign n14573 = n638 & n14572 ;
  assign n14574 = ~n14571 & ~n14573 ;
  assign n14575 = \b[42]  & n644 ;
  assign n14576 = \a[9]  & \b[41]  ;
  assign n14577 = n635 & n14576 ;
  assign n14578 = \a[11]  & ~n14577 ;
  assign n14579 = ~n14575 & n14578 ;
  assign n14580 = n14574 & n14579 ;
  assign n14581 = ~n14569 & n14580 ;
  assign n14582 = ~n14566 & n14581 ;
  assign n14583 = ~n14575 & ~n14577 ;
  assign n14584 = n14574 & n14583 ;
  assign n14585 = ~n14569 & n14584 ;
  assign n14586 = ~n14566 & n14585 ;
  assign n14587 = ~\a[11]  & ~n14586 ;
  assign n14588 = ~n14582 & ~n14587 ;
  assign n14589 = ~n14564 & n14588 ;
  assign n14590 = n14139 & n14589 ;
  assign n14591 = n14564 & n14588 ;
  assign n14592 = ~n14139 & n14591 ;
  assign n14593 = ~n14590 & ~n14592 ;
  assign n14594 = ~n14139 & n14564 ;
  assign n14595 = ~n13976 & ~n14564 ;
  assign n14596 = ~n14138 & n14595 ;
  assign n14597 = ~n14588 & ~n14596 ;
  assign n14598 = ~n14594 & n14597 ;
  assign n14599 = n14593 & ~n14598 ;
  assign n14600 = ~n13446 & n14004 ;
  assign n14601 = n14009 & ~n14600 ;
  assign n14602 = n13452 & n14009 ;
  assign n14603 = n13002 & n14602 ;
  assign n14604 = ~n14601 & ~n14603 ;
  assign n14605 = n14599 & ~n14604 ;
  assign n14606 = ~n14599 & n14604 ;
  assign n14607 = ~n14605 & ~n14606 ;
  assign n14608 = n430 & ~n11397 ;
  assign n14609 = ~n11395 & n14608 ;
  assign n14610 = \b[45]  & n428 ;
  assign n14611 = \a[6]  & \b[44]  ;
  assign n14612 = n419 & n14611 ;
  assign n14613 = ~n14610 & ~n14612 ;
  assign n14614 = \b[43]  & n486 ;
  assign n14615 = n483 & n14614 ;
  assign n14616 = ~\a[6]  & \b[44]  ;
  assign n14617 = n422 & n14616 ;
  assign n14618 = ~n14615 & ~n14617 ;
  assign n14619 = n14613 & n14618 ;
  assign n14620 = ~n14609 & n14619 ;
  assign n14621 = ~\a[8]  & ~n14620 ;
  assign n14622 = \a[8]  & n14619 ;
  assign n14623 = ~n14609 & n14622 ;
  assign n14624 = ~n14621 & ~n14623 ;
  assign n14625 = n14607 & ~n14624 ;
  assign n14626 = ~n14607 & n14624 ;
  assign n14627 = ~n14625 & ~n14626 ;
  assign n14628 = n14137 & ~n14627 ;
  assign n14629 = n14113 & n14628 ;
  assign n14630 = n14137 & n14627 ;
  assign n14631 = ~n14113 & n14630 ;
  assign n14632 = ~n14629 & ~n14631 ;
  assign n14633 = ~n14137 & ~n14627 ;
  assign n14634 = ~n14113 & n14633 ;
  assign n14635 = ~n14137 & n14627 ;
  assign n14636 = n14113 & n14635 ;
  assign n14637 = ~n14634 & ~n14636 ;
  assign n14638 = n14632 & n14637 ;
  assign n14639 = ~n14112 & ~n14638 ;
  assign n14640 = n14089 & n14639 ;
  assign n14641 = ~n14112 & n14638 ;
  assign n14642 = ~n14089 & n14641 ;
  assign n14643 = ~n14640 & ~n14642 ;
  assign n14644 = n14112 & ~n14638 ;
  assign n14645 = ~n14089 & n14644 ;
  assign n14646 = n14112 & n14638 ;
  assign n14647 = n14089 & n14646 ;
  assign n14648 = ~n14645 & ~n14647 ;
  assign n14649 = n14643 & n14648 ;
  assign n14650 = ~n14086 & n14649 ;
  assign n14651 = n14076 & ~n14649 ;
  assign n14652 = ~n14083 & n14651 ;
  assign n14653 = ~n14650 & ~n14652 ;
  assign n14654 = n14076 & n14643 ;
  assign n14655 = ~n14083 & n14654 ;
  assign n14656 = n14648 & ~n14655 ;
  assign n14657 = n14089 & n14638 ;
  assign n14658 = n14637 & ~n14657 ;
  assign n14659 = ~n14034 & ~n14625 ;
  assign n14660 = ~n14041 & n14659 ;
  assign n14661 = ~n14626 & ~n14660 ;
  assign n14662 = ~n14598 & ~n14605 ;
  assign n14663 = n430 & n11906 ;
  assign n14664 = ~n11903 & n14663 ;
  assign n14665 = n430 & n13483 ;
  assign n14666 = ~n11902 & n14665 ;
  assign n14667 = \b[44]  & n486 ;
  assign n14668 = n483 & n14667 ;
  assign n14669 = ~\a[6]  & \b[45]  ;
  assign n14670 = n422 & n14669 ;
  assign n14671 = ~n14668 & ~n14670 ;
  assign n14672 = \b[46]  & n428 ;
  assign n14673 = \a[6]  & \b[45]  ;
  assign n14674 = n419 & n14673 ;
  assign n14675 = \a[8]  & ~n14674 ;
  assign n14676 = ~n14672 & n14675 ;
  assign n14677 = n14671 & n14676 ;
  assign n14678 = ~n14666 & n14677 ;
  assign n14679 = ~n14664 & n14678 ;
  assign n14680 = ~n14672 & ~n14674 ;
  assign n14681 = n14671 & n14680 ;
  assign n14682 = ~n14666 & n14681 ;
  assign n14683 = ~n14664 & n14682 ;
  assign n14684 = ~\a[8]  & ~n14683 ;
  assign n14685 = ~n14679 & ~n14684 ;
  assign n14686 = ~n13976 & ~n14558 ;
  assign n14687 = ~n14138 & n14686 ;
  assign n14688 = n14563 & ~n14687 ;
  assign n14689 = n14530 & ~n14539 ;
  assign n14690 = n13925 & n14519 ;
  assign n14691 = ~n13927 & n14690 ;
  assign n14692 = n14524 & ~n14691 ;
  assign n14693 = n14170 & n14497 ;
  assign n14694 = n14491 & ~n14693 ;
  assign n14695 = ~n13908 & ~n14480 ;
  assign n14696 = ~n13910 & n14695 ;
  assign n14697 = n14485 & ~n14696 ;
  assign n14698 = n14454 & ~n14458 ;
  assign n14699 = n13864 & ~n14418 ;
  assign n14700 = ~n13873 & n14699 ;
  assign n14701 = ~n14419 & ~n14700 ;
  assign n14702 = ~n14384 & ~n14391 ;
  assign n14703 = n2768 & n5211 ;
  assign n14704 = ~n2765 & n14703 ;
  assign n14705 = n5211 & n6462 ;
  assign n14706 = ~n2764 & n14705 ;
  assign n14707 = \b[20]  & n5595 ;
  assign n14708 = n5592 & n14707 ;
  assign n14709 = ~\a[30]  & \b[21]  ;
  assign n14710 = n5203 & n14709 ;
  assign n14711 = ~n14708 & ~n14710 ;
  assign n14712 = \b[22]  & n5209 ;
  assign n14713 = \a[30]  & \b[21]  ;
  assign n14714 = n5200 & n14713 ;
  assign n14715 = \a[32]  & ~n14714 ;
  assign n14716 = ~n14712 & n14715 ;
  assign n14717 = n14711 & n14716 ;
  assign n14718 = ~n14706 & n14717 ;
  assign n14719 = ~n14704 & n14718 ;
  assign n14720 = ~n14712 & ~n14714 ;
  assign n14721 = n14711 & n14720 ;
  assign n14722 = ~n14706 & n14721 ;
  assign n14723 = ~n14704 & n14722 ;
  assign n14724 = ~\a[32]  & ~n14723 ;
  assign n14725 = ~n14719 & ~n14724 ;
  assign n14726 = n13842 & n14350 ;
  assign n14727 = n14355 & ~n14726 ;
  assign n14728 = n13848 & n14355 ;
  assign n14729 = n13692 & n14728 ;
  assign n14730 = ~n14727 & ~n14729 ;
  assign n14731 = n14207 & n14345 ;
  assign n14732 = n14339 & ~n14731 ;
  assign n14733 = ~n13808 & ~n14333 ;
  assign n14734 = ~n13811 & n14733 ;
  assign n14735 = ~n14332 & ~n14734 ;
  assign n14736 = ~n948 & n8759 ;
  assign n14737 = ~n908 & n8759 ;
  assign n14738 = ~n912 & n14737 ;
  assign n14739 = ~n14736 & ~n14738 ;
  assign n14740 = ~n951 & ~n14739 ;
  assign n14741 = \b[11]  & n9301 ;
  assign n14742 = n9298 & n14741 ;
  assign n14743 = ~\a[39]  & \b[12]  ;
  assign n14744 = n8751 & n14743 ;
  assign n14745 = ~n14742 & ~n14744 ;
  assign n14746 = \b[13]  & n8757 ;
  assign n14747 = \a[39]  & \b[12]  ;
  assign n14748 = n8748 & n14747 ;
  assign n14749 = \a[41]  & ~n14748 ;
  assign n14750 = ~n14746 & n14749 ;
  assign n14751 = n14745 & n14750 ;
  assign n14752 = ~n14740 & n14751 ;
  assign n14753 = ~n14746 & ~n14748 ;
  assign n14754 = n14745 & n14753 ;
  assign n14755 = ~\a[41]  & ~n14754 ;
  assign n14756 = ~\a[41]  & ~n951 ;
  assign n14757 = ~n14739 & n14756 ;
  assign n14758 = ~n14755 & ~n14757 ;
  assign n14759 = ~n14752 & n14758 ;
  assign n14760 = ~n14309 & ~n14313 ;
  assign n14761 = ~n14279 & ~n14282 ;
  assign n14762 = n222 & n13125 ;
  assign n14763 = \b[4]  & n13123 ;
  assign n14764 = \a[47]  & \b[3]  ;
  assign n14765 = n13114 & n14764 ;
  assign n14766 = ~\a[48]  & \b[3]  ;
  assign n14767 = n13117 & n14766 ;
  assign n14768 = ~n14765 & ~n14767 ;
  assign n14769 = ~n14763 & n14768 ;
  assign n14770 = \b[2]  & n13794 ;
  assign n14771 = n13792 & n14770 ;
  assign n14772 = \a[50]  & ~n14771 ;
  assign n14773 = n14769 & n14772 ;
  assign n14774 = ~n14762 & n14773 ;
  assign n14775 = n14769 & ~n14771 ;
  assign n14776 = ~n14762 & n14775 ;
  assign n14777 = ~\a[50]  & ~n14776 ;
  assign n14778 = ~n14774 & ~n14777 ;
  assign n14779 = \a[53]  & \b[0]  ;
  assign n14780 = ~n14276 & n14779 ;
  assign n14781 = \a[51]  & \b[0]  ;
  assign n14782 = \a[50]  & ~\a[52]  ;
  assign n14783 = n14781 & n14782 ;
  assign n14784 = ~\a[51]  & \b[0]  ;
  assign n14785 = ~\a[50]  & \a[52]  ;
  assign n14786 = n14784 & n14785 ;
  assign n14787 = ~n14783 & ~n14786 ;
  assign n14788 = \a[52]  & ~\a[53]  ;
  assign n14789 = ~\a[52]  & \a[53]  ;
  assign n14790 = ~n14788 & ~n14789 ;
  assign n14791 = ~n14276 & n14790 ;
  assign n14792 = \b[1]  & n14791 ;
  assign n14793 = ~n14276 & ~n14790 ;
  assign n14794 = ~n137 & n14793 ;
  assign n14795 = ~n14792 & ~n14794 ;
  assign n14796 = n14787 & n14795 ;
  assign n14797 = n14780 & ~n14796 ;
  assign n14798 = ~n14780 & n14787 ;
  assign n14799 = n14795 & n14798 ;
  assign n14800 = ~n14797 & ~n14799 ;
  assign n14801 = n14778 & ~n14800 ;
  assign n14802 = ~n14778 & n14800 ;
  assign n14803 = ~n14801 & ~n14802 ;
  assign n14804 = ~n14761 & n14803 ;
  assign n14805 = n14761 & ~n14803 ;
  assign n14806 = ~n14804 & ~n14805 ;
  assign n14807 = ~n383 & n11572 ;
  assign n14808 = ~n381 & n14807 ;
  assign n14809 = \b[5]  & n12159 ;
  assign n14810 = n12156 & n14809 ;
  assign n14811 = ~\a[45]  & \b[6]  ;
  assign n14812 = n11564 & n14811 ;
  assign n14813 = ~n14810 & ~n14812 ;
  assign n14814 = \b[7]  & n11570 ;
  assign n14815 = \a[45]  & \b[6]  ;
  assign n14816 = n11561 & n14815 ;
  assign n14817 = \a[47]  & ~n14816 ;
  assign n14818 = ~n14814 & n14817 ;
  assign n14819 = n14813 & n14818 ;
  assign n14820 = ~n14808 & n14819 ;
  assign n14821 = ~n14814 & ~n14816 ;
  assign n14822 = n14813 & n14821 ;
  assign n14823 = ~n14808 & n14822 ;
  assign n14824 = ~\a[47]  & ~n14823 ;
  assign n14825 = ~n14820 & ~n14824 ;
  assign n14826 = n14806 & ~n14825 ;
  assign n14827 = ~n14806 & n14825 ;
  assign n14828 = ~n14826 & ~n14827 ;
  assign n14829 = n685 & n10082 ;
  assign n14830 = ~n682 & n14829 ;
  assign n14831 = ~n685 & n10082 ;
  assign n14832 = ~n584 & n14831 ;
  assign n14833 = ~n681 & n14832 ;
  assign n14834 = \b[8]  & n10681 ;
  assign n14835 = n10678 & n14834 ;
  assign n14836 = \b[10]  & n10080 ;
  assign n14837 = \a[41]  & \b[9]  ;
  assign n14838 = n10679 & n14837 ;
  assign n14839 = ~\a[42]  & \b[9]  ;
  assign n14840 = n10074 & n14839 ;
  assign n14841 = ~n14838 & ~n14840 ;
  assign n14842 = ~n14836 & n14841 ;
  assign n14843 = ~n14835 & n14842 ;
  assign n14844 = ~n14833 & n14843 ;
  assign n14845 = ~n14830 & n14844 ;
  assign n14846 = ~\a[44]  & ~n14845 ;
  assign n14847 = \a[44]  & n14843 ;
  assign n14848 = ~n14833 & n14847 ;
  assign n14849 = ~n14830 & n14848 ;
  assign n14850 = ~n14846 & ~n14849 ;
  assign n14851 = ~n14828 & ~n14850 ;
  assign n14852 = ~n14760 & n14851 ;
  assign n14853 = n14828 & ~n14850 ;
  assign n14854 = n14760 & n14853 ;
  assign n14855 = ~n14852 & ~n14854 ;
  assign n14856 = ~n14828 & n14850 ;
  assign n14857 = n14760 & n14856 ;
  assign n14858 = n14828 & n14850 ;
  assign n14859 = ~n14760 & n14858 ;
  assign n14860 = ~n14857 & ~n14859 ;
  assign n14861 = n14855 & n14860 ;
  assign n14862 = n14759 & ~n14861 ;
  assign n14863 = ~n14735 & n14862 ;
  assign n14864 = n14759 & n14861 ;
  assign n14865 = n14735 & n14864 ;
  assign n14866 = ~n14863 & ~n14865 ;
  assign n14867 = ~n14759 & ~n14861 ;
  assign n14868 = n14735 & n14867 ;
  assign n14869 = ~n14759 & n14861 ;
  assign n14870 = ~n14735 & n14869 ;
  assign n14871 = ~n14868 & ~n14870 ;
  assign n14872 = n14866 & n14871 ;
  assign n14873 = ~n14732 & n14872 ;
  assign n14874 = n14339 & ~n14872 ;
  assign n14875 = ~n14731 & n14874 ;
  assign n14876 = n1512 & n7534 ;
  assign n14877 = ~n1509 & n14876 ;
  assign n14878 = n7534 & n10165 ;
  assign n14879 = ~n1508 & n14878 ;
  assign n14880 = \b[14]  & n7973 ;
  assign n14881 = n7970 & n14880 ;
  assign n14882 = \b[16]  & n7532 ;
  assign n14883 = \a[36]  & \b[15]  ;
  assign n14884 = n7523 & n14883 ;
  assign n14885 = ~\a[36]  & \b[15]  ;
  assign n14886 = n7526 & n14885 ;
  assign n14887 = ~n14884 & ~n14886 ;
  assign n14888 = ~n14882 & n14887 ;
  assign n14889 = ~n14881 & n14888 ;
  assign n14890 = ~n14879 & n14889 ;
  assign n14891 = ~n14877 & n14890 ;
  assign n14892 = ~\a[38]  & ~n14891 ;
  assign n14893 = \a[38]  & n14889 ;
  assign n14894 = ~n14879 & n14893 ;
  assign n14895 = ~n14877 & n14894 ;
  assign n14896 = ~n14892 & ~n14895 ;
  assign n14897 = ~n14875 & ~n14896 ;
  assign n14898 = ~n14873 & n14897 ;
  assign n14899 = ~n14872 & n14896 ;
  assign n14900 = n14732 & n14899 ;
  assign n14901 = n14872 & n14896 ;
  assign n14902 = ~n14732 & n14901 ;
  assign n14903 = ~n14900 & ~n14902 ;
  assign n14904 = ~n14898 & n14903 ;
  assign n14905 = n14730 & ~n14904 ;
  assign n14906 = ~n14730 & n14904 ;
  assign n14907 = ~n14905 & ~n14906 ;
  assign n14908 = ~n2076 & n6309 ;
  assign n14909 = ~n1874 & n6309 ;
  assign n14910 = ~n1878 & n14909 ;
  assign n14911 = ~n14908 & ~n14910 ;
  assign n14912 = ~n2079 & ~n14911 ;
  assign n14913 = \b[17]  & n6778 ;
  assign n14914 = n6775 & n14913 ;
  assign n14915 = ~\a[33]  & \b[18]  ;
  assign n14916 = n6301 & n14915 ;
  assign n14917 = ~n14914 & ~n14916 ;
  assign n14918 = \b[19]  & n6307 ;
  assign n14919 = \a[33]  & \b[18]  ;
  assign n14920 = n6298 & n14919 ;
  assign n14921 = \a[35]  & ~n14920 ;
  assign n14922 = ~n14918 & n14921 ;
  assign n14923 = n14917 & n14922 ;
  assign n14924 = ~n14912 & n14923 ;
  assign n14925 = ~n14918 & ~n14920 ;
  assign n14926 = n14917 & n14925 ;
  assign n14927 = ~\a[35]  & ~n14926 ;
  assign n14928 = ~\a[35]  & ~n2079 ;
  assign n14929 = ~n14911 & n14928 ;
  assign n14930 = ~n14927 & ~n14929 ;
  assign n14931 = ~n14924 & n14930 ;
  assign n14932 = n14907 & ~n14931 ;
  assign n14933 = ~n14907 & n14931 ;
  assign n14934 = ~n14932 & ~n14933 ;
  assign n14935 = ~n14725 & ~n14934 ;
  assign n14936 = ~n14702 & n14935 ;
  assign n14937 = ~n14725 & n14934 ;
  assign n14938 = n14702 & n14937 ;
  assign n14939 = ~n14936 & ~n14938 ;
  assign n14940 = n14725 & ~n14934 ;
  assign n14941 = n14702 & n14940 ;
  assign n14942 = n14725 & n14934 ;
  assign n14943 = ~n14702 & n14942 ;
  assign n14944 = ~n14941 & ~n14943 ;
  assign n14945 = n14939 & n14944 ;
  assign n14946 = ~n3567 & n4249 ;
  assign n14947 = ~n3565 & n14946 ;
  assign n14948 = \b[25]  & n4247 ;
  assign n14949 = \a[27]  & \b[24]  ;
  assign n14950 = n4238 & n14949 ;
  assign n14951 = ~n14948 & ~n14950 ;
  assign n14952 = \b[23]  & n4647 ;
  assign n14953 = n4644 & n14952 ;
  assign n14954 = ~\a[27]  & \b[24]  ;
  assign n14955 = n4241 & n14954 ;
  assign n14956 = ~n14953 & ~n14955 ;
  assign n14957 = n14951 & n14956 ;
  assign n14958 = ~n14947 & n14957 ;
  assign n14959 = ~\a[29]  & ~n14958 ;
  assign n14960 = \a[29]  & n14957 ;
  assign n14961 = ~n14947 & n14960 ;
  assign n14962 = ~n14959 & ~n14961 ;
  assign n14963 = ~n14945 & ~n14962 ;
  assign n14964 = n14701 & n14963 ;
  assign n14965 = n14945 & ~n14962 ;
  assign n14966 = ~n14701 & n14965 ;
  assign n14967 = ~n14964 & ~n14966 ;
  assign n14968 = ~n14945 & n14962 ;
  assign n14969 = ~n14701 & n14968 ;
  assign n14970 = n14945 & n14962 ;
  assign n14971 = n14701 & n14970 ;
  assign n14972 = ~n14969 & ~n14971 ;
  assign n14973 = n14967 & n14972 ;
  assign n14974 = ~n14698 & n14973 ;
  assign n14975 = n3402 & n4456 ;
  assign n14976 = ~n4453 & n14975 ;
  assign n14977 = n3402 & ~n4456 ;
  assign n14978 = ~n4143 & n14977 ;
  assign n14979 = ~n4452 & n14978 ;
  assign n14980 = \b[26]  & n3733 ;
  assign n14981 = n3730 & n14980 ;
  assign n14982 = ~\a[24]  & \b[27]  ;
  assign n14983 = n3394 & n14982 ;
  assign n14984 = ~n14981 & ~n14983 ;
  assign n14985 = \b[28]  & n3400 ;
  assign n14986 = \a[24]  & \b[27]  ;
  assign n14987 = n3391 & n14986 ;
  assign n14988 = \a[26]  & ~n14987 ;
  assign n14989 = ~n14985 & n14988 ;
  assign n14990 = n14984 & n14989 ;
  assign n14991 = ~n14979 & n14990 ;
  assign n14992 = ~n14976 & n14991 ;
  assign n14993 = ~n14985 & ~n14987 ;
  assign n14994 = n14984 & n14993 ;
  assign n14995 = ~n14979 & n14994 ;
  assign n14996 = ~n14976 & n14995 ;
  assign n14997 = ~\a[26]  & ~n14996 ;
  assign n14998 = ~n14992 & ~n14997 ;
  assign n14999 = n14454 & ~n14973 ;
  assign n15000 = ~n14458 & n14999 ;
  assign n15001 = ~n14998 & ~n15000 ;
  assign n15002 = ~n14974 & n15001 ;
  assign n15003 = ~n14973 & n14998 ;
  assign n15004 = n14698 & n15003 ;
  assign n15005 = n14973 & n14998 ;
  assign n15006 = ~n14698 & n15005 ;
  assign n15007 = ~n15004 & ~n15006 ;
  assign n15008 = ~n15002 & n15007 ;
  assign n15009 = n2622 & ~n5462 ;
  assign n15010 = ~n5460 & n15009 ;
  assign n15011 = \b[31]  & n2620 ;
  assign n15012 = \a[21]  & \b[30]  ;
  assign n15013 = n2611 & n15012 ;
  assign n15014 = ~n15011 & ~n15013 ;
  assign n15015 = \b[29]  & n2912 ;
  assign n15016 = n2909 & n15015 ;
  assign n15017 = ~\a[21]  & \b[30]  ;
  assign n15018 = n2614 & n15017 ;
  assign n15019 = ~n15016 & ~n15018 ;
  assign n15020 = n15014 & n15019 ;
  assign n15021 = ~n15010 & n15020 ;
  assign n15022 = ~\a[23]  & ~n15021 ;
  assign n15023 = \a[23]  & n15020 ;
  assign n15024 = ~n15010 & n15023 ;
  assign n15025 = ~n15022 & ~n15024 ;
  assign n15026 = ~n15008 & ~n15025 ;
  assign n15027 = n14697 & n15026 ;
  assign n15028 = n15008 & ~n15025 ;
  assign n15029 = ~n14697 & n15028 ;
  assign n15030 = ~n15027 & ~n15029 ;
  assign n15031 = ~n15008 & n15025 ;
  assign n15032 = ~n14697 & n15031 ;
  assign n15033 = n15008 & n15025 ;
  assign n15034 = n14697 & n15033 ;
  assign n15035 = ~n15032 & ~n15034 ;
  assign n15036 = n15030 & n15035 ;
  assign n15037 = ~n14694 & n15036 ;
  assign n15038 = n14491 & ~n15036 ;
  assign n15039 = ~n14693 & n15038 ;
  assign n15040 = n1965 & n6565 ;
  assign n15041 = ~n6562 & n15040 ;
  assign n15042 = n1965 & ~n6565 ;
  assign n15043 = ~n5850 & n15042 ;
  assign n15044 = ~n6561 & n15043 ;
  assign n15045 = \b[32]  & n2218 ;
  assign n15046 = n2216 & n15045 ;
  assign n15047 = ~\a[18]  & \b[33]  ;
  assign n15048 = n1957 & n15047 ;
  assign n15049 = ~n15046 & ~n15048 ;
  assign n15050 = \b[34]  & n1963 ;
  assign n15051 = \a[18]  & \b[33]  ;
  assign n15052 = n2210 & n15051 ;
  assign n15053 = \a[20]  & ~n15052 ;
  assign n15054 = ~n15050 & n15053 ;
  assign n15055 = n15049 & n15054 ;
  assign n15056 = ~n15044 & n15055 ;
  assign n15057 = ~n15041 & n15056 ;
  assign n15058 = ~n15050 & ~n15052 ;
  assign n15059 = n15049 & n15058 ;
  assign n15060 = ~n15044 & n15059 ;
  assign n15061 = ~n15041 & n15060 ;
  assign n15062 = ~\a[20]  & ~n15061 ;
  assign n15063 = ~n15057 & ~n15062 ;
  assign n15064 = ~n15039 & ~n15063 ;
  assign n15065 = ~n15037 & n15064 ;
  assign n15066 = ~n15036 & n15063 ;
  assign n15067 = n14694 & n15066 ;
  assign n15068 = n15036 & n15063 ;
  assign n15069 = ~n14694 & n15068 ;
  assign n15070 = ~n15067 & ~n15069 ;
  assign n15071 = ~n15065 & n15070 ;
  assign n15072 = ~n14692 & ~n15071 ;
  assign n15073 = n14692 & n15071 ;
  assign n15074 = ~n15072 & ~n15073 ;
  assign n15075 = n1467 & ~n7761 ;
  assign n15076 = ~n7759 & n15075 ;
  assign n15077 = \b[37]  & n1465 ;
  assign n15078 = \a[15]  & \b[36]  ;
  assign n15079 = n1456 & n15078 ;
  assign n15080 = ~n15077 & ~n15079 ;
  assign n15081 = \b[35]  & n1652 ;
  assign n15082 = n1649 & n15081 ;
  assign n15083 = ~\a[15]  & \b[36]  ;
  assign n15084 = n1459 & n15083 ;
  assign n15085 = ~n15082 & ~n15084 ;
  assign n15086 = n15080 & n15085 ;
  assign n15087 = ~n15076 & n15086 ;
  assign n15088 = ~\a[17]  & ~n15087 ;
  assign n15089 = \a[17]  & n15086 ;
  assign n15090 = ~n15076 & n15089 ;
  assign n15091 = ~n15088 & ~n15090 ;
  assign n15092 = n15074 & ~n15091 ;
  assign n15093 = ~n15074 & n15091 ;
  assign n15094 = ~n15092 & ~n15093 ;
  assign n15095 = n999 & n9044 ;
  assign n15096 = ~n9041 & n15095 ;
  assign n15097 = n999 & ~n9044 ;
  assign n15098 = ~n8597 & n15097 ;
  assign n15099 = ~n9040 & n15098 ;
  assign n15100 = \b[38]  & n1182 ;
  assign n15101 = n1179 & n15100 ;
  assign n15102 = \b[40]  & n997 ;
  assign n15103 = \a[11]  & \b[39]  ;
  assign n15104 = n1180 & n15103 ;
  assign n15105 = ~\a[12]  & \b[39]  ;
  assign n15106 = n7674 & n15105 ;
  assign n15107 = ~n15104 & ~n15106 ;
  assign n15108 = ~n15102 & n15107 ;
  assign n15109 = ~n15101 & n15108 ;
  assign n15110 = ~n15099 & n15109 ;
  assign n15111 = ~n15096 & n15110 ;
  assign n15112 = ~\a[14]  & ~n15111 ;
  assign n15113 = \a[14]  & n15109 ;
  assign n15114 = ~n15099 & n15113 ;
  assign n15115 = ~n15096 & n15114 ;
  assign n15116 = ~n15112 & ~n15115 ;
  assign n15117 = ~n15094 & ~n15116 ;
  assign n15118 = ~n14689 & n15117 ;
  assign n15119 = n15094 & ~n15116 ;
  assign n15120 = n14689 & n15119 ;
  assign n15121 = ~n15118 & ~n15120 ;
  assign n15122 = ~n15094 & n15116 ;
  assign n15123 = n14689 & n15122 ;
  assign n15124 = n15094 & n15116 ;
  assign n15125 = ~n14689 & n15124 ;
  assign n15126 = ~n15123 & ~n15125 ;
  assign n15127 = n15121 & n15126 ;
  assign n15128 = ~n14688 & ~n15127 ;
  assign n15129 = n14563 & n15127 ;
  assign n15130 = ~n14687 & n15129 ;
  assign n15131 = n646 & ~n10409 ;
  assign n15132 = ~n10407 & n15131 ;
  assign n15133 = \b[43]  & n644 ;
  assign n15134 = \a[9]  & \b[42]  ;
  assign n15135 = n635 & n15134 ;
  assign n15136 = ~n15133 & ~n15135 ;
  assign n15137 = \b[41]  & n796 ;
  assign n15138 = n793 & n15137 ;
  assign n15139 = ~\a[9]  & \b[42]  ;
  assign n15140 = n638 & n15139 ;
  assign n15141 = ~n15138 & ~n15140 ;
  assign n15142 = n15136 & n15141 ;
  assign n15143 = ~n15132 & n15142 ;
  assign n15144 = ~\a[11]  & ~n15143 ;
  assign n15145 = \a[11]  & n15142 ;
  assign n15146 = ~n15132 & n15145 ;
  assign n15147 = ~n15144 & ~n15146 ;
  assign n15148 = ~n15130 & ~n15147 ;
  assign n15149 = ~n15128 & n15148 ;
  assign n15150 = ~n15127 & n15147 ;
  assign n15151 = ~n14688 & n15150 ;
  assign n15152 = n15127 & n15147 ;
  assign n15153 = n14688 & n15152 ;
  assign n15154 = ~n15151 & ~n15153 ;
  assign n15155 = ~n15149 & n15154 ;
  assign n15156 = ~n14685 & ~n15155 ;
  assign n15157 = ~n14662 & n15156 ;
  assign n15158 = ~n14685 & n15155 ;
  assign n15159 = n14662 & n15158 ;
  assign n15160 = ~n15157 & ~n15159 ;
  assign n15161 = n14685 & ~n15155 ;
  assign n15162 = n14662 & n15161 ;
  assign n15163 = n14685 & n15155 ;
  assign n15164 = ~n14662 & n15163 ;
  assign n15165 = ~n15162 & ~n15164 ;
  assign n15166 = n15160 & n15165 ;
  assign n15167 = n252 & ~n13524 ;
  assign n15168 = ~n13522 & n15167 ;
  assign n15169 = \b[49]  & n250 ;
  assign n15170 = \a[3]  & \b[48]  ;
  assign n15171 = n241 & n15170 ;
  assign n15172 = ~n15169 & ~n15171 ;
  assign n15173 = \b[47]  & n303 ;
  assign n15174 = n300 & n15173 ;
  assign n15175 = ~\a[3]  & \b[48]  ;
  assign n15176 = n244 & n15175 ;
  assign n15177 = ~n15174 & ~n15176 ;
  assign n15178 = n15172 & n15177 ;
  assign n15179 = ~n15168 & n15178 ;
  assign n15180 = ~\a[5]  & ~n15179 ;
  assign n15181 = \a[5]  & n15178 ;
  assign n15182 = ~n15168 & n15181 ;
  assign n15183 = ~n15180 & ~n15182 ;
  assign n15184 = ~n15166 & ~n15183 ;
  assign n15185 = n14661 & n15184 ;
  assign n15186 = n15166 & ~n15183 ;
  assign n15187 = ~n14661 & n15186 ;
  assign n15188 = ~n15185 & ~n15187 ;
  assign n15189 = ~n15166 & n15183 ;
  assign n15190 = ~n14661 & n15189 ;
  assign n15191 = n15166 & n15183 ;
  assign n15192 = n14661 & n15191 ;
  assign n15193 = ~n15190 & ~n15192 ;
  assign n15194 = n15188 & n15193 ;
  assign n15195 = ~n14658 & n15194 ;
  assign n15196 = ~n14051 & ~n14094 ;
  assign n15197 = ~n14091 & n15196 ;
  assign n15198 = ~n14093 & ~n15197 ;
  assign n15199 = ~\b[51]  & ~\b[52]  ;
  assign n15200 = \b[51]  & \b[52]  ;
  assign n15201 = ~n15199 & ~n15200 ;
  assign n15202 = n134 & n15201 ;
  assign n15203 = ~n15198 & n15202 ;
  assign n15204 = n134 & ~n15201 ;
  assign n15205 = ~n14093 & n15204 ;
  assign n15206 = ~n15197 & n15205 ;
  assign n15207 = \a[0]  & \b[52]  ;
  assign n15208 = n133 & n15207 ;
  assign n15209 = \b[51]  & n141 ;
  assign n15210 = ~\a[1]  & \b[50]  ;
  assign n15211 = n10416 & n15210 ;
  assign n15212 = ~n15209 & ~n15211 ;
  assign n15213 = ~n15208 & n15212 ;
  assign n15214 = \a[2]  & n15213 ;
  assign n15215 = ~n15206 & n15214 ;
  assign n15216 = ~n15203 & n15215 ;
  assign n15217 = ~n15206 & n15213 ;
  assign n15218 = ~n15203 & n15217 ;
  assign n15219 = ~\a[2]  & ~n15218 ;
  assign n15220 = ~n15216 & ~n15219 ;
  assign n15221 = n14637 & ~n15194 ;
  assign n15222 = ~n14657 & n15221 ;
  assign n15223 = ~n15220 & ~n15222 ;
  assign n15224 = ~n15195 & n15223 ;
  assign n15225 = ~n15194 & n15220 ;
  assign n15226 = n14658 & n15225 ;
  assign n15227 = n15194 & n15220 ;
  assign n15228 = ~n14658 & n15227 ;
  assign n15229 = ~n15226 & ~n15228 ;
  assign n15230 = ~n15224 & n15229 ;
  assign n15231 = n14656 & n15230 ;
  assign n15232 = ~n14656 & ~n15230 ;
  assign n15233 = ~n15231 & ~n15232 ;
  assign n15234 = ~n15224 & ~n15231 ;
  assign n15235 = n14637 & n15188 ;
  assign n15236 = ~n14657 & n15235 ;
  assign n15237 = n15193 & ~n15236 ;
  assign n15238 = ~n14093 & n15201 ;
  assign n15239 = ~n15197 & n15238 ;
  assign n15240 = ~n15200 & ~n15239 ;
  assign n15241 = ~\b[52]  & ~\b[53]  ;
  assign n15242 = \b[52]  & \b[53]  ;
  assign n15243 = ~n15241 & ~n15242 ;
  assign n15244 = ~n15240 & n15243 ;
  assign n15245 = ~n15200 & ~n15243 ;
  assign n15246 = ~n15239 & n15245 ;
  assign n15247 = n134 & ~n15246 ;
  assign n15248 = ~n15244 & n15247 ;
  assign n15249 = \a[0]  & \b[53]  ;
  assign n15250 = n133 & n15249 ;
  assign n15251 = \b[52]  & n141 ;
  assign n15252 = ~\a[1]  & \b[51]  ;
  assign n15253 = n10416 & n15252 ;
  assign n15254 = ~n15251 & ~n15253 ;
  assign n15255 = ~n15250 & n15254 ;
  assign n15256 = ~n15248 & n15255 ;
  assign n15257 = ~\a[2]  & ~n15256 ;
  assign n15258 = \a[2]  & n15255 ;
  assign n15259 = ~n15248 & n15258 ;
  assign n15260 = ~n15257 & ~n15259 ;
  assign n15261 = n14661 & n15166 ;
  assign n15262 = n15160 & ~n15261 ;
  assign n15263 = ~n14598 & ~n15149 ;
  assign n15264 = ~n14605 & n15263 ;
  assign n15265 = n15154 & ~n15264 ;
  assign n15266 = n430 & ~n12438 ;
  assign n15267 = ~n12436 & n15266 ;
  assign n15268 = \b[47]  & n428 ;
  assign n15269 = \a[6]  & \b[46]  ;
  assign n15270 = n419 & n15269 ;
  assign n15271 = ~n15268 & ~n15270 ;
  assign n15272 = \b[45]  & n486 ;
  assign n15273 = n483 & n15272 ;
  assign n15274 = ~\a[6]  & \b[46]  ;
  assign n15275 = n422 & n15274 ;
  assign n15276 = ~n15273 & ~n15275 ;
  assign n15277 = n15271 & n15276 ;
  assign n15278 = ~n15267 & n15277 ;
  assign n15279 = ~\a[8]  & ~n15278 ;
  assign n15280 = \a[8]  & n15277 ;
  assign n15281 = ~n15267 & n15280 ;
  assign n15282 = ~n15279 & ~n15281 ;
  assign n15283 = n15121 & ~n15130 ;
  assign n15284 = n14530 & ~n15092 ;
  assign n15285 = ~n14539 & n15284 ;
  assign n15286 = ~n15093 & ~n15285 ;
  assign n15287 = ~n15065 & ~n15073 ;
  assign n15288 = n14491 & n15030 ;
  assign n15289 = ~n14693 & n15288 ;
  assign n15290 = n15035 & ~n15289 ;
  assign n15291 = n14697 & n15008 ;
  assign n15292 = ~n15002 & ~n15291 ;
  assign n15293 = n2622 & n5810 ;
  assign n15294 = ~n5807 & n15293 ;
  assign n15295 = n2622 & ~n5810 ;
  assign n15296 = ~n5457 & n15295 ;
  assign n15297 = ~n5806 & n15296 ;
  assign n15298 = \b[30]  & n2912 ;
  assign n15299 = n2909 & n15298 ;
  assign n15300 = ~\a[21]  & \b[31]  ;
  assign n15301 = n2614 & n15300 ;
  assign n15302 = ~n15299 & ~n15301 ;
  assign n15303 = \b[32]  & n2620 ;
  assign n15304 = \a[21]  & \b[31]  ;
  assign n15305 = n2611 & n15304 ;
  assign n15306 = \a[23]  & ~n15305 ;
  assign n15307 = ~n15303 & n15306 ;
  assign n15308 = n15302 & n15307 ;
  assign n15309 = ~n15297 & n15308 ;
  assign n15310 = ~n15294 & n15309 ;
  assign n15311 = ~n15303 & ~n15305 ;
  assign n15312 = n15302 & n15311 ;
  assign n15313 = ~n15297 & n15312 ;
  assign n15314 = ~n15294 & n15313 ;
  assign n15315 = ~\a[23]  & ~n15314 ;
  assign n15316 = ~n15310 & ~n15315 ;
  assign n15317 = n14454 & n14967 ;
  assign n15318 = ~n14458 & n15317 ;
  assign n15319 = n14972 & ~n15318 ;
  assign n15320 = n3402 & ~n4502 ;
  assign n15321 = ~n4500 & n15320 ;
  assign n15322 = \b[29]  & n3400 ;
  assign n15323 = \a[24]  & \b[28]  ;
  assign n15324 = n3391 & n15323 ;
  assign n15325 = ~n15322 & ~n15324 ;
  assign n15326 = \b[27]  & n3733 ;
  assign n15327 = n3730 & n15326 ;
  assign n15328 = ~\a[24]  & \b[28]  ;
  assign n15329 = n3394 & n15328 ;
  assign n15330 = ~n15327 & ~n15329 ;
  assign n15331 = n15325 & n15330 ;
  assign n15332 = ~n15321 & n15331 ;
  assign n15333 = ~\a[26]  & ~n15332 ;
  assign n15334 = \a[26]  & n15331 ;
  assign n15335 = ~n15321 & n15334 ;
  assign n15336 = ~n15333 & ~n15335 ;
  assign n15337 = n14701 & n14945 ;
  assign n15338 = n14939 & ~n15337 ;
  assign n15339 = n3604 & n4249 ;
  assign n15340 = ~n3601 & n15339 ;
  assign n15341 = n4249 & n12021 ;
  assign n15342 = ~n3600 & n15341 ;
  assign n15343 = \b[24]  & n4647 ;
  assign n15344 = n4644 & n15343 ;
  assign n15345 = ~\a[27]  & \b[25]  ;
  assign n15346 = n4241 & n15345 ;
  assign n15347 = ~n15344 & ~n15346 ;
  assign n15348 = \b[26]  & n4247 ;
  assign n15349 = \a[27]  & \b[25]  ;
  assign n15350 = n4238 & n15349 ;
  assign n15351 = \a[29]  & ~n15350 ;
  assign n15352 = ~n15348 & n15351 ;
  assign n15353 = n15347 & n15352 ;
  assign n15354 = ~n15342 & n15353 ;
  assign n15355 = ~n15340 & n15354 ;
  assign n15356 = ~n15348 & ~n15350 ;
  assign n15357 = n15347 & n15356 ;
  assign n15358 = ~n15342 & n15357 ;
  assign n15359 = ~n15340 & n15358 ;
  assign n15360 = ~\a[29]  & ~n15359 ;
  assign n15361 = ~n15355 & ~n15360 ;
  assign n15362 = ~n14384 & ~n14932 ;
  assign n15363 = ~n14391 & n15362 ;
  assign n15364 = ~n14933 & ~n15363 ;
  assign n15365 = ~n3022 & n5211 ;
  assign n15366 = ~n3020 & n15365 ;
  assign n15367 = \b[23]  & n5209 ;
  assign n15368 = \a[30]  & \b[22]  ;
  assign n15369 = n5200 & n15368 ;
  assign n15370 = ~n15367 & ~n15369 ;
  assign n15371 = \b[21]  & n5595 ;
  assign n15372 = n5592 & n15371 ;
  assign n15373 = ~\a[30]  & \b[22]  ;
  assign n15374 = n5203 & n15373 ;
  assign n15375 = ~n15372 & ~n15374 ;
  assign n15376 = n15370 & n15375 ;
  assign n15377 = ~n15366 & n15376 ;
  assign n15378 = ~\a[32]  & ~n15377 ;
  assign n15379 = \a[32]  & n15376 ;
  assign n15380 = ~n15366 & n15379 ;
  assign n15381 = ~n15378 & ~n15380 ;
  assign n15382 = ~n14898 & ~n14906 ;
  assign n15383 = n2293 & n6309 ;
  assign n15384 = ~n2290 & n15383 ;
  assign n15385 = n5705 & n6309 ;
  assign n15386 = ~n2289 & n15385 ;
  assign n15387 = \b[18]  & n6778 ;
  assign n15388 = n6775 & n15387 ;
  assign n15389 = ~\a[33]  & \b[19]  ;
  assign n15390 = n6301 & n15389 ;
  assign n15391 = ~n15388 & ~n15390 ;
  assign n15392 = \b[20]  & n6307 ;
  assign n15393 = \a[33]  & \b[19]  ;
  assign n15394 = n6298 & n15393 ;
  assign n15395 = \a[35]  & ~n15394 ;
  assign n15396 = ~n15392 & n15395 ;
  assign n15397 = n15391 & n15396 ;
  assign n15398 = ~n15386 & n15397 ;
  assign n15399 = ~n15384 & n15398 ;
  assign n15400 = ~n15392 & ~n15394 ;
  assign n15401 = n15391 & n15400 ;
  assign n15402 = ~n15386 & n15401 ;
  assign n15403 = ~n15384 & n15402 ;
  assign n15404 = ~\a[35]  & ~n15403 ;
  assign n15405 = ~n15399 & ~n15404 ;
  assign n15406 = n14339 & n14871 ;
  assign n15407 = ~n14731 & n15406 ;
  assign n15408 = n14866 & ~n15407 ;
  assign n15409 = ~n1691 & n7534 ;
  assign n15410 = ~n1511 & n7534 ;
  assign n15411 = ~n1515 & n15410 ;
  assign n15412 = ~n15409 & ~n15411 ;
  assign n15413 = ~n1694 & ~n15412 ;
  assign n15414 = \b[15]  & n7973 ;
  assign n15415 = n7970 & n15414 ;
  assign n15416 = \b[17]  & n7532 ;
  assign n15417 = \a[36]  & \b[16]  ;
  assign n15418 = n7523 & n15417 ;
  assign n15419 = ~\a[36]  & \b[16]  ;
  assign n15420 = n7526 & n15419 ;
  assign n15421 = ~n15418 & ~n15420 ;
  assign n15422 = ~n15416 & n15421 ;
  assign n15423 = ~n15415 & n15422 ;
  assign n15424 = ~\a[38]  & n15423 ;
  assign n15425 = ~n15413 & n15424 ;
  assign n15426 = \a[38]  & ~n15423 ;
  assign n15427 = \a[38]  & ~n1694 ;
  assign n15428 = ~n15412 & n15427 ;
  assign n15429 = ~n15426 & ~n15428 ;
  assign n15430 = ~n15425 & n15429 ;
  assign n15431 = n14735 & n14861 ;
  assign n15432 = n14855 & ~n15431 ;
  assign n15433 = ~n728 & n10082 ;
  assign n15434 = ~n726 & n15433 ;
  assign n15435 = \b[9]  & n10681 ;
  assign n15436 = n10678 & n15435 ;
  assign n15437 = \b[11]  & n10080 ;
  assign n15438 = \a[41]  & \b[10]  ;
  assign n15439 = n10679 & n15438 ;
  assign n15440 = ~\a[42]  & \b[10]  ;
  assign n15441 = n10074 & n15440 ;
  assign n15442 = ~n15439 & ~n15441 ;
  assign n15443 = ~n15437 & n15442 ;
  assign n15444 = ~n15436 & n15443 ;
  assign n15445 = ~n15434 & n15444 ;
  assign n15446 = ~\a[44]  & ~n15445 ;
  assign n15447 = \a[44]  & n15444 ;
  assign n15448 = ~n15434 & n15447 ;
  assign n15449 = ~n15446 & ~n15448 ;
  assign n15450 = ~n14309 & ~n14826 ;
  assign n15451 = ~n14313 & n15450 ;
  assign n15452 = ~n14827 & ~n15451 ;
  assign n15453 = ~n505 & ~n10988 ;
  assign n15454 = ~n11569 & n15453 ;
  assign n15455 = n502 & n15454 ;
  assign n15456 = n505 & ~n10988 ;
  assign n15457 = ~n11569 & n15456 ;
  assign n15458 = ~n502 & n15457 ;
  assign n15459 = ~n15455 & ~n15458 ;
  assign n15460 = \b[6]  & n12159 ;
  assign n15461 = n12156 & n15460 ;
  assign n15462 = ~\a[45]  & \b[7]  ;
  assign n15463 = n11564 & n15462 ;
  assign n15464 = ~n15461 & ~n15463 ;
  assign n15465 = \b[8]  & n11570 ;
  assign n15466 = \a[45]  & \b[7]  ;
  assign n15467 = n11561 & n15466 ;
  assign n15468 = \a[47]  & ~n15467 ;
  assign n15469 = ~n15465 & n15468 ;
  assign n15470 = n15464 & n15469 ;
  assign n15471 = n15459 & n15470 ;
  assign n15472 = ~n15465 & ~n15467 ;
  assign n15473 = n15464 & n15472 ;
  assign n15474 = n15459 & n15473 ;
  assign n15475 = ~\a[47]  & ~n15474 ;
  assign n15476 = ~n15471 & ~n15475 ;
  assign n15477 = ~n14802 & ~n14804 ;
  assign n15478 = ~n270 & n13125 ;
  assign n15479 = ~n218 & n13125 ;
  assign n15480 = ~n220 & n15479 ;
  assign n15481 = ~n15478 & ~n15480 ;
  assign n15482 = ~n273 & ~n15481 ;
  assign n15483 = \b[3]  & n13794 ;
  assign n15484 = n13792 & n15483 ;
  assign n15485 = ~\a[47]  & \b[4]  ;
  assign n15486 = n13793 & n15485 ;
  assign n15487 = ~n15484 & ~n15486 ;
  assign n15488 = \b[5]  & n13123 ;
  assign n15489 = \a[48]  & \b[4]  ;
  assign n15490 = n13786 & n15489 ;
  assign n15491 = \a[50]  & ~n15490 ;
  assign n15492 = ~n15488 & n15491 ;
  assign n15493 = n15487 & n15492 ;
  assign n15494 = ~n15482 & n15493 ;
  assign n15495 = ~n15488 & ~n15490 ;
  assign n15496 = n15487 & n15495 ;
  assign n15497 = ~\a[50]  & ~n15496 ;
  assign n15498 = ~\a[50]  & ~n273 ;
  assign n15499 = ~n15481 & n15498 ;
  assign n15500 = ~n15497 & ~n15499 ;
  assign n15501 = ~n15494 & n15500 ;
  assign n15502 = \a[53]  & ~n14277 ;
  assign n15503 = n14787 & n15502 ;
  assign n15504 = n14795 & n15503 ;
  assign n15505 = \a[53]  & ~n15504 ;
  assign n15506 = \b[2]  & n14791 ;
  assign n15507 = ~\a[51]  & \b[1]  ;
  assign n15508 = n14785 & n15507 ;
  assign n15509 = \a[51]  & \b[1]  ;
  assign n15510 = n14782 & n15509 ;
  assign n15511 = ~n15508 & ~n15510 ;
  assign n15512 = ~n15506 & n15511 ;
  assign n15513 = n157 & n14793 ;
  assign n15514 = n14276 & ~n14790 ;
  assign n15515 = \a[51]  & ~\a[52]  ;
  assign n15516 = ~\a[51]  & \a[52]  ;
  assign n15517 = ~n15515 & ~n15516 ;
  assign n15518 = \b[0]  & n15517 ;
  assign n15519 = n15514 & n15518 ;
  assign n15520 = ~n15513 & ~n15519 ;
  assign n15521 = n15512 & n15520 ;
  assign n15522 = ~n15505 & ~n15521 ;
  assign n15523 = n15505 & n15521 ;
  assign n15524 = ~n15522 & ~n15523 ;
  assign n15525 = ~n15501 & ~n15524 ;
  assign n15526 = n15501 & n15524 ;
  assign n15527 = ~n15525 & ~n15526 ;
  assign n15528 = ~n15477 & n15527 ;
  assign n15529 = ~n14802 & ~n15527 ;
  assign n15530 = ~n14804 & n15529 ;
  assign n15531 = ~n15528 & ~n15530 ;
  assign n15532 = n15476 & ~n15531 ;
  assign n15533 = ~n15476 & ~n15530 ;
  assign n15534 = ~n15528 & n15533 ;
  assign n15535 = ~n15532 & ~n15534 ;
  assign n15536 = n15452 & n15535 ;
  assign n15537 = ~n15452 & ~n15535 ;
  assign n15538 = ~n15536 & ~n15537 ;
  assign n15539 = n15449 & ~n15538 ;
  assign n15540 = ~n15449 & n15538 ;
  assign n15541 = ~n15539 & ~n15540 ;
  assign n15542 = n1087 & n8759 ;
  assign n15543 = ~n1084 & n15542 ;
  assign n15544 = n1552 & n8759 ;
  assign n15545 = ~n1083 & n15544 ;
  assign n15546 = \b[12]  & n9301 ;
  assign n15547 = n9298 & n15546 ;
  assign n15548 = ~\a[39]  & \b[13]  ;
  assign n15549 = n8751 & n15548 ;
  assign n15550 = ~n15547 & ~n15549 ;
  assign n15551 = \b[14]  & n8757 ;
  assign n15552 = \a[39]  & \b[13]  ;
  assign n15553 = n8748 & n15552 ;
  assign n15554 = \a[41]  & ~n15553 ;
  assign n15555 = ~n15551 & n15554 ;
  assign n15556 = n15550 & n15555 ;
  assign n15557 = ~n15545 & n15556 ;
  assign n15558 = ~n15543 & n15557 ;
  assign n15559 = ~n15551 & ~n15553 ;
  assign n15560 = n15550 & n15559 ;
  assign n15561 = ~n15545 & n15560 ;
  assign n15562 = ~n15543 & n15561 ;
  assign n15563 = ~\a[41]  & ~n15562 ;
  assign n15564 = ~n15558 & ~n15563 ;
  assign n15565 = ~n15541 & ~n15564 ;
  assign n15566 = ~n15432 & n15565 ;
  assign n15567 = n15541 & ~n15564 ;
  assign n15568 = n15432 & n15567 ;
  assign n15569 = ~n15566 & ~n15568 ;
  assign n15570 = ~n15541 & n15564 ;
  assign n15571 = n15432 & n15570 ;
  assign n15572 = n15541 & n15564 ;
  assign n15573 = ~n15432 & n15572 ;
  assign n15574 = ~n15571 & ~n15573 ;
  assign n15575 = n15569 & n15574 ;
  assign n15576 = n15430 & ~n15575 ;
  assign n15577 = n15408 & n15576 ;
  assign n15578 = n15430 & n15575 ;
  assign n15579 = ~n15408 & n15578 ;
  assign n15580 = ~n15577 & ~n15579 ;
  assign n15581 = ~n15430 & ~n15575 ;
  assign n15582 = ~n15408 & n15581 ;
  assign n15583 = ~n15430 & n15575 ;
  assign n15584 = n15408 & n15583 ;
  assign n15585 = ~n15582 & ~n15584 ;
  assign n15586 = n15580 & n15585 ;
  assign n15587 = ~n15405 & ~n15586 ;
  assign n15588 = ~n15382 & n15587 ;
  assign n15589 = ~n15405 & n15586 ;
  assign n15590 = n15382 & n15589 ;
  assign n15591 = ~n15588 & ~n15590 ;
  assign n15592 = n15405 & ~n15586 ;
  assign n15593 = n15382 & n15592 ;
  assign n15594 = n15405 & n15586 ;
  assign n15595 = ~n15382 & n15594 ;
  assign n15596 = ~n15593 & ~n15595 ;
  assign n15597 = n15591 & n15596 ;
  assign n15598 = ~n15381 & ~n15597 ;
  assign n15599 = n15364 & n15598 ;
  assign n15600 = ~n15381 & n15597 ;
  assign n15601 = ~n15364 & n15600 ;
  assign n15602 = ~n15599 & ~n15601 ;
  assign n15603 = n15381 & ~n15597 ;
  assign n15604 = ~n15364 & n15603 ;
  assign n15605 = n15381 & n15597 ;
  assign n15606 = n15364 & n15605 ;
  assign n15607 = ~n15604 & ~n15606 ;
  assign n15608 = n15602 & n15607 ;
  assign n15609 = n15361 & ~n15608 ;
  assign n15610 = n15338 & n15609 ;
  assign n15611 = n15361 & n15608 ;
  assign n15612 = ~n15338 & n15611 ;
  assign n15613 = ~n15610 & ~n15612 ;
  assign n15614 = ~n15338 & n15608 ;
  assign n15615 = n14939 & ~n15608 ;
  assign n15616 = ~n15337 & n15615 ;
  assign n15617 = ~n15361 & ~n15616 ;
  assign n15618 = ~n15614 & n15617 ;
  assign n15619 = n15613 & ~n15618 ;
  assign n15620 = n15336 & ~n15619 ;
  assign n15621 = ~n15319 & n15620 ;
  assign n15622 = n15336 & n15619 ;
  assign n15623 = n15319 & n15622 ;
  assign n15624 = ~n15621 & ~n15623 ;
  assign n15625 = ~n15336 & ~n15619 ;
  assign n15626 = n15319 & n15625 ;
  assign n15627 = ~n15336 & n15619 ;
  assign n15628 = ~n15319 & n15627 ;
  assign n15629 = ~n15626 & ~n15628 ;
  assign n15630 = n15624 & n15629 ;
  assign n15631 = n15316 & ~n15630 ;
  assign n15632 = n15292 & n15631 ;
  assign n15633 = n15316 & n15630 ;
  assign n15634 = ~n15292 & n15633 ;
  assign n15635 = ~n15632 & ~n15634 ;
  assign n15636 = ~n15292 & n15630 ;
  assign n15637 = ~n15002 & ~n15630 ;
  assign n15638 = ~n15291 & n15637 ;
  assign n15639 = ~n15316 & ~n15638 ;
  assign n15640 = ~n15636 & n15639 ;
  assign n15641 = n15635 & ~n15640 ;
  assign n15642 = n1965 & ~n6610 ;
  assign n15643 = ~n6608 & n15642 ;
  assign n15644 = \b[35]  & n1963 ;
  assign n15645 = \a[18]  & \b[34]  ;
  assign n15646 = n2210 & n15645 ;
  assign n15647 = ~n15644 & ~n15646 ;
  assign n15648 = \b[33]  & n2218 ;
  assign n15649 = n2216 & n15648 ;
  assign n15650 = ~\a[18]  & \b[34]  ;
  assign n15651 = n1957 & n15650 ;
  assign n15652 = ~n15649 & ~n15651 ;
  assign n15653 = n15647 & n15652 ;
  assign n15654 = ~n15643 & n15653 ;
  assign n15655 = ~\a[20]  & ~n15654 ;
  assign n15656 = \a[20]  & n15653 ;
  assign n15657 = ~n15643 & n15656 ;
  assign n15658 = ~n15655 & ~n15657 ;
  assign n15659 = ~n15641 & ~n15658 ;
  assign n15660 = n15290 & n15659 ;
  assign n15661 = n15641 & ~n15658 ;
  assign n15662 = ~n15290 & n15661 ;
  assign n15663 = ~n15660 & ~n15662 ;
  assign n15664 = ~n15641 & n15658 ;
  assign n15665 = ~n15290 & n15664 ;
  assign n15666 = n15641 & n15658 ;
  assign n15667 = n15290 & n15666 ;
  assign n15668 = ~n15665 & ~n15667 ;
  assign n15669 = n15663 & n15668 ;
  assign n15670 = n1467 & n8175 ;
  assign n15671 = ~n8172 & n15670 ;
  assign n15672 = n1467 & ~n8175 ;
  assign n15673 = ~n7756 & n15672 ;
  assign n15674 = ~n8171 & n15673 ;
  assign n15675 = \b[36]  & n1652 ;
  assign n15676 = n1649 & n15675 ;
  assign n15677 = ~\a[15]  & \b[37]  ;
  assign n15678 = n1459 & n15677 ;
  assign n15679 = ~n15676 & ~n15678 ;
  assign n15680 = \b[38]  & n1465 ;
  assign n15681 = \a[15]  & \b[37]  ;
  assign n15682 = n1456 & n15681 ;
  assign n15683 = \a[17]  & ~n15682 ;
  assign n15684 = ~n15680 & n15683 ;
  assign n15685 = n15679 & n15684 ;
  assign n15686 = ~n15674 & n15685 ;
  assign n15687 = ~n15671 & n15686 ;
  assign n15688 = ~n15680 & ~n15682 ;
  assign n15689 = n15679 & n15688 ;
  assign n15690 = ~n15674 & n15689 ;
  assign n15691 = ~n15671 & n15690 ;
  assign n15692 = ~\a[17]  & ~n15691 ;
  assign n15693 = ~n15687 & ~n15692 ;
  assign n15694 = ~n15669 & ~n15693 ;
  assign n15695 = ~n15287 & n15694 ;
  assign n15696 = n15669 & ~n15693 ;
  assign n15697 = n15287 & n15696 ;
  assign n15698 = ~n15695 & ~n15697 ;
  assign n15699 = ~n15669 & n15693 ;
  assign n15700 = n15287 & n15699 ;
  assign n15701 = n15669 & n15693 ;
  assign n15702 = ~n15287 & n15701 ;
  assign n15703 = ~n15700 & ~n15702 ;
  assign n15704 = n15698 & n15703 ;
  assign n15705 = n999 & ~n9482 ;
  assign n15706 = ~n9480 & n15705 ;
  assign n15707 = \b[39]  & n1182 ;
  assign n15708 = n1179 & n15707 ;
  assign n15709 = \b[41]  & n997 ;
  assign n15710 = \a[11]  & \b[40]  ;
  assign n15711 = n1180 & n15710 ;
  assign n15712 = ~\a[12]  & \b[40]  ;
  assign n15713 = n7674 & n15712 ;
  assign n15714 = ~n15711 & ~n15713 ;
  assign n15715 = ~n15709 & n15714 ;
  assign n15716 = ~n15708 & n15715 ;
  assign n15717 = ~n15706 & n15716 ;
  assign n15718 = ~\a[14]  & ~n15717 ;
  assign n15719 = \a[14]  & n15716 ;
  assign n15720 = ~n15706 & n15719 ;
  assign n15721 = ~n15718 & ~n15720 ;
  assign n15722 = ~n15704 & ~n15721 ;
  assign n15723 = n15286 & n15722 ;
  assign n15724 = n15704 & ~n15721 ;
  assign n15725 = ~n15286 & n15724 ;
  assign n15726 = ~n15723 & ~n15725 ;
  assign n15727 = ~n15704 & n15721 ;
  assign n15728 = ~n15286 & n15727 ;
  assign n15729 = n15704 & n15721 ;
  assign n15730 = n15286 & n15729 ;
  assign n15731 = ~n15728 & ~n15730 ;
  assign n15732 = n15726 & n15731 ;
  assign n15733 = ~n15283 & n15732 ;
  assign n15734 = n15121 & ~n15732 ;
  assign n15735 = ~n15130 & n15734 ;
  assign n15736 = n646 & ~n10892 ;
  assign n15737 = ~n10890 & n15736 ;
  assign n15738 = \b[42]  & n796 ;
  assign n15739 = n793 & n15738 ;
  assign n15740 = ~\a[9]  & \b[43]  ;
  assign n15741 = n638 & n15740 ;
  assign n15742 = ~n15739 & ~n15741 ;
  assign n15743 = \b[44]  & n644 ;
  assign n15744 = \a[9]  & \b[43]  ;
  assign n15745 = n635 & n15744 ;
  assign n15746 = \a[11]  & ~n15745 ;
  assign n15747 = ~n15743 & n15746 ;
  assign n15748 = n15742 & n15747 ;
  assign n15749 = ~n15737 & n15748 ;
  assign n15750 = ~n15743 & ~n15745 ;
  assign n15751 = n15742 & n15750 ;
  assign n15752 = ~n15737 & n15751 ;
  assign n15753 = ~\a[11]  & ~n15752 ;
  assign n15754 = ~n15749 & ~n15753 ;
  assign n15755 = ~n15735 & ~n15754 ;
  assign n15756 = ~n15733 & n15755 ;
  assign n15757 = ~n15732 & n15754 ;
  assign n15758 = n15283 & n15757 ;
  assign n15759 = n15732 & n15754 ;
  assign n15760 = ~n15283 & n15759 ;
  assign n15761 = ~n15758 & ~n15760 ;
  assign n15762 = ~n15756 & n15761 ;
  assign n15763 = ~n15282 & ~n15762 ;
  assign n15764 = n15265 & n15763 ;
  assign n15765 = ~n15282 & n15762 ;
  assign n15766 = ~n15265 & n15765 ;
  assign n15767 = ~n15764 & ~n15766 ;
  assign n15768 = n15282 & ~n15762 ;
  assign n15769 = ~n15265 & n15768 ;
  assign n15770 = n15282 & n15762 ;
  assign n15771 = n15265 & n15770 ;
  assign n15772 = ~n15769 & ~n15771 ;
  assign n15773 = n15767 & n15772 ;
  assign n15774 = ~n15262 & n15773 ;
  assign n15775 = n15160 & ~n15773 ;
  assign n15776 = ~n15261 & n15775 ;
  assign n15777 = n252 & n14052 ;
  assign n15778 = ~n14049 & n15777 ;
  assign n15779 = ~n13519 & ~n14052 ;
  assign n15780 = n252 & n15779 ;
  assign n15781 = ~n14048 & n15780 ;
  assign n15782 = \b[48]  & n303 ;
  assign n15783 = n300 & n15782 ;
  assign n15784 = ~\a[3]  & \b[49]  ;
  assign n15785 = n244 & n15784 ;
  assign n15786 = ~n15783 & ~n15785 ;
  assign n15787 = \b[50]  & n250 ;
  assign n15788 = \a[3]  & \b[49]  ;
  assign n15789 = n241 & n15788 ;
  assign n15790 = \a[5]  & ~n15789 ;
  assign n15791 = ~n15787 & n15790 ;
  assign n15792 = n15786 & n15791 ;
  assign n15793 = ~n15781 & n15792 ;
  assign n15794 = ~n15778 & n15793 ;
  assign n15795 = ~n15787 & ~n15789 ;
  assign n15796 = n15786 & n15795 ;
  assign n15797 = ~n15781 & n15796 ;
  assign n15798 = ~n15778 & n15797 ;
  assign n15799 = ~\a[5]  & ~n15798 ;
  assign n15800 = ~n15794 & ~n15799 ;
  assign n15801 = ~n15776 & ~n15800 ;
  assign n15802 = ~n15774 & n15801 ;
  assign n15803 = ~n15773 & n15800 ;
  assign n15804 = n15262 & n15803 ;
  assign n15805 = n15773 & n15800 ;
  assign n15806 = ~n15262 & n15805 ;
  assign n15807 = ~n15804 & ~n15806 ;
  assign n15808 = ~n15802 & n15807 ;
  assign n15809 = ~n15260 & ~n15808 ;
  assign n15810 = n15237 & n15809 ;
  assign n15811 = ~n15260 & n15808 ;
  assign n15812 = ~n15237 & n15811 ;
  assign n15813 = ~n15810 & ~n15812 ;
  assign n15814 = n15260 & ~n15808 ;
  assign n15815 = ~n15237 & n15814 ;
  assign n15816 = n15260 & n15808 ;
  assign n15817 = n15237 & n15816 ;
  assign n15818 = ~n15815 & ~n15817 ;
  assign n15819 = n15813 & n15818 ;
  assign n15820 = ~n15234 & n15819 ;
  assign n15821 = ~n15224 & ~n15819 ;
  assign n15822 = ~n15231 & n15821 ;
  assign n15823 = ~n15820 & ~n15822 ;
  assign n15824 = ~n15224 & n15813 ;
  assign n15825 = ~n15231 & n15824 ;
  assign n15826 = n15818 & ~n15825 ;
  assign n15827 = n15237 & n15808 ;
  assign n15828 = ~n15802 & ~n15827 ;
  assign n15829 = n15160 & n15767 ;
  assign n15830 = ~n15261 & n15829 ;
  assign n15831 = n15772 & ~n15830 ;
  assign n15832 = n15265 & n15762 ;
  assign n15833 = ~n15756 & ~n15832 ;
  assign n15834 = n15121 & n15726 ;
  assign n15835 = ~n15130 & n15834 ;
  assign n15836 = n15731 & ~n15835 ;
  assign n15837 = n646 & ~n11397 ;
  assign n15838 = ~n11395 & n15837 ;
  assign n15839 = \b[45]  & n644 ;
  assign n15840 = \a[9]  & \b[44]  ;
  assign n15841 = n635 & n15840 ;
  assign n15842 = ~n15839 & ~n15841 ;
  assign n15843 = \b[43]  & n796 ;
  assign n15844 = n793 & n15843 ;
  assign n15845 = ~\a[9]  & \b[44]  ;
  assign n15846 = n638 & n15845 ;
  assign n15847 = ~n15844 & ~n15846 ;
  assign n15848 = n15842 & n15847 ;
  assign n15849 = ~n15838 & n15848 ;
  assign n15850 = ~\a[11]  & ~n15849 ;
  assign n15851 = \a[11]  & n15848 ;
  assign n15852 = ~n15838 & n15851 ;
  assign n15853 = ~n15850 & ~n15852 ;
  assign n15854 = n15286 & n15704 ;
  assign n15855 = n15698 & ~n15854 ;
  assign n15856 = ~n15065 & n15663 ;
  assign n15857 = ~n15073 & n15856 ;
  assign n15858 = n15668 & ~n15857 ;
  assign n15859 = n15290 & n15641 ;
  assign n15860 = ~n15640 & ~n15859 ;
  assign n15861 = ~n15002 & n15629 ;
  assign n15862 = ~n15291 & n15861 ;
  assign n15863 = n15624 & ~n15862 ;
  assign n15864 = n15319 & n15619 ;
  assign n15865 = ~n15618 & ~n15864 ;
  assign n15866 = n14939 & n15602 ;
  assign n15867 = ~n15337 & n15866 ;
  assign n15868 = n15607 & ~n15867 ;
  assign n15869 = ~n4148 & n4249 ;
  assign n15870 = ~n4146 & n15869 ;
  assign n15871 = \b[25]  & n4647 ;
  assign n15872 = n4644 & n15871 ;
  assign n15873 = ~\a[27]  & \b[26]  ;
  assign n15874 = n4241 & n15873 ;
  assign n15875 = ~n15872 & ~n15874 ;
  assign n15876 = \b[27]  & n4247 ;
  assign n15877 = \a[27]  & \b[26]  ;
  assign n15878 = n4238 & n15877 ;
  assign n15879 = \a[29]  & ~n15878 ;
  assign n15880 = ~n15876 & n15879 ;
  assign n15881 = n15875 & n15880 ;
  assign n15882 = ~n15870 & n15881 ;
  assign n15883 = ~n15876 & ~n15878 ;
  assign n15884 = n15875 & n15883 ;
  assign n15885 = ~n15870 & n15884 ;
  assign n15886 = ~\a[29]  & ~n15885 ;
  assign n15887 = ~n15882 & ~n15886 ;
  assign n15888 = n15364 & n15597 ;
  assign n15889 = n15591 & ~n15888 ;
  assign n15890 = n3283 & n5211 ;
  assign n15891 = ~n3280 & n15890 ;
  assign n15892 = ~n3283 & n5211 ;
  assign n15893 = ~n3017 & n15892 ;
  assign n15894 = ~n3279 & n15893 ;
  assign n15895 = \b[22]  & n5595 ;
  assign n15896 = n5592 & n15895 ;
  assign n15897 = ~\a[30]  & \b[23]  ;
  assign n15898 = n5203 & n15897 ;
  assign n15899 = ~n15896 & ~n15898 ;
  assign n15900 = \b[24]  & n5209 ;
  assign n15901 = \a[30]  & \b[23]  ;
  assign n15902 = n5200 & n15901 ;
  assign n15903 = \a[32]  & ~n15902 ;
  assign n15904 = ~n15900 & n15903 ;
  assign n15905 = n15899 & n15904 ;
  assign n15906 = ~n15894 & n15905 ;
  assign n15907 = ~n15891 & n15906 ;
  assign n15908 = ~n15900 & ~n15902 ;
  assign n15909 = n15899 & n15908 ;
  assign n15910 = ~n15894 & n15909 ;
  assign n15911 = ~n15891 & n15910 ;
  assign n15912 = ~\a[32]  & ~n15911 ;
  assign n15913 = ~n15907 & ~n15912 ;
  assign n15914 = ~n2520 & n6309 ;
  assign n15915 = ~n2292 & n6309 ;
  assign n15916 = ~n2516 & n15915 ;
  assign n15917 = ~n15914 & ~n15916 ;
  assign n15918 = ~n2523 & ~n15917 ;
  assign n15919 = \b[19]  & n6778 ;
  assign n15920 = n6775 & n15919 ;
  assign n15921 = ~\a[33]  & \b[20]  ;
  assign n15922 = n6301 & n15921 ;
  assign n15923 = ~n15920 & ~n15922 ;
  assign n15924 = \b[21]  & n6307 ;
  assign n15925 = \a[33]  & \b[20]  ;
  assign n15926 = n6298 & n15925 ;
  assign n15927 = \a[35]  & ~n15926 ;
  assign n15928 = ~n15924 & n15927 ;
  assign n15929 = n15923 & n15928 ;
  assign n15930 = ~n15918 & n15929 ;
  assign n15931 = ~n15924 & ~n15926 ;
  assign n15932 = n15923 & n15931 ;
  assign n15933 = ~\a[35]  & ~n15932 ;
  assign n15934 = ~\a[35]  & ~n2523 ;
  assign n15935 = ~n15917 & n15934 ;
  assign n15936 = ~n15933 & ~n15935 ;
  assign n15937 = ~n15930 & n15936 ;
  assign n15938 = ~n14898 & n15580 ;
  assign n15939 = ~n14906 & n15938 ;
  assign n15940 = n15585 & ~n15939 ;
  assign n15941 = n15408 & n15575 ;
  assign n15942 = n15569 & ~n15941 ;
  assign n15943 = n14855 & ~n15540 ;
  assign n15944 = ~n15431 & n15943 ;
  assign n15945 = ~n15539 & ~n15944 ;
  assign n15946 = ~n1230 & n8759 ;
  assign n15947 = ~n1086 & n8759 ;
  assign n15948 = ~n1226 & n15947 ;
  assign n15949 = ~n15946 & ~n15948 ;
  assign n15950 = ~n1233 & ~n15949 ;
  assign n15951 = \b[13]  & n9301 ;
  assign n15952 = n9298 & n15951 ;
  assign n15953 = ~\a[39]  & \b[14]  ;
  assign n15954 = n8751 & n15953 ;
  assign n15955 = ~n15952 & ~n15954 ;
  assign n15956 = \b[15]  & n8757 ;
  assign n15957 = \a[39]  & \b[14]  ;
  assign n15958 = n8748 & n15957 ;
  assign n15959 = \a[41]  & ~n15958 ;
  assign n15960 = ~n15956 & n15959 ;
  assign n15961 = n15955 & n15960 ;
  assign n15962 = ~n15950 & n15961 ;
  assign n15963 = ~n15956 & ~n15958 ;
  assign n15964 = n15955 & n15963 ;
  assign n15965 = ~\a[41]  & ~n15964 ;
  assign n15966 = ~\a[41]  & ~n1233 ;
  assign n15967 = ~n15949 & n15966 ;
  assign n15968 = ~n15965 & ~n15967 ;
  assign n15969 = ~n15962 & n15968 ;
  assign n15970 = ~n15534 & ~n15536 ;
  assign n15971 = ~n14802 & ~n15525 ;
  assign n15972 = ~n14804 & n15971 ;
  assign n15973 = ~n15526 & ~n15972 ;
  assign n15974 = ~n586 & n11572 ;
  assign n15975 = ~n504 & n11572 ;
  assign n15976 = ~n508 & n15975 ;
  assign n15977 = ~n15974 & ~n15976 ;
  assign n15978 = ~n589 & ~n15977 ;
  assign n15979 = \b[7]  & n12159 ;
  assign n15980 = n12156 & n15979 ;
  assign n15981 = ~\a[45]  & \b[8]  ;
  assign n15982 = n11564 & n15981 ;
  assign n15983 = ~n15980 & ~n15982 ;
  assign n15984 = \b[9]  & n11570 ;
  assign n15985 = \a[45]  & \b[8]  ;
  assign n15986 = n11561 & n15985 ;
  assign n15987 = \a[47]  & ~n15986 ;
  assign n15988 = ~n15984 & n15987 ;
  assign n15989 = n15983 & n15988 ;
  assign n15990 = ~n15978 & n15989 ;
  assign n15991 = ~n15984 & ~n15986 ;
  assign n15992 = n15983 & n15991 ;
  assign n15993 = ~\a[47]  & ~n15992 ;
  assign n15994 = ~\a[47]  & ~n589 ;
  assign n15995 = ~n15977 & n15994 ;
  assign n15996 = ~n15993 & ~n15995 ;
  assign n15997 = ~n15990 & n15996 ;
  assign n15998 = n177 & n14793 ;
  assign n15999 = \b[3]  & n14791 ;
  assign n16000 = \a[50]  & \b[2]  ;
  assign n16001 = n15515 & n16000 ;
  assign n16002 = ~\a[51]  & \b[2]  ;
  assign n16003 = n14785 & n16002 ;
  assign n16004 = ~n16001 & ~n16003 ;
  assign n16005 = ~n15999 & n16004 ;
  assign n16006 = ~n15998 & n16005 ;
  assign n16007 = \b[1]  & n15517 ;
  assign n16008 = n15514 & n16007 ;
  assign n16009 = ~\a[53]  & ~n16008 ;
  assign n16010 = n16006 & n16009 ;
  assign n16011 = n16006 & ~n16008 ;
  assign n16012 = \a[53]  & ~n16011 ;
  assign n16013 = ~n16010 & ~n16012 ;
  assign n16014 = \a[53]  & ~\a[54]  ;
  assign n16015 = ~\a[53]  & \a[54]  ;
  assign n16016 = ~n16014 & ~n16015 ;
  assign n16017 = \b[0]  & ~n16016 ;
  assign n16018 = n15504 & n15521 ;
  assign n16019 = n16017 & n16018 ;
  assign n16020 = ~n16017 & ~n16018 ;
  assign n16021 = ~n16019 & ~n16020 ;
  assign n16022 = n16013 & n16021 ;
  assign n16023 = ~n16013 & ~n16021 ;
  assign n16024 = ~n16022 & ~n16023 ;
  assign n16025 = ~n323 & ~n12606 ;
  assign n16026 = ~n13122 & n16025 ;
  assign n16027 = n320 & n16026 ;
  assign n16028 = n323 & ~n12606 ;
  assign n16029 = ~n13122 & n16028 ;
  assign n16030 = ~n320 & n16029 ;
  assign n16031 = ~n16027 & ~n16030 ;
  assign n16032 = \b[4]  & n13794 ;
  assign n16033 = n13792 & n16032 ;
  assign n16034 = \b[6]  & n13123 ;
  assign n16035 = \a[48]  & \b[5]  ;
  assign n16036 = n13786 & n16035 ;
  assign n16037 = ~\a[48]  & \b[5]  ;
  assign n16038 = n13117 & n16037 ;
  assign n16039 = ~n16036 & ~n16038 ;
  assign n16040 = ~n16034 & n16039 ;
  assign n16041 = ~n16033 & n16040 ;
  assign n16042 = n16031 & n16041 ;
  assign n16043 = ~\a[50]  & ~n16042 ;
  assign n16044 = \a[50]  & n16041 ;
  assign n16045 = n16031 & n16044 ;
  assign n16046 = ~n16043 & ~n16045 ;
  assign n16047 = n16024 & ~n16046 ;
  assign n16048 = ~n16024 & n16046 ;
  assign n16049 = ~n16047 & ~n16048 ;
  assign n16050 = ~n15997 & ~n16049 ;
  assign n16051 = n15973 & n16050 ;
  assign n16052 = ~n15997 & n16049 ;
  assign n16053 = ~n15973 & n16052 ;
  assign n16054 = ~n16051 & ~n16053 ;
  assign n16055 = n15997 & ~n16049 ;
  assign n16056 = ~n15973 & n16055 ;
  assign n16057 = n15997 & n16049 ;
  assign n16058 = n15973 & n16057 ;
  assign n16059 = ~n16056 & ~n16058 ;
  assign n16060 = n16054 & n16059 ;
  assign n16061 = ~n15970 & n16060 ;
  assign n16062 = ~n909 & ~n9646 ;
  assign n16063 = ~n10079 & n16062 ;
  assign n16064 = n906 & n16063 ;
  assign n16065 = n909 & ~n9646 ;
  assign n16066 = ~n10079 & n16065 ;
  assign n16067 = ~n906 & n16066 ;
  assign n16068 = ~n16064 & ~n16067 ;
  assign n16069 = \b[10]  & n10681 ;
  assign n16070 = n10678 & n16069 ;
  assign n16071 = ~\a[42]  & \b[11]  ;
  assign n16072 = n10074 & n16071 ;
  assign n16073 = ~n16070 & ~n16072 ;
  assign n16074 = \b[12]  & n10080 ;
  assign n16075 = \a[42]  & \b[11]  ;
  assign n16076 = n10071 & n16075 ;
  assign n16077 = \a[44]  & ~n16076 ;
  assign n16078 = ~n16074 & n16077 ;
  assign n16079 = n16073 & n16078 ;
  assign n16080 = n16068 & n16079 ;
  assign n16081 = ~n16074 & ~n16076 ;
  assign n16082 = n16073 & n16081 ;
  assign n16083 = n16068 & n16082 ;
  assign n16084 = ~\a[44]  & ~n16083 ;
  assign n16085 = ~n16080 & ~n16084 ;
  assign n16086 = ~n15534 & ~n16060 ;
  assign n16087 = ~n15536 & n16086 ;
  assign n16088 = ~n16085 & ~n16087 ;
  assign n16089 = ~n16061 & n16088 ;
  assign n16090 = ~n16060 & n16085 ;
  assign n16091 = n15970 & n16090 ;
  assign n16092 = n16060 & n16085 ;
  assign n16093 = ~n15970 & n16092 ;
  assign n16094 = ~n16091 & ~n16093 ;
  assign n16095 = ~n16089 & n16094 ;
  assign n16096 = ~n15969 & ~n16095 ;
  assign n16097 = n15945 & n16096 ;
  assign n16098 = ~n15969 & n16095 ;
  assign n16099 = ~n15945 & n16098 ;
  assign n16100 = ~n16097 & ~n16099 ;
  assign n16101 = n15969 & ~n16095 ;
  assign n16102 = ~n15945 & n16101 ;
  assign n16103 = n15969 & n16095 ;
  assign n16104 = n15945 & n16103 ;
  assign n16105 = ~n16102 & ~n16104 ;
  assign n16106 = n16100 & n16105 ;
  assign n16107 = ~n15942 & n16106 ;
  assign n16108 = n1875 & n7534 ;
  assign n16109 = ~n1872 & n16108 ;
  assign n16110 = n5000 & n7534 ;
  assign n16111 = ~n1871 & n16110 ;
  assign n16112 = \b[16]  & n7973 ;
  assign n16113 = n7970 & n16112 ;
  assign n16114 = \b[18]  & n7532 ;
  assign n16115 = \a[36]  & \b[17]  ;
  assign n16116 = n7523 & n16115 ;
  assign n16117 = ~\a[36]  & \b[17]  ;
  assign n16118 = n7526 & n16117 ;
  assign n16119 = ~n16116 & ~n16118 ;
  assign n16120 = ~n16114 & n16119 ;
  assign n16121 = ~n16113 & n16120 ;
  assign n16122 = ~n16111 & n16121 ;
  assign n16123 = ~n16109 & n16122 ;
  assign n16124 = ~\a[38]  & ~n16123 ;
  assign n16125 = \a[38]  & n16121 ;
  assign n16126 = ~n16111 & n16125 ;
  assign n16127 = ~n16109 & n16126 ;
  assign n16128 = ~n16124 & ~n16127 ;
  assign n16129 = n15569 & ~n16106 ;
  assign n16130 = ~n15941 & n16129 ;
  assign n16131 = ~n16128 & ~n16130 ;
  assign n16132 = ~n16107 & n16131 ;
  assign n16133 = ~n16106 & n16128 ;
  assign n16134 = n15942 & n16133 ;
  assign n16135 = n16106 & n16128 ;
  assign n16136 = ~n15942 & n16135 ;
  assign n16137 = ~n16134 & ~n16136 ;
  assign n16138 = ~n16132 & n16137 ;
  assign n16139 = n15940 & n16138 ;
  assign n16140 = ~n15940 & ~n16138 ;
  assign n16141 = ~n16139 & ~n16140 ;
  assign n16142 = ~n15937 & n16141 ;
  assign n16143 = n15937 & ~n16141 ;
  assign n16144 = ~n16142 & ~n16143 ;
  assign n16145 = ~n15913 & ~n16144 ;
  assign n16146 = ~n15889 & n16145 ;
  assign n16147 = ~n15913 & n16144 ;
  assign n16148 = n15889 & n16147 ;
  assign n16149 = ~n16146 & ~n16148 ;
  assign n16150 = n15913 & ~n16144 ;
  assign n16151 = n15889 & n16150 ;
  assign n16152 = n15913 & n16144 ;
  assign n16153 = ~n15889 & n16152 ;
  assign n16154 = ~n16151 & ~n16153 ;
  assign n16155 = n16149 & n16154 ;
  assign n16156 = ~n15887 & ~n16155 ;
  assign n16157 = n15868 & n16156 ;
  assign n16158 = ~n15887 & n16155 ;
  assign n16159 = ~n15868 & n16158 ;
  assign n16160 = ~n16157 & ~n16159 ;
  assign n16161 = n15887 & ~n16155 ;
  assign n16162 = ~n15868 & n16161 ;
  assign n16163 = n15887 & n16155 ;
  assign n16164 = n15868 & n16163 ;
  assign n16165 = ~n16162 & ~n16164 ;
  assign n16166 = n16160 & n16165 ;
  assign n16167 = ~n15865 & n16166 ;
  assign n16168 = n3402 & n5105 ;
  assign n16169 = ~n5102 & n16168 ;
  assign n16170 = n3402 & ~n5105 ;
  assign n16171 = ~n4497 & n16170 ;
  assign n16172 = ~n5101 & n16171 ;
  assign n16173 = \b[28]  & n3733 ;
  assign n16174 = n3730 & n16173 ;
  assign n16175 = ~\a[24]  & \b[29]  ;
  assign n16176 = n3394 & n16175 ;
  assign n16177 = ~n16174 & ~n16176 ;
  assign n16178 = \b[30]  & n3400 ;
  assign n16179 = \a[24]  & \b[29]  ;
  assign n16180 = n3391 & n16179 ;
  assign n16181 = \a[26]  & ~n16180 ;
  assign n16182 = ~n16178 & n16181 ;
  assign n16183 = n16177 & n16182 ;
  assign n16184 = ~n16172 & n16183 ;
  assign n16185 = ~n16169 & n16184 ;
  assign n16186 = ~n16178 & ~n16180 ;
  assign n16187 = n16177 & n16186 ;
  assign n16188 = ~n16172 & n16187 ;
  assign n16189 = ~n16169 & n16188 ;
  assign n16190 = ~\a[26]  & ~n16189 ;
  assign n16191 = ~n16185 & ~n16190 ;
  assign n16192 = ~n15618 & ~n16166 ;
  assign n16193 = ~n15864 & n16192 ;
  assign n16194 = ~n16191 & ~n16193 ;
  assign n16195 = ~n16167 & n16194 ;
  assign n16196 = ~n16166 & n16191 ;
  assign n16197 = n15865 & n16196 ;
  assign n16198 = n16166 & n16191 ;
  assign n16199 = ~n15865 & n16198 ;
  assign n16200 = ~n16197 & ~n16199 ;
  assign n16201 = ~n16195 & n16200 ;
  assign n16202 = n2622 & ~n5855 ;
  assign n16203 = ~n5853 & n16202 ;
  assign n16204 = \b[33]  & n2620 ;
  assign n16205 = \a[21]  & \b[32]  ;
  assign n16206 = n2611 & n16205 ;
  assign n16207 = ~n16204 & ~n16206 ;
  assign n16208 = \b[31]  & n2912 ;
  assign n16209 = n2909 & n16208 ;
  assign n16210 = ~\a[21]  & \b[32]  ;
  assign n16211 = n2614 & n16210 ;
  assign n16212 = ~n16209 & ~n16211 ;
  assign n16213 = n16207 & n16212 ;
  assign n16214 = ~n16203 & n16213 ;
  assign n16215 = ~\a[23]  & ~n16214 ;
  assign n16216 = \a[23]  & n16213 ;
  assign n16217 = ~n16203 & n16216 ;
  assign n16218 = ~n16215 & ~n16217 ;
  assign n16219 = ~n16201 & ~n16218 ;
  assign n16220 = n15863 & n16219 ;
  assign n16221 = n16201 & ~n16218 ;
  assign n16222 = ~n15863 & n16221 ;
  assign n16223 = ~n16220 & ~n16222 ;
  assign n16224 = ~n16201 & n16218 ;
  assign n16225 = ~n15863 & n16224 ;
  assign n16226 = n16201 & n16218 ;
  assign n16227 = n15863 & n16226 ;
  assign n16228 = ~n16225 & ~n16227 ;
  assign n16229 = n16223 & n16228 ;
  assign n16230 = ~n15860 & n16229 ;
  assign n16231 = n1965 & n7337 ;
  assign n16232 = ~n7334 & n16231 ;
  assign n16233 = n1965 & ~n7337 ;
  assign n16234 = ~n6605 & n16233 ;
  assign n16235 = ~n7333 & n16234 ;
  assign n16236 = \b[34]  & n2218 ;
  assign n16237 = n2216 & n16236 ;
  assign n16238 = ~\a[18]  & \b[35]  ;
  assign n16239 = n1957 & n16238 ;
  assign n16240 = ~n16237 & ~n16239 ;
  assign n16241 = \b[36]  & n1963 ;
  assign n16242 = \a[18]  & \b[35]  ;
  assign n16243 = n2210 & n16242 ;
  assign n16244 = \a[20]  & ~n16243 ;
  assign n16245 = ~n16241 & n16244 ;
  assign n16246 = n16240 & n16245 ;
  assign n16247 = ~n16235 & n16246 ;
  assign n16248 = ~n16232 & n16247 ;
  assign n16249 = ~n16241 & ~n16243 ;
  assign n16250 = n16240 & n16249 ;
  assign n16251 = ~n16235 & n16250 ;
  assign n16252 = ~n16232 & n16251 ;
  assign n16253 = ~\a[20]  & ~n16252 ;
  assign n16254 = ~n16248 & ~n16253 ;
  assign n16255 = ~n15640 & ~n16229 ;
  assign n16256 = ~n15859 & n16255 ;
  assign n16257 = ~n16254 & ~n16256 ;
  assign n16258 = ~n16230 & n16257 ;
  assign n16259 = ~n16229 & n16254 ;
  assign n16260 = n15860 & n16259 ;
  assign n16261 = n16229 & n16254 ;
  assign n16262 = ~n15860 & n16261 ;
  assign n16263 = ~n16260 & ~n16262 ;
  assign n16264 = ~n16258 & n16263 ;
  assign n16265 = ~n15858 & ~n16264 ;
  assign n16266 = n15858 & n16264 ;
  assign n16267 = ~n16265 & ~n16266 ;
  assign n16268 = n1467 & ~n8602 ;
  assign n16269 = ~n8600 & n16268 ;
  assign n16270 = \b[39]  & n1465 ;
  assign n16271 = \a[15]  & \b[38]  ;
  assign n16272 = n1456 & n16271 ;
  assign n16273 = ~n16270 & ~n16272 ;
  assign n16274 = \b[37]  & n1652 ;
  assign n16275 = n1649 & n16274 ;
  assign n16276 = ~\a[15]  & \b[38]  ;
  assign n16277 = n1459 & n16276 ;
  assign n16278 = ~n16275 & ~n16277 ;
  assign n16279 = n16273 & n16278 ;
  assign n16280 = ~n16269 & n16279 ;
  assign n16281 = ~\a[17]  & ~n16280 ;
  assign n16282 = \a[17]  & n16279 ;
  assign n16283 = ~n16269 & n16282 ;
  assign n16284 = ~n16281 & ~n16283 ;
  assign n16285 = n16267 & ~n16284 ;
  assign n16286 = ~n16267 & n16284 ;
  assign n16287 = ~n16285 & ~n16286 ;
  assign n16288 = n999 & n9930 ;
  assign n16289 = ~n9927 & n16288 ;
  assign n16290 = n999 & ~n9930 ;
  assign n16291 = ~n9477 & n16290 ;
  assign n16292 = ~n9926 & n16291 ;
  assign n16293 = \b[40]  & n1182 ;
  assign n16294 = n1179 & n16293 ;
  assign n16295 = \b[42]  & n997 ;
  assign n16296 = \a[11]  & \b[41]  ;
  assign n16297 = n1180 & n16296 ;
  assign n16298 = ~\a[12]  & \b[41]  ;
  assign n16299 = n7674 & n16298 ;
  assign n16300 = ~n16297 & ~n16299 ;
  assign n16301 = ~n16295 & n16300 ;
  assign n16302 = ~n16294 & n16301 ;
  assign n16303 = ~n16292 & n16302 ;
  assign n16304 = ~n16289 & n16303 ;
  assign n16305 = ~\a[14]  & ~n16304 ;
  assign n16306 = \a[14]  & n16302 ;
  assign n16307 = ~n16292 & n16306 ;
  assign n16308 = ~n16289 & n16307 ;
  assign n16309 = ~n16305 & ~n16308 ;
  assign n16310 = ~n16287 & n16309 ;
  assign n16311 = n15855 & n16310 ;
  assign n16312 = n16287 & n16309 ;
  assign n16313 = ~n15855 & n16312 ;
  assign n16314 = ~n16311 & ~n16313 ;
  assign n16315 = ~n16287 & ~n16309 ;
  assign n16316 = ~n15855 & n16315 ;
  assign n16317 = n16287 & ~n16309 ;
  assign n16318 = n15855 & n16317 ;
  assign n16319 = ~n16316 & ~n16318 ;
  assign n16320 = n16314 & n16319 ;
  assign n16321 = ~n15853 & ~n16320 ;
  assign n16322 = n15836 & n16321 ;
  assign n16323 = ~n15853 & n16320 ;
  assign n16324 = ~n15836 & n16323 ;
  assign n16325 = ~n16322 & ~n16324 ;
  assign n16326 = n15853 & ~n16320 ;
  assign n16327 = ~n15836 & n16326 ;
  assign n16328 = n15853 & n16320 ;
  assign n16329 = n15836 & n16328 ;
  assign n16330 = ~n16327 & ~n16329 ;
  assign n16331 = n16325 & n16330 ;
  assign n16332 = ~n15833 & n16331 ;
  assign n16333 = n430 & n12478 ;
  assign n16334 = ~n12475 & n16333 ;
  assign n16335 = n430 & ~n12478 ;
  assign n16336 = ~n12433 & n16335 ;
  assign n16337 = ~n12474 & n16336 ;
  assign n16338 = \b[46]  & n486 ;
  assign n16339 = n483 & n16338 ;
  assign n16340 = ~\a[6]  & \b[47]  ;
  assign n16341 = n422 & n16340 ;
  assign n16342 = ~n16339 & ~n16341 ;
  assign n16343 = \b[48]  & n428 ;
  assign n16344 = \a[6]  & \b[47]  ;
  assign n16345 = n419 & n16344 ;
  assign n16346 = \a[8]  & ~n16345 ;
  assign n16347 = ~n16343 & n16346 ;
  assign n16348 = n16342 & n16347 ;
  assign n16349 = ~n16337 & n16348 ;
  assign n16350 = ~n16334 & n16349 ;
  assign n16351 = ~n16343 & ~n16345 ;
  assign n16352 = n16342 & n16351 ;
  assign n16353 = ~n16337 & n16352 ;
  assign n16354 = ~n16334 & n16353 ;
  assign n16355 = ~\a[8]  & ~n16354 ;
  assign n16356 = ~n16350 & ~n16355 ;
  assign n16357 = ~n15756 & ~n16331 ;
  assign n16358 = ~n15832 & n16357 ;
  assign n16359 = ~n16356 & ~n16358 ;
  assign n16360 = ~n16332 & n16359 ;
  assign n16361 = ~n16331 & n16356 ;
  assign n16362 = n15833 & n16361 ;
  assign n16363 = n16331 & n16356 ;
  assign n16364 = ~n15833 & n16363 ;
  assign n16365 = ~n16362 & ~n16364 ;
  assign n16366 = ~n16360 & n16365 ;
  assign n16367 = n252 & ~n14098 ;
  assign n16368 = ~n14096 & n16367 ;
  assign n16369 = \b[51]  & n250 ;
  assign n16370 = \a[3]  & \b[50]  ;
  assign n16371 = n241 & n16370 ;
  assign n16372 = ~n16369 & ~n16371 ;
  assign n16373 = \b[49]  & n303 ;
  assign n16374 = n300 & n16373 ;
  assign n16375 = ~\a[3]  & \b[50]  ;
  assign n16376 = n244 & n16375 ;
  assign n16377 = ~n16374 & ~n16376 ;
  assign n16378 = n16372 & n16377 ;
  assign n16379 = ~n16368 & n16378 ;
  assign n16380 = ~\a[5]  & ~n16379 ;
  assign n16381 = \a[5]  & n16378 ;
  assign n16382 = ~n16368 & n16381 ;
  assign n16383 = ~n16380 & ~n16382 ;
  assign n16384 = ~n16366 & n16383 ;
  assign n16385 = ~n15831 & n16384 ;
  assign n16386 = n16366 & n16383 ;
  assign n16387 = n15831 & n16386 ;
  assign n16388 = ~n16385 & ~n16387 ;
  assign n16389 = ~n16366 & ~n16383 ;
  assign n16390 = n15831 & n16389 ;
  assign n16391 = n16366 & ~n16383 ;
  assign n16392 = ~n15831 & n16391 ;
  assign n16393 = ~n16390 & ~n16392 ;
  assign n16394 = n16388 & n16393 ;
  assign n16395 = ~n15828 & n16394 ;
  assign n16396 = ~\b[53]  & ~\b[54]  ;
  assign n16397 = \b[53]  & \b[54]  ;
  assign n16398 = ~n16396 & ~n16397 ;
  assign n16399 = n15241 & ~n16398 ;
  assign n16400 = ~n15200 & ~n15242 ;
  assign n16401 = ~n16398 & n16400 ;
  assign n16402 = ~n15239 & n16401 ;
  assign n16403 = ~n16399 & ~n16402 ;
  assign n16404 = ~n15239 & n16400 ;
  assign n16405 = ~n15241 & n16398 ;
  assign n16406 = ~n16404 & n16405 ;
  assign n16407 = n16403 & ~n16406 ;
  assign n16408 = n134 & n16407 ;
  assign n16409 = \a[0]  & \b[54]  ;
  assign n16410 = n133 & n16409 ;
  assign n16411 = \b[53]  & n141 ;
  assign n16412 = ~\a[1]  & \b[52]  ;
  assign n16413 = n10416 & n16412 ;
  assign n16414 = ~n16411 & ~n16413 ;
  assign n16415 = ~n16410 & n16414 ;
  assign n16416 = \a[2]  & n16415 ;
  assign n16417 = ~n16408 & n16416 ;
  assign n16418 = ~\a[2]  & ~n16415 ;
  assign n16419 = ~\a[2]  & n134 ;
  assign n16420 = n16407 & n16419 ;
  assign n16421 = ~n16418 & ~n16420 ;
  assign n16422 = ~n16417 & n16421 ;
  assign n16423 = ~n15802 & ~n16394 ;
  assign n16424 = ~n15827 & n16423 ;
  assign n16425 = ~n16422 & ~n16424 ;
  assign n16426 = ~n16395 & n16425 ;
  assign n16427 = ~n16394 & n16422 ;
  assign n16428 = n15828 & n16427 ;
  assign n16429 = n16394 & n16422 ;
  assign n16430 = ~n15828 & n16429 ;
  assign n16431 = ~n16428 & ~n16430 ;
  assign n16432 = ~n16426 & n16431 ;
  assign n16433 = n15826 & n16432 ;
  assign n16434 = ~n15826 & ~n16432 ;
  assign n16435 = ~n16433 & ~n16434 ;
  assign n16436 = ~n16426 & ~n16433 ;
  assign n16437 = ~n15802 & n16393 ;
  assign n16438 = ~n15827 & n16437 ;
  assign n16439 = n16388 & ~n16438 ;
  assign n16440 = ~n16397 & ~n16406 ;
  assign n16441 = ~\b[54]  & ~\b[55]  ;
  assign n16442 = \b[54]  & \b[55]  ;
  assign n16443 = ~n16441 & ~n16442 ;
  assign n16444 = ~n16440 & n16443 ;
  assign n16445 = ~n16397 & ~n16443 ;
  assign n16446 = ~n16406 & n16445 ;
  assign n16447 = n134 & ~n16446 ;
  assign n16448 = ~n16444 & n16447 ;
  assign n16449 = \a[0]  & \b[55]  ;
  assign n16450 = n133 & n16449 ;
  assign n16451 = \b[54]  & n141 ;
  assign n16452 = ~\a[1]  & \b[53]  ;
  assign n16453 = n10416 & n16452 ;
  assign n16454 = ~n16451 & ~n16453 ;
  assign n16455 = ~n16450 & n16454 ;
  assign n16456 = ~n16448 & n16455 ;
  assign n16457 = ~\a[2]  & ~n16456 ;
  assign n16458 = \a[2]  & n16455 ;
  assign n16459 = ~n16448 & n16458 ;
  assign n16460 = ~n16457 & ~n16459 ;
  assign n16461 = n15831 & n16366 ;
  assign n16462 = ~n16360 & ~n16461 ;
  assign n16463 = ~n15756 & n16325 ;
  assign n16464 = ~n15832 & n16463 ;
  assign n16465 = n16330 & ~n16464 ;
  assign n16466 = n430 & ~n13524 ;
  assign n16467 = ~n13522 & n16466 ;
  assign n16468 = \b[49]  & n428 ;
  assign n16469 = \a[6]  & \b[48]  ;
  assign n16470 = n419 & n16469 ;
  assign n16471 = ~n16468 & ~n16470 ;
  assign n16472 = \b[47]  & n486 ;
  assign n16473 = n483 & n16472 ;
  assign n16474 = ~\a[6]  & \b[48]  ;
  assign n16475 = n422 & n16474 ;
  assign n16476 = ~n16473 & ~n16475 ;
  assign n16477 = n16471 & n16476 ;
  assign n16478 = ~n16467 & n16477 ;
  assign n16479 = ~\a[8]  & ~n16478 ;
  assign n16480 = \a[8]  & n16477 ;
  assign n16481 = ~n16467 & n16480 ;
  assign n16482 = ~n16479 & ~n16481 ;
  assign n16483 = n15836 & n16320 ;
  assign n16484 = n16319 & ~n16483 ;
  assign n16485 = n646 & n11906 ;
  assign n16486 = ~n11903 & n16485 ;
  assign n16487 = n646 & n13483 ;
  assign n16488 = ~n11902 & n16487 ;
  assign n16489 = \b[44]  & n796 ;
  assign n16490 = n793 & n16489 ;
  assign n16491 = ~\a[9]  & \b[45]  ;
  assign n16492 = n638 & n16491 ;
  assign n16493 = ~n16490 & ~n16492 ;
  assign n16494 = \b[46]  & n644 ;
  assign n16495 = \a[9]  & \b[45]  ;
  assign n16496 = n635 & n16495 ;
  assign n16497 = \a[11]  & ~n16496 ;
  assign n16498 = ~n16494 & n16497 ;
  assign n16499 = n16493 & n16498 ;
  assign n16500 = ~n16488 & n16499 ;
  assign n16501 = ~n16486 & n16500 ;
  assign n16502 = ~n16494 & ~n16496 ;
  assign n16503 = n16493 & n16502 ;
  assign n16504 = ~n16488 & n16503 ;
  assign n16505 = ~n16486 & n16504 ;
  assign n16506 = ~\a[11]  & ~n16505 ;
  assign n16507 = ~n16501 & ~n16506 ;
  assign n16508 = n15698 & ~n16285 ;
  assign n16509 = ~n15854 & n16508 ;
  assign n16510 = ~n16286 & ~n16509 ;
  assign n16511 = ~n16258 & ~n16266 ;
  assign n16512 = ~n15640 & n16223 ;
  assign n16513 = ~n15859 & n16512 ;
  assign n16514 = n16228 & ~n16513 ;
  assign n16515 = n15863 & n16201 ;
  assign n16516 = ~n16195 & ~n16515 ;
  assign n16517 = ~n15618 & n16160 ;
  assign n16518 = ~n15864 & n16517 ;
  assign n16519 = n16165 & ~n16518 ;
  assign n16520 = n15868 & n16155 ;
  assign n16521 = n16149 & ~n16520 ;
  assign n16522 = n15591 & ~n16142 ;
  assign n16523 = ~n15888 & n16522 ;
  assign n16524 = ~n16143 & ~n16523 ;
  assign n16525 = ~n16132 & ~n16139 ;
  assign n16526 = n2768 & n6309 ;
  assign n16527 = ~n2765 & n16526 ;
  assign n16528 = n6309 & n6462 ;
  assign n16529 = ~n2764 & n16528 ;
  assign n16530 = \b[20]  & n6778 ;
  assign n16531 = n6775 & n16530 ;
  assign n16532 = ~\a[33]  & \b[21]  ;
  assign n16533 = n6301 & n16532 ;
  assign n16534 = ~n16531 & ~n16533 ;
  assign n16535 = \b[22]  & n6307 ;
  assign n16536 = \a[33]  & \b[21]  ;
  assign n16537 = n6298 & n16536 ;
  assign n16538 = \a[35]  & ~n16537 ;
  assign n16539 = ~n16535 & n16538 ;
  assign n16540 = n16534 & n16539 ;
  assign n16541 = ~n16529 & n16540 ;
  assign n16542 = ~n16527 & n16541 ;
  assign n16543 = ~n16535 & ~n16537 ;
  assign n16544 = n16534 & n16543 ;
  assign n16545 = ~n16529 & n16544 ;
  assign n16546 = ~n16527 & n16545 ;
  assign n16547 = ~\a[35]  & ~n16546 ;
  assign n16548 = ~n16542 & ~n16547 ;
  assign n16549 = n15569 & n16100 ;
  assign n16550 = ~n15941 & n16549 ;
  assign n16551 = n16105 & ~n16550 ;
  assign n16552 = n15945 & n16095 ;
  assign n16553 = ~n16089 & ~n16552 ;
  assign n16554 = ~n15534 & n16054 ;
  assign n16555 = ~n15536 & n16554 ;
  assign n16556 = n16059 & ~n16555 ;
  assign n16557 = ~n948 & n10082 ;
  assign n16558 = ~n908 & n10082 ;
  assign n16559 = ~n912 & n16558 ;
  assign n16560 = ~n16557 & ~n16559 ;
  assign n16561 = ~n951 & ~n16560 ;
  assign n16562 = \b[11]  & n10681 ;
  assign n16563 = n10678 & n16562 ;
  assign n16564 = ~\a[42]  & \b[12]  ;
  assign n16565 = n10074 & n16564 ;
  assign n16566 = ~n16563 & ~n16565 ;
  assign n16567 = \b[13]  & n10080 ;
  assign n16568 = \a[42]  & \b[12]  ;
  assign n16569 = n10071 & n16568 ;
  assign n16570 = \a[44]  & ~n16569 ;
  assign n16571 = ~n16567 & n16570 ;
  assign n16572 = n16566 & n16571 ;
  assign n16573 = ~n16561 & n16572 ;
  assign n16574 = ~n16567 & ~n16569 ;
  assign n16575 = n16566 & n16574 ;
  assign n16576 = ~\a[44]  & ~n16575 ;
  assign n16577 = ~\a[44]  & ~n951 ;
  assign n16578 = ~n16560 & n16577 ;
  assign n16579 = ~n16576 & ~n16578 ;
  assign n16580 = ~n16573 & n16579 ;
  assign n16581 = n15973 & n16049 ;
  assign n16582 = ~n16047 & ~n16581 ;
  assign n16583 = n685 & n11572 ;
  assign n16584 = ~n682 & n16583 ;
  assign n16585 = n11572 & n11610 ;
  assign n16586 = ~n681 & n16585 ;
  assign n16587 = \b[8]  & n12159 ;
  assign n16588 = n12156 & n16587 ;
  assign n16589 = ~\a[45]  & \b[9]  ;
  assign n16590 = n11564 & n16589 ;
  assign n16591 = ~n16588 & ~n16590 ;
  assign n16592 = \b[10]  & n11570 ;
  assign n16593 = \a[45]  & \b[9]  ;
  assign n16594 = n11561 & n16593 ;
  assign n16595 = \a[47]  & ~n16594 ;
  assign n16596 = ~n16592 & n16595 ;
  assign n16597 = n16591 & n16596 ;
  assign n16598 = ~n16586 & n16597 ;
  assign n16599 = ~n16584 & n16598 ;
  assign n16600 = ~n16592 & ~n16594 ;
  assign n16601 = n16591 & n16600 ;
  assign n16602 = ~n16586 & n16601 ;
  assign n16603 = ~n16584 & n16602 ;
  assign n16604 = ~\a[47]  & ~n16603 ;
  assign n16605 = ~n16599 & ~n16604 ;
  assign n16606 = ~n383 & n13125 ;
  assign n16607 = ~n381 & n16606 ;
  assign n16608 = \b[5]  & n13794 ;
  assign n16609 = n13792 & n16608 ;
  assign n16610 = \b[7]  & n13123 ;
  assign n16611 = \a[48]  & \b[6]  ;
  assign n16612 = n13786 & n16611 ;
  assign n16613 = ~\a[48]  & \b[6]  ;
  assign n16614 = n13117 & n16613 ;
  assign n16615 = ~n16612 & ~n16614 ;
  assign n16616 = ~n16610 & n16615 ;
  assign n16617 = ~n16609 & n16616 ;
  assign n16618 = ~\a[50]  & n16617 ;
  assign n16619 = ~n16607 & n16618 ;
  assign n16620 = ~n16607 & n16617 ;
  assign n16621 = \a[50]  & ~n16620 ;
  assign n16622 = ~n16619 & ~n16621 ;
  assign n16623 = ~n16019 & ~n16022 ;
  assign n16624 = n222 & n14793 ;
  assign n16625 = \b[4]  & n14791 ;
  assign n16626 = \a[50]  & \b[3]  ;
  assign n16627 = n15515 & n16626 ;
  assign n16628 = ~\a[51]  & \b[3]  ;
  assign n16629 = n14785 & n16628 ;
  assign n16630 = ~n16627 & ~n16629 ;
  assign n16631 = ~n16625 & n16630 ;
  assign n16632 = \b[2]  & n15517 ;
  assign n16633 = n15514 & n16632 ;
  assign n16634 = \a[53]  & ~n16633 ;
  assign n16635 = n16631 & n16634 ;
  assign n16636 = ~n16624 & n16635 ;
  assign n16637 = n16631 & ~n16633 ;
  assign n16638 = ~n16624 & n16637 ;
  assign n16639 = ~\a[53]  & ~n16638 ;
  assign n16640 = ~n16636 & ~n16639 ;
  assign n16641 = \a[56]  & \b[0]  ;
  assign n16642 = ~n16016 & n16641 ;
  assign n16643 = \a[54]  & \b[0]  ;
  assign n16644 = \a[53]  & ~\a[55]  ;
  assign n16645 = n16643 & n16644 ;
  assign n16646 = ~\a[54]  & \b[0]  ;
  assign n16647 = ~\a[53]  & \a[55]  ;
  assign n16648 = n16646 & n16647 ;
  assign n16649 = ~n16645 & ~n16648 ;
  assign n16650 = \a[55]  & ~\a[56]  ;
  assign n16651 = ~\a[55]  & \a[56]  ;
  assign n16652 = ~n16650 & ~n16651 ;
  assign n16653 = ~n16016 & n16652 ;
  assign n16654 = \b[1]  & n16653 ;
  assign n16655 = ~n16016 & ~n16652 ;
  assign n16656 = ~n137 & n16655 ;
  assign n16657 = ~n16654 & ~n16656 ;
  assign n16658 = n16649 & n16657 ;
  assign n16659 = n16642 & ~n16658 ;
  assign n16660 = ~n16642 & n16649 ;
  assign n16661 = n16657 & n16660 ;
  assign n16662 = ~n16659 & ~n16661 ;
  assign n16663 = n16640 & ~n16662 ;
  assign n16664 = ~n16640 & n16662 ;
  assign n16665 = ~n16663 & ~n16664 ;
  assign n16666 = ~n16623 & n16665 ;
  assign n16667 = n16623 & ~n16665 ;
  assign n16668 = ~n16666 & ~n16667 ;
  assign n16669 = ~n16622 & ~n16668 ;
  assign n16670 = n16622 & n16668 ;
  assign n16671 = ~n16669 & ~n16670 ;
  assign n16672 = n16605 & ~n16671 ;
  assign n16673 = n16582 & n16672 ;
  assign n16674 = n16605 & n16671 ;
  assign n16675 = ~n16582 & n16674 ;
  assign n16676 = ~n16673 & ~n16675 ;
  assign n16677 = ~n16605 & ~n16671 ;
  assign n16678 = ~n16582 & n16677 ;
  assign n16679 = ~n16605 & n16671 ;
  assign n16680 = n16582 & n16679 ;
  assign n16681 = ~n16678 & ~n16680 ;
  assign n16682 = n16676 & n16681 ;
  assign n16683 = n16580 & ~n16682 ;
  assign n16684 = ~n16556 & n16683 ;
  assign n16685 = n16580 & n16682 ;
  assign n16686 = n16556 & n16685 ;
  assign n16687 = ~n16684 & ~n16686 ;
  assign n16688 = ~n16580 & ~n16682 ;
  assign n16689 = n16556 & n16688 ;
  assign n16690 = ~n16580 & n16682 ;
  assign n16691 = ~n16556 & n16690 ;
  assign n16692 = ~n16689 & ~n16691 ;
  assign n16693 = n16687 & n16692 ;
  assign n16694 = ~n16553 & n16693 ;
  assign n16695 = ~n16089 & ~n16693 ;
  assign n16696 = ~n16552 & n16695 ;
  assign n16697 = n1512 & n8759 ;
  assign n16698 = ~n1509 & n16697 ;
  assign n16699 = n8759 & n10165 ;
  assign n16700 = ~n1508 & n16699 ;
  assign n16701 = \b[14]  & n9301 ;
  assign n16702 = n9298 & n16701 ;
  assign n16703 = ~\a[39]  & \b[15]  ;
  assign n16704 = n8751 & n16703 ;
  assign n16705 = ~n16702 & ~n16704 ;
  assign n16706 = \b[16]  & n8757 ;
  assign n16707 = \a[39]  & \b[15]  ;
  assign n16708 = n8748 & n16707 ;
  assign n16709 = \a[41]  & ~n16708 ;
  assign n16710 = ~n16706 & n16709 ;
  assign n16711 = n16705 & n16710 ;
  assign n16712 = ~n16700 & n16711 ;
  assign n16713 = ~n16698 & n16712 ;
  assign n16714 = ~n16706 & ~n16708 ;
  assign n16715 = n16705 & n16714 ;
  assign n16716 = ~n16700 & n16715 ;
  assign n16717 = ~n16698 & n16716 ;
  assign n16718 = ~\a[41]  & ~n16717 ;
  assign n16719 = ~n16713 & ~n16718 ;
  assign n16720 = ~n16696 & ~n16719 ;
  assign n16721 = ~n16694 & n16720 ;
  assign n16722 = ~n16693 & n16719 ;
  assign n16723 = n16553 & n16722 ;
  assign n16724 = n16693 & n16719 ;
  assign n16725 = ~n16553 & n16724 ;
  assign n16726 = ~n16723 & ~n16725 ;
  assign n16727 = ~n16721 & n16726 ;
  assign n16728 = ~n2076 & n7534 ;
  assign n16729 = ~n1874 & n7534 ;
  assign n16730 = ~n1878 & n16729 ;
  assign n16731 = ~n16728 & ~n16730 ;
  assign n16732 = ~n2079 & ~n16731 ;
  assign n16733 = \b[17]  & n7973 ;
  assign n16734 = n7970 & n16733 ;
  assign n16735 = \b[19]  & n7532 ;
  assign n16736 = \a[36]  & \b[18]  ;
  assign n16737 = n7523 & n16736 ;
  assign n16738 = ~\a[36]  & \b[18]  ;
  assign n16739 = n7526 & n16738 ;
  assign n16740 = ~n16737 & ~n16739 ;
  assign n16741 = ~n16735 & n16740 ;
  assign n16742 = ~n16734 & n16741 ;
  assign n16743 = ~\a[38]  & n16742 ;
  assign n16744 = ~n16732 & n16743 ;
  assign n16745 = \a[38]  & ~n16742 ;
  assign n16746 = \a[38]  & ~n2079 ;
  assign n16747 = ~n16731 & n16746 ;
  assign n16748 = ~n16745 & ~n16747 ;
  assign n16749 = ~n16744 & n16748 ;
  assign n16750 = ~n16727 & n16749 ;
  assign n16751 = n16551 & n16750 ;
  assign n16752 = n16727 & n16749 ;
  assign n16753 = ~n16551 & n16752 ;
  assign n16754 = ~n16751 & ~n16753 ;
  assign n16755 = ~n16727 & ~n16749 ;
  assign n16756 = ~n16551 & n16755 ;
  assign n16757 = n16727 & ~n16749 ;
  assign n16758 = n16551 & n16757 ;
  assign n16759 = ~n16756 & ~n16758 ;
  assign n16760 = n16754 & n16759 ;
  assign n16761 = ~n16548 & ~n16760 ;
  assign n16762 = ~n16525 & n16761 ;
  assign n16763 = ~n16548 & n16760 ;
  assign n16764 = n16525 & n16763 ;
  assign n16765 = ~n16762 & ~n16764 ;
  assign n16766 = n16548 & ~n16760 ;
  assign n16767 = n16525 & n16766 ;
  assign n16768 = n16548 & n16760 ;
  assign n16769 = ~n16525 & n16768 ;
  assign n16770 = ~n16767 & ~n16769 ;
  assign n16771 = n16765 & n16770 ;
  assign n16772 = ~n3567 & n5211 ;
  assign n16773 = ~n3565 & n16772 ;
  assign n16774 = \b[25]  & n5209 ;
  assign n16775 = \a[30]  & \b[24]  ;
  assign n16776 = n5200 & n16775 ;
  assign n16777 = ~n16774 & ~n16776 ;
  assign n16778 = \b[23]  & n5595 ;
  assign n16779 = n5592 & n16778 ;
  assign n16780 = ~\a[30]  & \b[24]  ;
  assign n16781 = n5203 & n16780 ;
  assign n16782 = ~n16779 & ~n16781 ;
  assign n16783 = n16777 & n16782 ;
  assign n16784 = ~n16773 & n16783 ;
  assign n16785 = ~\a[32]  & ~n16784 ;
  assign n16786 = \a[32]  & n16783 ;
  assign n16787 = ~n16773 & n16786 ;
  assign n16788 = ~n16785 & ~n16787 ;
  assign n16789 = ~n16771 & ~n16788 ;
  assign n16790 = n16524 & n16789 ;
  assign n16791 = n16771 & ~n16788 ;
  assign n16792 = ~n16524 & n16791 ;
  assign n16793 = ~n16790 & ~n16792 ;
  assign n16794 = ~n16771 & n16788 ;
  assign n16795 = ~n16524 & n16794 ;
  assign n16796 = n16771 & n16788 ;
  assign n16797 = n16524 & n16796 ;
  assign n16798 = ~n16795 & ~n16797 ;
  assign n16799 = n16793 & n16798 ;
  assign n16800 = ~n16521 & n16799 ;
  assign n16801 = n16149 & ~n16799 ;
  assign n16802 = ~n16520 & n16801 ;
  assign n16803 = n4249 & n4456 ;
  assign n16804 = ~n4453 & n16803 ;
  assign n16805 = ~n4143 & ~n4456 ;
  assign n16806 = n4249 & n16805 ;
  assign n16807 = ~n4452 & n16806 ;
  assign n16808 = \b[26]  & n4647 ;
  assign n16809 = n4644 & n16808 ;
  assign n16810 = ~\a[27]  & \b[27]  ;
  assign n16811 = n4241 & n16810 ;
  assign n16812 = ~n16809 & ~n16811 ;
  assign n16813 = \b[28]  & n4247 ;
  assign n16814 = \a[27]  & \b[27]  ;
  assign n16815 = n4238 & n16814 ;
  assign n16816 = \a[29]  & ~n16815 ;
  assign n16817 = ~n16813 & n16816 ;
  assign n16818 = n16812 & n16817 ;
  assign n16819 = ~n16807 & n16818 ;
  assign n16820 = ~n16804 & n16819 ;
  assign n16821 = ~n16813 & ~n16815 ;
  assign n16822 = n16812 & n16821 ;
  assign n16823 = ~n16807 & n16822 ;
  assign n16824 = ~n16804 & n16823 ;
  assign n16825 = ~\a[29]  & ~n16824 ;
  assign n16826 = ~n16820 & ~n16825 ;
  assign n16827 = ~n16802 & ~n16826 ;
  assign n16828 = ~n16800 & n16827 ;
  assign n16829 = ~n16799 & n16826 ;
  assign n16830 = n16521 & n16829 ;
  assign n16831 = n16799 & n16826 ;
  assign n16832 = ~n16521 & n16831 ;
  assign n16833 = ~n16830 & ~n16832 ;
  assign n16834 = ~n16828 & n16833 ;
  assign n16835 = n3402 & ~n5462 ;
  assign n16836 = ~n5460 & n16835 ;
  assign n16837 = \b[31]  & n3400 ;
  assign n16838 = \a[24]  & \b[30]  ;
  assign n16839 = n3391 & n16838 ;
  assign n16840 = ~n16837 & ~n16839 ;
  assign n16841 = \b[29]  & n3733 ;
  assign n16842 = n3730 & n16841 ;
  assign n16843 = ~\a[24]  & \b[30]  ;
  assign n16844 = n3394 & n16843 ;
  assign n16845 = ~n16842 & ~n16844 ;
  assign n16846 = n16840 & n16845 ;
  assign n16847 = ~n16836 & n16846 ;
  assign n16848 = ~\a[26]  & ~n16847 ;
  assign n16849 = \a[26]  & n16846 ;
  assign n16850 = ~n16836 & n16849 ;
  assign n16851 = ~n16848 & ~n16850 ;
  assign n16852 = ~n16834 & ~n16851 ;
  assign n16853 = n16519 & n16852 ;
  assign n16854 = n16834 & ~n16851 ;
  assign n16855 = ~n16519 & n16854 ;
  assign n16856 = ~n16853 & ~n16855 ;
  assign n16857 = ~n16834 & n16851 ;
  assign n16858 = ~n16519 & n16857 ;
  assign n16859 = n16834 & n16851 ;
  assign n16860 = n16519 & n16859 ;
  assign n16861 = ~n16858 & ~n16860 ;
  assign n16862 = n16856 & n16861 ;
  assign n16863 = ~n16516 & n16862 ;
  assign n16864 = ~n16195 & ~n16862 ;
  assign n16865 = ~n16515 & n16864 ;
  assign n16866 = n2622 & n6565 ;
  assign n16867 = ~n6562 & n16866 ;
  assign n16868 = n2622 & ~n6565 ;
  assign n16869 = ~n5850 & n16868 ;
  assign n16870 = ~n6561 & n16869 ;
  assign n16871 = \b[32]  & n2912 ;
  assign n16872 = n2909 & n16871 ;
  assign n16873 = ~\a[21]  & \b[33]  ;
  assign n16874 = n2614 & n16873 ;
  assign n16875 = ~n16872 & ~n16874 ;
  assign n16876 = \b[34]  & n2620 ;
  assign n16877 = \a[21]  & \b[33]  ;
  assign n16878 = n2611 & n16877 ;
  assign n16879 = \a[23]  & ~n16878 ;
  assign n16880 = ~n16876 & n16879 ;
  assign n16881 = n16875 & n16880 ;
  assign n16882 = ~n16870 & n16881 ;
  assign n16883 = ~n16867 & n16882 ;
  assign n16884 = ~n16876 & ~n16878 ;
  assign n16885 = n16875 & n16884 ;
  assign n16886 = ~n16870 & n16885 ;
  assign n16887 = ~n16867 & n16886 ;
  assign n16888 = ~\a[23]  & ~n16887 ;
  assign n16889 = ~n16883 & ~n16888 ;
  assign n16890 = ~n16865 & ~n16889 ;
  assign n16891 = ~n16863 & n16890 ;
  assign n16892 = ~n16862 & n16889 ;
  assign n16893 = n16516 & n16892 ;
  assign n16894 = n16862 & n16889 ;
  assign n16895 = ~n16516 & n16894 ;
  assign n16896 = ~n16893 & ~n16895 ;
  assign n16897 = ~n16891 & n16896 ;
  assign n16898 = n1965 & ~n7761 ;
  assign n16899 = ~n7759 & n16898 ;
  assign n16900 = \b[37]  & n1963 ;
  assign n16901 = \a[18]  & \b[36]  ;
  assign n16902 = n2210 & n16901 ;
  assign n16903 = ~n16900 & ~n16902 ;
  assign n16904 = \b[35]  & n2218 ;
  assign n16905 = n2216 & n16904 ;
  assign n16906 = ~\a[18]  & \b[36]  ;
  assign n16907 = n1957 & n16906 ;
  assign n16908 = ~n16905 & ~n16907 ;
  assign n16909 = n16903 & n16908 ;
  assign n16910 = ~n16899 & n16909 ;
  assign n16911 = ~\a[20]  & ~n16910 ;
  assign n16912 = \a[20]  & n16909 ;
  assign n16913 = ~n16899 & n16912 ;
  assign n16914 = ~n16911 & ~n16913 ;
  assign n16915 = ~n16897 & ~n16914 ;
  assign n16916 = n16514 & n16915 ;
  assign n16917 = n16897 & ~n16914 ;
  assign n16918 = ~n16514 & n16917 ;
  assign n16919 = ~n16916 & ~n16918 ;
  assign n16920 = ~n16897 & n16914 ;
  assign n16921 = ~n16514 & n16920 ;
  assign n16922 = n16897 & n16914 ;
  assign n16923 = n16514 & n16922 ;
  assign n16924 = ~n16921 & ~n16923 ;
  assign n16925 = n16919 & n16924 ;
  assign n16926 = n1467 & n9044 ;
  assign n16927 = ~n9041 & n16926 ;
  assign n16928 = n1467 & ~n9044 ;
  assign n16929 = ~n8597 & n16928 ;
  assign n16930 = ~n9040 & n16929 ;
  assign n16931 = \b[38]  & n1652 ;
  assign n16932 = n1649 & n16931 ;
  assign n16933 = ~\a[15]  & \b[39]  ;
  assign n16934 = n1459 & n16933 ;
  assign n16935 = ~n16932 & ~n16934 ;
  assign n16936 = \b[40]  & n1465 ;
  assign n16937 = \a[15]  & \b[39]  ;
  assign n16938 = n1456 & n16937 ;
  assign n16939 = \a[17]  & ~n16938 ;
  assign n16940 = ~n16936 & n16939 ;
  assign n16941 = n16935 & n16940 ;
  assign n16942 = ~n16930 & n16941 ;
  assign n16943 = ~n16927 & n16942 ;
  assign n16944 = ~n16936 & ~n16938 ;
  assign n16945 = n16935 & n16944 ;
  assign n16946 = ~n16930 & n16945 ;
  assign n16947 = ~n16927 & n16946 ;
  assign n16948 = ~\a[17]  & ~n16947 ;
  assign n16949 = ~n16943 & ~n16948 ;
  assign n16950 = ~n16925 & ~n16949 ;
  assign n16951 = ~n16511 & n16950 ;
  assign n16952 = n16925 & ~n16949 ;
  assign n16953 = n16511 & n16952 ;
  assign n16954 = ~n16951 & ~n16953 ;
  assign n16955 = ~n16925 & n16949 ;
  assign n16956 = n16511 & n16955 ;
  assign n16957 = n16925 & n16949 ;
  assign n16958 = ~n16511 & n16957 ;
  assign n16959 = ~n16956 & ~n16958 ;
  assign n16960 = n16954 & n16959 ;
  assign n16961 = n999 & ~n10409 ;
  assign n16962 = ~n10407 & n16961 ;
  assign n16963 = \b[41]  & n1182 ;
  assign n16964 = n1179 & n16963 ;
  assign n16965 = \b[43]  & n997 ;
  assign n16966 = \a[11]  & \b[42]  ;
  assign n16967 = n1180 & n16966 ;
  assign n16968 = ~\a[12]  & \b[42]  ;
  assign n16969 = n7674 & n16968 ;
  assign n16970 = ~n16967 & ~n16969 ;
  assign n16971 = ~n16965 & n16970 ;
  assign n16972 = ~n16964 & n16971 ;
  assign n16973 = ~n16962 & n16972 ;
  assign n16974 = ~\a[14]  & ~n16973 ;
  assign n16975 = \a[14]  & n16972 ;
  assign n16976 = ~n16962 & n16975 ;
  assign n16977 = ~n16974 & ~n16976 ;
  assign n16978 = ~n16960 & ~n16977 ;
  assign n16979 = n16510 & n16978 ;
  assign n16980 = n16960 & ~n16977 ;
  assign n16981 = ~n16510 & n16980 ;
  assign n16982 = ~n16979 & ~n16981 ;
  assign n16983 = ~n16960 & n16977 ;
  assign n16984 = ~n16510 & n16983 ;
  assign n16985 = n16960 & n16977 ;
  assign n16986 = n16510 & n16985 ;
  assign n16987 = ~n16984 & ~n16986 ;
  assign n16988 = n16982 & n16987 ;
  assign n16989 = n16507 & ~n16988 ;
  assign n16990 = n16484 & n16989 ;
  assign n16991 = n16507 & n16988 ;
  assign n16992 = ~n16484 & n16991 ;
  assign n16993 = ~n16990 & ~n16992 ;
  assign n16994 = ~n16484 & n16988 ;
  assign n16995 = n16319 & ~n16988 ;
  assign n16996 = ~n16483 & n16995 ;
  assign n16997 = ~n16507 & ~n16996 ;
  assign n16998 = ~n16994 & n16997 ;
  assign n16999 = n16993 & ~n16998 ;
  assign n17000 = n16482 & ~n16999 ;
  assign n17001 = ~n16465 & n17000 ;
  assign n17002 = n16482 & n16999 ;
  assign n17003 = n16465 & n17002 ;
  assign n17004 = ~n17001 & ~n17003 ;
  assign n17005 = ~n16482 & ~n16999 ;
  assign n17006 = n16465 & n17005 ;
  assign n17007 = ~n16482 & n16999 ;
  assign n17008 = ~n16465 & n17007 ;
  assign n17009 = ~n17006 & ~n17008 ;
  assign n17010 = n17004 & n17009 ;
  assign n17011 = ~n16462 & n17010 ;
  assign n17012 = ~n16360 & ~n17010 ;
  assign n17013 = ~n16461 & n17012 ;
  assign n17014 = n252 & n15201 ;
  assign n17015 = ~n15198 & n17014 ;
  assign n17016 = ~n14093 & ~n15201 ;
  assign n17017 = n252 & n17016 ;
  assign n17018 = ~n15197 & n17017 ;
  assign n17019 = \b[50]  & n303 ;
  assign n17020 = n300 & n17019 ;
  assign n17021 = ~\a[3]  & \b[51]  ;
  assign n17022 = n244 & n17021 ;
  assign n17023 = ~n17020 & ~n17022 ;
  assign n17024 = \b[52]  & n250 ;
  assign n17025 = \a[3]  & \b[51]  ;
  assign n17026 = n241 & n17025 ;
  assign n17027 = \a[5]  & ~n17026 ;
  assign n17028 = ~n17024 & n17027 ;
  assign n17029 = n17023 & n17028 ;
  assign n17030 = ~n17018 & n17029 ;
  assign n17031 = ~n17015 & n17030 ;
  assign n17032 = ~n17024 & ~n17026 ;
  assign n17033 = n17023 & n17032 ;
  assign n17034 = ~n17018 & n17033 ;
  assign n17035 = ~n17015 & n17034 ;
  assign n17036 = ~\a[5]  & ~n17035 ;
  assign n17037 = ~n17031 & ~n17036 ;
  assign n17038 = ~n17013 & ~n17037 ;
  assign n17039 = ~n17011 & n17038 ;
  assign n17040 = ~n17010 & n17037 ;
  assign n17041 = n16462 & n17040 ;
  assign n17042 = n17010 & n17037 ;
  assign n17043 = ~n16462 & n17042 ;
  assign n17044 = ~n17041 & ~n17043 ;
  assign n17045 = ~n17039 & n17044 ;
  assign n17046 = ~n16460 & ~n17045 ;
  assign n17047 = n16439 & n17046 ;
  assign n17048 = ~n16460 & n17045 ;
  assign n17049 = ~n16439 & n17048 ;
  assign n17050 = ~n17047 & ~n17049 ;
  assign n17051 = n16460 & ~n17045 ;
  assign n17052 = ~n16439 & n17051 ;
  assign n17053 = n16460 & n17045 ;
  assign n17054 = n16439 & n17053 ;
  assign n17055 = ~n17052 & ~n17054 ;
  assign n17056 = n17050 & n17055 ;
  assign n17057 = ~n16436 & n17056 ;
  assign n17058 = ~n16426 & ~n17056 ;
  assign n17059 = ~n16433 & n17058 ;
  assign n17060 = ~n17057 & ~n17059 ;
  assign n17061 = ~n16426 & n17050 ;
  assign n17062 = ~n16433 & n17061 ;
  assign n17063 = n17055 & ~n17062 ;
  assign n17064 = n16439 & n17045 ;
  assign n17065 = ~n17039 & ~n17064 ;
  assign n17066 = ~n16360 & n17009 ;
  assign n17067 = ~n16461 & n17066 ;
  assign n17068 = n17004 & ~n17067 ;
  assign n17069 = n252 & ~n15246 ;
  assign n17070 = ~n15244 & n17069 ;
  assign n17071 = \b[53]  & n250 ;
  assign n17072 = \a[3]  & \b[52]  ;
  assign n17073 = n241 & n17072 ;
  assign n17074 = ~n17071 & ~n17073 ;
  assign n17075 = \b[51]  & n303 ;
  assign n17076 = n300 & n17075 ;
  assign n17077 = ~\a[3]  & \b[52]  ;
  assign n17078 = n244 & n17077 ;
  assign n17079 = ~n17076 & ~n17078 ;
  assign n17080 = n17074 & n17079 ;
  assign n17081 = ~n17070 & n17080 ;
  assign n17082 = ~\a[5]  & ~n17081 ;
  assign n17083 = \a[5]  & n17080 ;
  assign n17084 = ~n17070 & n17083 ;
  assign n17085 = ~n17082 & ~n17084 ;
  assign n17086 = n16465 & n16999 ;
  assign n17087 = ~n16998 & ~n17086 ;
  assign n17088 = n16319 & n16982 ;
  assign n17089 = ~n16483 & n17088 ;
  assign n17090 = n16987 & ~n17089 ;
  assign n17091 = n646 & ~n12438 ;
  assign n17092 = ~n12436 & n17091 ;
  assign n17093 = \b[47]  & n644 ;
  assign n17094 = \a[9]  & \b[46]  ;
  assign n17095 = n635 & n17094 ;
  assign n17096 = ~n17093 & ~n17095 ;
  assign n17097 = \b[45]  & n796 ;
  assign n17098 = n793 & n17097 ;
  assign n17099 = ~\a[9]  & \b[46]  ;
  assign n17100 = n638 & n17099 ;
  assign n17101 = ~n17098 & ~n17100 ;
  assign n17102 = n17096 & n17101 ;
  assign n17103 = ~n17092 & n17102 ;
  assign n17104 = ~\a[11]  & ~n17103 ;
  assign n17105 = \a[11]  & n17102 ;
  assign n17106 = ~n17092 & n17105 ;
  assign n17107 = ~n17104 & ~n17106 ;
  assign n17108 = n16510 & n16960 ;
  assign n17109 = n16954 & ~n17108 ;
  assign n17110 = ~n16258 & n16919 ;
  assign n17111 = ~n16266 & n17110 ;
  assign n17112 = n16924 & ~n17111 ;
  assign n17113 = n16514 & n16897 ;
  assign n17114 = ~n16891 & ~n17113 ;
  assign n17115 = ~n16195 & n16856 ;
  assign n17116 = n16861 & ~n17115 ;
  assign n17117 = n16201 & n16861 ;
  assign n17118 = n15863 & n17117 ;
  assign n17119 = ~n17116 & ~n17118 ;
  assign n17120 = n16519 & n16834 ;
  assign n17121 = ~n16828 & ~n17120 ;
  assign n17122 = n3402 & n5810 ;
  assign n17123 = ~n5807 & n17122 ;
  assign n17124 = n3402 & ~n5810 ;
  assign n17125 = ~n5457 & n17124 ;
  assign n17126 = ~n5806 & n17125 ;
  assign n17127 = \b[30]  & n3733 ;
  assign n17128 = n3730 & n17127 ;
  assign n17129 = ~\a[24]  & \b[31]  ;
  assign n17130 = n3394 & n17129 ;
  assign n17131 = ~n17128 & ~n17130 ;
  assign n17132 = \b[32]  & n3400 ;
  assign n17133 = \a[24]  & \b[31]  ;
  assign n17134 = n3391 & n17133 ;
  assign n17135 = \a[26]  & ~n17134 ;
  assign n17136 = ~n17132 & n17135 ;
  assign n17137 = n17131 & n17136 ;
  assign n17138 = ~n17126 & n17137 ;
  assign n17139 = ~n17123 & n17138 ;
  assign n17140 = ~n17132 & ~n17134 ;
  assign n17141 = n17131 & n17140 ;
  assign n17142 = ~n17126 & n17141 ;
  assign n17143 = ~n17123 & n17142 ;
  assign n17144 = ~\a[26]  & ~n17143 ;
  assign n17145 = ~n17139 & ~n17144 ;
  assign n17146 = n16149 & n16793 ;
  assign n17147 = ~n16520 & n17146 ;
  assign n17148 = n16798 & ~n17147 ;
  assign n17149 = n4249 & ~n4502 ;
  assign n17150 = ~n4500 & n17149 ;
  assign n17151 = \b[27]  & n4647 ;
  assign n17152 = n4644 & n17151 ;
  assign n17153 = ~\a[27]  & \b[28]  ;
  assign n17154 = n4241 & n17153 ;
  assign n17155 = ~n17152 & ~n17154 ;
  assign n17156 = \b[29]  & n4247 ;
  assign n17157 = \a[27]  & \b[28]  ;
  assign n17158 = n4238 & n17157 ;
  assign n17159 = \a[29]  & ~n17158 ;
  assign n17160 = ~n17156 & n17159 ;
  assign n17161 = n17155 & n17160 ;
  assign n17162 = ~n17150 & n17161 ;
  assign n17163 = ~n17156 & ~n17158 ;
  assign n17164 = n17155 & n17163 ;
  assign n17165 = ~n17150 & n17164 ;
  assign n17166 = ~\a[29]  & ~n17165 ;
  assign n17167 = ~n17162 & ~n17166 ;
  assign n17168 = n16524 & n16771 ;
  assign n17169 = n16765 & ~n17168 ;
  assign n17170 = ~n3022 & n6309 ;
  assign n17171 = ~n3020 & n17170 ;
  assign n17172 = \b[23]  & n6307 ;
  assign n17173 = \a[33]  & \b[22]  ;
  assign n17174 = n6298 & n17173 ;
  assign n17175 = ~n17172 & ~n17174 ;
  assign n17176 = \b[21]  & n6778 ;
  assign n17177 = n6775 & n17176 ;
  assign n17178 = ~\a[33]  & \b[22]  ;
  assign n17179 = n6301 & n17178 ;
  assign n17180 = ~n17177 & ~n17179 ;
  assign n17181 = n17175 & n17180 ;
  assign n17182 = ~n17171 & n17181 ;
  assign n17183 = ~\a[35]  & ~n17182 ;
  assign n17184 = \a[35]  & n17181 ;
  assign n17185 = ~n17171 & n17184 ;
  assign n17186 = ~n17183 & ~n17185 ;
  assign n17187 = ~n16132 & n16754 ;
  assign n17188 = ~n16139 & n17187 ;
  assign n17189 = n16759 & ~n17188 ;
  assign n17190 = n16551 & n16727 ;
  assign n17191 = ~n16721 & ~n17190 ;
  assign n17192 = ~n16089 & n16692 ;
  assign n17193 = ~n16552 & n17192 ;
  assign n17194 = n16687 & ~n17193 ;
  assign n17195 = ~n1691 & n8759 ;
  assign n17196 = ~n1511 & n8759 ;
  assign n17197 = ~n1515 & n17196 ;
  assign n17198 = ~n17195 & ~n17197 ;
  assign n17199 = ~n1694 & ~n17198 ;
  assign n17200 = \b[15]  & n9301 ;
  assign n17201 = n9298 & n17200 ;
  assign n17202 = ~\a[39]  & \b[16]  ;
  assign n17203 = n8751 & n17202 ;
  assign n17204 = ~n17201 & ~n17203 ;
  assign n17205 = \b[17]  & n8757 ;
  assign n17206 = \a[39]  & \b[16]  ;
  assign n17207 = n8748 & n17206 ;
  assign n17208 = \a[41]  & ~n17207 ;
  assign n17209 = ~n17205 & n17208 ;
  assign n17210 = n17204 & n17209 ;
  assign n17211 = ~n17199 & n17210 ;
  assign n17212 = ~n17205 & ~n17207 ;
  assign n17213 = n17204 & n17212 ;
  assign n17214 = ~\a[41]  & ~n17213 ;
  assign n17215 = ~\a[41]  & ~n1694 ;
  assign n17216 = ~n17198 & n17215 ;
  assign n17217 = ~n17214 & ~n17216 ;
  assign n17218 = ~n17211 & n17217 ;
  assign n17219 = n16556 & n16682 ;
  assign n17220 = n16681 & ~n17219 ;
  assign n17221 = ~n725 & n11572 ;
  assign n17222 = ~n684 & n11572 ;
  assign n17223 = ~n721 & n17222 ;
  assign n17224 = ~n17221 & ~n17223 ;
  assign n17225 = ~n728 & ~n17224 ;
  assign n17226 = \b[9]  & n12159 ;
  assign n17227 = n12156 & n17226 ;
  assign n17228 = ~\a[45]  & \b[10]  ;
  assign n17229 = n11564 & n17228 ;
  assign n17230 = ~n17227 & ~n17229 ;
  assign n17231 = \b[11]  & n11570 ;
  assign n17232 = \a[45]  & \b[10]  ;
  assign n17233 = n11561 & n17232 ;
  assign n17234 = \a[47]  & ~n17233 ;
  assign n17235 = ~n17231 & n17234 ;
  assign n17236 = n17230 & n17235 ;
  assign n17237 = ~n17225 & n17236 ;
  assign n17238 = ~n17231 & ~n17233 ;
  assign n17239 = n17230 & n17238 ;
  assign n17240 = ~\a[47]  & ~n17239 ;
  assign n17241 = ~\a[47]  & ~n728 ;
  assign n17242 = ~n17224 & n17241 ;
  assign n17243 = ~n17240 & ~n17242 ;
  assign n17244 = ~n17237 & n17243 ;
  assign n17245 = ~n16047 & ~n16670 ;
  assign n17246 = ~n16581 & n17245 ;
  assign n17247 = ~n16669 & ~n17246 ;
  assign n17248 = ~n505 & ~n12606 ;
  assign n17249 = ~n13122 & n17248 ;
  assign n17250 = n502 & n17249 ;
  assign n17251 = n505 & ~n12606 ;
  assign n17252 = ~n13122 & n17251 ;
  assign n17253 = ~n502 & n17252 ;
  assign n17254 = ~n17250 & ~n17253 ;
  assign n17255 = \b[6]  & n13794 ;
  assign n17256 = n13792 & n17255 ;
  assign n17257 = \b[8]  & n13123 ;
  assign n17258 = \a[48]  & \b[7]  ;
  assign n17259 = n13786 & n17258 ;
  assign n17260 = ~\a[48]  & \b[7]  ;
  assign n17261 = n13117 & n17260 ;
  assign n17262 = ~n17259 & ~n17261 ;
  assign n17263 = ~n17257 & n17262 ;
  assign n17264 = ~n17256 & n17263 ;
  assign n17265 = n17254 & n17264 ;
  assign n17266 = ~\a[50]  & ~n17265 ;
  assign n17267 = \a[50]  & n17264 ;
  assign n17268 = n17254 & n17267 ;
  assign n17269 = ~n17266 & ~n17268 ;
  assign n17270 = ~n16664 & ~n16666 ;
  assign n17271 = ~n270 & n14793 ;
  assign n17272 = ~n218 & n14793 ;
  assign n17273 = ~n220 & n17272 ;
  assign n17274 = ~n17271 & ~n17273 ;
  assign n17275 = ~n273 & ~n17274 ;
  assign n17276 = \b[3]  & n15517 ;
  assign n17277 = n15514 & n17276 ;
  assign n17278 = \b[5]  & n14791 ;
  assign n17279 = \a[50]  & \b[4]  ;
  assign n17280 = n15515 & n17279 ;
  assign n17281 = ~\a[51]  & \b[4]  ;
  assign n17282 = n14785 & n17281 ;
  assign n17283 = ~n17280 & ~n17282 ;
  assign n17284 = ~n17278 & n17283 ;
  assign n17285 = ~n17277 & n17284 ;
  assign n17286 = ~\a[53]  & n17285 ;
  assign n17287 = ~n17275 & n17286 ;
  assign n17288 = \a[53]  & ~n17285 ;
  assign n17289 = \a[53]  & ~n273 ;
  assign n17290 = ~n17274 & n17289 ;
  assign n17291 = ~n17288 & ~n17290 ;
  assign n17292 = ~n17287 & n17291 ;
  assign n17293 = \a[56]  & ~n16017 ;
  assign n17294 = n16649 & n17293 ;
  assign n17295 = n16657 & n17294 ;
  assign n17296 = \a[56]  & ~n17295 ;
  assign n17297 = \b[2]  & n16653 ;
  assign n17298 = ~\a[54]  & \b[1]  ;
  assign n17299 = n16647 & n17298 ;
  assign n17300 = \a[54]  & \b[1]  ;
  assign n17301 = n16644 & n17300 ;
  assign n17302 = ~n17299 & ~n17301 ;
  assign n17303 = ~n17297 & n17302 ;
  assign n17304 = n157 & n16655 ;
  assign n17305 = n16016 & ~n16652 ;
  assign n17306 = \a[54]  & ~\a[55]  ;
  assign n17307 = ~\a[54]  & \a[55]  ;
  assign n17308 = ~n17306 & ~n17307 ;
  assign n17309 = \b[0]  & n17308 ;
  assign n17310 = n17305 & n17309 ;
  assign n17311 = ~n17304 & ~n17310 ;
  assign n17312 = n17303 & n17311 ;
  assign n17313 = ~n17296 & ~n17312 ;
  assign n17314 = n17296 & n17312 ;
  assign n17315 = ~n17313 & ~n17314 ;
  assign n17316 = n17292 & ~n17315 ;
  assign n17317 = ~n17292 & n17315 ;
  assign n17318 = ~n17316 & ~n17317 ;
  assign n17319 = ~n17270 & n17318 ;
  assign n17320 = ~n16664 & ~n17318 ;
  assign n17321 = ~n16666 & n17320 ;
  assign n17322 = ~n17319 & ~n17321 ;
  assign n17323 = n17269 & ~n17322 ;
  assign n17324 = ~n17269 & ~n17321 ;
  assign n17325 = ~n17319 & n17324 ;
  assign n17326 = ~n17323 & ~n17325 ;
  assign n17327 = n17247 & n17326 ;
  assign n17328 = ~n17247 & ~n17326 ;
  assign n17329 = ~n17327 & ~n17328 ;
  assign n17330 = n17244 & ~n17329 ;
  assign n17331 = ~n17244 & n17329 ;
  assign n17332 = ~n17330 & ~n17331 ;
  assign n17333 = n1087 & n10082 ;
  assign n17334 = ~n1084 & n17333 ;
  assign n17335 = n1552 & n10082 ;
  assign n17336 = ~n1083 & n17335 ;
  assign n17337 = \b[12]  & n10681 ;
  assign n17338 = n10678 & n17337 ;
  assign n17339 = ~\a[42]  & \b[13]  ;
  assign n17340 = n10074 & n17339 ;
  assign n17341 = ~n17338 & ~n17340 ;
  assign n17342 = \b[14]  & n10080 ;
  assign n17343 = \a[42]  & \b[13]  ;
  assign n17344 = n10071 & n17343 ;
  assign n17345 = \a[44]  & ~n17344 ;
  assign n17346 = ~n17342 & n17345 ;
  assign n17347 = n17341 & n17346 ;
  assign n17348 = ~n17336 & n17347 ;
  assign n17349 = ~n17334 & n17348 ;
  assign n17350 = ~n17342 & ~n17344 ;
  assign n17351 = n17341 & n17350 ;
  assign n17352 = ~n17336 & n17351 ;
  assign n17353 = ~n17334 & n17352 ;
  assign n17354 = ~\a[44]  & ~n17353 ;
  assign n17355 = ~n17349 & ~n17354 ;
  assign n17356 = ~n17332 & ~n17355 ;
  assign n17357 = ~n17220 & n17356 ;
  assign n17358 = n17332 & ~n17355 ;
  assign n17359 = n17220 & n17358 ;
  assign n17360 = ~n17357 & ~n17359 ;
  assign n17361 = ~n17332 & n17355 ;
  assign n17362 = n17220 & n17361 ;
  assign n17363 = n17332 & n17355 ;
  assign n17364 = ~n17220 & n17363 ;
  assign n17365 = ~n17362 & ~n17364 ;
  assign n17366 = n17360 & n17365 ;
  assign n17367 = ~n17218 & ~n17366 ;
  assign n17368 = n17194 & n17367 ;
  assign n17369 = ~n17218 & n17366 ;
  assign n17370 = ~n17194 & n17369 ;
  assign n17371 = ~n17368 & ~n17370 ;
  assign n17372 = n17218 & ~n17366 ;
  assign n17373 = ~n17194 & n17372 ;
  assign n17374 = n17218 & n17366 ;
  assign n17375 = n17194 & n17374 ;
  assign n17376 = ~n17373 & ~n17375 ;
  assign n17377 = n17371 & n17376 ;
  assign n17378 = ~n17191 & n17377 ;
  assign n17379 = n2293 & n7534 ;
  assign n17380 = ~n2290 & n17379 ;
  assign n17381 = n5705 & n7534 ;
  assign n17382 = ~n2289 & n17381 ;
  assign n17383 = \b[18]  & n7973 ;
  assign n17384 = n7970 & n17383 ;
  assign n17385 = \b[20]  & n7532 ;
  assign n17386 = \a[36]  & \b[19]  ;
  assign n17387 = n7523 & n17386 ;
  assign n17388 = ~\a[36]  & \b[19]  ;
  assign n17389 = n7526 & n17388 ;
  assign n17390 = ~n17387 & ~n17389 ;
  assign n17391 = ~n17385 & n17390 ;
  assign n17392 = ~n17384 & n17391 ;
  assign n17393 = ~n17382 & n17392 ;
  assign n17394 = ~n17380 & n17393 ;
  assign n17395 = ~\a[38]  & ~n17394 ;
  assign n17396 = \a[38]  & n17392 ;
  assign n17397 = ~n17382 & n17396 ;
  assign n17398 = ~n17380 & n17397 ;
  assign n17399 = ~n17395 & ~n17398 ;
  assign n17400 = ~n16721 & ~n17377 ;
  assign n17401 = ~n17190 & n17400 ;
  assign n17402 = ~n17399 & ~n17401 ;
  assign n17403 = ~n17378 & n17402 ;
  assign n17404 = ~n17377 & n17399 ;
  assign n17405 = n17191 & n17404 ;
  assign n17406 = n17377 & n17399 ;
  assign n17407 = ~n17191 & n17406 ;
  assign n17408 = ~n17405 & ~n17407 ;
  assign n17409 = ~n17403 & n17408 ;
  assign n17410 = n17189 & n17409 ;
  assign n17411 = ~n17189 & ~n17409 ;
  assign n17412 = ~n17410 & ~n17411 ;
  assign n17413 = ~n17186 & n17412 ;
  assign n17414 = n17186 & ~n17412 ;
  assign n17415 = ~n17413 & ~n17414 ;
  assign n17416 = n3604 & n5211 ;
  assign n17417 = ~n3601 & n17416 ;
  assign n17418 = ~n3604 & n5211 ;
  assign n17419 = ~n3562 & n17418 ;
  assign n17420 = ~n3600 & n17419 ;
  assign n17421 = \b[24]  & n5595 ;
  assign n17422 = n5592 & n17421 ;
  assign n17423 = ~\a[30]  & \b[25]  ;
  assign n17424 = n5203 & n17423 ;
  assign n17425 = ~n17422 & ~n17424 ;
  assign n17426 = \b[26]  & n5209 ;
  assign n17427 = \a[30]  & \b[25]  ;
  assign n17428 = n5200 & n17427 ;
  assign n17429 = \a[32]  & ~n17428 ;
  assign n17430 = ~n17426 & n17429 ;
  assign n17431 = n17425 & n17430 ;
  assign n17432 = ~n17420 & n17431 ;
  assign n17433 = ~n17417 & n17432 ;
  assign n17434 = ~n17426 & ~n17428 ;
  assign n17435 = n17425 & n17434 ;
  assign n17436 = ~n17420 & n17435 ;
  assign n17437 = ~n17417 & n17436 ;
  assign n17438 = ~\a[32]  & ~n17437 ;
  assign n17439 = ~n17433 & ~n17438 ;
  assign n17440 = ~n17415 & ~n17439 ;
  assign n17441 = ~n17169 & n17440 ;
  assign n17442 = n17415 & ~n17439 ;
  assign n17443 = n17169 & n17442 ;
  assign n17444 = ~n17441 & ~n17443 ;
  assign n17445 = ~n17415 & n17439 ;
  assign n17446 = n17169 & n17445 ;
  assign n17447 = n17415 & n17439 ;
  assign n17448 = ~n17169 & n17447 ;
  assign n17449 = ~n17446 & ~n17448 ;
  assign n17450 = n17444 & n17449 ;
  assign n17451 = n17167 & ~n17450 ;
  assign n17452 = ~n17148 & n17451 ;
  assign n17453 = n17167 & n17450 ;
  assign n17454 = n17148 & n17453 ;
  assign n17455 = ~n17452 & ~n17454 ;
  assign n17456 = ~n17167 & ~n17450 ;
  assign n17457 = n17148 & n17456 ;
  assign n17458 = ~n17167 & n17450 ;
  assign n17459 = ~n17148 & n17458 ;
  assign n17460 = ~n17457 & ~n17459 ;
  assign n17461 = n17455 & n17460 ;
  assign n17462 = n17145 & ~n17461 ;
  assign n17463 = n17121 & n17462 ;
  assign n17464 = n17145 & n17461 ;
  assign n17465 = ~n17121 & n17464 ;
  assign n17466 = ~n17463 & ~n17465 ;
  assign n17467 = ~n17121 & n17461 ;
  assign n17468 = ~n16828 & ~n17461 ;
  assign n17469 = ~n17120 & n17468 ;
  assign n17470 = ~n17145 & ~n17469 ;
  assign n17471 = ~n17467 & n17470 ;
  assign n17472 = n17466 & ~n17471 ;
  assign n17473 = ~n17119 & n17472 ;
  assign n17474 = n17119 & ~n17472 ;
  assign n17475 = ~n17473 & ~n17474 ;
  assign n17476 = n2622 & ~n6610 ;
  assign n17477 = ~n6608 & n17476 ;
  assign n17478 = \b[35]  & n2620 ;
  assign n17479 = \a[21]  & \b[34]  ;
  assign n17480 = n2611 & n17479 ;
  assign n17481 = ~n17478 & ~n17480 ;
  assign n17482 = \b[33]  & n2912 ;
  assign n17483 = n2909 & n17482 ;
  assign n17484 = ~\a[21]  & \b[34]  ;
  assign n17485 = n2614 & n17484 ;
  assign n17486 = ~n17483 & ~n17485 ;
  assign n17487 = n17481 & n17486 ;
  assign n17488 = ~n17477 & n17487 ;
  assign n17489 = ~\a[23]  & ~n17488 ;
  assign n17490 = \a[23]  & n17487 ;
  assign n17491 = ~n17477 & n17490 ;
  assign n17492 = ~n17489 & ~n17491 ;
  assign n17493 = n17475 & ~n17492 ;
  assign n17494 = ~n17475 & n17492 ;
  assign n17495 = ~n17493 & ~n17494 ;
  assign n17496 = ~n17114 & n17495 ;
  assign n17497 = ~n16891 & ~n17495 ;
  assign n17498 = ~n17113 & n17497 ;
  assign n17499 = n1965 & n8175 ;
  assign n17500 = ~n8172 & n17499 ;
  assign n17501 = n1965 & ~n8175 ;
  assign n17502 = ~n7756 & n17501 ;
  assign n17503 = ~n8171 & n17502 ;
  assign n17504 = \b[36]  & n2218 ;
  assign n17505 = n2216 & n17504 ;
  assign n17506 = ~\a[18]  & \b[37]  ;
  assign n17507 = n1957 & n17506 ;
  assign n17508 = ~n17505 & ~n17507 ;
  assign n17509 = \b[38]  & n1963 ;
  assign n17510 = \a[18]  & \b[37]  ;
  assign n17511 = n2210 & n17510 ;
  assign n17512 = \a[20]  & ~n17511 ;
  assign n17513 = ~n17509 & n17512 ;
  assign n17514 = n17508 & n17513 ;
  assign n17515 = ~n17503 & n17514 ;
  assign n17516 = ~n17500 & n17515 ;
  assign n17517 = ~n17509 & ~n17511 ;
  assign n17518 = n17508 & n17517 ;
  assign n17519 = ~n17503 & n17518 ;
  assign n17520 = ~n17500 & n17519 ;
  assign n17521 = ~\a[20]  & ~n17520 ;
  assign n17522 = ~n17516 & ~n17521 ;
  assign n17523 = ~n17498 & ~n17522 ;
  assign n17524 = ~n17496 & n17523 ;
  assign n17525 = ~n17495 & n17522 ;
  assign n17526 = n17114 & n17525 ;
  assign n17527 = n17495 & n17522 ;
  assign n17528 = ~n17114 & n17527 ;
  assign n17529 = ~n17526 & ~n17528 ;
  assign n17530 = ~n17524 & n17529 ;
  assign n17531 = ~n17112 & ~n17530 ;
  assign n17532 = n17112 & n17530 ;
  assign n17533 = ~n17531 & ~n17532 ;
  assign n17534 = n1467 & ~n9482 ;
  assign n17535 = ~n9480 & n17534 ;
  assign n17536 = \b[41]  & n1465 ;
  assign n17537 = \a[15]  & \b[40]  ;
  assign n17538 = n1456 & n17537 ;
  assign n17539 = ~n17536 & ~n17538 ;
  assign n17540 = \b[39]  & n1652 ;
  assign n17541 = n1649 & n17540 ;
  assign n17542 = ~\a[15]  & \b[40]  ;
  assign n17543 = n1459 & n17542 ;
  assign n17544 = ~n17541 & ~n17543 ;
  assign n17545 = n17539 & n17544 ;
  assign n17546 = ~n17535 & n17545 ;
  assign n17547 = ~\a[17]  & ~n17546 ;
  assign n17548 = \a[17]  & n17545 ;
  assign n17549 = ~n17535 & n17548 ;
  assign n17550 = ~n17547 & ~n17549 ;
  assign n17551 = n17533 & ~n17550 ;
  assign n17552 = ~n17533 & n17550 ;
  assign n17553 = ~n17551 & ~n17552 ;
  assign n17554 = n999 & ~n10892 ;
  assign n17555 = ~n10890 & n17554 ;
  assign n17556 = \b[42]  & n1182 ;
  assign n17557 = n1179 & n17556 ;
  assign n17558 = \b[44]  & n997 ;
  assign n17559 = \a[11]  & \b[43]  ;
  assign n17560 = n1180 & n17559 ;
  assign n17561 = ~\a[12]  & \b[43]  ;
  assign n17562 = n7674 & n17561 ;
  assign n17563 = ~n17560 & ~n17562 ;
  assign n17564 = ~n17558 & n17563 ;
  assign n17565 = ~n17557 & n17564 ;
  assign n17566 = ~n17555 & n17565 ;
  assign n17567 = ~\a[14]  & ~n17566 ;
  assign n17568 = \a[14]  & n17565 ;
  assign n17569 = ~n17555 & n17568 ;
  assign n17570 = ~n17567 & ~n17569 ;
  assign n17571 = ~n17553 & ~n17570 ;
  assign n17572 = ~n17109 & n17571 ;
  assign n17573 = n17553 & ~n17570 ;
  assign n17574 = n17109 & n17573 ;
  assign n17575 = ~n17572 & ~n17574 ;
  assign n17576 = ~n17553 & n17570 ;
  assign n17577 = n17109 & n17576 ;
  assign n17578 = n17553 & n17570 ;
  assign n17579 = ~n17109 & n17578 ;
  assign n17580 = ~n17577 & ~n17579 ;
  assign n17581 = n17575 & n17580 ;
  assign n17582 = ~n17107 & ~n17581 ;
  assign n17583 = n17090 & n17582 ;
  assign n17584 = ~n17107 & n17581 ;
  assign n17585 = ~n17090 & n17584 ;
  assign n17586 = ~n17583 & ~n17585 ;
  assign n17587 = n17107 & ~n17581 ;
  assign n17588 = ~n17090 & n17587 ;
  assign n17589 = n17107 & n17581 ;
  assign n17590 = n17090 & n17589 ;
  assign n17591 = ~n17588 & ~n17590 ;
  assign n17592 = n17586 & n17591 ;
  assign n17593 = ~n17087 & n17592 ;
  assign n17594 = ~n359 & ~n13519 ;
  assign n17595 = ~n14052 & n17594 ;
  assign n17596 = ~n14048 & n17595 ;
  assign n17597 = ~n427 & n17596 ;
  assign n17598 = n430 & n14052 ;
  assign n17599 = ~n14049 & n17598 ;
  assign n17600 = ~n17597 & ~n17599 ;
  assign n17601 = \b[48]  & n486 ;
  assign n17602 = n483 & n17601 ;
  assign n17603 = ~\a[6]  & \b[49]  ;
  assign n17604 = n422 & n17603 ;
  assign n17605 = ~n17602 & ~n17604 ;
  assign n17606 = \b[50]  & n428 ;
  assign n17607 = \a[6]  & \b[49]  ;
  assign n17608 = n419 & n17607 ;
  assign n17609 = \a[8]  & ~n17608 ;
  assign n17610 = ~n17606 & n17609 ;
  assign n17611 = n17605 & n17610 ;
  assign n17612 = n17600 & n17611 ;
  assign n17613 = ~n17606 & ~n17608 ;
  assign n17614 = n17605 & n17613 ;
  assign n17615 = n17600 & n17614 ;
  assign n17616 = ~\a[8]  & ~n17615 ;
  assign n17617 = ~n17612 & ~n17616 ;
  assign n17618 = ~n16998 & ~n17592 ;
  assign n17619 = ~n17086 & n17618 ;
  assign n17620 = ~n17617 & ~n17619 ;
  assign n17621 = ~n17593 & n17620 ;
  assign n17622 = ~n17592 & n17617 ;
  assign n17623 = n17087 & n17622 ;
  assign n17624 = n17592 & n17617 ;
  assign n17625 = ~n17087 & n17624 ;
  assign n17626 = ~n17623 & ~n17625 ;
  assign n17627 = ~n17621 & n17626 ;
  assign n17628 = n17085 & ~n17627 ;
  assign n17629 = ~n17068 & n17628 ;
  assign n17630 = n17085 & n17627 ;
  assign n17631 = n17068 & n17630 ;
  assign n17632 = ~n17629 & ~n17631 ;
  assign n17633 = ~n17085 & ~n17627 ;
  assign n17634 = n17068 & n17633 ;
  assign n17635 = ~n17085 & n17627 ;
  assign n17636 = ~n17068 & n17635 ;
  assign n17637 = ~n17634 & ~n17636 ;
  assign n17638 = n17632 & n17637 ;
  assign n17639 = ~n17065 & n17638 ;
  assign n17640 = ~n17039 & ~n17638 ;
  assign n17641 = ~n17064 & n17640 ;
  assign n17642 = ~n16397 & ~n16442 ;
  assign n17643 = ~n16406 & n17642 ;
  assign n17644 = ~n16441 & ~n17643 ;
  assign n17645 = ~\b[55]  & ~\b[56]  ;
  assign n17646 = \b[55]  & \b[56]  ;
  assign n17647 = ~n17645 & ~n17646 ;
  assign n17648 = n134 & n17647 ;
  assign n17649 = ~n17644 & n17648 ;
  assign n17650 = n134 & ~n17647 ;
  assign n17651 = ~n16441 & n17650 ;
  assign n17652 = ~n17643 & n17651 ;
  assign n17653 = \a[0]  & \b[56]  ;
  assign n17654 = n133 & n17653 ;
  assign n17655 = \b[55]  & n141 ;
  assign n17656 = ~\a[1]  & \b[54]  ;
  assign n17657 = n10416 & n17656 ;
  assign n17658 = ~n17655 & ~n17657 ;
  assign n17659 = ~n17654 & n17658 ;
  assign n17660 = \a[2]  & n17659 ;
  assign n17661 = ~n17652 & n17660 ;
  assign n17662 = ~n17649 & n17661 ;
  assign n17663 = ~n17652 & n17659 ;
  assign n17664 = ~n17649 & n17663 ;
  assign n17665 = ~\a[2]  & ~n17664 ;
  assign n17666 = ~n17662 & ~n17665 ;
  assign n17667 = ~n17641 & ~n17666 ;
  assign n17668 = ~n17639 & n17667 ;
  assign n17669 = ~n17638 & n17666 ;
  assign n17670 = n17065 & n17669 ;
  assign n17671 = n17638 & n17666 ;
  assign n17672 = ~n17065 & n17671 ;
  assign n17673 = ~n17670 & ~n17672 ;
  assign n17674 = ~n17668 & n17673 ;
  assign n17675 = n17063 & n17674 ;
  assign n17676 = ~n17063 & ~n17674 ;
  assign n17677 = ~n17675 & ~n17676 ;
  assign n17678 = ~n17668 & ~n17675 ;
  assign n17679 = ~n17039 & n17637 ;
  assign n17680 = ~n17064 & n17679 ;
  assign n17681 = n17632 & ~n17680 ;
  assign n17682 = ~n16441 & n17647 ;
  assign n17683 = ~n17643 & n17682 ;
  assign n17684 = ~n17646 & ~n17683 ;
  assign n17685 = ~\b[56]  & ~\b[57]  ;
  assign n17686 = \b[56]  & \b[57]  ;
  assign n17687 = ~n17685 & ~n17686 ;
  assign n17688 = ~n17684 & n17687 ;
  assign n17689 = ~n17646 & ~n17687 ;
  assign n17690 = ~n17683 & n17689 ;
  assign n17691 = n134 & ~n17690 ;
  assign n17692 = ~n17688 & n17691 ;
  assign n17693 = \a[0]  & \b[57]  ;
  assign n17694 = n133 & n17693 ;
  assign n17695 = \b[56]  & n141 ;
  assign n17696 = ~\a[1]  & \b[55]  ;
  assign n17697 = n10416 & n17696 ;
  assign n17698 = ~n17695 & ~n17697 ;
  assign n17699 = ~n17694 & n17698 ;
  assign n17700 = ~n17692 & n17699 ;
  assign n17701 = ~\a[2]  & ~n17700 ;
  assign n17702 = \a[2]  & n17699 ;
  assign n17703 = ~n17692 & n17702 ;
  assign n17704 = ~n17701 & ~n17703 ;
  assign n17705 = n17068 & n17627 ;
  assign n17706 = ~n17621 & ~n17705 ;
  assign n17707 = ~n16998 & n17586 ;
  assign n17708 = ~n17086 & n17707 ;
  assign n17709 = n17591 & ~n17708 ;
  assign n17710 = n430 & ~n14098 ;
  assign n17711 = ~n14096 & n17710 ;
  assign n17712 = \b[51]  & n428 ;
  assign n17713 = \a[6]  & \b[50]  ;
  assign n17714 = n419 & n17713 ;
  assign n17715 = ~n17712 & ~n17714 ;
  assign n17716 = \b[49]  & n486 ;
  assign n17717 = n483 & n17716 ;
  assign n17718 = ~\a[6]  & \b[50]  ;
  assign n17719 = n422 & n17718 ;
  assign n17720 = ~n17717 & ~n17719 ;
  assign n17721 = n17715 & n17720 ;
  assign n17722 = ~n17711 & n17721 ;
  assign n17723 = ~\a[8]  & ~n17722 ;
  assign n17724 = \a[8]  & n17721 ;
  assign n17725 = ~n17711 & n17724 ;
  assign n17726 = ~n17723 & ~n17725 ;
  assign n17727 = n17090 & n17581 ;
  assign n17728 = n17575 & ~n17727 ;
  assign n17729 = n16954 & ~n17551 ;
  assign n17730 = ~n17108 & n17729 ;
  assign n17731 = ~n17552 & ~n17730 ;
  assign n17732 = n999 & ~n11397 ;
  assign n17733 = ~n11395 & n17732 ;
  assign n17734 = \b[43]  & n1182 ;
  assign n17735 = n1179 & n17734 ;
  assign n17736 = \b[45]  & n997 ;
  assign n17737 = \a[11]  & \b[44]  ;
  assign n17738 = n1180 & n17737 ;
  assign n17739 = ~\a[12]  & \b[44]  ;
  assign n17740 = n7674 & n17739 ;
  assign n17741 = ~n17738 & ~n17740 ;
  assign n17742 = ~n17736 & n17741 ;
  assign n17743 = ~n17735 & n17742 ;
  assign n17744 = ~n17733 & n17743 ;
  assign n17745 = ~\a[14]  & ~n17744 ;
  assign n17746 = \a[14]  & n17743 ;
  assign n17747 = ~n17733 & n17746 ;
  assign n17748 = ~n17745 & ~n17747 ;
  assign n17749 = ~n17524 & ~n17532 ;
  assign n17750 = ~n16891 & ~n17493 ;
  assign n17751 = ~n17113 & n17750 ;
  assign n17752 = ~n17494 & ~n17751 ;
  assign n17753 = ~n17471 & ~n17473 ;
  assign n17754 = n2622 & n7337 ;
  assign n17755 = ~n7334 & n17754 ;
  assign n17756 = n2622 & ~n7337 ;
  assign n17757 = ~n6605 & n17756 ;
  assign n17758 = ~n7333 & n17757 ;
  assign n17759 = \b[34]  & n2912 ;
  assign n17760 = n2909 & n17759 ;
  assign n17761 = ~\a[21]  & \b[35]  ;
  assign n17762 = n2614 & n17761 ;
  assign n17763 = ~n17760 & ~n17762 ;
  assign n17764 = \b[36]  & n2620 ;
  assign n17765 = \a[21]  & \b[35]  ;
  assign n17766 = n2611 & n17765 ;
  assign n17767 = \a[23]  & ~n17766 ;
  assign n17768 = ~n17764 & n17767 ;
  assign n17769 = n17763 & n17768 ;
  assign n17770 = ~n17758 & n17769 ;
  assign n17771 = ~n17755 & n17770 ;
  assign n17772 = ~n17764 & ~n17766 ;
  assign n17773 = n17763 & n17772 ;
  assign n17774 = ~n17758 & n17773 ;
  assign n17775 = ~n17755 & n17774 ;
  assign n17776 = ~\a[23]  & ~n17775 ;
  assign n17777 = ~n17771 & ~n17776 ;
  assign n17778 = ~n16828 & n17460 ;
  assign n17779 = ~n17120 & n17778 ;
  assign n17780 = n17455 & ~n17779 ;
  assign n17781 = n17148 & n17450 ;
  assign n17782 = n17444 & ~n17781 ;
  assign n17783 = n16765 & ~n17413 ;
  assign n17784 = ~n17168 & n17783 ;
  assign n17785 = ~n17414 & ~n17784 ;
  assign n17786 = ~n17403 & ~n17410 ;
  assign n17787 = ~n16721 & n17371 ;
  assign n17788 = ~n17190 & n17787 ;
  assign n17789 = n17376 & ~n17788 ;
  assign n17790 = ~n2520 & n7534 ;
  assign n17791 = ~n2292 & n7534 ;
  assign n17792 = ~n2516 & n17791 ;
  assign n17793 = ~n17790 & ~n17792 ;
  assign n17794 = ~n2523 & ~n17793 ;
  assign n17795 = \b[19]  & n7973 ;
  assign n17796 = n7970 & n17795 ;
  assign n17797 = ~\a[35]  & \b[20]  ;
  assign n17798 = n7972 & n17797 ;
  assign n17799 = ~n17796 & ~n17798 ;
  assign n17800 = \b[21]  & n7532 ;
  assign n17801 = \a[35]  & ~\a[37]  ;
  assign n17802 = \a[36]  & \b[20]  ;
  assign n17803 = n17801 & n17802 ;
  assign n17804 = \a[38]  & ~n17803 ;
  assign n17805 = ~n17800 & n17804 ;
  assign n17806 = n17799 & n17805 ;
  assign n17807 = ~n17794 & n17806 ;
  assign n17808 = ~n17800 & ~n17803 ;
  assign n17809 = n17799 & n17808 ;
  assign n17810 = ~\a[38]  & ~n17809 ;
  assign n17811 = ~\a[38]  & ~n2523 ;
  assign n17812 = ~n17793 & n17811 ;
  assign n17813 = ~n17810 & ~n17812 ;
  assign n17814 = ~n17807 & n17813 ;
  assign n17815 = n17194 & n17366 ;
  assign n17816 = n17360 & ~n17815 ;
  assign n17817 = n16681 & ~n17331 ;
  assign n17818 = ~n17219 & n17817 ;
  assign n17819 = ~n17330 & ~n17818 ;
  assign n17820 = ~n1230 & n10082 ;
  assign n17821 = ~n1086 & n10082 ;
  assign n17822 = ~n1226 & n17821 ;
  assign n17823 = ~n17820 & ~n17822 ;
  assign n17824 = ~n1233 & ~n17823 ;
  assign n17825 = \b[13]  & n10681 ;
  assign n17826 = n10678 & n17825 ;
  assign n17827 = ~\a[42]  & \b[14]  ;
  assign n17828 = n10074 & n17827 ;
  assign n17829 = ~n17826 & ~n17828 ;
  assign n17830 = \b[15]  & n10080 ;
  assign n17831 = \a[42]  & \b[14]  ;
  assign n17832 = n10071 & n17831 ;
  assign n17833 = \a[44]  & ~n17832 ;
  assign n17834 = ~n17830 & n17833 ;
  assign n17835 = n17829 & n17834 ;
  assign n17836 = ~n17824 & n17835 ;
  assign n17837 = ~n17830 & ~n17832 ;
  assign n17838 = n17829 & n17837 ;
  assign n17839 = ~\a[44]  & ~n17838 ;
  assign n17840 = ~\a[44]  & ~n1233 ;
  assign n17841 = ~n17823 & n17840 ;
  assign n17842 = ~n17839 & ~n17841 ;
  assign n17843 = ~n17836 & n17842 ;
  assign n17844 = ~n17325 & ~n17327 ;
  assign n17845 = ~n909 & ~n10988 ;
  assign n17846 = ~n11569 & n17845 ;
  assign n17847 = n906 & n17846 ;
  assign n17848 = n909 & ~n10988 ;
  assign n17849 = ~n11569 & n17848 ;
  assign n17850 = ~n906 & n17849 ;
  assign n17851 = ~n17847 & ~n17850 ;
  assign n17852 = \b[10]  & n12159 ;
  assign n17853 = n12156 & n17852 ;
  assign n17854 = ~\a[45]  & \b[11]  ;
  assign n17855 = n11564 & n17854 ;
  assign n17856 = ~n17853 & ~n17855 ;
  assign n17857 = \b[12]  & n11570 ;
  assign n17858 = \a[45]  & \b[11]  ;
  assign n17859 = n11561 & n17858 ;
  assign n17860 = \a[47]  & ~n17859 ;
  assign n17861 = ~n17857 & n17860 ;
  assign n17862 = n17856 & n17861 ;
  assign n17863 = n17851 & n17862 ;
  assign n17864 = ~n17857 & ~n17859 ;
  assign n17865 = n17856 & n17864 ;
  assign n17866 = n17851 & n17865 ;
  assign n17867 = ~\a[47]  & ~n17866 ;
  assign n17868 = ~n17863 & ~n17867 ;
  assign n17869 = ~n16664 & ~n17316 ;
  assign n17870 = ~n16666 & n17869 ;
  assign n17871 = ~n17317 & ~n17870 ;
  assign n17872 = ~n586 & n13125 ;
  assign n17873 = ~n504 & n13125 ;
  assign n17874 = ~n508 & n17873 ;
  assign n17875 = ~n17872 & ~n17874 ;
  assign n17876 = ~n589 & ~n17875 ;
  assign n17877 = \b[7]  & n13794 ;
  assign n17878 = n13792 & n17877 ;
  assign n17879 = \b[9]  & n13123 ;
  assign n17880 = \a[48]  & \b[8]  ;
  assign n17881 = n13786 & n17880 ;
  assign n17882 = ~\a[48]  & \b[8]  ;
  assign n17883 = n13117 & n17882 ;
  assign n17884 = ~n17881 & ~n17883 ;
  assign n17885 = ~n17879 & n17884 ;
  assign n17886 = ~n17878 & n17885 ;
  assign n17887 = ~\a[50]  & n17886 ;
  assign n17888 = ~n17876 & n17887 ;
  assign n17889 = \a[50]  & ~n17886 ;
  assign n17890 = \a[50]  & ~n589 ;
  assign n17891 = ~n17875 & n17890 ;
  assign n17892 = ~n17889 & ~n17891 ;
  assign n17893 = ~n17888 & n17892 ;
  assign n17894 = n177 & n16655 ;
  assign n17895 = \b[3]  & n16653 ;
  assign n17896 = \a[53]  & \b[2]  ;
  assign n17897 = n17306 & n17896 ;
  assign n17898 = ~\a[54]  & \b[2]  ;
  assign n17899 = n16647 & n17898 ;
  assign n17900 = ~n17897 & ~n17899 ;
  assign n17901 = ~n17895 & n17900 ;
  assign n17902 = ~n17894 & n17901 ;
  assign n17903 = \b[1]  & n17308 ;
  assign n17904 = n17305 & n17903 ;
  assign n17905 = ~\a[56]  & ~n17904 ;
  assign n17906 = n17902 & n17905 ;
  assign n17907 = n17902 & ~n17904 ;
  assign n17908 = \a[56]  & ~n17907 ;
  assign n17909 = ~n17906 & ~n17908 ;
  assign n17910 = \a[56]  & ~\a[57]  ;
  assign n17911 = ~\a[56]  & \a[57]  ;
  assign n17912 = ~n17910 & ~n17911 ;
  assign n17913 = \b[0]  & ~n17912 ;
  assign n17914 = n17295 & n17312 ;
  assign n17915 = n17913 & n17914 ;
  assign n17916 = ~n17913 & ~n17914 ;
  assign n17917 = ~n17915 & ~n17916 ;
  assign n17918 = n17909 & n17917 ;
  assign n17919 = ~n17909 & ~n17917 ;
  assign n17920 = ~n17918 & ~n17919 ;
  assign n17921 = ~n323 & ~n14276 ;
  assign n17922 = ~n14790 & n17921 ;
  assign n17923 = n320 & n17922 ;
  assign n17924 = n323 & ~n14276 ;
  assign n17925 = ~n14790 & n17924 ;
  assign n17926 = ~n320 & n17925 ;
  assign n17927 = ~n17923 & ~n17926 ;
  assign n17928 = \b[4]  & n15517 ;
  assign n17929 = n15514 & n17928 ;
  assign n17930 = \b[6]  & n14791 ;
  assign n17931 = \a[50]  & \b[5]  ;
  assign n17932 = n15515 & n17931 ;
  assign n17933 = ~\a[51]  & \b[5]  ;
  assign n17934 = n14785 & n17933 ;
  assign n17935 = ~n17932 & ~n17934 ;
  assign n17936 = ~n17930 & n17935 ;
  assign n17937 = ~n17929 & n17936 ;
  assign n17938 = n17927 & n17937 ;
  assign n17939 = ~\a[53]  & ~n17938 ;
  assign n17940 = \a[53]  & n17937 ;
  assign n17941 = n17927 & n17940 ;
  assign n17942 = ~n17939 & ~n17941 ;
  assign n17943 = n17920 & ~n17942 ;
  assign n17944 = ~n17920 & n17942 ;
  assign n17945 = ~n17943 & ~n17944 ;
  assign n17946 = n17893 & ~n17945 ;
  assign n17947 = n17871 & n17946 ;
  assign n17948 = n17893 & n17945 ;
  assign n17949 = ~n17871 & n17948 ;
  assign n17950 = ~n17947 & ~n17949 ;
  assign n17951 = ~n17893 & ~n17945 ;
  assign n17952 = ~n17871 & n17951 ;
  assign n17953 = ~n17893 & n17945 ;
  assign n17954 = n17871 & n17953 ;
  assign n17955 = ~n17952 & ~n17954 ;
  assign n17956 = n17950 & n17955 ;
  assign n17957 = n17868 & ~n17956 ;
  assign n17958 = n17844 & n17957 ;
  assign n17959 = n17868 & n17956 ;
  assign n17960 = ~n17844 & n17959 ;
  assign n17961 = ~n17958 & ~n17960 ;
  assign n17962 = ~n17844 & n17956 ;
  assign n17963 = ~n17325 & ~n17956 ;
  assign n17964 = ~n17327 & n17963 ;
  assign n17965 = ~n17868 & ~n17964 ;
  assign n17966 = ~n17962 & n17965 ;
  assign n17967 = n17961 & ~n17966 ;
  assign n17968 = ~n17843 & ~n17967 ;
  assign n17969 = n17819 & n17968 ;
  assign n17970 = ~n17843 & n17967 ;
  assign n17971 = ~n17819 & n17970 ;
  assign n17972 = ~n17969 & ~n17971 ;
  assign n17973 = n17843 & ~n17967 ;
  assign n17974 = ~n17819 & n17973 ;
  assign n17975 = n17843 & n17967 ;
  assign n17976 = n17819 & n17975 ;
  assign n17977 = ~n17974 & ~n17976 ;
  assign n17978 = n17972 & n17977 ;
  assign n17979 = ~n17816 & n17978 ;
  assign n17980 = n1875 & n8759 ;
  assign n17981 = ~n1872 & n17980 ;
  assign n17982 = n5000 & n8759 ;
  assign n17983 = ~n1871 & n17982 ;
  assign n17984 = \b[16]  & n9301 ;
  assign n17985 = n9298 & n17984 ;
  assign n17986 = ~\a[39]  & \b[17]  ;
  assign n17987 = n8751 & n17986 ;
  assign n17988 = ~n17985 & ~n17987 ;
  assign n17989 = \b[18]  & n8757 ;
  assign n17990 = \a[39]  & \b[17]  ;
  assign n17991 = n8748 & n17990 ;
  assign n17992 = \a[41]  & ~n17991 ;
  assign n17993 = ~n17989 & n17992 ;
  assign n17994 = n17988 & n17993 ;
  assign n17995 = ~n17983 & n17994 ;
  assign n17996 = ~n17981 & n17995 ;
  assign n17997 = ~n17989 & ~n17991 ;
  assign n17998 = n17988 & n17997 ;
  assign n17999 = ~n17983 & n17998 ;
  assign n18000 = ~n17981 & n17999 ;
  assign n18001 = ~\a[41]  & ~n18000 ;
  assign n18002 = ~n17996 & ~n18001 ;
  assign n18003 = n17360 & ~n17978 ;
  assign n18004 = ~n17815 & n18003 ;
  assign n18005 = ~n18002 & ~n18004 ;
  assign n18006 = ~n17979 & n18005 ;
  assign n18007 = ~n17978 & n18002 ;
  assign n18008 = n17816 & n18007 ;
  assign n18009 = n17978 & n18002 ;
  assign n18010 = ~n17816 & n18009 ;
  assign n18011 = ~n18008 & ~n18010 ;
  assign n18012 = ~n18006 & n18011 ;
  assign n18013 = ~n17814 & ~n18012 ;
  assign n18014 = n17789 & n18013 ;
  assign n18015 = ~n17814 & n18012 ;
  assign n18016 = ~n17789 & n18015 ;
  assign n18017 = ~n18014 & ~n18016 ;
  assign n18018 = n17814 & ~n18012 ;
  assign n18019 = ~n17789 & n18018 ;
  assign n18020 = n17814 & n18012 ;
  assign n18021 = n17789 & n18020 ;
  assign n18022 = ~n18019 & ~n18021 ;
  assign n18023 = n18017 & n18022 ;
  assign n18024 = n3283 & n6309 ;
  assign n18025 = ~n3280 & n18024 ;
  assign n18026 = ~n3283 & n6309 ;
  assign n18027 = ~n3017 & n18026 ;
  assign n18028 = ~n3279 & n18027 ;
  assign n18029 = \b[22]  & n6778 ;
  assign n18030 = n6775 & n18029 ;
  assign n18031 = ~\a[33]  & \b[23]  ;
  assign n18032 = n6301 & n18031 ;
  assign n18033 = ~n18030 & ~n18032 ;
  assign n18034 = \b[24]  & n6307 ;
  assign n18035 = \a[33]  & \b[23]  ;
  assign n18036 = n6298 & n18035 ;
  assign n18037 = \a[35]  & ~n18036 ;
  assign n18038 = ~n18034 & n18037 ;
  assign n18039 = n18033 & n18038 ;
  assign n18040 = ~n18028 & n18039 ;
  assign n18041 = ~n18025 & n18040 ;
  assign n18042 = ~n18034 & ~n18036 ;
  assign n18043 = n18033 & n18042 ;
  assign n18044 = ~n18028 & n18043 ;
  assign n18045 = ~n18025 & n18044 ;
  assign n18046 = ~\a[35]  & ~n18045 ;
  assign n18047 = ~n18041 & ~n18046 ;
  assign n18048 = ~n18023 & ~n18047 ;
  assign n18049 = ~n17786 & n18048 ;
  assign n18050 = n18023 & ~n18047 ;
  assign n18051 = n17786 & n18050 ;
  assign n18052 = ~n18049 & ~n18051 ;
  assign n18053 = ~n18023 & n18047 ;
  assign n18054 = n17786 & n18053 ;
  assign n18055 = n18023 & n18047 ;
  assign n18056 = ~n17786 & n18055 ;
  assign n18057 = ~n18054 & ~n18056 ;
  assign n18058 = n18052 & n18057 ;
  assign n18059 = ~n4148 & n5211 ;
  assign n18060 = ~n4146 & n18059 ;
  assign n18061 = \b[25]  & n5595 ;
  assign n18062 = n5592 & n18061 ;
  assign n18063 = ~\a[30]  & \b[26]  ;
  assign n18064 = n5203 & n18063 ;
  assign n18065 = ~n18062 & ~n18064 ;
  assign n18066 = \b[27]  & n5209 ;
  assign n18067 = \a[30]  & \b[26]  ;
  assign n18068 = n5200 & n18067 ;
  assign n18069 = \a[32]  & ~n18068 ;
  assign n18070 = ~n18066 & n18069 ;
  assign n18071 = n18065 & n18070 ;
  assign n18072 = ~n18060 & n18071 ;
  assign n18073 = ~n18066 & ~n18068 ;
  assign n18074 = n18065 & n18073 ;
  assign n18075 = ~n18060 & n18074 ;
  assign n18076 = ~\a[32]  & ~n18075 ;
  assign n18077 = ~n18072 & ~n18076 ;
  assign n18078 = ~n18058 & n18077 ;
  assign n18079 = ~n17785 & n18078 ;
  assign n18080 = n18058 & n18077 ;
  assign n18081 = n17785 & n18080 ;
  assign n18082 = ~n18079 & ~n18081 ;
  assign n18083 = ~n18058 & ~n18077 ;
  assign n18084 = n17785 & n18083 ;
  assign n18085 = n18058 & ~n18077 ;
  assign n18086 = ~n17785 & n18085 ;
  assign n18087 = ~n18084 & ~n18086 ;
  assign n18088 = n18082 & n18087 ;
  assign n18089 = ~n17782 & n18088 ;
  assign n18090 = n4249 & n5105 ;
  assign n18091 = ~n5102 & n18090 ;
  assign n18092 = ~n4497 & ~n5105 ;
  assign n18093 = n4249 & n18092 ;
  assign n18094 = ~n5101 & n18093 ;
  assign n18095 = \b[28]  & n4647 ;
  assign n18096 = n4644 & n18095 ;
  assign n18097 = ~\a[27]  & \b[29]  ;
  assign n18098 = n4241 & n18097 ;
  assign n18099 = ~n18096 & ~n18098 ;
  assign n18100 = \b[30]  & n4247 ;
  assign n18101 = \a[27]  & \b[29]  ;
  assign n18102 = n4238 & n18101 ;
  assign n18103 = \a[29]  & ~n18102 ;
  assign n18104 = ~n18100 & n18103 ;
  assign n18105 = n18099 & n18104 ;
  assign n18106 = ~n18094 & n18105 ;
  assign n18107 = ~n18091 & n18106 ;
  assign n18108 = ~n18100 & ~n18102 ;
  assign n18109 = n18099 & n18108 ;
  assign n18110 = ~n18094 & n18109 ;
  assign n18111 = ~n18091 & n18110 ;
  assign n18112 = ~\a[29]  & ~n18111 ;
  assign n18113 = ~n18107 & ~n18112 ;
  assign n18114 = n17444 & ~n18088 ;
  assign n18115 = ~n17781 & n18114 ;
  assign n18116 = ~n18113 & ~n18115 ;
  assign n18117 = ~n18089 & n18116 ;
  assign n18118 = ~n18088 & n18113 ;
  assign n18119 = n17782 & n18118 ;
  assign n18120 = n18088 & n18113 ;
  assign n18121 = ~n17782 & n18120 ;
  assign n18122 = ~n18119 & ~n18121 ;
  assign n18123 = ~n18117 & n18122 ;
  assign n18124 = n3402 & ~n5855 ;
  assign n18125 = ~n5853 & n18124 ;
  assign n18126 = \b[33]  & n3400 ;
  assign n18127 = \a[24]  & \b[32]  ;
  assign n18128 = n3391 & n18127 ;
  assign n18129 = ~n18126 & ~n18128 ;
  assign n18130 = \b[31]  & n3733 ;
  assign n18131 = n3730 & n18130 ;
  assign n18132 = ~\a[24]  & \b[32]  ;
  assign n18133 = n3394 & n18132 ;
  assign n18134 = ~n18131 & ~n18133 ;
  assign n18135 = n18129 & n18134 ;
  assign n18136 = ~n18125 & n18135 ;
  assign n18137 = ~\a[26]  & ~n18136 ;
  assign n18138 = \a[26]  & n18135 ;
  assign n18139 = ~n18125 & n18138 ;
  assign n18140 = ~n18137 & ~n18139 ;
  assign n18141 = ~n18123 & ~n18140 ;
  assign n18142 = n17780 & n18141 ;
  assign n18143 = n18123 & ~n18140 ;
  assign n18144 = ~n17780 & n18143 ;
  assign n18145 = ~n18142 & ~n18144 ;
  assign n18146 = ~n18123 & n18140 ;
  assign n18147 = ~n17780 & n18146 ;
  assign n18148 = n18123 & n18140 ;
  assign n18149 = n17780 & n18148 ;
  assign n18150 = ~n18147 & ~n18149 ;
  assign n18151 = n18145 & n18150 ;
  assign n18152 = ~n17777 & ~n18151 ;
  assign n18153 = ~n17753 & n18152 ;
  assign n18154 = ~n17777 & n18151 ;
  assign n18155 = n17753 & n18154 ;
  assign n18156 = ~n18153 & ~n18155 ;
  assign n18157 = n17777 & ~n18151 ;
  assign n18158 = n17753 & n18157 ;
  assign n18159 = n17777 & n18151 ;
  assign n18160 = ~n17753 & n18159 ;
  assign n18161 = ~n18158 & ~n18160 ;
  assign n18162 = n18156 & n18161 ;
  assign n18163 = ~n17752 & ~n18162 ;
  assign n18164 = ~n17494 & n18162 ;
  assign n18165 = ~n17751 & n18164 ;
  assign n18166 = n1965 & ~n8602 ;
  assign n18167 = ~n8600 & n18166 ;
  assign n18168 = \b[39]  & n1963 ;
  assign n18169 = \a[18]  & \b[38]  ;
  assign n18170 = n2210 & n18169 ;
  assign n18171 = ~n18168 & ~n18170 ;
  assign n18172 = \b[37]  & n2218 ;
  assign n18173 = n2216 & n18172 ;
  assign n18174 = ~\a[18]  & \b[38]  ;
  assign n18175 = n1957 & n18174 ;
  assign n18176 = ~n18173 & ~n18175 ;
  assign n18177 = n18171 & n18176 ;
  assign n18178 = ~n18167 & n18177 ;
  assign n18179 = ~\a[20]  & ~n18178 ;
  assign n18180 = \a[20]  & n18177 ;
  assign n18181 = ~n18167 & n18180 ;
  assign n18182 = ~n18179 & ~n18181 ;
  assign n18183 = ~n18165 & ~n18182 ;
  assign n18184 = ~n18163 & n18183 ;
  assign n18185 = ~n18162 & n18182 ;
  assign n18186 = ~n17752 & n18185 ;
  assign n18187 = n18162 & n18182 ;
  assign n18188 = n17752 & n18187 ;
  assign n18189 = ~n18186 & ~n18188 ;
  assign n18190 = ~n18184 & n18189 ;
  assign n18191 = n1467 & n9930 ;
  assign n18192 = ~n9927 & n18191 ;
  assign n18193 = n1467 & ~n9930 ;
  assign n18194 = ~n9477 & n18193 ;
  assign n18195 = ~n9926 & n18194 ;
  assign n18196 = \b[40]  & n1652 ;
  assign n18197 = n1649 & n18196 ;
  assign n18198 = \b[42]  & n1465 ;
  assign n18199 = \a[15]  & \b[41]  ;
  assign n18200 = n1456 & n18199 ;
  assign n18201 = ~\a[15]  & \b[41]  ;
  assign n18202 = n1459 & n18201 ;
  assign n18203 = ~n18200 & ~n18202 ;
  assign n18204 = ~n18198 & n18203 ;
  assign n18205 = ~n18197 & n18204 ;
  assign n18206 = ~n18195 & n18205 ;
  assign n18207 = ~n18192 & n18206 ;
  assign n18208 = ~\a[17]  & ~n18207 ;
  assign n18209 = \a[17]  & n18205 ;
  assign n18210 = ~n18195 & n18209 ;
  assign n18211 = ~n18192 & n18210 ;
  assign n18212 = ~n18208 & ~n18211 ;
  assign n18213 = ~n18190 & n18212 ;
  assign n18214 = n17749 & n18213 ;
  assign n18215 = n18190 & n18212 ;
  assign n18216 = ~n17749 & n18215 ;
  assign n18217 = ~n18214 & ~n18216 ;
  assign n18218 = ~n18190 & ~n18212 ;
  assign n18219 = ~n17749 & n18218 ;
  assign n18220 = n18190 & ~n18212 ;
  assign n18221 = n17749 & n18220 ;
  assign n18222 = ~n18219 & ~n18221 ;
  assign n18223 = n18217 & n18222 ;
  assign n18224 = ~n17748 & ~n18223 ;
  assign n18225 = n17731 & n18224 ;
  assign n18226 = ~n17748 & n18223 ;
  assign n18227 = ~n17731 & n18226 ;
  assign n18228 = ~n18225 & ~n18227 ;
  assign n18229 = n17748 & ~n18223 ;
  assign n18230 = ~n17731 & n18229 ;
  assign n18231 = n17748 & n18223 ;
  assign n18232 = n17731 & n18231 ;
  assign n18233 = ~n18230 & ~n18232 ;
  assign n18234 = n18228 & n18233 ;
  assign n18235 = ~n17728 & n18234 ;
  assign n18236 = n646 & n12478 ;
  assign n18237 = ~n12475 & n18236 ;
  assign n18238 = n646 & ~n12478 ;
  assign n18239 = ~n12433 & n18238 ;
  assign n18240 = ~n12474 & n18239 ;
  assign n18241 = \b[46]  & n796 ;
  assign n18242 = n793 & n18241 ;
  assign n18243 = ~\a[9]  & \b[47]  ;
  assign n18244 = n638 & n18243 ;
  assign n18245 = ~n18242 & ~n18244 ;
  assign n18246 = \b[48]  & n644 ;
  assign n18247 = \a[9]  & \b[47]  ;
  assign n18248 = n635 & n18247 ;
  assign n18249 = \a[11]  & ~n18248 ;
  assign n18250 = ~n18246 & n18249 ;
  assign n18251 = n18245 & n18250 ;
  assign n18252 = ~n18240 & n18251 ;
  assign n18253 = ~n18237 & n18252 ;
  assign n18254 = ~n18246 & ~n18248 ;
  assign n18255 = n18245 & n18254 ;
  assign n18256 = ~n18240 & n18255 ;
  assign n18257 = ~n18237 & n18256 ;
  assign n18258 = ~\a[11]  & ~n18257 ;
  assign n18259 = ~n18253 & ~n18258 ;
  assign n18260 = n17575 & ~n18234 ;
  assign n18261 = ~n17727 & n18260 ;
  assign n18262 = ~n18259 & ~n18261 ;
  assign n18263 = ~n18235 & n18262 ;
  assign n18264 = ~n18234 & n18259 ;
  assign n18265 = n17728 & n18264 ;
  assign n18266 = n18234 & n18259 ;
  assign n18267 = ~n17728 & n18266 ;
  assign n18268 = ~n18265 & ~n18267 ;
  assign n18269 = ~n18263 & n18268 ;
  assign n18270 = ~n17726 & ~n18269 ;
  assign n18271 = n17709 & n18270 ;
  assign n18272 = ~n17726 & n18269 ;
  assign n18273 = ~n17709 & n18272 ;
  assign n18274 = ~n18271 & ~n18273 ;
  assign n18275 = n17726 & ~n18269 ;
  assign n18276 = ~n17709 & n18275 ;
  assign n18277 = n17726 & n18269 ;
  assign n18278 = n17709 & n18277 ;
  assign n18279 = ~n18276 & ~n18278 ;
  assign n18280 = n18274 & n18279 ;
  assign n18281 = ~n17706 & n18280 ;
  assign n18282 = n252 & n16407 ;
  assign n18283 = \b[52]  & n303 ;
  assign n18284 = n300 & n18283 ;
  assign n18285 = ~\a[3]  & \b[53]  ;
  assign n18286 = n244 & n18285 ;
  assign n18287 = ~n18284 & ~n18286 ;
  assign n18288 = \b[54]  & n250 ;
  assign n18289 = \a[3]  & \b[53]  ;
  assign n18290 = n241 & n18289 ;
  assign n18291 = \a[5]  & ~n18290 ;
  assign n18292 = ~n18288 & n18291 ;
  assign n18293 = n18287 & n18292 ;
  assign n18294 = ~n18282 & n18293 ;
  assign n18295 = ~n18288 & ~n18290 ;
  assign n18296 = n18287 & n18295 ;
  assign n18297 = ~\a[5]  & ~n18296 ;
  assign n18298 = ~\a[5]  & n252 ;
  assign n18299 = n16407 & n18298 ;
  assign n18300 = ~n18297 & ~n18299 ;
  assign n18301 = ~n18294 & n18300 ;
  assign n18302 = ~n17621 & ~n18280 ;
  assign n18303 = ~n17705 & n18302 ;
  assign n18304 = ~n18301 & ~n18303 ;
  assign n18305 = ~n18281 & n18304 ;
  assign n18306 = ~n18280 & n18301 ;
  assign n18307 = n17706 & n18306 ;
  assign n18308 = n18280 & n18301 ;
  assign n18309 = ~n17706 & n18308 ;
  assign n18310 = ~n18307 & ~n18309 ;
  assign n18311 = ~n18305 & n18310 ;
  assign n18312 = ~n17704 & ~n18311 ;
  assign n18313 = n17681 & n18312 ;
  assign n18314 = ~n17704 & n18311 ;
  assign n18315 = ~n17681 & n18314 ;
  assign n18316 = ~n18313 & ~n18315 ;
  assign n18317 = n17704 & ~n18311 ;
  assign n18318 = ~n17681 & n18317 ;
  assign n18319 = n17704 & n18311 ;
  assign n18320 = n17681 & n18319 ;
  assign n18321 = ~n18318 & ~n18320 ;
  assign n18322 = n18316 & n18321 ;
  assign n18323 = ~n17678 & n18322 ;
  assign n18324 = ~n17668 & ~n18322 ;
  assign n18325 = ~n17675 & n18324 ;
  assign n18326 = ~n18323 & ~n18325 ;
  assign n18327 = ~n17668 & n18316 ;
  assign n18328 = n18321 & ~n18327 ;
  assign n18329 = n17674 & n18321 ;
  assign n18330 = n17063 & n18329 ;
  assign n18331 = ~n18328 & ~n18330 ;
  assign n18332 = n17681 & n18311 ;
  assign n18333 = ~n18305 & ~n18332 ;
  assign n18334 = ~n17621 & n18274 ;
  assign n18335 = ~n17705 & n18334 ;
  assign n18336 = n18279 & ~n18335 ;
  assign n18337 = n252 & ~n16446 ;
  assign n18338 = ~n16444 & n18337 ;
  assign n18339 = \b[53]  & n303 ;
  assign n18340 = n300 & n18339 ;
  assign n18341 = \b[55]  & n250 ;
  assign n18342 = \a[2]  & \b[54]  ;
  assign n18343 = n301 & n18342 ;
  assign n18344 = ~\a[3]  & \b[54]  ;
  assign n18345 = n244 & n18344 ;
  assign n18346 = ~n18343 & ~n18345 ;
  assign n18347 = ~n18341 & n18346 ;
  assign n18348 = ~n18340 & n18347 ;
  assign n18349 = ~\a[5]  & n18348 ;
  assign n18350 = ~n18338 & n18349 ;
  assign n18351 = ~n18338 & n18348 ;
  assign n18352 = \a[5]  & ~n18351 ;
  assign n18353 = ~n18350 & ~n18352 ;
  assign n18354 = n17709 & n18269 ;
  assign n18355 = ~n18263 & ~n18354 ;
  assign n18356 = ~n15198 & ~n15201 ;
  assign n18357 = n430 & ~n15239 ;
  assign n18358 = ~n18356 & n18357 ;
  assign n18359 = \b[50]  & n486 ;
  assign n18360 = n483 & n18359 ;
  assign n18361 = \b[52]  & n428 ;
  assign n18362 = \a[5]  & \b[51]  ;
  assign n18363 = n484 & n18362 ;
  assign n18364 = ~\a[6]  & \b[51]  ;
  assign n18365 = n422 & n18364 ;
  assign n18366 = ~n18363 & ~n18365 ;
  assign n18367 = ~n18361 & n18366 ;
  assign n18368 = ~n18360 & n18367 ;
  assign n18369 = ~n18358 & n18368 ;
  assign n18370 = ~\a[8]  & ~n18369 ;
  assign n18371 = \a[8]  & n18368 ;
  assign n18372 = ~n18358 & n18371 ;
  assign n18373 = ~n18370 & ~n18372 ;
  assign n18374 = n17575 & n18228 ;
  assign n18375 = ~n17727 & n18374 ;
  assign n18376 = n18233 & ~n18375 ;
  assign n18377 = n646 & ~n13524 ;
  assign n18378 = ~n13522 & n18377 ;
  assign n18379 = \b[47]  & n796 ;
  assign n18380 = n793 & n18379 ;
  assign n18381 = \b[49]  & n644 ;
  assign n18382 = \a[8]  & \b[48]  ;
  assign n18383 = n794 & n18382 ;
  assign n18384 = ~\a[9]  & \b[48]  ;
  assign n18385 = n638 & n18384 ;
  assign n18386 = ~n18383 & ~n18385 ;
  assign n18387 = ~n18381 & n18386 ;
  assign n18388 = ~n18380 & n18387 ;
  assign n18389 = ~n18378 & n18388 ;
  assign n18390 = ~\a[11]  & ~n18389 ;
  assign n18391 = \a[11]  & n18388 ;
  assign n18392 = ~n18378 & n18391 ;
  assign n18393 = ~n18390 & ~n18392 ;
  assign n18394 = n17731 & n18223 ;
  assign n18395 = n18222 & ~n18394 ;
  assign n18396 = ~n847 & ~n11392 ;
  assign n18397 = ~n11906 & n18396 ;
  assign n18398 = ~n11902 & n18397 ;
  assign n18399 = ~n996 & n18398 ;
  assign n18400 = n999 & n11906 ;
  assign n18401 = ~n11903 & n18400 ;
  assign n18402 = ~n18399 & ~n18401 ;
  assign n18403 = \b[44]  & n1182 ;
  assign n18404 = n1179 & n18403 ;
  assign n18405 = \a[11]  & \b[45]  ;
  assign n18406 = n1180 & n18405 ;
  assign n18407 = ~\a[12]  & \b[45]  ;
  assign n18408 = n7674 & n18407 ;
  assign n18409 = ~n18406 & ~n18408 ;
  assign n18410 = ~n18404 & n18409 ;
  assign n18411 = \b[46]  & n997 ;
  assign n18412 = \a[14]  & ~n18411 ;
  assign n18413 = n18410 & n18412 ;
  assign n18414 = n18402 & n18413 ;
  assign n18415 = n18410 & ~n18411 ;
  assign n18416 = n18402 & n18415 ;
  assign n18417 = ~\a[14]  & ~n18416 ;
  assign n18418 = ~n18414 & ~n18417 ;
  assign n18419 = ~n17524 & ~n18184 ;
  assign n18420 = ~n17532 & n18419 ;
  assign n18421 = n18189 & ~n18420 ;
  assign n18422 = n18156 & ~n18165 ;
  assign n18423 = ~n17471 & n18145 ;
  assign n18424 = ~n17473 & n18423 ;
  assign n18425 = n18150 & ~n18424 ;
  assign n18426 = n17780 & n18123 ;
  assign n18427 = ~n18117 & ~n18426 ;
  assign n18428 = n17444 & n18087 ;
  assign n18429 = ~n17781 & n18428 ;
  assign n18430 = n18082 & ~n18429 ;
  assign n18431 = n4249 & ~n5462 ;
  assign n18432 = ~n5460 & n18431 ;
  assign n18433 = \b[29]  & n4647 ;
  assign n18434 = n4644 & n18433 ;
  assign n18435 = ~\a[27]  & \b[30]  ;
  assign n18436 = n4241 & n18435 ;
  assign n18437 = ~n18434 & ~n18436 ;
  assign n18438 = \b[31]  & n4247 ;
  assign n18439 = \a[27]  & \b[30]  ;
  assign n18440 = n4238 & n18439 ;
  assign n18441 = \a[29]  & ~n18440 ;
  assign n18442 = ~n18438 & n18441 ;
  assign n18443 = n18437 & n18442 ;
  assign n18444 = ~n18432 & n18443 ;
  assign n18445 = ~n18438 & ~n18440 ;
  assign n18446 = n18437 & n18445 ;
  assign n18447 = ~n18432 & n18446 ;
  assign n18448 = ~\a[29]  & ~n18447 ;
  assign n18449 = ~n18444 & ~n18448 ;
  assign n18450 = n17785 & n18058 ;
  assign n18451 = n18052 & ~n18450 ;
  assign n18452 = ~n17403 & n18017 ;
  assign n18453 = ~n17410 & n18452 ;
  assign n18454 = n18022 & ~n18453 ;
  assign n18455 = n17789 & n18012 ;
  assign n18456 = ~n18006 & ~n18455 ;
  assign n18457 = n17360 & n17972 ;
  assign n18458 = ~n17815 & n18457 ;
  assign n18459 = n17977 & ~n18458 ;
  assign n18460 = n17819 & n17967 ;
  assign n18461 = ~n17966 & ~n18460 ;
  assign n18462 = ~n17325 & n17950 ;
  assign n18463 = ~n17327 & n18462 ;
  assign n18464 = n17955 & ~n18463 ;
  assign n18465 = n17871 & n17945 ;
  assign n18466 = ~n17943 & ~n18465 ;
  assign n18467 = ~n383 & n14793 ;
  assign n18468 = ~n381 & n18467 ;
  assign n18469 = \b[5]  & n15517 ;
  assign n18470 = n15514 & n18469 ;
  assign n18471 = \b[7]  & n14791 ;
  assign n18472 = \a[50]  & \b[6]  ;
  assign n18473 = n15515 & n18472 ;
  assign n18474 = ~\a[51]  & \b[6]  ;
  assign n18475 = n14785 & n18474 ;
  assign n18476 = ~n18473 & ~n18475 ;
  assign n18477 = ~n18471 & n18476 ;
  assign n18478 = ~n18470 & n18477 ;
  assign n18479 = ~\a[53]  & n18478 ;
  assign n18480 = ~n18468 & n18479 ;
  assign n18481 = ~n18468 & n18478 ;
  assign n18482 = \a[53]  & ~n18481 ;
  assign n18483 = ~n18480 & ~n18482 ;
  assign n18484 = ~n17915 & ~n17918 ;
  assign n18485 = n222 & n16655 ;
  assign n18486 = \b[4]  & n16653 ;
  assign n18487 = \a[53]  & \b[3]  ;
  assign n18488 = n17306 & n18487 ;
  assign n18489 = ~\a[54]  & \b[3]  ;
  assign n18490 = n16647 & n18489 ;
  assign n18491 = ~n18488 & ~n18490 ;
  assign n18492 = ~n18486 & n18491 ;
  assign n18493 = \b[2]  & n17308 ;
  assign n18494 = n17305 & n18493 ;
  assign n18495 = \a[56]  & ~n18494 ;
  assign n18496 = n18492 & n18495 ;
  assign n18497 = ~n18485 & n18496 ;
  assign n18498 = n18492 & ~n18494 ;
  assign n18499 = ~n18485 & n18498 ;
  assign n18500 = ~\a[56]  & ~n18499 ;
  assign n18501 = ~n18497 & ~n18500 ;
  assign n18502 = \a[59]  & \b[0]  ;
  assign n18503 = ~n17912 & n18502 ;
  assign n18504 = \a[57]  & \b[0]  ;
  assign n18505 = \a[56]  & ~\a[58]  ;
  assign n18506 = n18504 & n18505 ;
  assign n18507 = ~\a[57]  & \b[0]  ;
  assign n18508 = ~\a[56]  & \a[58]  ;
  assign n18509 = n18507 & n18508 ;
  assign n18510 = ~n18506 & ~n18509 ;
  assign n18511 = \a[58]  & ~\a[59]  ;
  assign n18512 = ~\a[58]  & \a[59]  ;
  assign n18513 = ~n18511 & ~n18512 ;
  assign n18514 = ~n17912 & n18513 ;
  assign n18515 = \b[1]  & n18514 ;
  assign n18516 = ~n17912 & ~n18513 ;
  assign n18517 = ~n137 & n18516 ;
  assign n18518 = ~n18515 & ~n18517 ;
  assign n18519 = n18510 & n18518 ;
  assign n18520 = n18503 & ~n18519 ;
  assign n18521 = ~n18503 & n18510 ;
  assign n18522 = n18518 & n18521 ;
  assign n18523 = ~n18520 & ~n18522 ;
  assign n18524 = n18501 & ~n18523 ;
  assign n18525 = ~n18501 & n18523 ;
  assign n18526 = ~n18524 & ~n18525 ;
  assign n18527 = ~n18484 & n18526 ;
  assign n18528 = n18484 & ~n18526 ;
  assign n18529 = ~n18527 & ~n18528 ;
  assign n18530 = ~n18483 & ~n18529 ;
  assign n18531 = n18483 & n18529 ;
  assign n18532 = ~n18530 & ~n18531 ;
  assign n18533 = ~n685 & ~n12606 ;
  assign n18534 = ~n13122 & n18533 ;
  assign n18535 = n682 & n18534 ;
  assign n18536 = n685 & ~n12606 ;
  assign n18537 = ~n13122 & n18536 ;
  assign n18538 = ~n682 & n18537 ;
  assign n18539 = ~n18535 & ~n18538 ;
  assign n18540 = \b[8]  & n13794 ;
  assign n18541 = n13792 & n18540 ;
  assign n18542 = ~\a[48]  & \b[9]  ;
  assign n18543 = n13117 & n18542 ;
  assign n18544 = ~n18541 & ~n18543 ;
  assign n18545 = \b[10]  & n13123 ;
  assign n18546 = \a[48]  & \b[9]  ;
  assign n18547 = n13786 & n18546 ;
  assign n18548 = \a[50]  & ~n18547 ;
  assign n18549 = ~n18545 & n18548 ;
  assign n18550 = n18544 & n18549 ;
  assign n18551 = n18539 & n18550 ;
  assign n18552 = ~n18545 & ~n18547 ;
  assign n18553 = n18544 & n18552 ;
  assign n18554 = n18539 & n18553 ;
  assign n18555 = ~\a[50]  & ~n18554 ;
  assign n18556 = ~n18551 & ~n18555 ;
  assign n18557 = ~n18532 & ~n18556 ;
  assign n18558 = ~n18466 & n18557 ;
  assign n18559 = n18532 & ~n18556 ;
  assign n18560 = n18466 & n18559 ;
  assign n18561 = ~n18558 & ~n18560 ;
  assign n18562 = ~n18532 & n18556 ;
  assign n18563 = n18466 & n18562 ;
  assign n18564 = n18532 & n18556 ;
  assign n18565 = ~n18466 & n18564 ;
  assign n18566 = ~n18563 & ~n18565 ;
  assign n18567 = n18561 & n18566 ;
  assign n18568 = ~n948 & n11572 ;
  assign n18569 = ~n908 & n11572 ;
  assign n18570 = ~n912 & n18569 ;
  assign n18571 = ~n18568 & ~n18570 ;
  assign n18572 = ~n951 & ~n18571 ;
  assign n18573 = \b[11]  & n12159 ;
  assign n18574 = n12156 & n18573 ;
  assign n18575 = \b[13]  & n11570 ;
  assign n18576 = \a[44]  & \b[12]  ;
  assign n18577 = n12157 & n18576 ;
  assign n18578 = ~\a[45]  & \b[12]  ;
  assign n18579 = n11564 & n18578 ;
  assign n18580 = ~n18577 & ~n18579 ;
  assign n18581 = ~n18575 & n18580 ;
  assign n18582 = ~n18574 & n18581 ;
  assign n18583 = ~\a[47]  & n18582 ;
  assign n18584 = ~n18572 & n18583 ;
  assign n18585 = \a[47]  & ~n18582 ;
  assign n18586 = \a[47]  & ~n951 ;
  assign n18587 = ~n18571 & n18586 ;
  assign n18588 = ~n18585 & ~n18587 ;
  assign n18589 = ~n18584 & n18588 ;
  assign n18590 = ~n18567 & n18589 ;
  assign n18591 = n18464 & n18590 ;
  assign n18592 = n18567 & n18589 ;
  assign n18593 = ~n18464 & n18592 ;
  assign n18594 = ~n18591 & ~n18593 ;
  assign n18595 = ~n18567 & ~n18589 ;
  assign n18596 = ~n18464 & n18595 ;
  assign n18597 = n18567 & ~n18589 ;
  assign n18598 = n18464 & n18597 ;
  assign n18599 = ~n18596 & ~n18598 ;
  assign n18600 = n18594 & n18599 ;
  assign n18601 = ~n18461 & n18600 ;
  assign n18602 = n1512 & n10082 ;
  assign n18603 = ~n1509 & n18602 ;
  assign n18604 = ~n1512 & n10082 ;
  assign n18605 = ~n1228 & n18604 ;
  assign n18606 = ~n1508 & n18605 ;
  assign n18607 = \b[14]  & n10681 ;
  assign n18608 = n10678 & n18607 ;
  assign n18609 = \b[16]  & n10080 ;
  assign n18610 = \a[41]  & \b[15]  ;
  assign n18611 = n10679 & n18610 ;
  assign n18612 = ~\a[42]  & \b[15]  ;
  assign n18613 = n10074 & n18612 ;
  assign n18614 = ~n18611 & ~n18613 ;
  assign n18615 = ~n18609 & n18614 ;
  assign n18616 = ~n18608 & n18615 ;
  assign n18617 = ~n18606 & n18616 ;
  assign n18618 = ~n18603 & n18617 ;
  assign n18619 = ~\a[44]  & ~n18618 ;
  assign n18620 = \a[44]  & n18616 ;
  assign n18621 = ~n18606 & n18620 ;
  assign n18622 = ~n18603 & n18621 ;
  assign n18623 = ~n18619 & ~n18622 ;
  assign n18624 = ~n17966 & ~n18600 ;
  assign n18625 = ~n18460 & n18624 ;
  assign n18626 = ~n18623 & ~n18625 ;
  assign n18627 = ~n18601 & n18626 ;
  assign n18628 = ~n18600 & n18623 ;
  assign n18629 = n18461 & n18628 ;
  assign n18630 = n18600 & n18623 ;
  assign n18631 = ~n18461 & n18630 ;
  assign n18632 = ~n18629 & ~n18631 ;
  assign n18633 = ~n18627 & n18632 ;
  assign n18634 = ~n2079 & n8759 ;
  assign n18635 = ~n2077 & n18634 ;
  assign n18636 = \b[17]  & n9301 ;
  assign n18637 = n9298 & n18636 ;
  assign n18638 = ~\a[39]  & \b[18]  ;
  assign n18639 = n8751 & n18638 ;
  assign n18640 = ~n18637 & ~n18639 ;
  assign n18641 = \b[19]  & n8757 ;
  assign n18642 = \a[39]  & \b[18]  ;
  assign n18643 = n8748 & n18642 ;
  assign n18644 = \a[41]  & ~n18643 ;
  assign n18645 = ~n18641 & n18644 ;
  assign n18646 = n18640 & n18645 ;
  assign n18647 = ~n18635 & n18646 ;
  assign n18648 = ~n18641 & ~n18643 ;
  assign n18649 = n18640 & n18648 ;
  assign n18650 = ~n18635 & n18649 ;
  assign n18651 = ~\a[41]  & ~n18650 ;
  assign n18652 = ~n18647 & ~n18651 ;
  assign n18653 = ~n18633 & ~n18652 ;
  assign n18654 = n18459 & n18653 ;
  assign n18655 = n18633 & ~n18652 ;
  assign n18656 = ~n18459 & n18655 ;
  assign n18657 = ~n18654 & ~n18656 ;
  assign n18658 = ~n18633 & n18652 ;
  assign n18659 = ~n18459 & n18658 ;
  assign n18660 = n18633 & n18652 ;
  assign n18661 = n18459 & n18660 ;
  assign n18662 = ~n18659 & ~n18661 ;
  assign n18663 = n18657 & n18662 ;
  assign n18664 = ~n18456 & n18663 ;
  assign n18665 = n2768 & n7534 ;
  assign n18666 = ~n2765 & n18665 ;
  assign n18667 = ~n2768 & n7534 ;
  assign n18668 = ~n2518 & n18667 ;
  assign n18669 = ~n2764 & n18668 ;
  assign n18670 = \b[20]  & n7973 ;
  assign n18671 = n7970 & n18670 ;
  assign n18672 = ~\a[36]  & \b[21]  ;
  assign n18673 = n7526 & n18672 ;
  assign n18674 = ~n18671 & ~n18673 ;
  assign n18675 = \b[22]  & n7532 ;
  assign n18676 = \a[36]  & \b[21]  ;
  assign n18677 = n17801 & n18676 ;
  assign n18678 = \a[38]  & ~n18677 ;
  assign n18679 = ~n18675 & n18678 ;
  assign n18680 = n18674 & n18679 ;
  assign n18681 = ~n18669 & n18680 ;
  assign n18682 = ~n18666 & n18681 ;
  assign n18683 = ~n18675 & ~n18677 ;
  assign n18684 = n18674 & n18683 ;
  assign n18685 = ~n18669 & n18684 ;
  assign n18686 = ~n18666 & n18685 ;
  assign n18687 = ~\a[38]  & ~n18686 ;
  assign n18688 = ~n18682 & ~n18687 ;
  assign n18689 = ~n18006 & ~n18663 ;
  assign n18690 = ~n18455 & n18689 ;
  assign n18691 = ~n18688 & ~n18690 ;
  assign n18692 = ~n18664 & n18691 ;
  assign n18693 = ~n18663 & n18688 ;
  assign n18694 = n18456 & n18693 ;
  assign n18695 = n18663 & n18688 ;
  assign n18696 = ~n18456 & n18695 ;
  assign n18697 = ~n18694 & ~n18696 ;
  assign n18698 = ~n18692 & n18697 ;
  assign n18699 = ~n18454 & ~n18698 ;
  assign n18700 = n18454 & n18698 ;
  assign n18701 = ~n18699 & ~n18700 ;
  assign n18702 = ~n3567 & n6309 ;
  assign n18703 = ~n3565 & n18702 ;
  assign n18704 = \b[25]  & n6307 ;
  assign n18705 = \a[33]  & \b[24]  ;
  assign n18706 = n6298 & n18705 ;
  assign n18707 = ~n18704 & ~n18706 ;
  assign n18708 = \b[23]  & n6778 ;
  assign n18709 = n6775 & n18708 ;
  assign n18710 = ~\a[33]  & \b[24]  ;
  assign n18711 = n6301 & n18710 ;
  assign n18712 = ~n18709 & ~n18711 ;
  assign n18713 = n18707 & n18712 ;
  assign n18714 = ~n18703 & n18713 ;
  assign n18715 = ~\a[35]  & ~n18714 ;
  assign n18716 = \a[35]  & n18713 ;
  assign n18717 = ~n18703 & n18716 ;
  assign n18718 = ~n18715 & ~n18717 ;
  assign n18719 = n18701 & ~n18718 ;
  assign n18720 = ~n18701 & n18718 ;
  assign n18721 = ~n18719 & ~n18720 ;
  assign n18722 = n4456 & n5211 ;
  assign n18723 = ~n4143 & ~n4452 ;
  assign n18724 = n18722 & ~n18723 ;
  assign n18725 = ~n4456 & n5211 ;
  assign n18726 = ~n4143 & n18725 ;
  assign n18727 = ~n4452 & n18726 ;
  assign n18728 = \b[26]  & n5595 ;
  assign n18729 = n5592 & n18728 ;
  assign n18730 = ~\a[30]  & \b[27]  ;
  assign n18731 = n5203 & n18730 ;
  assign n18732 = ~n18729 & ~n18731 ;
  assign n18733 = \b[28]  & n5209 ;
  assign n18734 = \a[30]  & \b[27]  ;
  assign n18735 = n5200 & n18734 ;
  assign n18736 = \a[32]  & ~n18735 ;
  assign n18737 = ~n18733 & n18736 ;
  assign n18738 = n18732 & n18737 ;
  assign n18739 = ~n18727 & n18738 ;
  assign n18740 = ~n18724 & n18739 ;
  assign n18741 = ~n18733 & ~n18735 ;
  assign n18742 = n18732 & n18741 ;
  assign n18743 = ~n18727 & n18742 ;
  assign n18744 = ~n18724 & n18743 ;
  assign n18745 = ~\a[32]  & ~n18744 ;
  assign n18746 = ~n18740 & ~n18745 ;
  assign n18747 = ~n18721 & ~n18746 ;
  assign n18748 = ~n18451 & n18747 ;
  assign n18749 = n18721 & ~n18746 ;
  assign n18750 = n18451 & n18749 ;
  assign n18751 = ~n18748 & ~n18750 ;
  assign n18752 = ~n18721 & n18746 ;
  assign n18753 = n18451 & n18752 ;
  assign n18754 = n18721 & n18746 ;
  assign n18755 = ~n18451 & n18754 ;
  assign n18756 = ~n18753 & ~n18755 ;
  assign n18757 = n18751 & n18756 ;
  assign n18758 = ~n18449 & ~n18757 ;
  assign n18759 = n18430 & n18758 ;
  assign n18760 = ~n18449 & n18757 ;
  assign n18761 = ~n18430 & n18760 ;
  assign n18762 = ~n18759 & ~n18761 ;
  assign n18763 = n18449 & ~n18757 ;
  assign n18764 = ~n18430 & n18763 ;
  assign n18765 = n18449 & n18757 ;
  assign n18766 = n18430 & n18765 ;
  assign n18767 = ~n18764 & ~n18766 ;
  assign n18768 = n18762 & n18767 ;
  assign n18769 = ~n18427 & n18768 ;
  assign n18770 = ~n18117 & ~n18768 ;
  assign n18771 = ~n18426 & n18770 ;
  assign n18772 = n3402 & n6565 ;
  assign n18773 = ~n6562 & n18772 ;
  assign n18774 = n3402 & ~n6565 ;
  assign n18775 = ~n5850 & n18774 ;
  assign n18776 = ~n6561 & n18775 ;
  assign n18777 = \b[32]  & n3733 ;
  assign n18778 = n3730 & n18777 ;
  assign n18779 = \b[34]  & n3400 ;
  assign n18780 = \a[23]  & \b[33]  ;
  assign n18781 = n3731 & n18780 ;
  assign n18782 = ~\a[24]  & \b[33]  ;
  assign n18783 = n3394 & n18782 ;
  assign n18784 = ~n18781 & ~n18783 ;
  assign n18785 = ~n18779 & n18784 ;
  assign n18786 = ~n18778 & n18785 ;
  assign n18787 = ~n18776 & n18786 ;
  assign n18788 = ~n18773 & n18787 ;
  assign n18789 = ~\a[26]  & ~n18788 ;
  assign n18790 = \a[26]  & n18786 ;
  assign n18791 = ~n18776 & n18790 ;
  assign n18792 = ~n18773 & n18791 ;
  assign n18793 = ~n18789 & ~n18792 ;
  assign n18794 = ~n18771 & ~n18793 ;
  assign n18795 = ~n18769 & n18794 ;
  assign n18796 = ~n18768 & n18793 ;
  assign n18797 = n18427 & n18796 ;
  assign n18798 = n18768 & n18793 ;
  assign n18799 = ~n18427 & n18798 ;
  assign n18800 = ~n18797 & ~n18799 ;
  assign n18801 = ~n18795 & n18800 ;
  assign n18802 = ~n18425 & ~n18801 ;
  assign n18803 = n18425 & n18801 ;
  assign n18804 = ~n18802 & ~n18803 ;
  assign n18805 = n2622 & ~n7761 ;
  assign n18806 = ~n7759 & n18805 ;
  assign n18807 = \b[35]  & n2912 ;
  assign n18808 = n2909 & n18807 ;
  assign n18809 = \b[37]  & n2620 ;
  assign n18810 = \a[20]  & \b[36]  ;
  assign n18811 = n2910 & n18810 ;
  assign n18812 = ~\a[21]  & \b[36]  ;
  assign n18813 = n2614 & n18812 ;
  assign n18814 = ~n18811 & ~n18813 ;
  assign n18815 = ~n18809 & n18814 ;
  assign n18816 = ~n18808 & n18815 ;
  assign n18817 = ~n18806 & n18816 ;
  assign n18818 = ~\a[23]  & ~n18817 ;
  assign n18819 = \a[23]  & n18816 ;
  assign n18820 = ~n18806 & n18819 ;
  assign n18821 = ~n18818 & ~n18820 ;
  assign n18822 = n18804 & ~n18821 ;
  assign n18823 = ~n18804 & n18821 ;
  assign n18824 = ~n18822 & ~n18823 ;
  assign n18825 = n1965 & n9044 ;
  assign n18826 = ~n9041 & n18825 ;
  assign n18827 = n1965 & ~n9044 ;
  assign n18828 = ~n8597 & n18827 ;
  assign n18829 = ~n9040 & n18828 ;
  assign n18830 = \b[38]  & n2218 ;
  assign n18831 = n2216 & n18830 ;
  assign n18832 = ~\a[18]  & \b[39]  ;
  assign n18833 = n1957 & n18832 ;
  assign n18834 = ~n18831 & ~n18833 ;
  assign n18835 = \b[40]  & n1963 ;
  assign n18836 = \a[18]  & \b[39]  ;
  assign n18837 = n2210 & n18836 ;
  assign n18838 = \a[20]  & ~n18837 ;
  assign n18839 = ~n18835 & n18838 ;
  assign n18840 = n18834 & n18839 ;
  assign n18841 = ~n18829 & n18840 ;
  assign n18842 = ~n18826 & n18841 ;
  assign n18843 = ~n18835 & ~n18837 ;
  assign n18844 = n18834 & n18843 ;
  assign n18845 = ~n18829 & n18844 ;
  assign n18846 = ~n18826 & n18845 ;
  assign n18847 = ~\a[20]  & ~n18846 ;
  assign n18848 = ~n18842 & ~n18847 ;
  assign n18849 = ~n18824 & ~n18848 ;
  assign n18850 = ~n18422 & n18849 ;
  assign n18851 = n18824 & ~n18848 ;
  assign n18852 = n18422 & n18851 ;
  assign n18853 = ~n18850 & ~n18852 ;
  assign n18854 = ~n18824 & n18848 ;
  assign n18855 = n18422 & n18854 ;
  assign n18856 = n18824 & n18848 ;
  assign n18857 = ~n18422 & n18856 ;
  assign n18858 = ~n18855 & ~n18857 ;
  assign n18859 = n18853 & n18858 ;
  assign n18860 = n1467 & ~n10409 ;
  assign n18861 = ~n10407 & n18860 ;
  assign n18862 = \b[43]  & n1465 ;
  assign n18863 = \a[15]  & \b[42]  ;
  assign n18864 = n1456 & n18863 ;
  assign n18865 = ~n18862 & ~n18864 ;
  assign n18866 = \b[41]  & n1652 ;
  assign n18867 = n1649 & n18866 ;
  assign n18868 = ~\a[15]  & \b[42]  ;
  assign n18869 = n1459 & n18868 ;
  assign n18870 = ~n18867 & ~n18869 ;
  assign n18871 = n18865 & n18870 ;
  assign n18872 = ~n18861 & n18871 ;
  assign n18873 = ~\a[17]  & ~n18872 ;
  assign n18874 = \a[17]  & n18871 ;
  assign n18875 = ~n18861 & n18874 ;
  assign n18876 = ~n18873 & ~n18875 ;
  assign n18877 = ~n18859 & ~n18876 ;
  assign n18878 = n18421 & n18877 ;
  assign n18879 = n18859 & ~n18876 ;
  assign n18880 = ~n18421 & n18879 ;
  assign n18881 = ~n18878 & ~n18880 ;
  assign n18882 = ~n18859 & n18876 ;
  assign n18883 = ~n18421 & n18882 ;
  assign n18884 = n18859 & n18876 ;
  assign n18885 = n18421 & n18884 ;
  assign n18886 = ~n18883 & ~n18885 ;
  assign n18887 = n18881 & n18886 ;
  assign n18888 = n18418 & ~n18887 ;
  assign n18889 = n18395 & n18888 ;
  assign n18890 = n18418 & n18887 ;
  assign n18891 = ~n18395 & n18890 ;
  assign n18892 = ~n18889 & ~n18891 ;
  assign n18893 = ~n18395 & n18887 ;
  assign n18894 = n18222 & ~n18887 ;
  assign n18895 = ~n18394 & n18894 ;
  assign n18896 = ~n18418 & ~n18895 ;
  assign n18897 = ~n18893 & n18896 ;
  assign n18898 = n18892 & ~n18897 ;
  assign n18899 = n18393 & ~n18898 ;
  assign n18900 = ~n18376 & n18899 ;
  assign n18901 = n18393 & n18898 ;
  assign n18902 = n18376 & n18901 ;
  assign n18903 = ~n18900 & ~n18902 ;
  assign n18904 = ~n18393 & ~n18898 ;
  assign n18905 = n18376 & n18904 ;
  assign n18906 = ~n18393 & n18898 ;
  assign n18907 = ~n18376 & n18906 ;
  assign n18908 = ~n18905 & ~n18907 ;
  assign n18909 = n18903 & n18908 ;
  assign n18910 = n18373 & ~n18909 ;
  assign n18911 = n18355 & n18910 ;
  assign n18912 = n18373 & n18909 ;
  assign n18913 = ~n18355 & n18912 ;
  assign n18914 = ~n18911 & ~n18913 ;
  assign n18915 = ~n18355 & n18909 ;
  assign n18916 = ~n18263 & ~n18909 ;
  assign n18917 = ~n18354 & n18916 ;
  assign n18918 = ~n18373 & ~n18917 ;
  assign n18919 = ~n18915 & n18918 ;
  assign n18920 = n18914 & ~n18919 ;
  assign n18921 = ~n18353 & ~n18920 ;
  assign n18922 = ~n18336 & n18921 ;
  assign n18923 = ~n18353 & n18920 ;
  assign n18924 = n18336 & n18923 ;
  assign n18925 = ~n18922 & ~n18924 ;
  assign n18926 = n18353 & ~n18920 ;
  assign n18927 = n18336 & n18926 ;
  assign n18928 = n18353 & n18920 ;
  assign n18929 = ~n18336 & n18928 ;
  assign n18930 = ~n18927 & ~n18929 ;
  assign n18931 = n18925 & n18930 ;
  assign n18932 = ~n18333 & n18931 ;
  assign n18933 = ~n18305 & ~n18931 ;
  assign n18934 = ~n18332 & n18933 ;
  assign n18935 = ~n17646 & ~n17686 ;
  assign n18936 = ~n17683 & n18935 ;
  assign n18937 = ~n17685 & ~n18936 ;
  assign n18938 = ~\b[57]  & ~\b[58]  ;
  assign n18939 = \b[57]  & \b[58]  ;
  assign n18940 = ~n18938 & ~n18939 ;
  assign n18941 = n134 & n18940 ;
  assign n18942 = ~n18937 & n18941 ;
  assign n18943 = n134 & ~n18940 ;
  assign n18944 = ~n17685 & n18943 ;
  assign n18945 = ~n18936 & n18944 ;
  assign n18946 = \a[0]  & \b[58]  ;
  assign n18947 = n133 & n18946 ;
  assign n18948 = \b[57]  & n141 ;
  assign n18949 = ~\a[1]  & \b[56]  ;
  assign n18950 = n10416 & n18949 ;
  assign n18951 = ~n18948 & ~n18950 ;
  assign n18952 = ~n18947 & n18951 ;
  assign n18953 = \a[2]  & n18952 ;
  assign n18954 = ~n18945 & n18953 ;
  assign n18955 = ~n18942 & n18954 ;
  assign n18956 = ~n18945 & n18952 ;
  assign n18957 = ~n18942 & n18956 ;
  assign n18958 = ~\a[2]  & ~n18957 ;
  assign n18959 = ~n18955 & ~n18958 ;
  assign n18960 = ~n18934 & ~n18959 ;
  assign n18961 = ~n18932 & n18960 ;
  assign n18962 = ~n18931 & n18959 ;
  assign n18963 = n18333 & n18962 ;
  assign n18964 = n18931 & n18959 ;
  assign n18965 = ~n18333 & n18964 ;
  assign n18966 = ~n18963 & ~n18965 ;
  assign n18967 = ~n18961 & n18966 ;
  assign n18968 = ~n18331 & n18967 ;
  assign n18969 = n18331 & ~n18967 ;
  assign n18970 = ~n18968 & ~n18969 ;
  assign n18971 = ~n18961 & ~n18968 ;
  assign n18972 = n18336 & n18920 ;
  assign n18973 = ~n18919 & ~n18972 ;
  assign n18974 = ~n18263 & n18908 ;
  assign n18975 = ~n18354 & n18974 ;
  assign n18976 = n18903 & ~n18975 ;
  assign n18977 = n430 & ~n15246 ;
  assign n18978 = ~n15244 & n18977 ;
  assign n18979 = \b[51]  & n486 ;
  assign n18980 = n483 & n18979 ;
  assign n18981 = \b[53]  & n428 ;
  assign n18982 = \a[5]  & \b[52]  ;
  assign n18983 = n484 & n18982 ;
  assign n18984 = ~\a[6]  & \b[52]  ;
  assign n18985 = n422 & n18984 ;
  assign n18986 = ~n18983 & ~n18985 ;
  assign n18987 = ~n18981 & n18986 ;
  assign n18988 = ~n18980 & n18987 ;
  assign n18989 = ~n18978 & n18988 ;
  assign n18990 = ~\a[8]  & ~n18989 ;
  assign n18991 = \a[8]  & n18988 ;
  assign n18992 = ~n18978 & n18991 ;
  assign n18993 = ~n18990 & ~n18992 ;
  assign n18994 = n18376 & n18898 ;
  assign n18995 = ~n18897 & ~n18994 ;
  assign n18996 = n18222 & n18881 ;
  assign n18997 = ~n18394 & n18996 ;
  assign n18998 = n18886 & ~n18997 ;
  assign n18999 = n999 & ~n12438 ;
  assign n19000 = ~n12436 & n18999 ;
  assign n19001 = \b[45]  & n1182 ;
  assign n19002 = n1179 & n19001 ;
  assign n19003 = \b[47]  & n997 ;
  assign n19004 = \a[11]  & \b[46]  ;
  assign n19005 = n1180 & n19004 ;
  assign n19006 = ~\a[12]  & \b[46]  ;
  assign n19007 = n7674 & n19006 ;
  assign n19008 = ~n19005 & ~n19007 ;
  assign n19009 = ~n19003 & n19008 ;
  assign n19010 = ~n19002 & n19009 ;
  assign n19011 = ~n19000 & n19010 ;
  assign n19012 = ~\a[14]  & ~n19011 ;
  assign n19013 = \a[14]  & n19010 ;
  assign n19014 = ~n19000 & n19013 ;
  assign n19015 = ~n19012 & ~n19014 ;
  assign n19016 = n18421 & n18859 ;
  assign n19017 = n18853 & ~n19016 ;
  assign n19018 = n18156 & ~n18822 ;
  assign n19019 = ~n18165 & n19018 ;
  assign n19020 = ~n18823 & ~n19019 ;
  assign n19021 = ~n18795 & ~n18803 ;
  assign n19022 = ~n18117 & n18762 ;
  assign n19023 = ~n18426 & n19022 ;
  assign n19024 = n18767 & ~n19023 ;
  assign n19025 = n18430 & n18757 ;
  assign n19026 = n18751 & ~n19025 ;
  assign n19027 = n4249 & n5810 ;
  assign n19028 = ~n5807 & n19027 ;
  assign n19029 = ~n5457 & ~n5810 ;
  assign n19030 = n4249 & n19029 ;
  assign n19031 = ~n5806 & n19030 ;
  assign n19032 = \b[30]  & n4647 ;
  assign n19033 = n4644 & n19032 ;
  assign n19034 = ~\a[27]  & \b[31]  ;
  assign n19035 = n4241 & n19034 ;
  assign n19036 = ~n19033 & ~n19035 ;
  assign n19037 = \b[32]  & n4247 ;
  assign n19038 = \a[27]  & \b[31]  ;
  assign n19039 = n4238 & n19038 ;
  assign n19040 = \a[29]  & ~n19039 ;
  assign n19041 = ~n19037 & n19040 ;
  assign n19042 = n19036 & n19041 ;
  assign n19043 = ~n19031 & n19042 ;
  assign n19044 = ~n19028 & n19043 ;
  assign n19045 = ~n19037 & ~n19039 ;
  assign n19046 = n19036 & n19045 ;
  assign n19047 = ~n19031 & n19046 ;
  assign n19048 = ~n19028 & n19047 ;
  assign n19049 = ~\a[29]  & ~n19048 ;
  assign n19050 = ~n19044 & ~n19049 ;
  assign n19051 = n18052 & ~n18719 ;
  assign n19052 = ~n18450 & n19051 ;
  assign n19053 = ~n18720 & ~n19052 ;
  assign n19054 = ~n18692 & ~n18700 ;
  assign n19055 = ~n18006 & n18657 ;
  assign n19056 = ~n18455 & n19055 ;
  assign n19057 = n18662 & ~n19056 ;
  assign n19058 = ~n3022 & n7534 ;
  assign n19059 = ~n3020 & n19058 ;
  assign n19060 = \b[23]  & n7532 ;
  assign n19061 = \a[36]  & \b[22]  ;
  assign n19062 = n17801 & n19061 ;
  assign n19063 = ~n19060 & ~n19062 ;
  assign n19064 = \b[21]  & n7973 ;
  assign n19065 = n7970 & n19064 ;
  assign n19066 = ~\a[36]  & \b[22]  ;
  assign n19067 = n7526 & n19066 ;
  assign n19068 = ~n19065 & ~n19067 ;
  assign n19069 = n19063 & n19068 ;
  assign n19070 = ~n19059 & n19069 ;
  assign n19071 = ~\a[38]  & ~n19070 ;
  assign n19072 = \a[38]  & n19069 ;
  assign n19073 = ~n19059 & n19072 ;
  assign n19074 = ~n19071 & ~n19073 ;
  assign n19075 = n18459 & n18633 ;
  assign n19076 = ~n18627 & ~n19075 ;
  assign n19077 = ~n1694 & n10082 ;
  assign n19078 = ~n1692 & n19077 ;
  assign n19079 = \b[15]  & n10681 ;
  assign n19080 = n10678 & n19079 ;
  assign n19081 = \b[17]  & n10080 ;
  assign n19082 = \a[41]  & \b[16]  ;
  assign n19083 = n10679 & n19082 ;
  assign n19084 = ~\a[42]  & \b[16]  ;
  assign n19085 = n10074 & n19084 ;
  assign n19086 = ~n19083 & ~n19085 ;
  assign n19087 = ~n19081 & n19086 ;
  assign n19088 = ~n19080 & n19087 ;
  assign n19089 = ~n19078 & n19088 ;
  assign n19090 = ~\a[44]  & ~n19089 ;
  assign n19091 = \a[44]  & n19088 ;
  assign n19092 = ~n19078 & n19091 ;
  assign n19093 = ~n19090 & ~n19092 ;
  assign n19094 = ~n17966 & n18594 ;
  assign n19095 = n18599 & ~n19094 ;
  assign n19096 = n17967 & n18599 ;
  assign n19097 = n17819 & n19096 ;
  assign n19098 = ~n19095 & ~n19097 ;
  assign n19099 = n18464 & n18567 ;
  assign n19100 = n18561 & ~n19099 ;
  assign n19101 = ~n725 & n13125 ;
  assign n19102 = ~n684 & n13125 ;
  assign n19103 = ~n721 & n19102 ;
  assign n19104 = ~n19101 & ~n19103 ;
  assign n19105 = ~n728 & ~n19104 ;
  assign n19106 = \b[9]  & n13794 ;
  assign n19107 = n13792 & n19106 ;
  assign n19108 = ~\a[48]  & \b[10]  ;
  assign n19109 = n13117 & n19108 ;
  assign n19110 = ~n19107 & ~n19109 ;
  assign n19111 = \b[11]  & n13123 ;
  assign n19112 = \a[48]  & \b[10]  ;
  assign n19113 = n13786 & n19112 ;
  assign n19114 = \a[50]  & ~n19113 ;
  assign n19115 = ~n19111 & n19114 ;
  assign n19116 = n19110 & n19115 ;
  assign n19117 = ~n19105 & n19116 ;
  assign n19118 = ~n19111 & ~n19113 ;
  assign n19119 = n19110 & n19118 ;
  assign n19120 = ~\a[50]  & ~n19119 ;
  assign n19121 = ~\a[50]  & ~n728 ;
  assign n19122 = ~n19104 & n19121 ;
  assign n19123 = ~n19120 & ~n19122 ;
  assign n19124 = ~n19117 & n19123 ;
  assign n19125 = ~n17943 & ~n18531 ;
  assign n19126 = ~n18465 & n19125 ;
  assign n19127 = ~n18530 & ~n19126 ;
  assign n19128 = ~n505 & ~n14276 ;
  assign n19129 = ~n14790 & n19128 ;
  assign n19130 = n502 & n19129 ;
  assign n19131 = n505 & ~n14276 ;
  assign n19132 = ~n14790 & n19131 ;
  assign n19133 = ~n502 & n19132 ;
  assign n19134 = ~n19130 & ~n19133 ;
  assign n19135 = \b[6]  & n15517 ;
  assign n19136 = n15514 & n19135 ;
  assign n19137 = \b[8]  & n14791 ;
  assign n19138 = \a[50]  & \b[7]  ;
  assign n19139 = n15515 & n19138 ;
  assign n19140 = ~\a[51]  & \b[7]  ;
  assign n19141 = n14785 & n19140 ;
  assign n19142 = ~n19139 & ~n19141 ;
  assign n19143 = ~n19137 & n19142 ;
  assign n19144 = ~n19136 & n19143 ;
  assign n19145 = n19134 & n19144 ;
  assign n19146 = ~\a[53]  & ~n19145 ;
  assign n19147 = \a[53]  & n19144 ;
  assign n19148 = n19134 & n19147 ;
  assign n19149 = ~n19146 & ~n19148 ;
  assign n19150 = ~n18525 & ~n18527 ;
  assign n19151 = ~n273 & n16655 ;
  assign n19152 = ~n271 & n19151 ;
  assign n19153 = \b[3]  & n17308 ;
  assign n19154 = n17305 & n19153 ;
  assign n19155 = \b[5]  & n16653 ;
  assign n19156 = \a[53]  & \b[4]  ;
  assign n19157 = n17306 & n19156 ;
  assign n19158 = ~\a[54]  & \b[4]  ;
  assign n19159 = n16647 & n19158 ;
  assign n19160 = ~n19157 & ~n19159 ;
  assign n19161 = ~n19155 & n19160 ;
  assign n19162 = ~n19154 & n19161 ;
  assign n19163 = ~\a[56]  & n19162 ;
  assign n19164 = ~n19152 & n19163 ;
  assign n19165 = ~n19152 & n19162 ;
  assign n19166 = \a[56]  & ~n19165 ;
  assign n19167 = ~n19164 & ~n19166 ;
  assign n19168 = \a[59]  & ~n17913 ;
  assign n19169 = n18510 & n19168 ;
  assign n19170 = n18518 & n19169 ;
  assign n19171 = \a[59]  & ~n19170 ;
  assign n19172 = \b[2]  & n18514 ;
  assign n19173 = ~\a[57]  & \b[1]  ;
  assign n19174 = n18508 & n19173 ;
  assign n19175 = \a[57]  & \b[1]  ;
  assign n19176 = n18505 & n19175 ;
  assign n19177 = ~n19174 & ~n19176 ;
  assign n19178 = ~n19172 & n19177 ;
  assign n19179 = n157 & n18516 ;
  assign n19180 = n17912 & ~n18513 ;
  assign n19181 = \a[57]  & ~\a[58]  ;
  assign n19182 = ~\a[57]  & \a[58]  ;
  assign n19183 = ~n19181 & ~n19182 ;
  assign n19184 = \b[0]  & n19183 ;
  assign n19185 = n19180 & n19184 ;
  assign n19186 = ~n19179 & ~n19185 ;
  assign n19187 = n19178 & n19186 ;
  assign n19188 = ~n19171 & ~n19187 ;
  assign n19189 = n19171 & n19187 ;
  assign n19190 = ~n19188 & ~n19189 ;
  assign n19191 = n19167 & ~n19190 ;
  assign n19192 = ~n19167 & n19190 ;
  assign n19193 = ~n19191 & ~n19192 ;
  assign n19194 = ~n19150 & n19193 ;
  assign n19195 = n19150 & ~n19193 ;
  assign n19196 = ~n19194 & ~n19195 ;
  assign n19197 = n19149 & ~n19196 ;
  assign n19198 = ~n19149 & n19196 ;
  assign n19199 = ~n19197 & ~n19198 ;
  assign n19200 = n19127 & n19199 ;
  assign n19201 = ~n19127 & ~n19199 ;
  assign n19202 = ~n19200 & ~n19201 ;
  assign n19203 = n19124 & ~n19202 ;
  assign n19204 = ~n19124 & n19202 ;
  assign n19205 = ~n19203 & ~n19204 ;
  assign n19206 = n1087 & n11572 ;
  assign n19207 = ~n1084 & n19206 ;
  assign n19208 = ~n1087 & n11572 ;
  assign n19209 = ~n946 & n19208 ;
  assign n19210 = ~n1083 & n19209 ;
  assign n19211 = \b[12]  & n12159 ;
  assign n19212 = n12156 & n19211 ;
  assign n19213 = \b[14]  & n11570 ;
  assign n19214 = \a[44]  & \b[13]  ;
  assign n19215 = n12157 & n19214 ;
  assign n19216 = ~\a[45]  & \b[13]  ;
  assign n19217 = n11564 & n19216 ;
  assign n19218 = ~n19215 & ~n19217 ;
  assign n19219 = ~n19213 & n19218 ;
  assign n19220 = ~n19212 & n19219 ;
  assign n19221 = ~n19210 & n19220 ;
  assign n19222 = ~n19207 & n19221 ;
  assign n19223 = ~\a[47]  & ~n19222 ;
  assign n19224 = \a[47]  & n19220 ;
  assign n19225 = ~n19210 & n19224 ;
  assign n19226 = ~n19207 & n19225 ;
  assign n19227 = ~n19223 & ~n19226 ;
  assign n19228 = ~n19205 & ~n19227 ;
  assign n19229 = ~n19100 & n19228 ;
  assign n19230 = n19205 & ~n19227 ;
  assign n19231 = n19100 & n19230 ;
  assign n19232 = ~n19229 & ~n19231 ;
  assign n19233 = ~n19205 & n19227 ;
  assign n19234 = n19100 & n19233 ;
  assign n19235 = n19205 & n19227 ;
  assign n19236 = ~n19100 & n19235 ;
  assign n19237 = ~n19234 & ~n19236 ;
  assign n19238 = n19232 & n19237 ;
  assign n19239 = ~n19098 & n19238 ;
  assign n19240 = n19098 & ~n19238 ;
  assign n19241 = ~n19239 & ~n19240 ;
  assign n19242 = ~n19093 & n19241 ;
  assign n19243 = n19093 & ~n19241 ;
  assign n19244 = ~n19242 & ~n19243 ;
  assign n19245 = ~n19076 & n19244 ;
  assign n19246 = n2293 & n8759 ;
  assign n19247 = ~n2074 & ~n2289 ;
  assign n19248 = n19246 & ~n19247 ;
  assign n19249 = n5705 & n8759 ;
  assign n19250 = ~n2289 & n19249 ;
  assign n19251 = \b[18]  & n9301 ;
  assign n19252 = n9298 & n19251 ;
  assign n19253 = ~\a[39]  & \b[19]  ;
  assign n19254 = n8751 & n19253 ;
  assign n19255 = ~n19252 & ~n19254 ;
  assign n19256 = \b[20]  & n8757 ;
  assign n19257 = \a[39]  & \b[19]  ;
  assign n19258 = n8748 & n19257 ;
  assign n19259 = \a[41]  & ~n19258 ;
  assign n19260 = ~n19256 & n19259 ;
  assign n19261 = n19255 & n19260 ;
  assign n19262 = ~n19250 & n19261 ;
  assign n19263 = ~n19248 & n19262 ;
  assign n19264 = ~n19256 & ~n19258 ;
  assign n19265 = n19255 & n19264 ;
  assign n19266 = ~n19250 & n19265 ;
  assign n19267 = ~n19248 & n19266 ;
  assign n19268 = ~\a[41]  & ~n19267 ;
  assign n19269 = ~n19263 & ~n19268 ;
  assign n19270 = ~n18627 & ~n19244 ;
  assign n19271 = ~n19075 & n19270 ;
  assign n19272 = ~n19269 & ~n19271 ;
  assign n19273 = ~n19245 & n19272 ;
  assign n19274 = ~n19244 & n19269 ;
  assign n19275 = n19076 & n19274 ;
  assign n19276 = n19244 & n19269 ;
  assign n19277 = ~n19076 & n19276 ;
  assign n19278 = ~n19275 & ~n19277 ;
  assign n19279 = ~n19273 & n19278 ;
  assign n19280 = ~n19074 & ~n19279 ;
  assign n19281 = n19057 & n19280 ;
  assign n19282 = ~n19074 & n19279 ;
  assign n19283 = ~n19057 & n19282 ;
  assign n19284 = ~n19281 & ~n19283 ;
  assign n19285 = n19074 & ~n19279 ;
  assign n19286 = ~n19057 & n19285 ;
  assign n19287 = n19074 & n19279 ;
  assign n19288 = n19057 & n19287 ;
  assign n19289 = ~n19286 & ~n19288 ;
  assign n19290 = n19284 & n19289 ;
  assign n19291 = n3604 & n6309 ;
  assign n19292 = ~n3562 & ~n3600 ;
  assign n19293 = n19291 & ~n19292 ;
  assign n19294 = ~n3604 & n6309 ;
  assign n19295 = ~n3562 & n19294 ;
  assign n19296 = ~n3600 & n19295 ;
  assign n19297 = \b[24]  & n6778 ;
  assign n19298 = n6775 & n19297 ;
  assign n19299 = ~\a[33]  & \b[25]  ;
  assign n19300 = n6301 & n19299 ;
  assign n19301 = ~n19298 & ~n19300 ;
  assign n19302 = \b[26]  & n6307 ;
  assign n19303 = \a[33]  & \b[25]  ;
  assign n19304 = n6298 & n19303 ;
  assign n19305 = \a[35]  & ~n19304 ;
  assign n19306 = ~n19302 & n19305 ;
  assign n19307 = n19301 & n19306 ;
  assign n19308 = ~n19296 & n19307 ;
  assign n19309 = ~n19293 & n19308 ;
  assign n19310 = ~n19302 & ~n19304 ;
  assign n19311 = n19301 & n19310 ;
  assign n19312 = ~n19296 & n19311 ;
  assign n19313 = ~n19293 & n19312 ;
  assign n19314 = ~\a[35]  & ~n19313 ;
  assign n19315 = ~n19309 & ~n19314 ;
  assign n19316 = ~n19290 & ~n19315 ;
  assign n19317 = ~n19054 & n19316 ;
  assign n19318 = n19290 & ~n19315 ;
  assign n19319 = n19054 & n19318 ;
  assign n19320 = ~n19317 & ~n19319 ;
  assign n19321 = ~n19290 & n19315 ;
  assign n19322 = n19054 & n19321 ;
  assign n19323 = n19290 & n19315 ;
  assign n19324 = ~n19054 & n19323 ;
  assign n19325 = ~n19322 & ~n19324 ;
  assign n19326 = n19320 & n19325 ;
  assign n19327 = ~n4502 & n5211 ;
  assign n19328 = ~n4500 & n19327 ;
  assign n19329 = \b[27]  & n5595 ;
  assign n19330 = n5592 & n19329 ;
  assign n19331 = ~\a[30]  & \b[28]  ;
  assign n19332 = n5203 & n19331 ;
  assign n19333 = ~n19330 & ~n19332 ;
  assign n19334 = \b[29]  & n5209 ;
  assign n19335 = \a[30]  & \b[28]  ;
  assign n19336 = n5200 & n19335 ;
  assign n19337 = \a[32]  & ~n19336 ;
  assign n19338 = ~n19334 & n19337 ;
  assign n19339 = n19333 & n19338 ;
  assign n19340 = ~n19328 & n19339 ;
  assign n19341 = ~n19334 & ~n19336 ;
  assign n19342 = n19333 & n19341 ;
  assign n19343 = ~n19328 & n19342 ;
  assign n19344 = ~\a[32]  & ~n19343 ;
  assign n19345 = ~n19340 & ~n19344 ;
  assign n19346 = ~n19326 & ~n19345 ;
  assign n19347 = n19053 & n19346 ;
  assign n19348 = n19326 & ~n19345 ;
  assign n19349 = ~n19053 & n19348 ;
  assign n19350 = ~n19347 & ~n19349 ;
  assign n19351 = ~n19326 & n19345 ;
  assign n19352 = ~n19053 & n19351 ;
  assign n19353 = n19326 & n19345 ;
  assign n19354 = n19053 & n19353 ;
  assign n19355 = ~n19352 & ~n19354 ;
  assign n19356 = n19350 & n19355 ;
  assign n19357 = n19050 & ~n19356 ;
  assign n19358 = n19026 & n19357 ;
  assign n19359 = n19050 & n19356 ;
  assign n19360 = ~n19026 & n19359 ;
  assign n19361 = ~n19358 & ~n19360 ;
  assign n19362 = ~n19026 & n19356 ;
  assign n19363 = n18751 & ~n19356 ;
  assign n19364 = ~n19025 & n19363 ;
  assign n19365 = ~n19050 & ~n19364 ;
  assign n19366 = ~n19362 & n19365 ;
  assign n19367 = n19361 & ~n19366 ;
  assign n19368 = n3402 & ~n6610 ;
  assign n19369 = ~n6608 & n19368 ;
  assign n19370 = \b[33]  & n3733 ;
  assign n19371 = n3730 & n19370 ;
  assign n19372 = \b[35]  & n3400 ;
  assign n19373 = \a[23]  & \b[34]  ;
  assign n19374 = n3731 & n19373 ;
  assign n19375 = ~\a[24]  & \b[34]  ;
  assign n19376 = n3394 & n19375 ;
  assign n19377 = ~n19374 & ~n19376 ;
  assign n19378 = ~n19372 & n19377 ;
  assign n19379 = ~n19371 & n19378 ;
  assign n19380 = ~n19369 & n19379 ;
  assign n19381 = ~\a[26]  & ~n19380 ;
  assign n19382 = \a[26]  & n19379 ;
  assign n19383 = ~n19369 & n19382 ;
  assign n19384 = ~n19381 & ~n19383 ;
  assign n19385 = ~n19367 & ~n19384 ;
  assign n19386 = n19024 & n19385 ;
  assign n19387 = n19367 & ~n19384 ;
  assign n19388 = ~n19024 & n19387 ;
  assign n19389 = ~n19386 & ~n19388 ;
  assign n19390 = ~n19367 & n19384 ;
  assign n19391 = ~n19024 & n19390 ;
  assign n19392 = n19367 & n19384 ;
  assign n19393 = n19024 & n19392 ;
  assign n19394 = ~n19391 & ~n19393 ;
  assign n19395 = n19389 & n19394 ;
  assign n19396 = n2622 & n8175 ;
  assign n19397 = ~n8172 & n19396 ;
  assign n19398 = n2622 & ~n8175 ;
  assign n19399 = ~n7756 & n19398 ;
  assign n19400 = ~n8171 & n19399 ;
  assign n19401 = \b[36]  & n2912 ;
  assign n19402 = n2909 & n19401 ;
  assign n19403 = \b[38]  & n2620 ;
  assign n19404 = \a[20]  & \b[37]  ;
  assign n19405 = n2910 & n19404 ;
  assign n19406 = ~\a[21]  & \b[37]  ;
  assign n19407 = n2614 & n19406 ;
  assign n19408 = ~n19405 & ~n19407 ;
  assign n19409 = ~n19403 & n19408 ;
  assign n19410 = ~n19402 & n19409 ;
  assign n19411 = ~n19400 & n19410 ;
  assign n19412 = ~n19397 & n19411 ;
  assign n19413 = ~\a[23]  & ~n19412 ;
  assign n19414 = \a[23]  & n19410 ;
  assign n19415 = ~n19400 & n19414 ;
  assign n19416 = ~n19397 & n19415 ;
  assign n19417 = ~n19413 & ~n19416 ;
  assign n19418 = ~n19395 & ~n19417 ;
  assign n19419 = ~n19021 & n19418 ;
  assign n19420 = n19395 & ~n19417 ;
  assign n19421 = n19021 & n19420 ;
  assign n19422 = ~n19419 & ~n19421 ;
  assign n19423 = ~n19395 & n19417 ;
  assign n19424 = n19021 & n19423 ;
  assign n19425 = n19395 & n19417 ;
  assign n19426 = ~n19021 & n19425 ;
  assign n19427 = ~n19424 & ~n19426 ;
  assign n19428 = n19422 & n19427 ;
  assign n19429 = n1965 & ~n9482 ;
  assign n19430 = ~n9480 & n19429 ;
  assign n19431 = \b[41]  & n1963 ;
  assign n19432 = \a[18]  & \b[40]  ;
  assign n19433 = n2210 & n19432 ;
  assign n19434 = ~n19431 & ~n19433 ;
  assign n19435 = \b[39]  & n2218 ;
  assign n19436 = n2216 & n19435 ;
  assign n19437 = ~\a[18]  & \b[40]  ;
  assign n19438 = n1957 & n19437 ;
  assign n19439 = ~n19436 & ~n19438 ;
  assign n19440 = n19434 & n19439 ;
  assign n19441 = ~n19430 & n19440 ;
  assign n19442 = ~\a[20]  & ~n19441 ;
  assign n19443 = \a[20]  & n19440 ;
  assign n19444 = ~n19430 & n19443 ;
  assign n19445 = ~n19442 & ~n19444 ;
  assign n19446 = ~n19428 & ~n19445 ;
  assign n19447 = n19020 & n19446 ;
  assign n19448 = n19428 & ~n19445 ;
  assign n19449 = ~n19020 & n19448 ;
  assign n19450 = ~n19447 & ~n19449 ;
  assign n19451 = ~n19428 & n19445 ;
  assign n19452 = ~n19020 & n19451 ;
  assign n19453 = n19428 & n19445 ;
  assign n19454 = n19020 & n19453 ;
  assign n19455 = ~n19452 & ~n19454 ;
  assign n19456 = n19450 & n19455 ;
  assign n19457 = ~n19017 & n19456 ;
  assign n19458 = n1467 & ~n10892 ;
  assign n19459 = ~n10890 & n19458 ;
  assign n19460 = \b[42]  & n1652 ;
  assign n19461 = n1649 & n19460 ;
  assign n19462 = ~\a[15]  & \b[43]  ;
  assign n19463 = n1459 & n19462 ;
  assign n19464 = ~n19461 & ~n19463 ;
  assign n19465 = \b[44]  & n1465 ;
  assign n19466 = \a[15]  & \b[43]  ;
  assign n19467 = n1456 & n19466 ;
  assign n19468 = \a[17]  & ~n19467 ;
  assign n19469 = ~n19465 & n19468 ;
  assign n19470 = n19464 & n19469 ;
  assign n19471 = ~n19459 & n19470 ;
  assign n19472 = ~n19465 & ~n19467 ;
  assign n19473 = n19464 & n19472 ;
  assign n19474 = ~n19459 & n19473 ;
  assign n19475 = ~\a[17]  & ~n19474 ;
  assign n19476 = ~n19471 & ~n19475 ;
  assign n19477 = n18853 & ~n19456 ;
  assign n19478 = ~n19016 & n19477 ;
  assign n19479 = ~n19476 & ~n19478 ;
  assign n19480 = ~n19457 & n19479 ;
  assign n19481 = ~n19456 & n19476 ;
  assign n19482 = n19017 & n19481 ;
  assign n19483 = n19456 & n19476 ;
  assign n19484 = ~n19017 & n19483 ;
  assign n19485 = ~n19482 & ~n19484 ;
  assign n19486 = ~n19480 & n19485 ;
  assign n19487 = ~n19015 & ~n19486 ;
  assign n19488 = n18998 & n19487 ;
  assign n19489 = ~n19015 & n19486 ;
  assign n19490 = ~n18998 & n19489 ;
  assign n19491 = ~n19488 & ~n19490 ;
  assign n19492 = n19015 & ~n19486 ;
  assign n19493 = ~n18998 & n19492 ;
  assign n19494 = n19015 & n19486 ;
  assign n19495 = n18998 & n19494 ;
  assign n19496 = ~n19493 & ~n19495 ;
  assign n19497 = n19491 & n19496 ;
  assign n19498 = ~n18995 & n19497 ;
  assign n19499 = ~n18897 & ~n19497 ;
  assign n19500 = ~n18994 & n19499 ;
  assign n19501 = n646 & n14052 ;
  assign n19502 = ~n14049 & n19501 ;
  assign n19503 = n646 & ~n14052 ;
  assign n19504 = ~n13519 & n19503 ;
  assign n19505 = ~n14048 & n19504 ;
  assign n19506 = \b[48]  & n796 ;
  assign n19507 = n793 & n19506 ;
  assign n19508 = \b[50]  & n644 ;
  assign n19509 = \a[8]  & \b[49]  ;
  assign n19510 = n794 & n19509 ;
  assign n19511 = ~\a[9]  & \b[49]  ;
  assign n19512 = n638 & n19511 ;
  assign n19513 = ~n19510 & ~n19512 ;
  assign n19514 = ~n19508 & n19513 ;
  assign n19515 = ~n19507 & n19514 ;
  assign n19516 = ~n19505 & n19515 ;
  assign n19517 = ~n19502 & n19516 ;
  assign n19518 = ~\a[11]  & ~n19517 ;
  assign n19519 = \a[11]  & n19515 ;
  assign n19520 = ~n19505 & n19519 ;
  assign n19521 = ~n19502 & n19520 ;
  assign n19522 = ~n19518 & ~n19521 ;
  assign n19523 = ~n19500 & ~n19522 ;
  assign n19524 = ~n19498 & n19523 ;
  assign n19525 = ~n19497 & n19522 ;
  assign n19526 = n18995 & n19525 ;
  assign n19527 = n19497 & n19522 ;
  assign n19528 = ~n18995 & n19527 ;
  assign n19529 = ~n19526 & ~n19528 ;
  assign n19530 = ~n19524 & n19529 ;
  assign n19531 = ~n18993 & ~n19530 ;
  assign n19532 = n18976 & n19531 ;
  assign n19533 = ~n18993 & n19530 ;
  assign n19534 = ~n18976 & n19533 ;
  assign n19535 = ~n19532 & ~n19534 ;
  assign n19536 = n18993 & ~n19530 ;
  assign n19537 = ~n18976 & n19536 ;
  assign n19538 = n18993 & n19530 ;
  assign n19539 = n18976 & n19538 ;
  assign n19540 = ~n19537 & ~n19539 ;
  assign n19541 = n19535 & n19540 ;
  assign n19542 = ~n17685 & n18940 ;
  assign n19543 = ~n18936 & n19542 ;
  assign n19544 = ~n18939 & ~n19543 ;
  assign n19545 = ~\b[58]  & ~\b[59]  ;
  assign n19546 = \b[58]  & \b[59]  ;
  assign n19547 = ~n19545 & ~n19546 ;
  assign n19548 = ~n19544 & n19547 ;
  assign n19549 = ~n18939 & ~n19547 ;
  assign n19550 = ~n19543 & n19549 ;
  assign n19551 = n134 & ~n19550 ;
  assign n19552 = ~n19548 & n19551 ;
  assign n19553 = \a[0]  & \b[59]  ;
  assign n19554 = n133 & n19553 ;
  assign n19555 = \b[58]  & n141 ;
  assign n19556 = ~\a[1]  & \b[57]  ;
  assign n19557 = n10416 & n19556 ;
  assign n19558 = ~n19555 & ~n19557 ;
  assign n19559 = ~n19554 & n19558 ;
  assign n19560 = \a[2]  & n19559 ;
  assign n19561 = ~n19552 & n19560 ;
  assign n19562 = ~n19552 & n19559 ;
  assign n19563 = ~\a[2]  & ~n19562 ;
  assign n19564 = ~n19561 & ~n19563 ;
  assign n19565 = n252 & n17647 ;
  assign n19566 = ~n17644 & n19565 ;
  assign n19567 = ~n16441 & ~n17647 ;
  assign n19568 = n252 & n19567 ;
  assign n19569 = ~n17643 & n19568 ;
  assign n19570 = \b[54]  & n303 ;
  assign n19571 = n300 & n19570 ;
  assign n19572 = ~\a[3]  & \b[55]  ;
  assign n19573 = n244 & n19572 ;
  assign n19574 = ~n19571 & ~n19573 ;
  assign n19575 = \b[56]  & n250 ;
  assign n19576 = \a[3]  & \b[55]  ;
  assign n19577 = n241 & n19576 ;
  assign n19578 = \a[5]  & ~n19577 ;
  assign n19579 = ~n19575 & n19578 ;
  assign n19580 = n19574 & n19579 ;
  assign n19581 = ~n19569 & n19580 ;
  assign n19582 = ~n19566 & n19581 ;
  assign n19583 = ~n19575 & ~n19577 ;
  assign n19584 = n19574 & n19583 ;
  assign n19585 = ~n19569 & n19584 ;
  assign n19586 = ~n19566 & n19585 ;
  assign n19587 = ~\a[5]  & ~n19586 ;
  assign n19588 = ~n19582 & ~n19587 ;
  assign n19589 = ~n19564 & n19588 ;
  assign n19590 = ~n19541 & n19589 ;
  assign n19591 = ~n18973 & n19590 ;
  assign n19592 = ~n19564 & ~n19588 ;
  assign n19593 = n19541 & n19592 ;
  assign n19594 = ~n18973 & n19593 ;
  assign n19595 = ~n19591 & ~n19594 ;
  assign n19596 = ~n19541 & n19592 ;
  assign n19597 = n18973 & n19596 ;
  assign n19598 = n19541 & n19589 ;
  assign n19599 = n18973 & n19598 ;
  assign n19600 = ~n19597 & ~n19599 ;
  assign n19601 = n19595 & n19600 ;
  assign n19602 = ~n18305 & n18930 ;
  assign n19603 = ~n18332 & n19602 ;
  assign n19604 = n18925 & ~n19603 ;
  assign n19605 = ~n19561 & ~n19588 ;
  assign n19606 = ~n19541 & n19605 ;
  assign n19607 = ~n18973 & n19606 ;
  assign n19608 = ~n19561 & n19588 ;
  assign n19609 = n19541 & n19608 ;
  assign n19610 = ~n18973 & n19609 ;
  assign n19611 = ~n19607 & ~n19610 ;
  assign n19612 = ~n19541 & n19608 ;
  assign n19613 = n18973 & n19612 ;
  assign n19614 = n19541 & n19605 ;
  assign n19615 = n18973 & n19614 ;
  assign n19616 = ~n19613 & ~n19615 ;
  assign n19617 = n19611 & n19616 ;
  assign n19618 = ~n19563 & ~n19617 ;
  assign n19619 = n19604 & ~n19618 ;
  assign n19620 = n19601 & n19619 ;
  assign n19621 = n19564 & ~n19588 ;
  assign n19622 = ~n19541 & n19621 ;
  assign n19623 = ~n18973 & n19622 ;
  assign n19624 = n19564 & n19588 ;
  assign n19625 = n19541 & n19624 ;
  assign n19626 = ~n18973 & n19625 ;
  assign n19627 = ~n19623 & ~n19626 ;
  assign n19628 = ~n19541 & n19624 ;
  assign n19629 = n18973 & n19628 ;
  assign n19630 = n19541 & n19621 ;
  assign n19631 = n18973 & n19630 ;
  assign n19632 = ~n19629 & ~n19631 ;
  assign n19633 = n19627 & n19632 ;
  assign n19634 = ~n19604 & ~n19633 ;
  assign n19635 = ~n18973 & n19541 ;
  assign n19636 = ~n18919 & ~n19541 ;
  assign n19637 = ~n18972 & n19636 ;
  assign n19638 = ~n19588 & ~n19637 ;
  assign n19639 = ~n19635 & n19638 ;
  assign n19640 = ~n19541 & n19588 ;
  assign n19641 = n18973 & n19640 ;
  assign n19642 = n19541 & n19588 ;
  assign n19643 = ~n18973 & n19642 ;
  assign n19644 = ~n19641 & ~n19643 ;
  assign n19645 = ~n19639 & n19644 ;
  assign n19646 = ~n19564 & n19645 ;
  assign n19647 = ~n19604 & n19646 ;
  assign n19648 = ~n19634 & ~n19647 ;
  assign n19649 = ~n19620 & n19648 ;
  assign n19650 = ~n18971 & n19649 ;
  assign n19651 = n18971 & ~n19649 ;
  assign n19652 = ~n19650 & ~n19651 ;
  assign n19653 = ~n19620 & ~n19649 ;
  assign n19654 = ~n18961 & ~n19620 ;
  assign n19655 = ~n18968 & n19654 ;
  assign n19656 = ~n19653 & ~n19655 ;
  assign n19657 = ~n18919 & n19535 ;
  assign n19658 = ~n18972 & n19657 ;
  assign n19659 = n19540 & ~n19658 ;
  assign n19660 = n18976 & n19530 ;
  assign n19661 = ~n19524 & ~n19660 ;
  assign n19662 = ~n18897 & n19491 ;
  assign n19663 = ~n18994 & n19662 ;
  assign n19664 = n19496 & ~n19663 ;
  assign n19665 = n646 & ~n14098 ;
  assign n19666 = ~n14096 & n19665 ;
  assign n19667 = \b[49]  & n796 ;
  assign n19668 = n793 & n19667 ;
  assign n19669 = \b[51]  & n644 ;
  assign n19670 = \a[8]  & \b[50]  ;
  assign n19671 = n794 & n19670 ;
  assign n19672 = ~\a[9]  & \b[50]  ;
  assign n19673 = n638 & n19672 ;
  assign n19674 = ~n19671 & ~n19673 ;
  assign n19675 = ~n19669 & n19674 ;
  assign n19676 = ~n19668 & n19675 ;
  assign n19677 = ~n19666 & n19676 ;
  assign n19678 = ~\a[11]  & ~n19677 ;
  assign n19679 = \a[11]  & n19676 ;
  assign n19680 = ~n19666 & n19679 ;
  assign n19681 = ~n19678 & ~n19680 ;
  assign n19682 = n18998 & n19486 ;
  assign n19683 = ~n19480 & ~n19682 ;
  assign n19684 = n18853 & n19450 ;
  assign n19685 = ~n19016 & n19684 ;
  assign n19686 = n19455 & ~n19685 ;
  assign n19687 = n1467 & ~n11397 ;
  assign n19688 = ~n11395 & n19687 ;
  assign n19689 = \b[45]  & n1465 ;
  assign n19690 = \a[15]  & \b[44]  ;
  assign n19691 = n1456 & n19690 ;
  assign n19692 = ~n19689 & ~n19691 ;
  assign n19693 = \b[43]  & n1652 ;
  assign n19694 = n1649 & n19693 ;
  assign n19695 = ~\a[15]  & \b[44]  ;
  assign n19696 = n1459 & n19695 ;
  assign n19697 = ~n19694 & ~n19696 ;
  assign n19698 = n19692 & n19697 ;
  assign n19699 = ~n19688 & n19698 ;
  assign n19700 = ~\a[17]  & ~n19699 ;
  assign n19701 = \a[17]  & n19698 ;
  assign n19702 = ~n19688 & n19701 ;
  assign n19703 = ~n19700 & ~n19702 ;
  assign n19704 = n19020 & n19428 ;
  assign n19705 = n19422 & ~n19704 ;
  assign n19706 = ~n18795 & n19389 ;
  assign n19707 = ~n18803 & n19706 ;
  assign n19708 = n19394 & ~n19707 ;
  assign n19709 = n19024 & n19367 ;
  assign n19710 = ~n19366 & ~n19709 ;
  assign n19711 = n18751 & n19350 ;
  assign n19712 = ~n19025 & n19711 ;
  assign n19713 = n19355 & ~n19712 ;
  assign n19714 = n19053 & n19326 ;
  assign n19715 = n19320 & ~n19714 ;
  assign n19716 = ~n18692 & n19284 ;
  assign n19717 = ~n18700 & n19716 ;
  assign n19718 = n19289 & ~n19717 ;
  assign n19719 = n19057 & n19279 ;
  assign n19720 = ~n19273 & ~n19719 ;
  assign n19721 = ~n18627 & ~n19242 ;
  assign n19722 = ~n19243 & ~n19721 ;
  assign n19723 = n18633 & ~n19243 ;
  assign n19724 = n18459 & n19723 ;
  assign n19725 = ~n19722 & ~n19724 ;
  assign n19726 = ~n2520 & n8759 ;
  assign n19727 = ~n2292 & n8759 ;
  assign n19728 = ~n2516 & n19727 ;
  assign n19729 = ~n19726 & ~n19728 ;
  assign n19730 = ~n2523 & ~n19729 ;
  assign n19731 = \b[19]  & n9301 ;
  assign n19732 = n9298 & n19731 ;
  assign n19733 = ~\a[39]  & \b[20]  ;
  assign n19734 = n8751 & n19733 ;
  assign n19735 = ~n19732 & ~n19734 ;
  assign n19736 = \b[21]  & n8757 ;
  assign n19737 = \a[39]  & \b[20]  ;
  assign n19738 = n8748 & n19737 ;
  assign n19739 = \a[41]  & ~n19738 ;
  assign n19740 = ~n19736 & n19739 ;
  assign n19741 = n19735 & n19740 ;
  assign n19742 = ~n19730 & n19741 ;
  assign n19743 = ~n19736 & ~n19738 ;
  assign n19744 = n19735 & n19743 ;
  assign n19745 = ~\a[41]  & ~n19744 ;
  assign n19746 = ~\a[41]  & ~n2523 ;
  assign n19747 = ~n19729 & n19746 ;
  assign n19748 = ~n19745 & ~n19747 ;
  assign n19749 = ~n19742 & n19748 ;
  assign n19750 = n19232 & ~n19239 ;
  assign n19751 = n1875 & n10082 ;
  assign n19752 = ~n1872 & n19751 ;
  assign n19753 = ~n1875 & n10082 ;
  assign n19754 = ~n1689 & n19753 ;
  assign n19755 = ~n1871 & n19754 ;
  assign n19756 = \b[16]  & n10681 ;
  assign n19757 = n10678 & n19756 ;
  assign n19758 = \b[18]  & n10080 ;
  assign n19759 = \a[41]  & \b[17]  ;
  assign n19760 = n10679 & n19759 ;
  assign n19761 = ~\a[42]  & \b[17]  ;
  assign n19762 = n10074 & n19761 ;
  assign n19763 = ~n19760 & ~n19762 ;
  assign n19764 = ~n19758 & n19763 ;
  assign n19765 = ~n19757 & n19764 ;
  assign n19766 = ~n19755 & n19765 ;
  assign n19767 = ~n19752 & n19766 ;
  assign n19768 = ~\a[44]  & ~n19767 ;
  assign n19769 = \a[44]  & n19765 ;
  assign n19770 = ~n19755 & n19769 ;
  assign n19771 = ~n19752 & n19770 ;
  assign n19772 = ~n19768 & ~n19771 ;
  assign n19773 = n18561 & ~n19204 ;
  assign n19774 = ~n19099 & n19773 ;
  assign n19775 = ~n19203 & ~n19774 ;
  assign n19776 = ~n1233 & n11572 ;
  assign n19777 = ~n1231 & n19776 ;
  assign n19778 = \b[13]  & n12159 ;
  assign n19779 = n12156 & n19778 ;
  assign n19780 = \b[15]  & n11570 ;
  assign n19781 = \a[44]  & \b[14]  ;
  assign n19782 = n12157 & n19781 ;
  assign n19783 = ~\a[45]  & \b[14]  ;
  assign n19784 = n11564 & n19783 ;
  assign n19785 = ~n19782 & ~n19784 ;
  assign n19786 = ~n19780 & n19785 ;
  assign n19787 = ~n19779 & n19786 ;
  assign n19788 = ~\a[47]  & n19787 ;
  assign n19789 = ~n19777 & n19788 ;
  assign n19790 = ~n19777 & n19787 ;
  assign n19791 = \a[47]  & ~n19790 ;
  assign n19792 = ~n19789 & ~n19791 ;
  assign n19793 = ~n19198 & ~n19200 ;
  assign n19794 = ~n909 & ~n12606 ;
  assign n19795 = ~n13122 & n19794 ;
  assign n19796 = n906 & n19795 ;
  assign n19797 = n909 & ~n12606 ;
  assign n19798 = ~n13122 & n19797 ;
  assign n19799 = ~n906 & n19798 ;
  assign n19800 = ~n19796 & ~n19799 ;
  assign n19801 = \b[10]  & n13794 ;
  assign n19802 = n13792 & n19801 ;
  assign n19803 = ~\a[48]  & \b[11]  ;
  assign n19804 = n13117 & n19803 ;
  assign n19805 = ~n19802 & ~n19804 ;
  assign n19806 = \b[12]  & n13123 ;
  assign n19807 = \a[48]  & \b[11]  ;
  assign n19808 = n13786 & n19807 ;
  assign n19809 = \a[50]  & ~n19808 ;
  assign n19810 = ~n19806 & n19809 ;
  assign n19811 = n19805 & n19810 ;
  assign n19812 = n19800 & n19811 ;
  assign n19813 = ~n19806 & ~n19808 ;
  assign n19814 = n19805 & n19813 ;
  assign n19815 = n19800 & n19814 ;
  assign n19816 = ~\a[50]  & ~n19815 ;
  assign n19817 = ~n19812 & ~n19816 ;
  assign n19818 = ~n18525 & ~n19191 ;
  assign n19819 = ~n18527 & n19818 ;
  assign n19820 = ~n19192 & ~n19819 ;
  assign n19821 = ~n586 & n14793 ;
  assign n19822 = ~n504 & n14793 ;
  assign n19823 = ~n508 & n19822 ;
  assign n19824 = ~n19821 & ~n19823 ;
  assign n19825 = ~n589 & ~n19824 ;
  assign n19826 = \b[7]  & n15517 ;
  assign n19827 = n15514 & n19826 ;
  assign n19828 = \b[9]  & n14791 ;
  assign n19829 = \a[50]  & \b[8]  ;
  assign n19830 = n15515 & n19829 ;
  assign n19831 = ~\a[51]  & \b[8]  ;
  assign n19832 = n14785 & n19831 ;
  assign n19833 = ~n19830 & ~n19832 ;
  assign n19834 = ~n19828 & n19833 ;
  assign n19835 = ~n19827 & n19834 ;
  assign n19836 = ~\a[53]  & n19835 ;
  assign n19837 = ~n19825 & n19836 ;
  assign n19838 = \a[53]  & ~n19835 ;
  assign n19839 = \a[53]  & ~n589 ;
  assign n19840 = ~n19824 & n19839 ;
  assign n19841 = ~n19838 & ~n19840 ;
  assign n19842 = ~n19837 & n19841 ;
  assign n19843 = n177 & n18516 ;
  assign n19844 = \b[3]  & n18514 ;
  assign n19845 = \a[56]  & \b[2]  ;
  assign n19846 = n19181 & n19845 ;
  assign n19847 = ~\a[57]  & \b[2]  ;
  assign n19848 = n18508 & n19847 ;
  assign n19849 = ~n19846 & ~n19848 ;
  assign n19850 = ~n19844 & n19849 ;
  assign n19851 = ~n19843 & n19850 ;
  assign n19852 = \b[1]  & n19183 ;
  assign n19853 = n19180 & n19852 ;
  assign n19854 = ~\a[59]  & ~n19853 ;
  assign n19855 = n19851 & n19854 ;
  assign n19856 = n19851 & ~n19853 ;
  assign n19857 = \a[59]  & ~n19856 ;
  assign n19858 = ~n19855 & ~n19857 ;
  assign n19859 = \a[59]  & ~\a[60]  ;
  assign n19860 = ~\a[59]  & \a[60]  ;
  assign n19861 = ~n19859 & ~n19860 ;
  assign n19862 = \b[0]  & ~n19861 ;
  assign n19863 = n19170 & n19187 ;
  assign n19864 = n19862 & n19863 ;
  assign n19865 = ~n19862 & ~n19863 ;
  assign n19866 = ~n19864 & ~n19865 ;
  assign n19867 = n19858 & n19866 ;
  assign n19868 = ~n19858 & ~n19866 ;
  assign n19869 = ~n19867 & ~n19868 ;
  assign n19870 = ~n323 & ~n16016 ;
  assign n19871 = ~n16652 & n19870 ;
  assign n19872 = n320 & n19871 ;
  assign n19873 = n323 & ~n16016 ;
  assign n19874 = ~n16652 & n19873 ;
  assign n19875 = ~n320 & n19874 ;
  assign n19876 = ~n19872 & ~n19875 ;
  assign n19877 = \b[4]  & n17308 ;
  assign n19878 = n17305 & n19877 ;
  assign n19879 = \b[6]  & n16653 ;
  assign n19880 = \a[53]  & \b[5]  ;
  assign n19881 = n17306 & n19880 ;
  assign n19882 = ~\a[54]  & \b[5]  ;
  assign n19883 = n16647 & n19882 ;
  assign n19884 = ~n19881 & ~n19883 ;
  assign n19885 = ~n19879 & n19884 ;
  assign n19886 = ~n19878 & n19885 ;
  assign n19887 = n19876 & n19886 ;
  assign n19888 = ~\a[56]  & ~n19887 ;
  assign n19889 = \a[56]  & n19886 ;
  assign n19890 = n19876 & n19889 ;
  assign n19891 = ~n19888 & ~n19890 ;
  assign n19892 = n19869 & ~n19891 ;
  assign n19893 = ~n19869 & n19891 ;
  assign n19894 = ~n19892 & ~n19893 ;
  assign n19895 = n19842 & ~n19894 ;
  assign n19896 = n19820 & n19895 ;
  assign n19897 = n19842 & n19894 ;
  assign n19898 = ~n19820 & n19897 ;
  assign n19899 = ~n19896 & ~n19898 ;
  assign n19900 = ~n19842 & ~n19894 ;
  assign n19901 = ~n19820 & n19900 ;
  assign n19902 = ~n19842 & n19894 ;
  assign n19903 = n19820 & n19902 ;
  assign n19904 = ~n19901 & ~n19903 ;
  assign n19905 = n19899 & n19904 ;
  assign n19906 = n19817 & ~n19905 ;
  assign n19907 = n19793 & n19906 ;
  assign n19908 = n19817 & n19905 ;
  assign n19909 = ~n19793 & n19908 ;
  assign n19910 = ~n19907 & ~n19909 ;
  assign n19911 = ~n19793 & n19905 ;
  assign n19912 = ~n19198 & ~n19905 ;
  assign n19913 = ~n19200 & n19912 ;
  assign n19914 = ~n19817 & ~n19913 ;
  assign n19915 = ~n19911 & n19914 ;
  assign n19916 = n19910 & ~n19915 ;
  assign n19917 = n19792 & ~n19916 ;
  assign n19918 = n19775 & n19917 ;
  assign n19919 = n19792 & n19916 ;
  assign n19920 = ~n19775 & n19919 ;
  assign n19921 = ~n19918 & ~n19920 ;
  assign n19922 = ~n19792 & ~n19916 ;
  assign n19923 = ~n19775 & n19922 ;
  assign n19924 = ~n19792 & n19916 ;
  assign n19925 = n19775 & n19924 ;
  assign n19926 = ~n19923 & ~n19925 ;
  assign n19927 = n19921 & n19926 ;
  assign n19928 = ~n19772 & ~n19927 ;
  assign n19929 = ~n19750 & n19928 ;
  assign n19930 = ~n19772 & n19927 ;
  assign n19931 = n19750 & n19930 ;
  assign n19932 = ~n19929 & ~n19931 ;
  assign n19933 = n19772 & ~n19927 ;
  assign n19934 = n19750 & n19933 ;
  assign n19935 = n19772 & n19927 ;
  assign n19936 = ~n19750 & n19935 ;
  assign n19937 = ~n19934 & ~n19936 ;
  assign n19938 = n19932 & n19937 ;
  assign n19939 = ~n19749 & ~n19938 ;
  assign n19940 = ~n19725 & n19939 ;
  assign n19941 = ~n19749 & n19938 ;
  assign n19942 = n19725 & n19941 ;
  assign n19943 = ~n19940 & ~n19942 ;
  assign n19944 = n19749 & ~n19938 ;
  assign n19945 = n19725 & n19944 ;
  assign n19946 = n19749 & n19938 ;
  assign n19947 = ~n19725 & n19946 ;
  assign n19948 = ~n19945 & ~n19947 ;
  assign n19949 = n19943 & n19948 ;
  assign n19950 = ~n19720 & n19949 ;
  assign n19951 = ~n19273 & ~n19949 ;
  assign n19952 = ~n19719 & n19951 ;
  assign n19953 = ~n3283 & ~n7098 ;
  assign n19954 = ~n7531 & n19953 ;
  assign n19955 = n3280 & n19954 ;
  assign n19956 = n3283 & ~n7098 ;
  assign n19957 = ~n7531 & n19956 ;
  assign n19958 = ~n3280 & n19957 ;
  assign n19959 = ~n19955 & ~n19958 ;
  assign n19960 = \b[22]  & n7973 ;
  assign n19961 = n7970 & n19960 ;
  assign n19962 = ~\a[36]  & \b[23]  ;
  assign n19963 = n7526 & n19962 ;
  assign n19964 = ~n19961 & ~n19963 ;
  assign n19965 = \b[24]  & n7532 ;
  assign n19966 = \a[36]  & \b[23]  ;
  assign n19967 = n17801 & n19966 ;
  assign n19968 = \a[38]  & ~n19967 ;
  assign n19969 = ~n19965 & n19968 ;
  assign n19970 = n19964 & n19969 ;
  assign n19971 = n19959 & n19970 ;
  assign n19972 = ~n19965 & ~n19967 ;
  assign n19973 = n19964 & n19972 ;
  assign n19974 = n19959 & n19973 ;
  assign n19975 = ~\a[38]  & ~n19974 ;
  assign n19976 = ~n19971 & ~n19975 ;
  assign n19977 = ~n19952 & ~n19976 ;
  assign n19978 = ~n19950 & n19977 ;
  assign n19979 = ~n19949 & n19976 ;
  assign n19980 = n19720 & n19979 ;
  assign n19981 = n19949 & n19976 ;
  assign n19982 = ~n19720 & n19981 ;
  assign n19983 = ~n19980 & ~n19982 ;
  assign n19984 = ~n19978 & n19983 ;
  assign n19985 = ~n19718 & ~n19984 ;
  assign n19986 = n19718 & n19984 ;
  assign n19987 = ~n19985 & ~n19986 ;
  assign n19988 = ~n4148 & n6309 ;
  assign n19989 = ~n4146 & n19988 ;
  assign n19990 = \b[25]  & n6778 ;
  assign n19991 = n6775 & n19990 ;
  assign n19992 = ~\a[33]  & \b[26]  ;
  assign n19993 = n6301 & n19992 ;
  assign n19994 = ~n19991 & ~n19993 ;
  assign n19995 = \b[27]  & n6307 ;
  assign n19996 = \a[33]  & \b[26]  ;
  assign n19997 = n6298 & n19996 ;
  assign n19998 = \a[35]  & ~n19997 ;
  assign n19999 = ~n19995 & n19998 ;
  assign n20000 = n19994 & n19999 ;
  assign n20001 = ~n19989 & n20000 ;
  assign n20002 = ~n19995 & ~n19997 ;
  assign n20003 = n19994 & n20002 ;
  assign n20004 = ~n19989 & n20003 ;
  assign n20005 = ~\a[35]  & ~n20004 ;
  assign n20006 = ~n20001 & ~n20005 ;
  assign n20007 = n19987 & ~n20006 ;
  assign n20008 = ~n19987 & n20006 ;
  assign n20009 = ~n20007 & ~n20008 ;
  assign n20010 = n5105 & n5211 ;
  assign n20011 = ~n5102 & n20010 ;
  assign n20012 = n5211 & n18092 ;
  assign n20013 = ~n5101 & n20012 ;
  assign n20014 = \b[28]  & n5595 ;
  assign n20015 = n5592 & n20014 ;
  assign n20016 = ~\a[30]  & \b[29]  ;
  assign n20017 = n5203 & n20016 ;
  assign n20018 = ~n20015 & ~n20017 ;
  assign n20019 = \b[30]  & n5209 ;
  assign n20020 = \a[30]  & \b[29]  ;
  assign n20021 = n5200 & n20020 ;
  assign n20022 = \a[32]  & ~n20021 ;
  assign n20023 = ~n20019 & n20022 ;
  assign n20024 = n20018 & n20023 ;
  assign n20025 = ~n20013 & n20024 ;
  assign n20026 = ~n20011 & n20025 ;
  assign n20027 = ~n20019 & ~n20021 ;
  assign n20028 = n20018 & n20027 ;
  assign n20029 = ~n20013 & n20028 ;
  assign n20030 = ~n20011 & n20029 ;
  assign n20031 = ~\a[32]  & ~n20030 ;
  assign n20032 = ~n20026 & ~n20031 ;
  assign n20033 = ~n20009 & n20032 ;
  assign n20034 = n19715 & n20033 ;
  assign n20035 = n20009 & n20032 ;
  assign n20036 = ~n19715 & n20035 ;
  assign n20037 = ~n20034 & ~n20036 ;
  assign n20038 = ~n20009 & ~n20032 ;
  assign n20039 = ~n19715 & n20038 ;
  assign n20040 = n20009 & ~n20032 ;
  assign n20041 = n19715 & n20040 ;
  assign n20042 = ~n20039 & ~n20041 ;
  assign n20043 = n20037 & n20042 ;
  assign n20044 = n4249 & ~n5855 ;
  assign n20045 = ~n5853 & n20044 ;
  assign n20046 = \b[33]  & n4247 ;
  assign n20047 = \a[27]  & \b[32]  ;
  assign n20048 = n4238 & n20047 ;
  assign n20049 = ~n20046 & ~n20048 ;
  assign n20050 = \b[31]  & n4647 ;
  assign n20051 = n4644 & n20050 ;
  assign n20052 = ~\a[27]  & \b[32]  ;
  assign n20053 = n4241 & n20052 ;
  assign n20054 = ~n20051 & ~n20053 ;
  assign n20055 = n20049 & n20054 ;
  assign n20056 = ~n20045 & n20055 ;
  assign n20057 = ~\a[29]  & ~n20056 ;
  assign n20058 = \a[29]  & n20055 ;
  assign n20059 = ~n20045 & n20058 ;
  assign n20060 = ~n20057 & ~n20059 ;
  assign n20061 = ~n20043 & ~n20060 ;
  assign n20062 = n19713 & n20061 ;
  assign n20063 = n20043 & ~n20060 ;
  assign n20064 = ~n19713 & n20063 ;
  assign n20065 = ~n20062 & ~n20064 ;
  assign n20066 = ~n20043 & n20060 ;
  assign n20067 = ~n19713 & n20066 ;
  assign n20068 = n20043 & n20060 ;
  assign n20069 = n19713 & n20068 ;
  assign n20070 = ~n20067 & ~n20069 ;
  assign n20071 = n20065 & n20070 ;
  assign n20072 = ~n19710 & n20071 ;
  assign n20073 = n3402 & n7337 ;
  assign n20074 = ~n7334 & n20073 ;
  assign n20075 = n3402 & ~n7337 ;
  assign n20076 = ~n6605 & n20075 ;
  assign n20077 = ~n7333 & n20076 ;
  assign n20078 = \b[34]  & n3733 ;
  assign n20079 = n3730 & n20078 ;
  assign n20080 = \b[36]  & n3400 ;
  assign n20081 = \a[23]  & \b[35]  ;
  assign n20082 = n3731 & n20081 ;
  assign n20083 = ~\a[24]  & \b[35]  ;
  assign n20084 = n3394 & n20083 ;
  assign n20085 = ~n20082 & ~n20084 ;
  assign n20086 = ~n20080 & n20085 ;
  assign n20087 = ~n20079 & n20086 ;
  assign n20088 = ~n20077 & n20087 ;
  assign n20089 = ~n20074 & n20088 ;
  assign n20090 = ~\a[26]  & ~n20089 ;
  assign n20091 = \a[26]  & n20087 ;
  assign n20092 = ~n20077 & n20091 ;
  assign n20093 = ~n20074 & n20092 ;
  assign n20094 = ~n20090 & ~n20093 ;
  assign n20095 = ~n19366 & ~n20071 ;
  assign n20096 = ~n19709 & n20095 ;
  assign n20097 = ~n20094 & ~n20096 ;
  assign n20098 = ~n20072 & n20097 ;
  assign n20099 = ~n20071 & n20094 ;
  assign n20100 = n19710 & n20099 ;
  assign n20101 = n20071 & n20094 ;
  assign n20102 = ~n19710 & n20101 ;
  assign n20103 = ~n20100 & ~n20102 ;
  assign n20104 = ~n20098 & n20103 ;
  assign n20105 = ~n19708 & ~n20104 ;
  assign n20106 = n19708 & n20104 ;
  assign n20107 = ~n20105 & ~n20106 ;
  assign n20108 = n2622 & ~n8602 ;
  assign n20109 = ~n8600 & n20108 ;
  assign n20110 = \b[37]  & n2912 ;
  assign n20111 = n2909 & n20110 ;
  assign n20112 = \b[39]  & n2620 ;
  assign n20113 = \a[20]  & \b[38]  ;
  assign n20114 = n2910 & n20113 ;
  assign n20115 = ~\a[21]  & \b[38]  ;
  assign n20116 = n2614 & n20115 ;
  assign n20117 = ~n20114 & ~n20116 ;
  assign n20118 = ~n20112 & n20117 ;
  assign n20119 = ~n20111 & n20118 ;
  assign n20120 = ~n20109 & n20119 ;
  assign n20121 = ~\a[23]  & ~n20120 ;
  assign n20122 = \a[23]  & n20119 ;
  assign n20123 = ~n20109 & n20122 ;
  assign n20124 = ~n20121 & ~n20123 ;
  assign n20125 = n20107 & ~n20124 ;
  assign n20126 = ~n20107 & n20124 ;
  assign n20127 = ~n20125 & ~n20126 ;
  assign n20128 = n1965 & n9930 ;
  assign n20129 = ~n9927 & n20128 ;
  assign n20130 = n1965 & ~n9930 ;
  assign n20131 = ~n9477 & n20130 ;
  assign n20132 = ~n9926 & n20131 ;
  assign n20133 = \b[40]  & n2218 ;
  assign n20134 = n2216 & n20133 ;
  assign n20135 = ~\a[18]  & \b[41]  ;
  assign n20136 = n1957 & n20135 ;
  assign n20137 = ~n20134 & ~n20136 ;
  assign n20138 = \b[42]  & n1963 ;
  assign n20139 = \a[18]  & \b[41]  ;
  assign n20140 = n2210 & n20139 ;
  assign n20141 = \a[20]  & ~n20140 ;
  assign n20142 = ~n20138 & n20141 ;
  assign n20143 = n20137 & n20142 ;
  assign n20144 = ~n20132 & n20143 ;
  assign n20145 = ~n20129 & n20144 ;
  assign n20146 = ~n20138 & ~n20140 ;
  assign n20147 = n20137 & n20146 ;
  assign n20148 = ~n20132 & n20147 ;
  assign n20149 = ~n20129 & n20148 ;
  assign n20150 = ~\a[20]  & ~n20149 ;
  assign n20151 = ~n20145 & ~n20150 ;
  assign n20152 = ~n20127 & n20151 ;
  assign n20153 = n19705 & n20152 ;
  assign n20154 = n20127 & n20151 ;
  assign n20155 = ~n19705 & n20154 ;
  assign n20156 = ~n20153 & ~n20155 ;
  assign n20157 = ~n20127 & ~n20151 ;
  assign n20158 = ~n19705 & n20157 ;
  assign n20159 = n20127 & ~n20151 ;
  assign n20160 = n19705 & n20159 ;
  assign n20161 = ~n20158 & ~n20160 ;
  assign n20162 = n20156 & n20161 ;
  assign n20163 = ~n19703 & ~n20162 ;
  assign n20164 = n19686 & n20163 ;
  assign n20165 = ~n19703 & n20162 ;
  assign n20166 = ~n19686 & n20165 ;
  assign n20167 = ~n20164 & ~n20166 ;
  assign n20168 = n19703 & ~n20162 ;
  assign n20169 = ~n19686 & n20168 ;
  assign n20170 = n19703 & n20162 ;
  assign n20171 = n19686 & n20170 ;
  assign n20172 = ~n20169 & ~n20171 ;
  assign n20173 = n20167 & n20172 ;
  assign n20174 = ~n19683 & n20173 ;
  assign n20175 = n999 & n12478 ;
  assign n20176 = ~n12475 & n20175 ;
  assign n20177 = n999 & ~n12478 ;
  assign n20178 = ~n12433 & n20177 ;
  assign n20179 = ~n12474 & n20178 ;
  assign n20180 = \b[46]  & n1182 ;
  assign n20181 = n1179 & n20180 ;
  assign n20182 = \b[48]  & n997 ;
  assign n20183 = \a[11]  & \b[47]  ;
  assign n20184 = n1180 & n20183 ;
  assign n20185 = ~\a[12]  & \b[47]  ;
  assign n20186 = n7674 & n20185 ;
  assign n20187 = ~n20184 & ~n20186 ;
  assign n20188 = ~n20182 & n20187 ;
  assign n20189 = ~n20181 & n20188 ;
  assign n20190 = ~n20179 & n20189 ;
  assign n20191 = ~n20176 & n20190 ;
  assign n20192 = ~\a[14]  & ~n20191 ;
  assign n20193 = \a[14]  & n20189 ;
  assign n20194 = ~n20179 & n20193 ;
  assign n20195 = ~n20176 & n20194 ;
  assign n20196 = ~n20192 & ~n20195 ;
  assign n20197 = ~n19480 & ~n20173 ;
  assign n20198 = ~n19682 & n20197 ;
  assign n20199 = ~n20196 & ~n20198 ;
  assign n20200 = ~n20174 & n20199 ;
  assign n20201 = ~n20173 & n20196 ;
  assign n20202 = n19683 & n20201 ;
  assign n20203 = n20173 & n20196 ;
  assign n20204 = ~n19683 & n20203 ;
  assign n20205 = ~n20202 & ~n20204 ;
  assign n20206 = ~n20200 & n20205 ;
  assign n20207 = ~n19681 & ~n20206 ;
  assign n20208 = n19664 & n20207 ;
  assign n20209 = ~n19681 & n20206 ;
  assign n20210 = ~n19664 & n20209 ;
  assign n20211 = ~n20208 & ~n20210 ;
  assign n20212 = n19681 & ~n20206 ;
  assign n20213 = ~n19664 & n20212 ;
  assign n20214 = n19681 & n20206 ;
  assign n20215 = n19664 & n20214 ;
  assign n20216 = ~n20213 & ~n20215 ;
  assign n20217 = n20211 & n20216 ;
  assign n20218 = ~n19661 & n20217 ;
  assign n20219 = n430 & ~n16398 ;
  assign n20220 = ~n15241 & n20219 ;
  assign n20221 = ~n16404 & n20220 ;
  assign n20222 = n430 & n16398 ;
  assign n20223 = n15241 & n20222 ;
  assign n20224 = n16400 & n20222 ;
  assign n20225 = ~n15239 & n20224 ;
  assign n20226 = ~n20223 & ~n20225 ;
  assign n20227 = ~n20221 & n20226 ;
  assign n20228 = \b[52]  & n486 ;
  assign n20229 = n483 & n20228 ;
  assign n20230 = ~\a[6]  & \b[53]  ;
  assign n20231 = n422 & n20230 ;
  assign n20232 = ~n20229 & ~n20231 ;
  assign n20233 = \b[54]  & n428 ;
  assign n20234 = \a[6]  & \b[53]  ;
  assign n20235 = n419 & n20234 ;
  assign n20236 = \a[8]  & ~n20235 ;
  assign n20237 = ~n20233 & n20236 ;
  assign n20238 = n20232 & n20237 ;
  assign n20239 = n20227 & n20238 ;
  assign n20240 = ~n20233 & ~n20235 ;
  assign n20241 = n20232 & n20240 ;
  assign n20242 = n20227 & n20241 ;
  assign n20243 = ~\a[8]  & ~n20242 ;
  assign n20244 = ~n20239 & ~n20243 ;
  assign n20245 = ~n19524 & ~n20217 ;
  assign n20246 = ~n19660 & n20245 ;
  assign n20247 = ~n20244 & ~n20246 ;
  assign n20248 = ~n20218 & n20247 ;
  assign n20249 = ~n20217 & n20244 ;
  assign n20250 = n19661 & n20249 ;
  assign n20251 = n20217 & n20244 ;
  assign n20252 = ~n19661 & n20251 ;
  assign n20253 = ~n20250 & ~n20252 ;
  assign n20254 = ~n20248 & n20253 ;
  assign n20255 = ~n18939 & ~n19546 ;
  assign n20256 = ~n19543 & n20255 ;
  assign n20257 = ~n19545 & ~n20256 ;
  assign n20258 = ~\b[59]  & ~\b[60]  ;
  assign n20259 = \b[59]  & \b[60]  ;
  assign n20260 = ~n20258 & ~n20259 ;
  assign n20261 = n134 & n20260 ;
  assign n20262 = ~n20257 & n20261 ;
  assign n20263 = n134 & ~n20260 ;
  assign n20264 = ~n19545 & n20263 ;
  assign n20265 = ~n20256 & n20264 ;
  assign n20266 = \a[0]  & \b[60]  ;
  assign n20267 = n133 & n20266 ;
  assign n20268 = \b[59]  & n141 ;
  assign n20269 = ~\a[1]  & \b[58]  ;
  assign n20270 = n10416 & n20269 ;
  assign n20271 = ~n20268 & ~n20270 ;
  assign n20272 = ~n20267 & n20271 ;
  assign n20273 = \a[2]  & n20272 ;
  assign n20274 = ~n20265 & n20273 ;
  assign n20275 = ~n20262 & n20274 ;
  assign n20276 = ~n20265 & n20272 ;
  assign n20277 = ~n20262 & n20276 ;
  assign n20278 = ~\a[2]  & ~n20277 ;
  assign n20279 = ~n20275 & ~n20278 ;
  assign n20280 = n252 & ~n17690 ;
  assign n20281 = ~n17688 & n20280 ;
  assign n20282 = \b[57]  & n250 ;
  assign n20283 = \a[3]  & \b[56]  ;
  assign n20284 = n241 & n20283 ;
  assign n20285 = ~n20282 & ~n20284 ;
  assign n20286 = \b[55]  & n303 ;
  assign n20287 = n300 & n20286 ;
  assign n20288 = ~\a[3]  & \b[56]  ;
  assign n20289 = n244 & n20288 ;
  assign n20290 = ~n20287 & ~n20289 ;
  assign n20291 = n20285 & n20290 ;
  assign n20292 = ~n20281 & n20291 ;
  assign n20293 = ~\a[5]  & ~n20292 ;
  assign n20294 = \a[5]  & n20291 ;
  assign n20295 = ~n20281 & n20294 ;
  assign n20296 = ~n20293 & ~n20295 ;
  assign n20297 = ~n20279 & ~n20296 ;
  assign n20298 = ~n20254 & n20297 ;
  assign n20299 = ~n19659 & n20298 ;
  assign n20300 = ~n20279 & n20296 ;
  assign n20301 = n20254 & n20300 ;
  assign n20302 = ~n19659 & n20301 ;
  assign n20303 = ~n20299 & ~n20302 ;
  assign n20304 = ~n20254 & n20300 ;
  assign n20305 = n19659 & n20304 ;
  assign n20306 = n20254 & n20297 ;
  assign n20307 = n19659 & n20306 ;
  assign n20308 = ~n20305 & ~n20307 ;
  assign n20309 = n20303 & n20308 ;
  assign n20310 = n20279 & n20296 ;
  assign n20311 = ~n20254 & n20310 ;
  assign n20312 = ~n19659 & n20311 ;
  assign n20313 = n20279 & ~n20296 ;
  assign n20314 = n20254 & n20313 ;
  assign n20315 = ~n19659 & n20314 ;
  assign n20316 = ~n20312 & ~n20315 ;
  assign n20317 = ~n20254 & n20313 ;
  assign n20318 = n19659 & n20317 ;
  assign n20319 = n20254 & n20310 ;
  assign n20320 = n19659 & n20319 ;
  assign n20321 = ~n20318 & ~n20320 ;
  assign n20322 = n20316 & n20321 ;
  assign n20323 = n19564 & ~n19639 ;
  assign n20324 = n19644 & ~n20323 ;
  assign n20325 = n20322 & n20324 ;
  assign n20326 = n20309 & n20325 ;
  assign n20327 = n20309 & n20322 ;
  assign n20328 = ~n20324 & ~n20327 ;
  assign n20329 = ~n20326 & ~n20328 ;
  assign n20330 = n19656 & n20329 ;
  assign n20331 = ~n19656 & ~n20329 ;
  assign n20332 = ~n20330 & ~n20331 ;
  assign n20333 = ~n20254 & n20296 ;
  assign n20334 = ~n19659 & n20333 ;
  assign n20335 = n20254 & n20296 ;
  assign n20336 = n19659 & n20335 ;
  assign n20337 = ~n20334 & ~n20336 ;
  assign n20338 = ~n20254 & ~n20296 ;
  assign n20339 = n19659 & n20338 ;
  assign n20340 = n20254 & ~n20296 ;
  assign n20341 = ~n19659 & n20340 ;
  assign n20342 = ~n20339 & ~n20341 ;
  assign n20343 = n20279 & n20342 ;
  assign n20344 = n20337 & ~n20343 ;
  assign n20345 = n19659 & n20254 ;
  assign n20346 = ~n20248 & ~n20345 ;
  assign n20347 = ~n19524 & n20211 ;
  assign n20348 = ~n19660 & n20347 ;
  assign n20349 = n20216 & ~n20348 ;
  assign n20350 = n19664 & n20206 ;
  assign n20351 = ~n20200 & ~n20350 ;
  assign n20352 = ~n551 & ~n14093 ;
  assign n20353 = ~n15201 & n20352 ;
  assign n20354 = ~n15197 & n20353 ;
  assign n20355 = ~n643 & n20354 ;
  assign n20356 = n646 & n15201 ;
  assign n20357 = ~n15198 & n20356 ;
  assign n20358 = ~n20355 & ~n20357 ;
  assign n20359 = \b[50]  & n796 ;
  assign n20360 = n793 & n20359 ;
  assign n20361 = \b[52]  & n644 ;
  assign n20362 = \a[8]  & \b[51]  ;
  assign n20363 = n794 & n20362 ;
  assign n20364 = ~\a[9]  & \b[51]  ;
  assign n20365 = n638 & n20364 ;
  assign n20366 = ~n20363 & ~n20365 ;
  assign n20367 = ~n20361 & n20366 ;
  assign n20368 = ~n20360 & n20367 ;
  assign n20369 = n20358 & n20368 ;
  assign n20370 = ~\a[11]  & ~n20369 ;
  assign n20371 = \a[11]  & n20368 ;
  assign n20372 = n20358 & n20371 ;
  assign n20373 = ~n20370 & ~n20372 ;
  assign n20374 = ~n19480 & n20167 ;
  assign n20375 = ~n19682 & n20374 ;
  assign n20376 = n20172 & ~n20375 ;
  assign n20377 = n999 & ~n13524 ;
  assign n20378 = ~n13522 & n20377 ;
  assign n20379 = \b[47]  & n1182 ;
  assign n20380 = n1179 & n20379 ;
  assign n20381 = \b[49]  & n997 ;
  assign n20382 = \a[11]  & \b[48]  ;
  assign n20383 = n1180 & n20382 ;
  assign n20384 = ~\a[12]  & \b[48]  ;
  assign n20385 = n7674 & n20384 ;
  assign n20386 = ~n20383 & ~n20385 ;
  assign n20387 = ~n20381 & n20386 ;
  assign n20388 = ~n20380 & n20387 ;
  assign n20389 = ~n20378 & n20388 ;
  assign n20390 = ~\a[14]  & ~n20389 ;
  assign n20391 = \a[14]  & n20388 ;
  assign n20392 = ~n20378 & n20391 ;
  assign n20393 = ~n20390 & ~n20392 ;
  assign n20394 = n19686 & n20162 ;
  assign n20395 = n20161 & ~n20394 ;
  assign n20396 = n1467 & n11906 ;
  assign n20397 = ~n11903 & n20396 ;
  assign n20398 = n1467 & ~n11906 ;
  assign n20399 = ~n11392 & n20398 ;
  assign n20400 = ~n11902 & n20399 ;
  assign n20401 = \b[44]  & n1652 ;
  assign n20402 = n1649 & n20401 ;
  assign n20403 = ~\a[15]  & \b[45]  ;
  assign n20404 = n1459 & n20403 ;
  assign n20405 = ~n20402 & ~n20404 ;
  assign n20406 = \b[46]  & n1465 ;
  assign n20407 = \a[15]  & \b[45]  ;
  assign n20408 = n1456 & n20407 ;
  assign n20409 = \a[17]  & ~n20408 ;
  assign n20410 = ~n20406 & n20409 ;
  assign n20411 = n20405 & n20410 ;
  assign n20412 = ~n20400 & n20411 ;
  assign n20413 = ~n20397 & n20412 ;
  assign n20414 = ~n20406 & ~n20408 ;
  assign n20415 = n20405 & n20414 ;
  assign n20416 = ~n20400 & n20415 ;
  assign n20417 = ~n20397 & n20416 ;
  assign n20418 = ~\a[17]  & ~n20417 ;
  assign n20419 = ~n20413 & ~n20418 ;
  assign n20420 = n19422 & ~n20125 ;
  assign n20421 = ~n19704 & n20420 ;
  assign n20422 = ~n20126 & ~n20421 ;
  assign n20423 = ~n20098 & ~n20106 ;
  assign n20424 = ~n19366 & n20065 ;
  assign n20425 = ~n19709 & n20424 ;
  assign n20426 = n20070 & ~n20425 ;
  assign n20427 = n19713 & n20043 ;
  assign n20428 = n20042 & ~n20427 ;
  assign n20429 = n19320 & ~n20007 ;
  assign n20430 = ~n19714 & n20429 ;
  assign n20431 = ~n20008 & ~n20430 ;
  assign n20432 = ~n19978 & ~n19986 ;
  assign n20433 = ~n19273 & n19943 ;
  assign n20434 = ~n19719 & n20433 ;
  assign n20435 = n19948 & ~n20434 ;
  assign n20436 = ~n19725 & n19938 ;
  assign n20437 = n19932 & ~n20436 ;
  assign n20438 = n2768 & n8759 ;
  assign n20439 = ~n2765 & n20438 ;
  assign n20440 = ~n2768 & n8759 ;
  assign n20441 = ~n2518 & n20440 ;
  assign n20442 = ~n2764 & n20441 ;
  assign n20443 = \b[20]  & n9301 ;
  assign n20444 = n9298 & n20443 ;
  assign n20445 = ~\a[39]  & \b[21]  ;
  assign n20446 = n8751 & n20445 ;
  assign n20447 = ~n20444 & ~n20446 ;
  assign n20448 = \b[22]  & n8757 ;
  assign n20449 = \a[39]  & \b[21]  ;
  assign n20450 = n8748 & n20449 ;
  assign n20451 = \a[41]  & ~n20450 ;
  assign n20452 = ~n20448 & n20451 ;
  assign n20453 = n20447 & n20452 ;
  assign n20454 = ~n20442 & n20453 ;
  assign n20455 = ~n20439 & n20454 ;
  assign n20456 = ~n20448 & ~n20450 ;
  assign n20457 = n20447 & n20456 ;
  assign n20458 = ~n20442 & n20457 ;
  assign n20459 = ~n20439 & n20458 ;
  assign n20460 = ~\a[41]  & ~n20459 ;
  assign n20461 = ~n20455 & ~n20460 ;
  assign n20462 = n19232 & n19921 ;
  assign n20463 = ~n19239 & n20462 ;
  assign n20464 = n19926 & ~n20463 ;
  assign n20465 = n19775 & n19916 ;
  assign n20466 = ~n19915 & ~n20465 ;
  assign n20467 = ~n19198 & n19899 ;
  assign n20468 = ~n19200 & n20467 ;
  assign n20469 = n19904 & ~n20468 ;
  assign n20470 = n19820 & n19894 ;
  assign n20471 = ~n19892 & ~n20470 ;
  assign n20472 = ~n383 & n16655 ;
  assign n20473 = ~n381 & n20472 ;
  assign n20474 = \b[5]  & n17308 ;
  assign n20475 = n17305 & n20474 ;
  assign n20476 = \b[7]  & n16653 ;
  assign n20477 = \a[53]  & \b[6]  ;
  assign n20478 = n17306 & n20477 ;
  assign n20479 = ~\a[54]  & \b[6]  ;
  assign n20480 = n16647 & n20479 ;
  assign n20481 = ~n20478 & ~n20480 ;
  assign n20482 = ~n20476 & n20481 ;
  assign n20483 = ~n20475 & n20482 ;
  assign n20484 = ~\a[56]  & n20483 ;
  assign n20485 = ~n20473 & n20484 ;
  assign n20486 = ~n20473 & n20483 ;
  assign n20487 = \a[56]  & ~n20486 ;
  assign n20488 = ~n20485 & ~n20487 ;
  assign n20489 = ~n19864 & ~n19867 ;
  assign n20490 = n222 & n18516 ;
  assign n20491 = \b[4]  & n18514 ;
  assign n20492 = \a[56]  & \b[3]  ;
  assign n20493 = n19181 & n20492 ;
  assign n20494 = ~\a[57]  & \b[3]  ;
  assign n20495 = n18508 & n20494 ;
  assign n20496 = ~n20493 & ~n20495 ;
  assign n20497 = ~n20491 & n20496 ;
  assign n20498 = \b[2]  & n19183 ;
  assign n20499 = n19180 & n20498 ;
  assign n20500 = \a[59]  & ~n20499 ;
  assign n20501 = n20497 & n20500 ;
  assign n20502 = ~n20490 & n20501 ;
  assign n20503 = n20497 & ~n20499 ;
  assign n20504 = ~n20490 & n20503 ;
  assign n20505 = ~\a[59]  & ~n20504 ;
  assign n20506 = ~n20502 & ~n20505 ;
  assign n20507 = \a[62]  & \b[0]  ;
  assign n20508 = ~n19861 & n20507 ;
  assign n20509 = \a[60]  & \b[0]  ;
  assign n20510 = \a[59]  & ~\a[61]  ;
  assign n20511 = n20509 & n20510 ;
  assign n20512 = ~\a[60]  & \b[0]  ;
  assign n20513 = ~\a[59]  & \a[61]  ;
  assign n20514 = n20512 & n20513 ;
  assign n20515 = ~n20511 & ~n20514 ;
  assign n20516 = \a[61]  & ~\a[62]  ;
  assign n20517 = ~\a[61]  & \a[62]  ;
  assign n20518 = ~n20516 & ~n20517 ;
  assign n20519 = ~n19861 & n20518 ;
  assign n20520 = \b[1]  & n20519 ;
  assign n20521 = ~n19861 & ~n20518 ;
  assign n20522 = ~n137 & n20521 ;
  assign n20523 = ~n20520 & ~n20522 ;
  assign n20524 = n20515 & n20523 ;
  assign n20525 = n20508 & ~n20524 ;
  assign n20526 = ~n20508 & n20515 ;
  assign n20527 = n20523 & n20526 ;
  assign n20528 = ~n20525 & ~n20527 ;
  assign n20529 = n20506 & ~n20528 ;
  assign n20530 = ~n20506 & n20528 ;
  assign n20531 = ~n20529 & ~n20530 ;
  assign n20532 = ~n20489 & n20531 ;
  assign n20533 = n20489 & ~n20531 ;
  assign n20534 = ~n20532 & ~n20533 ;
  assign n20535 = ~n20488 & ~n20534 ;
  assign n20536 = n20488 & n20534 ;
  assign n20537 = ~n20535 & ~n20536 ;
  assign n20538 = ~n685 & ~n14276 ;
  assign n20539 = ~n14790 & n20538 ;
  assign n20540 = n682 & n20539 ;
  assign n20541 = n685 & ~n14276 ;
  assign n20542 = ~n14790 & n20541 ;
  assign n20543 = ~n682 & n20542 ;
  assign n20544 = ~n20540 & ~n20543 ;
  assign n20545 = \b[8]  & n15517 ;
  assign n20546 = n15514 & n20545 ;
  assign n20547 = ~\a[51]  & \b[9]  ;
  assign n20548 = n14785 & n20547 ;
  assign n20549 = ~n20546 & ~n20548 ;
  assign n20550 = \b[10]  & n14791 ;
  assign n20551 = \a[51]  & \b[9]  ;
  assign n20552 = n14782 & n20551 ;
  assign n20553 = \a[53]  & ~n20552 ;
  assign n20554 = ~n20550 & n20553 ;
  assign n20555 = n20549 & n20554 ;
  assign n20556 = n20544 & n20555 ;
  assign n20557 = ~n20550 & ~n20552 ;
  assign n20558 = n20549 & n20557 ;
  assign n20559 = n20544 & n20558 ;
  assign n20560 = ~\a[53]  & ~n20559 ;
  assign n20561 = ~n20556 & ~n20560 ;
  assign n20562 = ~n20537 & ~n20561 ;
  assign n20563 = ~n20471 & n20562 ;
  assign n20564 = n20537 & ~n20561 ;
  assign n20565 = n20471 & n20564 ;
  assign n20566 = ~n20563 & ~n20565 ;
  assign n20567 = ~n20537 & n20561 ;
  assign n20568 = n20471 & n20567 ;
  assign n20569 = n20537 & n20561 ;
  assign n20570 = ~n20471 & n20569 ;
  assign n20571 = ~n20568 & ~n20570 ;
  assign n20572 = n20566 & n20571 ;
  assign n20573 = ~n948 & n13125 ;
  assign n20574 = ~n908 & n13125 ;
  assign n20575 = ~n912 & n20574 ;
  assign n20576 = ~n20573 & ~n20575 ;
  assign n20577 = ~n951 & ~n20576 ;
  assign n20578 = \b[11]  & n13794 ;
  assign n20579 = n13792 & n20578 ;
  assign n20580 = ~\a[48]  & \b[12]  ;
  assign n20581 = n13117 & n20580 ;
  assign n20582 = ~n20579 & ~n20581 ;
  assign n20583 = \b[13]  & n13123 ;
  assign n20584 = \a[48]  & \b[12]  ;
  assign n20585 = n13786 & n20584 ;
  assign n20586 = \a[50]  & ~n20585 ;
  assign n20587 = ~n20583 & n20586 ;
  assign n20588 = n20582 & n20587 ;
  assign n20589 = ~n20577 & n20588 ;
  assign n20590 = ~n20583 & ~n20585 ;
  assign n20591 = n20582 & n20590 ;
  assign n20592 = ~\a[50]  & ~n20591 ;
  assign n20593 = ~\a[50]  & ~n951 ;
  assign n20594 = ~n20576 & n20593 ;
  assign n20595 = ~n20592 & ~n20594 ;
  assign n20596 = ~n20589 & n20595 ;
  assign n20597 = ~n20572 & ~n20596 ;
  assign n20598 = n20469 & n20597 ;
  assign n20599 = n20572 & ~n20596 ;
  assign n20600 = ~n20469 & n20599 ;
  assign n20601 = ~n20598 & ~n20600 ;
  assign n20602 = ~n20572 & n20596 ;
  assign n20603 = ~n20469 & n20602 ;
  assign n20604 = n20572 & n20596 ;
  assign n20605 = n20469 & n20604 ;
  assign n20606 = ~n20603 & ~n20605 ;
  assign n20607 = n20601 & n20606 ;
  assign n20608 = ~n20466 & n20607 ;
  assign n20609 = n1512 & n11572 ;
  assign n20610 = ~n1509 & n20609 ;
  assign n20611 = ~n1512 & n11572 ;
  assign n20612 = ~n1228 & n20611 ;
  assign n20613 = ~n1508 & n20612 ;
  assign n20614 = \b[14]  & n12159 ;
  assign n20615 = n12156 & n20614 ;
  assign n20616 = \b[16]  & n11570 ;
  assign n20617 = \a[44]  & \b[15]  ;
  assign n20618 = n12157 & n20617 ;
  assign n20619 = ~\a[45]  & \b[15]  ;
  assign n20620 = n11564 & n20619 ;
  assign n20621 = ~n20618 & ~n20620 ;
  assign n20622 = ~n20616 & n20621 ;
  assign n20623 = ~n20615 & n20622 ;
  assign n20624 = ~n20613 & n20623 ;
  assign n20625 = ~n20610 & n20624 ;
  assign n20626 = ~\a[47]  & ~n20625 ;
  assign n20627 = \a[47]  & n20623 ;
  assign n20628 = ~n20613 & n20627 ;
  assign n20629 = ~n20610 & n20628 ;
  assign n20630 = ~n20626 & ~n20629 ;
  assign n20631 = ~n19915 & ~n20607 ;
  assign n20632 = ~n20465 & n20631 ;
  assign n20633 = ~n20630 & ~n20632 ;
  assign n20634 = ~n20608 & n20633 ;
  assign n20635 = ~n20607 & n20630 ;
  assign n20636 = n20466 & n20635 ;
  assign n20637 = n20607 & n20630 ;
  assign n20638 = ~n20466 & n20637 ;
  assign n20639 = ~n20636 & ~n20638 ;
  assign n20640 = ~n20634 & n20639 ;
  assign n20641 = ~n20464 & ~n20640 ;
  assign n20642 = n20464 & n20640 ;
  assign n20643 = ~n20641 & ~n20642 ;
  assign n20644 = ~n2079 & n10082 ;
  assign n20645 = ~n2077 & n20644 ;
  assign n20646 = \b[17]  & n10681 ;
  assign n20647 = n10678 & n20646 ;
  assign n20648 = \b[19]  & n10080 ;
  assign n20649 = \a[41]  & \b[18]  ;
  assign n20650 = n10679 & n20649 ;
  assign n20651 = ~\a[42]  & \b[18]  ;
  assign n20652 = n10074 & n20651 ;
  assign n20653 = ~n20650 & ~n20652 ;
  assign n20654 = ~n20648 & n20653 ;
  assign n20655 = ~n20647 & n20654 ;
  assign n20656 = ~n20645 & n20655 ;
  assign n20657 = ~\a[44]  & ~n20656 ;
  assign n20658 = \a[44]  & n20655 ;
  assign n20659 = ~n20645 & n20658 ;
  assign n20660 = ~n20657 & ~n20659 ;
  assign n20661 = n20643 & ~n20660 ;
  assign n20662 = ~n20643 & n20660 ;
  assign n20663 = ~n20661 & ~n20662 ;
  assign n20664 = ~n20461 & ~n20663 ;
  assign n20665 = ~n20437 & n20664 ;
  assign n20666 = ~n20461 & n20663 ;
  assign n20667 = n20437 & n20666 ;
  assign n20668 = ~n20665 & ~n20667 ;
  assign n20669 = n20461 & ~n20663 ;
  assign n20670 = n20437 & n20669 ;
  assign n20671 = n20461 & n20663 ;
  assign n20672 = ~n20437 & n20671 ;
  assign n20673 = ~n20670 & ~n20672 ;
  assign n20674 = n20668 & n20673 ;
  assign n20675 = ~n20435 & ~n20674 ;
  assign n20676 = n19948 & n20674 ;
  assign n20677 = ~n20434 & n20676 ;
  assign n20678 = ~n3564 & n7534 ;
  assign n20679 = ~n3282 & n7534 ;
  assign n20680 = ~n3560 & n20679 ;
  assign n20681 = ~n20678 & ~n20680 ;
  assign n20682 = ~n3567 & ~n20681 ;
  assign n20683 = \b[23]  & n7973 ;
  assign n20684 = n7970 & n20683 ;
  assign n20685 = ~\a[36]  & \b[24]  ;
  assign n20686 = n7526 & n20685 ;
  assign n20687 = ~n20684 & ~n20686 ;
  assign n20688 = \b[25]  & n7532 ;
  assign n20689 = \a[36]  & \b[24]  ;
  assign n20690 = n17801 & n20689 ;
  assign n20691 = \a[38]  & ~n20690 ;
  assign n20692 = ~n20688 & n20691 ;
  assign n20693 = n20687 & n20692 ;
  assign n20694 = ~n20682 & n20693 ;
  assign n20695 = ~n20688 & ~n20690 ;
  assign n20696 = n20687 & n20695 ;
  assign n20697 = ~\a[38]  & ~n20696 ;
  assign n20698 = ~\a[38]  & ~n3567 ;
  assign n20699 = ~n20681 & n20698 ;
  assign n20700 = ~n20697 & ~n20699 ;
  assign n20701 = ~n20694 & n20700 ;
  assign n20702 = ~n20677 & ~n20701 ;
  assign n20703 = ~n20675 & n20702 ;
  assign n20704 = ~n20674 & n20701 ;
  assign n20705 = ~n20435 & n20704 ;
  assign n20706 = n20674 & n20701 ;
  assign n20707 = n20435 & n20706 ;
  assign n20708 = ~n20705 & ~n20707 ;
  assign n20709 = ~n20703 & n20708 ;
  assign n20710 = n4456 & n6309 ;
  assign n20711 = ~n18723 & n20710 ;
  assign n20712 = ~n4456 & n6309 ;
  assign n20713 = ~n4143 & n20712 ;
  assign n20714 = ~n4452 & n20713 ;
  assign n20715 = \b[26]  & n6778 ;
  assign n20716 = n6775 & n20715 ;
  assign n20717 = ~\a[33]  & \b[27]  ;
  assign n20718 = n6301 & n20717 ;
  assign n20719 = ~n20716 & ~n20718 ;
  assign n20720 = \b[28]  & n6307 ;
  assign n20721 = \a[33]  & \b[27]  ;
  assign n20722 = n6298 & n20721 ;
  assign n20723 = \a[35]  & ~n20722 ;
  assign n20724 = ~n20720 & n20723 ;
  assign n20725 = n20719 & n20724 ;
  assign n20726 = ~n20714 & n20725 ;
  assign n20727 = ~n20711 & n20726 ;
  assign n20728 = ~n20720 & ~n20722 ;
  assign n20729 = n20719 & n20728 ;
  assign n20730 = ~n20714 & n20729 ;
  assign n20731 = ~n20711 & n20730 ;
  assign n20732 = ~\a[35]  & ~n20731 ;
  assign n20733 = ~n20727 & ~n20732 ;
  assign n20734 = ~n20709 & ~n20733 ;
  assign n20735 = ~n20432 & n20734 ;
  assign n20736 = n20709 & ~n20733 ;
  assign n20737 = n20432 & n20736 ;
  assign n20738 = ~n20735 & ~n20737 ;
  assign n20739 = ~n20709 & n20733 ;
  assign n20740 = n20432 & n20739 ;
  assign n20741 = n20709 & n20733 ;
  assign n20742 = ~n20432 & n20741 ;
  assign n20743 = ~n20740 & ~n20742 ;
  assign n20744 = n20738 & n20743 ;
  assign n20745 = n5211 & ~n5462 ;
  assign n20746 = ~n5460 & n20745 ;
  assign n20747 = \b[29]  & n5595 ;
  assign n20748 = n5592 & n20747 ;
  assign n20749 = ~\a[30]  & \b[30]  ;
  assign n20750 = n5203 & n20749 ;
  assign n20751 = ~n20748 & ~n20750 ;
  assign n20752 = \b[31]  & n5209 ;
  assign n20753 = \a[30]  & \b[30]  ;
  assign n20754 = n5200 & n20753 ;
  assign n20755 = \a[32]  & ~n20754 ;
  assign n20756 = ~n20752 & n20755 ;
  assign n20757 = n20751 & n20756 ;
  assign n20758 = ~n20746 & n20757 ;
  assign n20759 = ~n20752 & ~n20754 ;
  assign n20760 = n20751 & n20759 ;
  assign n20761 = ~n20746 & n20760 ;
  assign n20762 = ~\a[32]  & ~n20761 ;
  assign n20763 = ~n20758 & ~n20762 ;
  assign n20764 = ~n20744 & ~n20763 ;
  assign n20765 = n20431 & n20764 ;
  assign n20766 = n20744 & ~n20763 ;
  assign n20767 = ~n20431 & n20766 ;
  assign n20768 = ~n20765 & ~n20767 ;
  assign n20769 = ~n20744 & n20763 ;
  assign n20770 = ~n20431 & n20769 ;
  assign n20771 = n20744 & n20763 ;
  assign n20772 = n20431 & n20771 ;
  assign n20773 = ~n20770 & ~n20772 ;
  assign n20774 = n20768 & n20773 ;
  assign n20775 = ~n20428 & n20774 ;
  assign n20776 = n4249 & n6565 ;
  assign n20777 = ~n6562 & n20776 ;
  assign n20778 = n4249 & ~n6565 ;
  assign n20779 = ~n5850 & n20778 ;
  assign n20780 = ~n6561 & n20779 ;
  assign n20781 = \b[32]  & n4647 ;
  assign n20782 = n4644 & n20781 ;
  assign n20783 = ~\a[27]  & \b[33]  ;
  assign n20784 = n4241 & n20783 ;
  assign n20785 = ~n20782 & ~n20784 ;
  assign n20786 = \b[34]  & n4247 ;
  assign n20787 = \a[27]  & \b[33]  ;
  assign n20788 = n4238 & n20787 ;
  assign n20789 = \a[29]  & ~n20788 ;
  assign n20790 = ~n20786 & n20789 ;
  assign n20791 = n20785 & n20790 ;
  assign n20792 = ~n20780 & n20791 ;
  assign n20793 = ~n20777 & n20792 ;
  assign n20794 = ~n20786 & ~n20788 ;
  assign n20795 = n20785 & n20794 ;
  assign n20796 = ~n20780 & n20795 ;
  assign n20797 = ~n20777 & n20796 ;
  assign n20798 = ~\a[29]  & ~n20797 ;
  assign n20799 = ~n20793 & ~n20798 ;
  assign n20800 = n20042 & ~n20774 ;
  assign n20801 = ~n20427 & n20800 ;
  assign n20802 = ~n20799 & ~n20801 ;
  assign n20803 = ~n20775 & n20802 ;
  assign n20804 = ~n20774 & n20799 ;
  assign n20805 = n20428 & n20804 ;
  assign n20806 = n20774 & n20799 ;
  assign n20807 = ~n20428 & n20806 ;
  assign n20808 = ~n20805 & ~n20807 ;
  assign n20809 = ~n20803 & n20808 ;
  assign n20810 = n3402 & ~n7761 ;
  assign n20811 = ~n7759 & n20810 ;
  assign n20812 = \b[35]  & n3733 ;
  assign n20813 = n3730 & n20812 ;
  assign n20814 = \b[37]  & n3400 ;
  assign n20815 = \a[23]  & \b[36]  ;
  assign n20816 = n3731 & n20815 ;
  assign n20817 = ~\a[24]  & \b[36]  ;
  assign n20818 = n3394 & n20817 ;
  assign n20819 = ~n20816 & ~n20818 ;
  assign n20820 = ~n20814 & n20819 ;
  assign n20821 = ~n20813 & n20820 ;
  assign n20822 = ~n20811 & n20821 ;
  assign n20823 = ~\a[26]  & ~n20822 ;
  assign n20824 = \a[26]  & n20821 ;
  assign n20825 = ~n20811 & n20824 ;
  assign n20826 = ~n20823 & ~n20825 ;
  assign n20827 = ~n20809 & ~n20826 ;
  assign n20828 = n20426 & n20827 ;
  assign n20829 = n20809 & ~n20826 ;
  assign n20830 = ~n20426 & n20829 ;
  assign n20831 = ~n20828 & ~n20830 ;
  assign n20832 = ~n20809 & n20826 ;
  assign n20833 = ~n20426 & n20832 ;
  assign n20834 = n20809 & n20826 ;
  assign n20835 = n20426 & n20834 ;
  assign n20836 = ~n20833 & ~n20835 ;
  assign n20837 = n20831 & n20836 ;
  assign n20838 = n2622 & n9044 ;
  assign n20839 = ~n9041 & n20838 ;
  assign n20840 = n2622 & ~n9044 ;
  assign n20841 = ~n8597 & n20840 ;
  assign n20842 = ~n9040 & n20841 ;
  assign n20843 = \b[38]  & n2912 ;
  assign n20844 = n2909 & n20843 ;
  assign n20845 = ~\a[21]  & \b[39]  ;
  assign n20846 = n2614 & n20845 ;
  assign n20847 = ~n20844 & ~n20846 ;
  assign n20848 = \b[40]  & n2620 ;
  assign n20849 = \a[20]  & ~\a[22]  ;
  assign n20850 = \a[21]  & \b[39]  ;
  assign n20851 = n20849 & n20850 ;
  assign n20852 = \a[23]  & ~n20851 ;
  assign n20853 = ~n20848 & n20852 ;
  assign n20854 = n20847 & n20853 ;
  assign n20855 = ~n20842 & n20854 ;
  assign n20856 = ~n20839 & n20855 ;
  assign n20857 = ~n20848 & ~n20851 ;
  assign n20858 = n20847 & n20857 ;
  assign n20859 = ~n20842 & n20858 ;
  assign n20860 = ~n20839 & n20859 ;
  assign n20861 = ~\a[23]  & ~n20860 ;
  assign n20862 = ~n20856 & ~n20861 ;
  assign n20863 = ~n20837 & ~n20862 ;
  assign n20864 = ~n20423 & n20863 ;
  assign n20865 = n20837 & ~n20862 ;
  assign n20866 = n20423 & n20865 ;
  assign n20867 = ~n20864 & ~n20866 ;
  assign n20868 = ~n20837 & n20862 ;
  assign n20869 = n20423 & n20868 ;
  assign n20870 = n20837 & n20862 ;
  assign n20871 = ~n20423 & n20870 ;
  assign n20872 = ~n20869 & ~n20871 ;
  assign n20873 = n20867 & n20872 ;
  assign n20874 = n1965 & ~n10409 ;
  assign n20875 = ~n10407 & n20874 ;
  assign n20876 = \b[43]  & n1963 ;
  assign n20877 = \a[18]  & \b[42]  ;
  assign n20878 = n2210 & n20877 ;
  assign n20879 = ~n20876 & ~n20878 ;
  assign n20880 = \b[41]  & n2218 ;
  assign n20881 = n2216 & n20880 ;
  assign n20882 = ~\a[18]  & \b[42]  ;
  assign n20883 = n1957 & n20882 ;
  assign n20884 = ~n20881 & ~n20883 ;
  assign n20885 = n20879 & n20884 ;
  assign n20886 = ~n20875 & n20885 ;
  assign n20887 = ~\a[20]  & ~n20886 ;
  assign n20888 = \a[20]  & n20885 ;
  assign n20889 = ~n20875 & n20888 ;
  assign n20890 = ~n20887 & ~n20889 ;
  assign n20891 = ~n20873 & ~n20890 ;
  assign n20892 = n20422 & n20891 ;
  assign n20893 = n20873 & ~n20890 ;
  assign n20894 = ~n20422 & n20893 ;
  assign n20895 = ~n20892 & ~n20894 ;
  assign n20896 = ~n20873 & n20890 ;
  assign n20897 = ~n20422 & n20896 ;
  assign n20898 = n20873 & n20890 ;
  assign n20899 = n20422 & n20898 ;
  assign n20900 = ~n20897 & ~n20899 ;
  assign n20901 = n20895 & n20900 ;
  assign n20902 = n20419 & ~n20901 ;
  assign n20903 = n20395 & n20902 ;
  assign n20904 = n20419 & n20901 ;
  assign n20905 = ~n20395 & n20904 ;
  assign n20906 = ~n20903 & ~n20905 ;
  assign n20907 = ~n20395 & n20901 ;
  assign n20908 = n20161 & ~n20901 ;
  assign n20909 = ~n20394 & n20908 ;
  assign n20910 = ~n20419 & ~n20909 ;
  assign n20911 = ~n20907 & n20910 ;
  assign n20912 = n20906 & ~n20911 ;
  assign n20913 = n20393 & ~n20912 ;
  assign n20914 = ~n20376 & n20913 ;
  assign n20915 = n20393 & n20912 ;
  assign n20916 = n20376 & n20915 ;
  assign n20917 = ~n20914 & ~n20916 ;
  assign n20918 = ~n20393 & ~n20912 ;
  assign n20919 = n20376 & n20918 ;
  assign n20920 = ~n20393 & n20912 ;
  assign n20921 = ~n20376 & n20920 ;
  assign n20922 = ~n20919 & ~n20921 ;
  assign n20923 = n20917 & n20922 ;
  assign n20924 = n20373 & ~n20923 ;
  assign n20925 = n20351 & n20924 ;
  assign n20926 = n20373 & n20923 ;
  assign n20927 = ~n20351 & n20926 ;
  assign n20928 = ~n20925 & ~n20927 ;
  assign n20929 = ~n20351 & n20923 ;
  assign n20930 = ~n20200 & ~n20923 ;
  assign n20931 = ~n20350 & n20930 ;
  assign n20932 = ~n20373 & ~n20931 ;
  assign n20933 = ~n20929 & n20932 ;
  assign n20934 = n20928 & ~n20933 ;
  assign n20935 = n430 & ~n16446 ;
  assign n20936 = ~n16444 & n20935 ;
  assign n20937 = \b[55]  & n428 ;
  assign n20938 = \a[6]  & \b[54]  ;
  assign n20939 = n419 & n20938 ;
  assign n20940 = ~n20937 & ~n20939 ;
  assign n20941 = \b[53]  & n486 ;
  assign n20942 = n483 & n20941 ;
  assign n20943 = ~\a[6]  & \b[54]  ;
  assign n20944 = n422 & n20943 ;
  assign n20945 = ~n20942 & ~n20944 ;
  assign n20946 = n20940 & n20945 ;
  assign n20947 = ~n20936 & n20946 ;
  assign n20948 = ~\a[8]  & ~n20947 ;
  assign n20949 = \a[8]  & n20946 ;
  assign n20950 = ~n20936 & n20949 ;
  assign n20951 = ~n20948 & ~n20950 ;
  assign n20952 = ~n20934 & ~n20951 ;
  assign n20953 = n20349 & n20952 ;
  assign n20954 = n20934 & ~n20951 ;
  assign n20955 = ~n20349 & n20954 ;
  assign n20956 = ~n20953 & ~n20955 ;
  assign n20957 = ~n20934 & n20951 ;
  assign n20958 = ~n20349 & n20957 ;
  assign n20959 = n20934 & n20951 ;
  assign n20960 = n20349 & n20959 ;
  assign n20961 = ~n20958 & ~n20960 ;
  assign n20962 = n20956 & n20961 ;
  assign n20963 = ~n19545 & n20260 ;
  assign n20964 = ~n20256 & n20963 ;
  assign n20965 = ~n20259 & ~n20964 ;
  assign n20966 = ~\b[60]  & ~\b[61]  ;
  assign n20967 = \b[60]  & \b[61]  ;
  assign n20968 = ~n20966 & ~n20967 ;
  assign n20969 = ~n20965 & n20968 ;
  assign n20970 = ~n20259 & ~n20968 ;
  assign n20971 = ~n20964 & n20970 ;
  assign n20972 = n134 & ~n20971 ;
  assign n20973 = ~n20969 & n20972 ;
  assign n20974 = \a[0]  & \b[61]  ;
  assign n20975 = n133 & n20974 ;
  assign n20976 = \b[60]  & n141 ;
  assign n20977 = ~\a[1]  & \b[59]  ;
  assign n20978 = n10416 & n20977 ;
  assign n20979 = ~n20976 & ~n20978 ;
  assign n20980 = ~n20975 & n20979 ;
  assign n20981 = \a[2]  & n20980 ;
  assign n20982 = ~n20973 & n20981 ;
  assign n20983 = ~n20973 & n20980 ;
  assign n20984 = ~\a[2]  & ~n20983 ;
  assign n20985 = ~n20982 & ~n20984 ;
  assign n20986 = n252 & n18940 ;
  assign n20987 = ~n18937 & n20986 ;
  assign n20988 = ~n17685 & ~n18940 ;
  assign n20989 = n252 & n20988 ;
  assign n20990 = ~n18936 & n20989 ;
  assign n20991 = \b[56]  & n303 ;
  assign n20992 = n300 & n20991 ;
  assign n20993 = \b[58]  & n250 ;
  assign n20994 = \a[3]  & \b[57]  ;
  assign n20995 = n241 & n20994 ;
  assign n20996 = ~\a[3]  & \b[57]  ;
  assign n20997 = n244 & n20996 ;
  assign n20998 = ~n20995 & ~n20997 ;
  assign n20999 = ~n20993 & n20998 ;
  assign n21000 = ~n20992 & n20999 ;
  assign n21001 = ~n20990 & n21000 ;
  assign n21002 = ~n20987 & n21001 ;
  assign n21003 = ~\a[5]  & ~n21002 ;
  assign n21004 = \a[5]  & n21000 ;
  assign n21005 = ~n20990 & n21004 ;
  assign n21006 = ~n20987 & n21005 ;
  assign n21007 = ~n21003 & ~n21006 ;
  assign n21008 = ~n20985 & ~n21007 ;
  assign n21009 = ~n20962 & n21008 ;
  assign n21010 = n20346 & n21009 ;
  assign n21011 = ~n20985 & n21007 ;
  assign n21012 = ~n20962 & n21011 ;
  assign n21013 = ~n20346 & n21012 ;
  assign n21014 = ~n21010 & ~n21013 ;
  assign n21015 = n20962 & n21008 ;
  assign n21016 = ~n20346 & n21015 ;
  assign n21017 = n20962 & n21011 ;
  assign n21018 = n20346 & n21017 ;
  assign n21019 = ~n21016 & ~n21018 ;
  assign n21020 = n21014 & n21019 ;
  assign n21021 = n20985 & ~n21007 ;
  assign n21022 = ~n20962 & n21021 ;
  assign n21023 = ~n20346 & n21022 ;
  assign n21024 = n20985 & n21007 ;
  assign n21025 = ~n20962 & n21024 ;
  assign n21026 = n20346 & n21025 ;
  assign n21027 = ~n21023 & ~n21026 ;
  assign n21028 = n20962 & n21021 ;
  assign n21029 = n20346 & n21028 ;
  assign n21030 = n20962 & n21024 ;
  assign n21031 = ~n20346 & n21030 ;
  assign n21032 = ~n21029 & ~n21031 ;
  assign n21033 = n21027 & n21032 ;
  assign n21034 = n21020 & n21033 ;
  assign n21035 = n20344 & n21034 ;
  assign n21036 = ~n20962 & n21007 ;
  assign n21037 = n20346 & n21036 ;
  assign n21038 = n20962 & n21007 ;
  assign n21039 = ~n20346 & n21038 ;
  assign n21040 = ~n21037 & ~n21039 ;
  assign n21041 = ~n20346 & n20962 ;
  assign n21042 = ~n20248 & ~n20962 ;
  assign n21043 = ~n20345 & n21042 ;
  assign n21044 = ~n21007 & ~n21043 ;
  assign n21045 = ~n21041 & n21044 ;
  assign n21046 = n21040 & ~n21045 ;
  assign n21047 = ~n20344 & n20985 ;
  assign n21048 = ~n21046 & n21047 ;
  assign n21049 = ~n20344 & ~n20985 ;
  assign n21050 = n21046 & n21049 ;
  assign n21051 = ~n21048 & ~n21050 ;
  assign n21052 = ~n21035 & n21051 ;
  assign n21053 = ~n20326 & ~n20330 ;
  assign n21054 = n21052 & ~n21053 ;
  assign n21055 = ~n20326 & ~n21052 ;
  assign n21056 = ~n20330 & n21055 ;
  assign n21057 = ~n21054 & ~n21056 ;
  assign n21058 = ~n20326 & ~n21035 ;
  assign n21059 = ~n20330 & n21058 ;
  assign n21060 = ~n20248 & n20956 ;
  assign n21061 = ~n20345 & n21060 ;
  assign n21062 = n20961 & ~n21061 ;
  assign n21063 = n20349 & n20934 ;
  assign n21064 = ~n20933 & ~n21063 ;
  assign n21065 = ~n20200 & n20922 ;
  assign n21066 = ~n20350 & n21065 ;
  assign n21067 = n20917 & ~n21066 ;
  assign n21068 = n646 & ~n15246 ;
  assign n21069 = ~n15244 & n21068 ;
  assign n21070 = \b[51]  & n796 ;
  assign n21071 = n793 & n21070 ;
  assign n21072 = \b[53]  & n644 ;
  assign n21073 = \a[8]  & \b[52]  ;
  assign n21074 = n794 & n21073 ;
  assign n21075 = ~\a[9]  & \b[52]  ;
  assign n21076 = n638 & n21075 ;
  assign n21077 = ~n21074 & ~n21076 ;
  assign n21078 = ~n21072 & n21077 ;
  assign n21079 = ~n21071 & n21078 ;
  assign n21080 = ~n21069 & n21079 ;
  assign n21081 = ~\a[11]  & ~n21080 ;
  assign n21082 = \a[11]  & n21079 ;
  assign n21083 = ~n21069 & n21082 ;
  assign n21084 = ~n21081 & ~n21083 ;
  assign n21085 = n20376 & n20912 ;
  assign n21086 = ~n20911 & ~n21085 ;
  assign n21087 = n20161 & n20895 ;
  assign n21088 = ~n20394 & n21087 ;
  assign n21089 = n20900 & ~n21088 ;
  assign n21090 = n1467 & ~n12438 ;
  assign n21091 = ~n12436 & n21090 ;
  assign n21092 = \b[47]  & n1465 ;
  assign n21093 = \a[15]  & \b[46]  ;
  assign n21094 = n1456 & n21093 ;
  assign n21095 = ~n21092 & ~n21094 ;
  assign n21096 = \b[45]  & n1652 ;
  assign n21097 = n1649 & n21096 ;
  assign n21098 = ~\a[15]  & \b[46]  ;
  assign n21099 = n1459 & n21098 ;
  assign n21100 = ~n21097 & ~n21099 ;
  assign n21101 = n21095 & n21100 ;
  assign n21102 = ~n21091 & n21101 ;
  assign n21103 = ~\a[17]  & ~n21102 ;
  assign n21104 = \a[17]  & n21101 ;
  assign n21105 = ~n21091 & n21104 ;
  assign n21106 = ~n21103 & ~n21105 ;
  assign n21107 = n20422 & n20873 ;
  assign n21108 = n20867 & ~n21107 ;
  assign n21109 = n1965 & ~n10892 ;
  assign n21110 = ~n10890 & n21109 ;
  assign n21111 = \b[42]  & n2218 ;
  assign n21112 = n2216 & n21111 ;
  assign n21113 = ~\a[18]  & \b[43]  ;
  assign n21114 = n1957 & n21113 ;
  assign n21115 = ~n21112 & ~n21114 ;
  assign n21116 = \b[44]  & n1963 ;
  assign n21117 = \a[18]  & \b[43]  ;
  assign n21118 = n2210 & n21117 ;
  assign n21119 = \a[20]  & ~n21118 ;
  assign n21120 = ~n21116 & n21119 ;
  assign n21121 = n21115 & n21120 ;
  assign n21122 = ~n21110 & n21121 ;
  assign n21123 = ~n21116 & ~n21118 ;
  assign n21124 = n21115 & n21123 ;
  assign n21125 = ~n21110 & n21124 ;
  assign n21126 = ~\a[20]  & ~n21125 ;
  assign n21127 = ~n21122 & ~n21126 ;
  assign n21128 = ~n20098 & n20831 ;
  assign n21129 = ~n20106 & n21128 ;
  assign n21130 = n20836 & ~n21129 ;
  assign n21131 = n20426 & n20809 ;
  assign n21132 = ~n20803 & ~n21131 ;
  assign n21133 = n20042 & n20768 ;
  assign n21134 = ~n20427 & n21133 ;
  assign n21135 = n20773 & ~n21134 ;
  assign n21136 = n4249 & ~n6610 ;
  assign n21137 = ~n6608 & n21136 ;
  assign n21138 = \b[35]  & n4247 ;
  assign n21139 = \a[27]  & \b[34]  ;
  assign n21140 = n4238 & n21139 ;
  assign n21141 = ~n21138 & ~n21140 ;
  assign n21142 = \b[33]  & n4647 ;
  assign n21143 = n4644 & n21142 ;
  assign n21144 = ~\a[27]  & \b[34]  ;
  assign n21145 = n4241 & n21144 ;
  assign n21146 = ~n21143 & ~n21145 ;
  assign n21147 = n21141 & n21146 ;
  assign n21148 = ~n21137 & n21147 ;
  assign n21149 = ~\a[29]  & ~n21148 ;
  assign n21150 = \a[29]  & n21147 ;
  assign n21151 = ~n21137 & n21150 ;
  assign n21152 = ~n21149 & ~n21151 ;
  assign n21153 = n20431 & n20744 ;
  assign n21154 = n20738 & ~n21153 ;
  assign n21155 = ~n19978 & ~n20703 ;
  assign n21156 = ~n19986 & n21155 ;
  assign n21157 = n20708 & ~n21156 ;
  assign n21158 = n20668 & ~n20677 ;
  assign n21159 = n19932 & ~n20661 ;
  assign n21160 = ~n20436 & n21159 ;
  assign n21161 = ~n20662 & ~n21160 ;
  assign n21162 = ~n3022 & n8759 ;
  assign n21163 = ~n3020 & n21162 ;
  assign n21164 = \b[23]  & n8757 ;
  assign n21165 = \a[39]  & \b[22]  ;
  assign n21166 = n8748 & n21165 ;
  assign n21167 = ~n21164 & ~n21166 ;
  assign n21168 = \b[21]  & n9301 ;
  assign n21169 = n9298 & n21168 ;
  assign n21170 = ~\a[39]  & \b[22]  ;
  assign n21171 = n8751 & n21170 ;
  assign n21172 = ~n21169 & ~n21171 ;
  assign n21173 = n21167 & n21172 ;
  assign n21174 = ~n21163 & n21173 ;
  assign n21175 = ~\a[41]  & ~n21174 ;
  assign n21176 = \a[41]  & n21173 ;
  assign n21177 = ~n21163 & n21176 ;
  assign n21178 = ~n21175 & ~n21177 ;
  assign n21179 = ~n20634 & ~n20642 ;
  assign n21180 = n2293 & n10082 ;
  assign n21181 = ~n19247 & n21180 ;
  assign n21182 = ~n2293 & n10082 ;
  assign n21183 = ~n2074 & n21182 ;
  assign n21184 = ~n2289 & n21183 ;
  assign n21185 = \b[18]  & n10681 ;
  assign n21186 = n10678 & n21185 ;
  assign n21187 = \b[20]  & n10080 ;
  assign n21188 = \a[42]  & \b[19]  ;
  assign n21189 = n10071 & n21188 ;
  assign n21190 = ~\a[42]  & \b[19]  ;
  assign n21191 = n10074 & n21190 ;
  assign n21192 = ~n21189 & ~n21191 ;
  assign n21193 = ~n21187 & n21192 ;
  assign n21194 = ~n21186 & n21193 ;
  assign n21195 = ~n21184 & n21194 ;
  assign n21196 = ~n21181 & n21195 ;
  assign n21197 = ~\a[44]  & ~n21196 ;
  assign n21198 = \a[44]  & n21194 ;
  assign n21199 = ~n21184 & n21198 ;
  assign n21200 = ~n21181 & n21199 ;
  assign n21201 = ~n21197 & ~n21200 ;
  assign n21202 = ~n19915 & n20601 ;
  assign n21203 = ~n20465 & n21202 ;
  assign n21204 = n20606 & ~n21203 ;
  assign n21205 = ~n1691 & n11572 ;
  assign n21206 = ~n1511 & n11572 ;
  assign n21207 = ~n1515 & n21206 ;
  assign n21208 = ~n21205 & ~n21207 ;
  assign n21209 = ~n1694 & ~n21208 ;
  assign n21210 = \b[15]  & n12159 ;
  assign n21211 = n12156 & n21210 ;
  assign n21212 = ~\a[45]  & \b[16]  ;
  assign n21213 = n11564 & n21212 ;
  assign n21214 = ~n21211 & ~n21213 ;
  assign n21215 = \b[17]  & n11570 ;
  assign n21216 = \a[45]  & \b[16]  ;
  assign n21217 = n11561 & n21216 ;
  assign n21218 = \a[47]  & ~n21217 ;
  assign n21219 = ~n21215 & n21218 ;
  assign n21220 = n21214 & n21219 ;
  assign n21221 = ~n21209 & n21220 ;
  assign n21222 = ~n21215 & ~n21217 ;
  assign n21223 = n21214 & n21222 ;
  assign n21224 = ~\a[47]  & ~n21223 ;
  assign n21225 = ~\a[47]  & ~n1694 ;
  assign n21226 = ~n21208 & n21225 ;
  assign n21227 = ~n21224 & ~n21226 ;
  assign n21228 = ~n21221 & n21227 ;
  assign n21229 = n20469 & n20572 ;
  assign n21230 = n20566 & ~n21229 ;
  assign n21231 = ~n725 & n14793 ;
  assign n21232 = ~n684 & n14793 ;
  assign n21233 = ~n721 & n21232 ;
  assign n21234 = ~n21231 & ~n21233 ;
  assign n21235 = ~n728 & ~n21234 ;
  assign n21236 = \b[9]  & n15517 ;
  assign n21237 = n15514 & n21236 ;
  assign n21238 = ~\a[51]  & \b[10]  ;
  assign n21239 = n14785 & n21238 ;
  assign n21240 = ~n21237 & ~n21239 ;
  assign n21241 = \b[11]  & n14791 ;
  assign n21242 = \a[51]  & \b[10]  ;
  assign n21243 = n14782 & n21242 ;
  assign n21244 = \a[53]  & ~n21243 ;
  assign n21245 = ~n21241 & n21244 ;
  assign n21246 = n21240 & n21245 ;
  assign n21247 = ~n21235 & n21246 ;
  assign n21248 = ~n21241 & ~n21243 ;
  assign n21249 = n21240 & n21248 ;
  assign n21250 = ~\a[53]  & ~n21249 ;
  assign n21251 = ~\a[53]  & ~n728 ;
  assign n21252 = ~n21234 & n21251 ;
  assign n21253 = ~n21250 & ~n21252 ;
  assign n21254 = ~n21247 & n21253 ;
  assign n21255 = ~n19892 & ~n20536 ;
  assign n21256 = ~n20470 & n21255 ;
  assign n21257 = ~n20535 & ~n21256 ;
  assign n21258 = ~n505 & ~n16016 ;
  assign n21259 = ~n16652 & n21258 ;
  assign n21260 = n502 & n21259 ;
  assign n21261 = n505 & ~n16016 ;
  assign n21262 = ~n16652 & n21261 ;
  assign n21263 = ~n502 & n21262 ;
  assign n21264 = ~n21260 & ~n21263 ;
  assign n21265 = \b[6]  & n17308 ;
  assign n21266 = n17305 & n21265 ;
  assign n21267 = ~\a[54]  & \b[7]  ;
  assign n21268 = n16647 & n21267 ;
  assign n21269 = ~n21266 & ~n21268 ;
  assign n21270 = \b[8]  & n16653 ;
  assign n21271 = \a[54]  & \b[7]  ;
  assign n21272 = n16644 & n21271 ;
  assign n21273 = \a[56]  & ~n21272 ;
  assign n21274 = ~n21270 & n21273 ;
  assign n21275 = n21269 & n21274 ;
  assign n21276 = n21264 & n21275 ;
  assign n21277 = ~n21270 & ~n21272 ;
  assign n21278 = n21269 & n21277 ;
  assign n21279 = n21264 & n21278 ;
  assign n21280 = ~\a[56]  & ~n21279 ;
  assign n21281 = ~n21276 & ~n21280 ;
  assign n21282 = ~n20530 & ~n20532 ;
  assign n21283 = ~n273 & n18516 ;
  assign n21284 = ~n271 & n21283 ;
  assign n21285 = \b[3]  & n19183 ;
  assign n21286 = n19180 & n21285 ;
  assign n21287 = \b[5]  & n18514 ;
  assign n21288 = \a[56]  & \b[4]  ;
  assign n21289 = n19181 & n21288 ;
  assign n21290 = ~\a[57]  & \b[4]  ;
  assign n21291 = n18508 & n21290 ;
  assign n21292 = ~n21289 & ~n21291 ;
  assign n21293 = ~n21287 & n21292 ;
  assign n21294 = ~n21286 & n21293 ;
  assign n21295 = ~\a[59]  & n21294 ;
  assign n21296 = ~n21284 & n21295 ;
  assign n21297 = ~n21284 & n21294 ;
  assign n21298 = \a[59]  & ~n21297 ;
  assign n21299 = ~n21296 & ~n21298 ;
  assign n21300 = \a[62]  & ~n19862 ;
  assign n21301 = n20515 & n21300 ;
  assign n21302 = n20523 & n21301 ;
  assign n21303 = \a[62]  & ~n21302 ;
  assign n21304 = \b[2]  & n20519 ;
  assign n21305 = ~\a[60]  & \b[1]  ;
  assign n21306 = n20513 & n21305 ;
  assign n21307 = \a[60]  & \b[1]  ;
  assign n21308 = n20510 & n21307 ;
  assign n21309 = ~n21306 & ~n21308 ;
  assign n21310 = ~n21304 & n21309 ;
  assign n21311 = n157 & n20521 ;
  assign n21312 = n19861 & ~n20518 ;
  assign n21313 = \a[60]  & ~\a[61]  ;
  assign n21314 = ~\a[60]  & \a[61]  ;
  assign n21315 = ~n21313 & ~n21314 ;
  assign n21316 = \b[0]  & n21315 ;
  assign n21317 = n21312 & n21316 ;
  assign n21318 = ~n21311 & ~n21317 ;
  assign n21319 = n21310 & n21318 ;
  assign n21320 = ~n21303 & ~n21319 ;
  assign n21321 = n21303 & n21319 ;
  assign n21322 = ~n21320 & ~n21321 ;
  assign n21323 = n21299 & ~n21322 ;
  assign n21324 = ~n21299 & n21322 ;
  assign n21325 = ~n21323 & ~n21324 ;
  assign n21326 = ~n21282 & n21325 ;
  assign n21327 = n21282 & ~n21325 ;
  assign n21328 = ~n21326 & ~n21327 ;
  assign n21329 = n21281 & ~n21328 ;
  assign n21330 = ~n21281 & n21328 ;
  assign n21331 = ~n21329 & ~n21330 ;
  assign n21332 = n21257 & n21331 ;
  assign n21333 = ~n21257 & ~n21331 ;
  assign n21334 = ~n21332 & ~n21333 ;
  assign n21335 = n21254 & ~n21334 ;
  assign n21336 = ~n21254 & n21334 ;
  assign n21337 = ~n21335 & ~n21336 ;
  assign n21338 = n1087 & n13125 ;
  assign n21339 = ~n1084 & n21338 ;
  assign n21340 = ~n946 & ~n1087 ;
  assign n21341 = n13125 & n21340 ;
  assign n21342 = ~n1083 & n21341 ;
  assign n21343 = \b[12]  & n13794 ;
  assign n21344 = n13792 & n21343 ;
  assign n21345 = ~\a[48]  & \b[13]  ;
  assign n21346 = n13117 & n21345 ;
  assign n21347 = ~n21344 & ~n21346 ;
  assign n21348 = \b[14]  & n13123 ;
  assign n21349 = \a[48]  & \b[13]  ;
  assign n21350 = n13786 & n21349 ;
  assign n21351 = \a[50]  & ~n21350 ;
  assign n21352 = ~n21348 & n21351 ;
  assign n21353 = n21347 & n21352 ;
  assign n21354 = ~n21342 & n21353 ;
  assign n21355 = ~n21339 & n21354 ;
  assign n21356 = ~n21348 & ~n21350 ;
  assign n21357 = n21347 & n21356 ;
  assign n21358 = ~n21342 & n21357 ;
  assign n21359 = ~n21339 & n21358 ;
  assign n21360 = ~\a[50]  & ~n21359 ;
  assign n21361 = ~n21355 & ~n21360 ;
  assign n21362 = ~n21337 & ~n21361 ;
  assign n21363 = ~n21230 & n21362 ;
  assign n21364 = n21337 & ~n21361 ;
  assign n21365 = n21230 & n21364 ;
  assign n21366 = ~n21363 & ~n21365 ;
  assign n21367 = ~n21337 & n21361 ;
  assign n21368 = n21230 & n21367 ;
  assign n21369 = n21337 & n21361 ;
  assign n21370 = ~n21230 & n21369 ;
  assign n21371 = ~n21368 & ~n21370 ;
  assign n21372 = n21366 & n21371 ;
  assign n21373 = ~n21228 & ~n21372 ;
  assign n21374 = n21204 & n21373 ;
  assign n21375 = ~n21228 & n21372 ;
  assign n21376 = ~n21204 & n21375 ;
  assign n21377 = ~n21374 & ~n21376 ;
  assign n21378 = n21228 & ~n21372 ;
  assign n21379 = ~n21204 & n21378 ;
  assign n21380 = n21228 & n21372 ;
  assign n21381 = n21204 & n21380 ;
  assign n21382 = ~n21379 & ~n21381 ;
  assign n21383 = n21377 & n21382 ;
  assign n21384 = ~n21201 & ~n21383 ;
  assign n21385 = ~n21179 & n21384 ;
  assign n21386 = ~n21201 & n21383 ;
  assign n21387 = n21179 & n21386 ;
  assign n21388 = ~n21385 & ~n21387 ;
  assign n21389 = n21201 & ~n21383 ;
  assign n21390 = n21179 & n21389 ;
  assign n21391 = n21201 & n21383 ;
  assign n21392 = ~n21179 & n21391 ;
  assign n21393 = ~n21390 & ~n21392 ;
  assign n21394 = n21388 & n21393 ;
  assign n21395 = ~n21178 & ~n21394 ;
  assign n21396 = n21161 & n21395 ;
  assign n21397 = ~n21178 & n21394 ;
  assign n21398 = ~n21161 & n21397 ;
  assign n21399 = ~n21396 & ~n21398 ;
  assign n21400 = n21178 & ~n21394 ;
  assign n21401 = ~n21161 & n21400 ;
  assign n21402 = n21178 & n21394 ;
  assign n21403 = n21161 & n21402 ;
  assign n21404 = ~n21401 & ~n21403 ;
  assign n21405 = n21399 & n21404 ;
  assign n21406 = ~n21158 & n21405 ;
  assign n21407 = n20668 & ~n21405 ;
  assign n21408 = ~n20677 & n21407 ;
  assign n21409 = n3604 & n7534 ;
  assign n21410 = ~n19292 & n21409 ;
  assign n21411 = n7534 & n12021 ;
  assign n21412 = ~n3600 & n21411 ;
  assign n21413 = \b[24]  & n7973 ;
  assign n21414 = n7970 & n21413 ;
  assign n21415 = ~\a[36]  & \b[25]  ;
  assign n21416 = n7526 & n21415 ;
  assign n21417 = ~n21414 & ~n21416 ;
  assign n21418 = \b[26]  & n7532 ;
  assign n21419 = \a[36]  & \b[25]  ;
  assign n21420 = n17801 & n21419 ;
  assign n21421 = \a[38]  & ~n21420 ;
  assign n21422 = ~n21418 & n21421 ;
  assign n21423 = n21417 & n21422 ;
  assign n21424 = ~n21412 & n21423 ;
  assign n21425 = ~n21410 & n21424 ;
  assign n21426 = ~n21418 & ~n21420 ;
  assign n21427 = n21417 & n21426 ;
  assign n21428 = ~n21412 & n21427 ;
  assign n21429 = ~n21410 & n21428 ;
  assign n21430 = ~\a[38]  & ~n21429 ;
  assign n21431 = ~n21425 & ~n21430 ;
  assign n21432 = ~n21408 & ~n21431 ;
  assign n21433 = ~n21406 & n21432 ;
  assign n21434 = ~n21405 & n21431 ;
  assign n21435 = n21158 & n21434 ;
  assign n21436 = n21405 & n21431 ;
  assign n21437 = ~n21158 & n21436 ;
  assign n21438 = ~n21435 & ~n21437 ;
  assign n21439 = ~n21433 & n21438 ;
  assign n21440 = ~n4502 & n6309 ;
  assign n21441 = ~n4500 & n21440 ;
  assign n21442 = \b[27]  & n6778 ;
  assign n21443 = n6775 & n21442 ;
  assign n21444 = ~\a[33]  & \b[28]  ;
  assign n21445 = n6301 & n21444 ;
  assign n21446 = ~n21443 & ~n21445 ;
  assign n21447 = \b[29]  & n6307 ;
  assign n21448 = \a[33]  & \b[28]  ;
  assign n21449 = n6298 & n21448 ;
  assign n21450 = \a[35]  & ~n21449 ;
  assign n21451 = ~n21447 & n21450 ;
  assign n21452 = n21446 & n21451 ;
  assign n21453 = ~n21441 & n21452 ;
  assign n21454 = ~n21447 & ~n21449 ;
  assign n21455 = n21446 & n21454 ;
  assign n21456 = ~n21441 & n21455 ;
  assign n21457 = ~\a[35]  & ~n21456 ;
  assign n21458 = ~n21453 & ~n21457 ;
  assign n21459 = ~n21439 & ~n21458 ;
  assign n21460 = n21157 & n21459 ;
  assign n21461 = n21439 & ~n21458 ;
  assign n21462 = ~n21157 & n21461 ;
  assign n21463 = ~n21460 & ~n21462 ;
  assign n21464 = ~n21439 & n21458 ;
  assign n21465 = ~n21157 & n21464 ;
  assign n21466 = n21439 & n21458 ;
  assign n21467 = n21157 & n21466 ;
  assign n21468 = ~n21465 & ~n21467 ;
  assign n21469 = n21463 & n21468 ;
  assign n21470 = ~n21154 & n21469 ;
  assign n21471 = n20738 & ~n21469 ;
  assign n21472 = ~n21153 & n21471 ;
  assign n21473 = n5211 & n5810 ;
  assign n21474 = ~n5807 & n21473 ;
  assign n21475 = n5211 & n19029 ;
  assign n21476 = ~n5806 & n21475 ;
  assign n21477 = \b[30]  & n5595 ;
  assign n21478 = n5592 & n21477 ;
  assign n21479 = ~\a[30]  & \b[31]  ;
  assign n21480 = n5203 & n21479 ;
  assign n21481 = ~n21478 & ~n21480 ;
  assign n21482 = \b[32]  & n5209 ;
  assign n21483 = \a[30]  & \b[31]  ;
  assign n21484 = n5200 & n21483 ;
  assign n21485 = \a[32]  & ~n21484 ;
  assign n21486 = ~n21482 & n21485 ;
  assign n21487 = n21481 & n21486 ;
  assign n21488 = ~n21476 & n21487 ;
  assign n21489 = ~n21474 & n21488 ;
  assign n21490 = ~n21482 & ~n21484 ;
  assign n21491 = n21481 & n21490 ;
  assign n21492 = ~n21476 & n21491 ;
  assign n21493 = ~n21474 & n21492 ;
  assign n21494 = ~\a[32]  & ~n21493 ;
  assign n21495 = ~n21489 & ~n21494 ;
  assign n21496 = ~n21472 & ~n21495 ;
  assign n21497 = ~n21470 & n21496 ;
  assign n21498 = ~n21469 & n21495 ;
  assign n21499 = n21154 & n21498 ;
  assign n21500 = n21469 & n21495 ;
  assign n21501 = ~n21154 & n21500 ;
  assign n21502 = ~n21499 & ~n21501 ;
  assign n21503 = ~n21497 & n21502 ;
  assign n21504 = ~n21152 & ~n21503 ;
  assign n21505 = n21135 & n21504 ;
  assign n21506 = ~n21152 & n21503 ;
  assign n21507 = ~n21135 & n21506 ;
  assign n21508 = ~n21505 & ~n21507 ;
  assign n21509 = n21152 & ~n21503 ;
  assign n21510 = ~n21135 & n21509 ;
  assign n21511 = n21152 & n21503 ;
  assign n21512 = n21135 & n21511 ;
  assign n21513 = ~n21510 & ~n21512 ;
  assign n21514 = n21508 & n21513 ;
  assign n21515 = ~n21132 & n21514 ;
  assign n21516 = ~n20803 & ~n21514 ;
  assign n21517 = ~n21131 & n21516 ;
  assign n21518 = n3402 & n8175 ;
  assign n21519 = ~n8172 & n21518 ;
  assign n21520 = n3402 & ~n8175 ;
  assign n21521 = ~n7756 & n21520 ;
  assign n21522 = ~n8171 & n21521 ;
  assign n21523 = \b[36]  & n3733 ;
  assign n21524 = n3730 & n21523 ;
  assign n21525 = \b[38]  & n3400 ;
  assign n21526 = \a[23]  & \b[37]  ;
  assign n21527 = n3731 & n21526 ;
  assign n21528 = ~\a[24]  & \b[37]  ;
  assign n21529 = n3394 & n21528 ;
  assign n21530 = ~n21527 & ~n21529 ;
  assign n21531 = ~n21525 & n21530 ;
  assign n21532 = ~n21524 & n21531 ;
  assign n21533 = ~n21522 & n21532 ;
  assign n21534 = ~n21519 & n21533 ;
  assign n21535 = ~\a[26]  & ~n21534 ;
  assign n21536 = \a[26]  & n21532 ;
  assign n21537 = ~n21522 & n21536 ;
  assign n21538 = ~n21519 & n21537 ;
  assign n21539 = ~n21535 & ~n21538 ;
  assign n21540 = ~n21517 & ~n21539 ;
  assign n21541 = ~n21515 & n21540 ;
  assign n21542 = ~n21514 & n21539 ;
  assign n21543 = n21132 & n21542 ;
  assign n21544 = n21514 & n21539 ;
  assign n21545 = ~n21132 & n21544 ;
  assign n21546 = ~n21543 & ~n21545 ;
  assign n21547 = ~n21541 & n21546 ;
  assign n21548 = ~n21130 & ~n21547 ;
  assign n21549 = n21130 & n21547 ;
  assign n21550 = ~n21548 & ~n21549 ;
  assign n21551 = n2622 & ~n9482 ;
  assign n21552 = ~n9480 & n21551 ;
  assign n21553 = \b[41]  & n2620 ;
  assign n21554 = \a[21]  & \b[40]  ;
  assign n21555 = n20849 & n21554 ;
  assign n21556 = ~n21553 & ~n21555 ;
  assign n21557 = \b[39]  & n2912 ;
  assign n21558 = n2909 & n21557 ;
  assign n21559 = ~\a[21]  & \b[40]  ;
  assign n21560 = n2614 & n21559 ;
  assign n21561 = ~n21558 & ~n21560 ;
  assign n21562 = n21556 & n21561 ;
  assign n21563 = ~n21552 & n21562 ;
  assign n21564 = ~\a[23]  & ~n21563 ;
  assign n21565 = \a[23]  & n21562 ;
  assign n21566 = ~n21552 & n21565 ;
  assign n21567 = ~n21564 & ~n21566 ;
  assign n21568 = n21550 & ~n21567 ;
  assign n21569 = ~n21550 & n21567 ;
  assign n21570 = ~n21568 & ~n21569 ;
  assign n21571 = ~n21127 & ~n21570 ;
  assign n21572 = ~n21108 & n21571 ;
  assign n21573 = ~n21127 & n21570 ;
  assign n21574 = n21108 & n21573 ;
  assign n21575 = ~n21572 & ~n21574 ;
  assign n21576 = n21127 & ~n21570 ;
  assign n21577 = n21108 & n21576 ;
  assign n21578 = n21127 & n21570 ;
  assign n21579 = ~n21108 & n21578 ;
  assign n21580 = ~n21577 & ~n21579 ;
  assign n21581 = n21575 & n21580 ;
  assign n21582 = ~n21106 & ~n21581 ;
  assign n21583 = n21089 & n21582 ;
  assign n21584 = ~n21106 & n21581 ;
  assign n21585 = ~n21089 & n21584 ;
  assign n21586 = ~n21583 & ~n21585 ;
  assign n21587 = n21106 & ~n21581 ;
  assign n21588 = ~n21089 & n21587 ;
  assign n21589 = n21106 & n21581 ;
  assign n21590 = n21089 & n21589 ;
  assign n21591 = ~n21588 & ~n21590 ;
  assign n21592 = n21586 & n21591 ;
  assign n21593 = ~n21086 & n21592 ;
  assign n21594 = ~n20911 & ~n21592 ;
  assign n21595 = ~n21085 & n21594 ;
  assign n21596 = n999 & n14052 ;
  assign n21597 = ~n14049 & n21596 ;
  assign n21598 = n999 & ~n14052 ;
  assign n21599 = ~n13519 & n21598 ;
  assign n21600 = ~n14048 & n21599 ;
  assign n21601 = \b[48]  & n1182 ;
  assign n21602 = n1179 & n21601 ;
  assign n21603 = \b[50]  & n997 ;
  assign n21604 = \a[11]  & \b[49]  ;
  assign n21605 = n1180 & n21604 ;
  assign n21606 = ~\a[12]  & \b[49]  ;
  assign n21607 = n7674 & n21606 ;
  assign n21608 = ~n21605 & ~n21607 ;
  assign n21609 = ~n21603 & n21608 ;
  assign n21610 = ~n21602 & n21609 ;
  assign n21611 = ~n21600 & n21610 ;
  assign n21612 = ~n21597 & n21611 ;
  assign n21613 = ~\a[14]  & ~n21612 ;
  assign n21614 = \a[14]  & n21610 ;
  assign n21615 = ~n21600 & n21614 ;
  assign n21616 = ~n21597 & n21615 ;
  assign n21617 = ~n21613 & ~n21616 ;
  assign n21618 = ~n21595 & ~n21617 ;
  assign n21619 = ~n21593 & n21618 ;
  assign n21620 = ~n21592 & n21617 ;
  assign n21621 = n21086 & n21620 ;
  assign n21622 = n21592 & n21617 ;
  assign n21623 = ~n21086 & n21622 ;
  assign n21624 = ~n21621 & ~n21623 ;
  assign n21625 = ~n21619 & n21624 ;
  assign n21626 = ~n21084 & ~n21625 ;
  assign n21627 = n21067 & n21626 ;
  assign n21628 = ~n21084 & n21625 ;
  assign n21629 = ~n21067 & n21628 ;
  assign n21630 = ~n21627 & ~n21629 ;
  assign n21631 = n21084 & ~n21625 ;
  assign n21632 = ~n21067 & n21631 ;
  assign n21633 = n21084 & n21625 ;
  assign n21634 = n21067 & n21633 ;
  assign n21635 = ~n21632 & ~n21634 ;
  assign n21636 = n21630 & n21635 ;
  assign n21637 = ~n359 & ~n16441 ;
  assign n21638 = ~n17647 & n21637 ;
  assign n21639 = ~n17643 & n21638 ;
  assign n21640 = ~n427 & n21639 ;
  assign n21641 = n430 & n17647 ;
  assign n21642 = ~n17644 & n21641 ;
  assign n21643 = ~n21640 & ~n21642 ;
  assign n21644 = \b[54]  & n486 ;
  assign n21645 = n483 & n21644 ;
  assign n21646 = ~\a[6]  & \b[55]  ;
  assign n21647 = n422 & n21646 ;
  assign n21648 = ~n21645 & ~n21647 ;
  assign n21649 = \b[56]  & n428 ;
  assign n21650 = \a[6]  & \b[55]  ;
  assign n21651 = n419 & n21650 ;
  assign n21652 = \a[8]  & ~n21651 ;
  assign n21653 = ~n21649 & n21652 ;
  assign n21654 = n21648 & n21653 ;
  assign n21655 = n21643 & n21654 ;
  assign n21656 = ~n21649 & ~n21651 ;
  assign n21657 = n21648 & n21656 ;
  assign n21658 = n21643 & n21657 ;
  assign n21659 = ~\a[8]  & ~n21658 ;
  assign n21660 = ~n21655 & ~n21659 ;
  assign n21661 = ~n21636 & n21660 ;
  assign n21662 = n21064 & n21661 ;
  assign n21663 = n21636 & n21660 ;
  assign n21664 = ~n21064 & n21663 ;
  assign n21665 = ~n21662 & ~n21664 ;
  assign n21666 = ~n21064 & n21636 ;
  assign n21667 = ~n20933 & ~n21636 ;
  assign n21668 = ~n21063 & n21667 ;
  assign n21669 = ~n21660 & ~n21668 ;
  assign n21670 = ~n21666 & n21669 ;
  assign n21671 = n21665 & ~n21670 ;
  assign n21672 = n252 & ~n19550 ;
  assign n21673 = ~n19548 & n21672 ;
  assign n21674 = \b[57]  & n303 ;
  assign n21675 = n300 & n21674 ;
  assign n21676 = ~\a[3]  & \b[58]  ;
  assign n21677 = n244 & n21676 ;
  assign n21678 = ~n21675 & ~n21677 ;
  assign n21679 = \b[59]  & n250 ;
  assign n21680 = \a[3]  & \b[58]  ;
  assign n21681 = n241 & n21680 ;
  assign n21682 = \a[5]  & ~n21681 ;
  assign n21683 = ~n21679 & n21682 ;
  assign n21684 = n21678 & n21683 ;
  assign n21685 = ~n21673 & n21684 ;
  assign n21686 = ~n21679 & ~n21681 ;
  assign n21687 = n21678 & n21686 ;
  assign n21688 = ~n21673 & n21687 ;
  assign n21689 = ~\a[5]  & ~n21688 ;
  assign n21690 = ~n21685 & ~n21689 ;
  assign n21691 = ~n20259 & ~n20967 ;
  assign n21692 = ~n20964 & n21691 ;
  assign n21693 = ~n20966 & ~n21692 ;
  assign n21694 = ~\b[61]  & ~\b[62]  ;
  assign n21695 = \b[61]  & \b[62]  ;
  assign n21696 = ~n21694 & ~n21695 ;
  assign n21697 = ~n21693 & ~n21696 ;
  assign n21698 = ~n20966 & n21696 ;
  assign n21699 = ~n21692 & n21698 ;
  assign n21700 = n134 & ~n21699 ;
  assign n21701 = ~n21697 & n21700 ;
  assign n21702 = \a[0]  & \b[62]  ;
  assign n21703 = n133 & n21702 ;
  assign n21704 = \b[61]  & n141 ;
  assign n21705 = ~\a[1]  & \b[60]  ;
  assign n21706 = n10416 & n21705 ;
  assign n21707 = ~n21704 & ~n21706 ;
  assign n21708 = ~n21703 & n21707 ;
  assign n21709 = \a[2]  & n21708 ;
  assign n21710 = ~n21701 & n21709 ;
  assign n21711 = ~n21701 & n21708 ;
  assign n21712 = ~\a[2]  & ~n21711 ;
  assign n21713 = ~n21710 & ~n21712 ;
  assign n21714 = n21690 & ~n21713 ;
  assign n21715 = ~n21671 & n21714 ;
  assign n21716 = ~n21062 & n21715 ;
  assign n21717 = ~n21690 & ~n21713 ;
  assign n21718 = n21671 & n21717 ;
  assign n21719 = ~n21062 & n21718 ;
  assign n21720 = ~n21716 & ~n21719 ;
  assign n21721 = ~n21671 & n21717 ;
  assign n21722 = n21062 & n21721 ;
  assign n21723 = n21671 & n21714 ;
  assign n21724 = n21062 & n21723 ;
  assign n21725 = ~n21722 & ~n21724 ;
  assign n21726 = n21720 & n21725 ;
  assign n21727 = n21671 & ~n21690 ;
  assign n21728 = ~n21062 & n21727 ;
  assign n21729 = ~n21671 & n21690 ;
  assign n21730 = ~n21062 & n21729 ;
  assign n21731 = ~n21728 & ~n21730 ;
  assign n21732 = ~n21660 & ~n21690 ;
  assign n21733 = ~n21636 & n21732 ;
  assign n21734 = n21064 & n21733 ;
  assign n21735 = n21660 & ~n21690 ;
  assign n21736 = ~n21636 & n21735 ;
  assign n21737 = ~n21064 & n21736 ;
  assign n21738 = ~n21734 & ~n21737 ;
  assign n21739 = n21636 & n21732 ;
  assign n21740 = ~n21064 & n21739 ;
  assign n21741 = n21636 & n21735 ;
  assign n21742 = n21064 & n21741 ;
  assign n21743 = ~n21740 & ~n21742 ;
  assign n21744 = n21738 & n21743 ;
  assign n21745 = ~n21660 & n21690 ;
  assign n21746 = ~n21636 & n21745 ;
  assign n21747 = ~n21064 & n21746 ;
  assign n21748 = n21660 & n21690 ;
  assign n21749 = ~n21636 & n21748 ;
  assign n21750 = n21064 & n21749 ;
  assign n21751 = ~n21747 & ~n21750 ;
  assign n21752 = n21636 & n21745 ;
  assign n21753 = n21064 & n21752 ;
  assign n21754 = n21636 & n21748 ;
  assign n21755 = ~n21064 & n21754 ;
  assign n21756 = ~n21753 & ~n21755 ;
  assign n21757 = n21751 & n21756 ;
  assign n21758 = n21744 & n21757 ;
  assign n21759 = n21062 & n21758 ;
  assign n21760 = n21713 & ~n21759 ;
  assign n21761 = n21731 & n21760 ;
  assign n21762 = n21726 & ~n21761 ;
  assign n21763 = \a[2]  & ~n20983 ;
  assign n21764 = ~\a[2]  & n20983 ;
  assign n21765 = ~n21763 & ~n21764 ;
  assign n21766 = n21040 & n21765 ;
  assign n21767 = ~n21045 & ~n21766 ;
  assign n21768 = ~n21762 & ~n21767 ;
  assign n21769 = n21762 & n21767 ;
  assign n21770 = ~n21768 & ~n21769 ;
  assign n21771 = n21051 & n21770 ;
  assign n21772 = ~n21059 & n21771 ;
  assign n21773 = n21051 & ~n21059 ;
  assign n21774 = ~n21770 & ~n21773 ;
  assign n21775 = ~n21772 & ~n21774 ;
  assign n21776 = \a[5]  & ~n21688 ;
  assign n21777 = ~\a[5]  & n21688 ;
  assign n21778 = ~n21776 & ~n21777 ;
  assign n21779 = n21665 & n21778 ;
  assign n21780 = ~n21670 & ~n21779 ;
  assign n21781 = ~n20933 & n21630 ;
  assign n21782 = ~n21063 & n21781 ;
  assign n21783 = n21635 & ~n21782 ;
  assign n21784 = n21067 & n21625 ;
  assign n21785 = ~n21619 & ~n21784 ;
  assign n21786 = ~n20911 & n21586 ;
  assign n21787 = ~n21085 & n21786 ;
  assign n21788 = n21591 & ~n21787 ;
  assign n21789 = n999 & ~n14098 ;
  assign n21790 = ~n14096 & n21789 ;
  assign n21791 = \b[49]  & n1182 ;
  assign n21792 = n1179 & n21791 ;
  assign n21793 = \b[51]  & n997 ;
  assign n21794 = \a[11]  & \b[50]  ;
  assign n21795 = n1180 & n21794 ;
  assign n21796 = ~\a[12]  & \b[50]  ;
  assign n21797 = n7674 & n21796 ;
  assign n21798 = ~n21795 & ~n21797 ;
  assign n21799 = ~n21793 & n21798 ;
  assign n21800 = ~n21792 & n21799 ;
  assign n21801 = ~n21790 & n21800 ;
  assign n21802 = ~\a[14]  & ~n21801 ;
  assign n21803 = \a[14]  & n21800 ;
  assign n21804 = ~n21790 & n21803 ;
  assign n21805 = ~n21802 & ~n21804 ;
  assign n21806 = n21089 & n21581 ;
  assign n21807 = n21575 & ~n21806 ;
  assign n21808 = n20867 & ~n21568 ;
  assign n21809 = ~n21107 & n21808 ;
  assign n21810 = ~n21569 & ~n21809 ;
  assign n21811 = n1965 & ~n11397 ;
  assign n21812 = ~n11395 & n21811 ;
  assign n21813 = \b[45]  & n1963 ;
  assign n21814 = \a[18]  & \b[44]  ;
  assign n21815 = n2210 & n21814 ;
  assign n21816 = ~n21813 & ~n21815 ;
  assign n21817 = \b[43]  & n2218 ;
  assign n21818 = n2216 & n21817 ;
  assign n21819 = ~\a[18]  & \b[44]  ;
  assign n21820 = n1957 & n21819 ;
  assign n21821 = ~n21818 & ~n21820 ;
  assign n21822 = n21816 & n21821 ;
  assign n21823 = ~n21812 & n21822 ;
  assign n21824 = ~\a[20]  & ~n21823 ;
  assign n21825 = \a[20]  & n21822 ;
  assign n21826 = ~n21812 & n21825 ;
  assign n21827 = ~n21824 & ~n21826 ;
  assign n21828 = ~n21541 & ~n21549 ;
  assign n21829 = n2622 & n9930 ;
  assign n21830 = ~n9927 & n21829 ;
  assign n21831 = n2622 & ~n9930 ;
  assign n21832 = ~n9477 & n21831 ;
  assign n21833 = ~n9926 & n21832 ;
  assign n21834 = \b[40]  & n2912 ;
  assign n21835 = n2909 & n21834 ;
  assign n21836 = ~\a[21]  & \b[41]  ;
  assign n21837 = n2614 & n21836 ;
  assign n21838 = ~n21835 & ~n21837 ;
  assign n21839 = \b[42]  & n2620 ;
  assign n21840 = \a[21]  & \b[41]  ;
  assign n21841 = n20849 & n21840 ;
  assign n21842 = \a[23]  & ~n21841 ;
  assign n21843 = ~n21839 & n21842 ;
  assign n21844 = n21838 & n21843 ;
  assign n21845 = ~n21833 & n21844 ;
  assign n21846 = ~n21830 & n21845 ;
  assign n21847 = ~n21839 & ~n21841 ;
  assign n21848 = n21838 & n21847 ;
  assign n21849 = ~n21833 & n21848 ;
  assign n21850 = ~n21830 & n21849 ;
  assign n21851 = ~\a[23]  & ~n21850 ;
  assign n21852 = ~n21846 & ~n21851 ;
  assign n21853 = ~n20803 & n21508 ;
  assign n21854 = ~n21131 & n21853 ;
  assign n21855 = n21513 & ~n21854 ;
  assign n21856 = n21135 & n21503 ;
  assign n21857 = ~n21497 & ~n21856 ;
  assign n21858 = n21157 & n21439 ;
  assign n21859 = ~n21433 & ~n21858 ;
  assign n21860 = n20668 & n21399 ;
  assign n21861 = ~n20677 & n21860 ;
  assign n21862 = n21404 & ~n21861 ;
  assign n21863 = n21161 & n21394 ;
  assign n21864 = n21388 & ~n21863 ;
  assign n21865 = ~n2523 & n10082 ;
  assign n21866 = ~n2521 & n21865 ;
  assign n21867 = \b[19]  & n10681 ;
  assign n21868 = n10678 & n21867 ;
  assign n21869 = \b[21]  & n10080 ;
  assign n21870 = \a[42]  & \b[20]  ;
  assign n21871 = n10071 & n21870 ;
  assign n21872 = ~\a[42]  & \b[20]  ;
  assign n21873 = n10074 & n21872 ;
  assign n21874 = ~n21871 & ~n21873 ;
  assign n21875 = ~n21869 & n21874 ;
  assign n21876 = ~n21868 & n21875 ;
  assign n21877 = ~n21866 & n21876 ;
  assign n21878 = ~\a[44]  & ~n21877 ;
  assign n21879 = \a[44]  & n21876 ;
  assign n21880 = ~n21866 & n21879 ;
  assign n21881 = ~n21878 & ~n21880 ;
  assign n21882 = ~n20634 & n21377 ;
  assign n21883 = ~n20642 & n21882 ;
  assign n21884 = n21382 & ~n21883 ;
  assign n21885 = n21204 & n21372 ;
  assign n21886 = n21366 & ~n21885 ;
  assign n21887 = n20566 & ~n21336 ;
  assign n21888 = ~n21229 & n21887 ;
  assign n21889 = ~n21335 & ~n21888 ;
  assign n21890 = ~n21330 & ~n21332 ;
  assign n21891 = ~n909 & ~n14276 ;
  assign n21892 = ~n14790 & n21891 ;
  assign n21893 = n906 & n21892 ;
  assign n21894 = n909 & ~n14276 ;
  assign n21895 = ~n14790 & n21894 ;
  assign n21896 = ~n906 & n21895 ;
  assign n21897 = ~n21893 & ~n21896 ;
  assign n21898 = \b[10]  & n15517 ;
  assign n21899 = n15514 & n21898 ;
  assign n21900 = ~\a[51]  & \b[11]  ;
  assign n21901 = n14785 & n21900 ;
  assign n21902 = ~n21899 & ~n21901 ;
  assign n21903 = \b[12]  & n14791 ;
  assign n21904 = \a[51]  & \b[11]  ;
  assign n21905 = n14782 & n21904 ;
  assign n21906 = \a[53]  & ~n21905 ;
  assign n21907 = ~n21903 & n21906 ;
  assign n21908 = n21902 & n21907 ;
  assign n21909 = n21897 & n21908 ;
  assign n21910 = ~n21903 & ~n21905 ;
  assign n21911 = n21902 & n21910 ;
  assign n21912 = n21897 & n21911 ;
  assign n21913 = ~\a[53]  & ~n21912 ;
  assign n21914 = ~n21909 & ~n21913 ;
  assign n21915 = ~n20530 & ~n21323 ;
  assign n21916 = ~n20532 & n21915 ;
  assign n21917 = ~n21324 & ~n21916 ;
  assign n21918 = ~n323 & ~n17912 ;
  assign n21919 = ~n18513 & n21918 ;
  assign n21920 = n320 & n21919 ;
  assign n21921 = n323 & ~n17912 ;
  assign n21922 = ~n18513 & n21921 ;
  assign n21923 = ~n320 & n21922 ;
  assign n21924 = ~n21920 & ~n21923 ;
  assign n21925 = \b[4]  & n19183 ;
  assign n21926 = n19180 & n21925 ;
  assign n21927 = \b[6]  & n18514 ;
  assign n21928 = \a[56]  & \b[5]  ;
  assign n21929 = n19181 & n21928 ;
  assign n21930 = ~\a[57]  & \b[5]  ;
  assign n21931 = n18508 & n21930 ;
  assign n21932 = ~n21929 & ~n21931 ;
  assign n21933 = ~n21927 & n21932 ;
  assign n21934 = ~n21926 & n21933 ;
  assign n21935 = n21924 & n21934 ;
  assign n21936 = ~\a[59]  & ~n21935 ;
  assign n21937 = \a[59]  & n21934 ;
  assign n21938 = n21924 & n21937 ;
  assign n21939 = ~n21936 & ~n21938 ;
  assign n21940 = n177 & n20521 ;
  assign n21941 = \b[3]  & n20519 ;
  assign n21942 = \a[59]  & \b[2]  ;
  assign n21943 = n21313 & n21942 ;
  assign n21944 = ~\a[60]  & \b[2]  ;
  assign n21945 = n20513 & n21944 ;
  assign n21946 = ~n21943 & ~n21945 ;
  assign n21947 = ~n21941 & n21946 ;
  assign n21948 = ~n21940 & n21947 ;
  assign n21949 = \b[1]  & n21315 ;
  assign n21950 = n21312 & n21949 ;
  assign n21951 = ~\a[62]  & ~n21950 ;
  assign n21952 = n21948 & n21951 ;
  assign n21953 = n21948 & ~n21950 ;
  assign n21954 = \a[62]  & ~n21953 ;
  assign n21955 = ~n21952 & ~n21954 ;
  assign n21956 = ~\a[62]  & ~\a[63]  ;
  assign n21957 = \a[62]  & \a[63]  ;
  assign n21958 = ~n21956 & ~n21957 ;
  assign n21959 = \b[0]  & n21958 ;
  assign n21960 = n21302 & n21319 ;
  assign n21961 = n21959 & n21960 ;
  assign n21962 = ~n21959 & ~n21960 ;
  assign n21963 = ~n21961 & ~n21962 ;
  assign n21964 = n21955 & n21963 ;
  assign n21965 = ~n21955 & ~n21963 ;
  assign n21966 = ~n21964 & ~n21965 ;
  assign n21967 = n21939 & ~n21966 ;
  assign n21968 = ~n21939 & n21966 ;
  assign n21969 = ~n21967 & ~n21968 ;
  assign n21970 = ~n586 & n16655 ;
  assign n21971 = ~n504 & n16655 ;
  assign n21972 = ~n508 & n21971 ;
  assign n21973 = ~n21970 & ~n21972 ;
  assign n21974 = ~n589 & ~n21973 ;
  assign n21975 = \b[7]  & n17308 ;
  assign n21976 = n17305 & n21975 ;
  assign n21977 = ~\a[54]  & \b[8]  ;
  assign n21978 = n16647 & n21977 ;
  assign n21979 = ~n21976 & ~n21978 ;
  assign n21980 = \b[9]  & n16653 ;
  assign n21981 = \a[54]  & \b[8]  ;
  assign n21982 = n16644 & n21981 ;
  assign n21983 = \a[56]  & ~n21982 ;
  assign n21984 = ~n21980 & n21983 ;
  assign n21985 = n21979 & n21984 ;
  assign n21986 = ~n21974 & n21985 ;
  assign n21987 = ~n21980 & ~n21982 ;
  assign n21988 = n21979 & n21987 ;
  assign n21989 = ~\a[56]  & ~n21988 ;
  assign n21990 = ~\a[56]  & ~n589 ;
  assign n21991 = ~n21973 & n21990 ;
  assign n21992 = ~n21989 & ~n21991 ;
  assign n21993 = ~n21986 & n21992 ;
  assign n21994 = ~n21969 & ~n21993 ;
  assign n21995 = n21917 & n21994 ;
  assign n21996 = n21969 & ~n21993 ;
  assign n21997 = ~n21917 & n21996 ;
  assign n21998 = ~n21995 & ~n21997 ;
  assign n21999 = ~n21969 & n21993 ;
  assign n22000 = ~n21917 & n21999 ;
  assign n22001 = n21969 & n21993 ;
  assign n22002 = n21917 & n22001 ;
  assign n22003 = ~n22000 & ~n22002 ;
  assign n22004 = n21998 & n22003 ;
  assign n22005 = n21914 & ~n22004 ;
  assign n22006 = n21890 & n22005 ;
  assign n22007 = n21914 & n22004 ;
  assign n22008 = ~n21890 & n22007 ;
  assign n22009 = ~n22006 & ~n22008 ;
  assign n22010 = ~n21890 & n22004 ;
  assign n22011 = ~n21330 & ~n22004 ;
  assign n22012 = ~n21332 & n22011 ;
  assign n22013 = ~n21914 & ~n22012 ;
  assign n22014 = ~n22010 & n22013 ;
  assign n22015 = n22009 & ~n22014 ;
  assign n22016 = ~n1233 & n13125 ;
  assign n22017 = ~n1231 & n22016 ;
  assign n22018 = \b[15]  & n13123 ;
  assign n22019 = \a[48]  & \b[14]  ;
  assign n22020 = n13786 & n22019 ;
  assign n22021 = ~n22018 & ~n22020 ;
  assign n22022 = \b[13]  & n13794 ;
  assign n22023 = n13792 & n22022 ;
  assign n22024 = ~\a[48]  & \b[14]  ;
  assign n22025 = n13117 & n22024 ;
  assign n22026 = ~n22023 & ~n22025 ;
  assign n22027 = n22021 & n22026 ;
  assign n22028 = ~n22017 & n22027 ;
  assign n22029 = ~\a[50]  & ~n22028 ;
  assign n22030 = \a[50]  & n22027 ;
  assign n22031 = ~n22017 & n22030 ;
  assign n22032 = ~n22029 & ~n22031 ;
  assign n22033 = ~n22015 & ~n22032 ;
  assign n22034 = n21889 & n22033 ;
  assign n22035 = n22015 & ~n22032 ;
  assign n22036 = ~n21889 & n22035 ;
  assign n22037 = ~n22034 & ~n22036 ;
  assign n22038 = ~n22015 & n22032 ;
  assign n22039 = ~n21889 & n22038 ;
  assign n22040 = n22015 & n22032 ;
  assign n22041 = n21889 & n22040 ;
  assign n22042 = ~n22039 & ~n22041 ;
  assign n22043 = n22037 & n22042 ;
  assign n22044 = n1875 & n11572 ;
  assign n22045 = ~n1872 & n22044 ;
  assign n22046 = n5000 & n11572 ;
  assign n22047 = ~n1871 & n22046 ;
  assign n22048 = \b[16]  & n12159 ;
  assign n22049 = n12156 & n22048 ;
  assign n22050 = ~\a[45]  & \b[17]  ;
  assign n22051 = n11564 & n22050 ;
  assign n22052 = ~n22049 & ~n22051 ;
  assign n22053 = \b[18]  & n11570 ;
  assign n22054 = \a[45]  & \b[17]  ;
  assign n22055 = n11561 & n22054 ;
  assign n22056 = \a[47]  & ~n22055 ;
  assign n22057 = ~n22053 & n22056 ;
  assign n22058 = n22052 & n22057 ;
  assign n22059 = ~n22047 & n22058 ;
  assign n22060 = ~n22045 & n22059 ;
  assign n22061 = ~n22053 & ~n22055 ;
  assign n22062 = n22052 & n22061 ;
  assign n22063 = ~n22047 & n22062 ;
  assign n22064 = ~n22045 & n22063 ;
  assign n22065 = ~\a[47]  & ~n22064 ;
  assign n22066 = ~n22060 & ~n22065 ;
  assign n22067 = ~n22043 & n22066 ;
  assign n22068 = n21886 & n22067 ;
  assign n22069 = n22043 & n22066 ;
  assign n22070 = ~n21886 & n22069 ;
  assign n22071 = ~n22068 & ~n22070 ;
  assign n22072 = ~n21886 & n22043 ;
  assign n22073 = n21366 & ~n22043 ;
  assign n22074 = ~n21885 & n22073 ;
  assign n22075 = ~n22066 & ~n22074 ;
  assign n22076 = ~n22072 & n22075 ;
  assign n22077 = n22071 & ~n22076 ;
  assign n22078 = n21884 & n22077 ;
  assign n22079 = ~n21884 & ~n22077 ;
  assign n22080 = ~n22078 & ~n22079 ;
  assign n22081 = ~n21881 & n22080 ;
  assign n22082 = n21881 & ~n22080 ;
  assign n22083 = ~n22081 & ~n22082 ;
  assign n22084 = ~n3283 & ~n8272 ;
  assign n22085 = ~n8756 & n22084 ;
  assign n22086 = n3280 & n22085 ;
  assign n22087 = n3283 & ~n8272 ;
  assign n22088 = ~n8756 & n22087 ;
  assign n22089 = ~n3280 & n22088 ;
  assign n22090 = ~n22086 & ~n22089 ;
  assign n22091 = \b[22]  & n9301 ;
  assign n22092 = n9298 & n22091 ;
  assign n22093 = ~\a[39]  & \b[23]  ;
  assign n22094 = n8751 & n22093 ;
  assign n22095 = ~n22092 & ~n22094 ;
  assign n22096 = \b[24]  & n8757 ;
  assign n22097 = \a[39]  & \b[23]  ;
  assign n22098 = n8748 & n22097 ;
  assign n22099 = \a[41]  & ~n22098 ;
  assign n22100 = ~n22096 & n22099 ;
  assign n22101 = n22095 & n22100 ;
  assign n22102 = n22090 & n22101 ;
  assign n22103 = ~n22096 & ~n22098 ;
  assign n22104 = n22095 & n22103 ;
  assign n22105 = n22090 & n22104 ;
  assign n22106 = ~\a[41]  & ~n22105 ;
  assign n22107 = ~n22102 & ~n22106 ;
  assign n22108 = ~n22083 & ~n22107 ;
  assign n22109 = ~n21864 & n22108 ;
  assign n22110 = n22083 & ~n22107 ;
  assign n22111 = n21864 & n22110 ;
  assign n22112 = ~n22109 & ~n22111 ;
  assign n22113 = ~n22083 & n22107 ;
  assign n22114 = n21864 & n22113 ;
  assign n22115 = n22083 & n22107 ;
  assign n22116 = ~n21864 & n22115 ;
  assign n22117 = ~n22114 & ~n22116 ;
  assign n22118 = n22112 & n22117 ;
  assign n22119 = ~n4148 & n7534 ;
  assign n22120 = ~n4146 & n22119 ;
  assign n22121 = \b[25]  & n7973 ;
  assign n22122 = n7970 & n22121 ;
  assign n22123 = ~\a[36]  & \b[26]  ;
  assign n22124 = n7526 & n22123 ;
  assign n22125 = ~n22122 & ~n22124 ;
  assign n22126 = \b[27]  & n7532 ;
  assign n22127 = \a[36]  & \b[26]  ;
  assign n22128 = n17801 & n22127 ;
  assign n22129 = \a[38]  & ~n22128 ;
  assign n22130 = ~n22126 & n22129 ;
  assign n22131 = n22125 & n22130 ;
  assign n22132 = ~n22120 & n22131 ;
  assign n22133 = ~n22126 & ~n22128 ;
  assign n22134 = n22125 & n22133 ;
  assign n22135 = ~n22120 & n22134 ;
  assign n22136 = ~\a[38]  & ~n22135 ;
  assign n22137 = ~n22132 & ~n22136 ;
  assign n22138 = ~n22118 & ~n22137 ;
  assign n22139 = n21862 & n22138 ;
  assign n22140 = n22118 & ~n22137 ;
  assign n22141 = ~n21862 & n22140 ;
  assign n22142 = ~n22139 & ~n22141 ;
  assign n22143 = ~n22118 & n22137 ;
  assign n22144 = ~n21862 & n22143 ;
  assign n22145 = n22118 & n22137 ;
  assign n22146 = n21862 & n22145 ;
  assign n22147 = ~n22144 & ~n22146 ;
  assign n22148 = n22142 & n22147 ;
  assign n22149 = ~n5105 & ~n5952 ;
  assign n22150 = ~n6306 & n22149 ;
  assign n22151 = n5102 & n22150 ;
  assign n22152 = n5105 & ~n5952 ;
  assign n22153 = ~n6306 & n22152 ;
  assign n22154 = ~n5102 & n22153 ;
  assign n22155 = ~n22151 & ~n22154 ;
  assign n22156 = \b[28]  & n6778 ;
  assign n22157 = n6775 & n22156 ;
  assign n22158 = ~\a[33]  & \b[29]  ;
  assign n22159 = n6301 & n22158 ;
  assign n22160 = ~n22157 & ~n22159 ;
  assign n22161 = \b[30]  & n6307 ;
  assign n22162 = \a[33]  & \b[29]  ;
  assign n22163 = n6298 & n22162 ;
  assign n22164 = \a[35]  & ~n22163 ;
  assign n22165 = ~n22161 & n22164 ;
  assign n22166 = n22160 & n22165 ;
  assign n22167 = n22155 & n22166 ;
  assign n22168 = ~n22161 & ~n22163 ;
  assign n22169 = n22160 & n22168 ;
  assign n22170 = n22155 & n22169 ;
  assign n22171 = ~\a[35]  & ~n22170 ;
  assign n22172 = ~n22167 & ~n22171 ;
  assign n22173 = ~n22148 & n22172 ;
  assign n22174 = n21859 & n22173 ;
  assign n22175 = n22148 & n22172 ;
  assign n22176 = ~n21859 & n22175 ;
  assign n22177 = ~n22174 & ~n22176 ;
  assign n22178 = ~n21859 & n22148 ;
  assign n22179 = ~n21433 & ~n22148 ;
  assign n22180 = ~n21858 & n22179 ;
  assign n22181 = ~n22172 & ~n22180 ;
  assign n22182 = ~n22178 & n22181 ;
  assign n22183 = n22177 & ~n22182 ;
  assign n22184 = n20738 & n21463 ;
  assign n22185 = n21468 & ~n22184 ;
  assign n22186 = n20744 & n21468 ;
  assign n22187 = n20431 & n22186 ;
  assign n22188 = ~n22185 & ~n22187 ;
  assign n22189 = n22183 & ~n22188 ;
  assign n22190 = ~n22183 & n22188 ;
  assign n22191 = ~n22189 & ~n22190 ;
  assign n22192 = n5211 & ~n5855 ;
  assign n22193 = ~n5853 & n22192 ;
  assign n22194 = \b[31]  & n5595 ;
  assign n22195 = n5592 & n22194 ;
  assign n22196 = ~\a[30]  & \b[32]  ;
  assign n22197 = n5203 & n22196 ;
  assign n22198 = ~n22195 & ~n22197 ;
  assign n22199 = \b[33]  & n5209 ;
  assign n22200 = \a[30]  & \b[32]  ;
  assign n22201 = n5200 & n22200 ;
  assign n22202 = \a[32]  & ~n22201 ;
  assign n22203 = ~n22199 & n22202 ;
  assign n22204 = n22198 & n22203 ;
  assign n22205 = ~n22193 & n22204 ;
  assign n22206 = ~n22199 & ~n22201 ;
  assign n22207 = n22198 & n22206 ;
  assign n22208 = ~n22193 & n22207 ;
  assign n22209 = ~\a[32]  & ~n22208 ;
  assign n22210 = ~n22205 & ~n22209 ;
  assign n22211 = n22191 & ~n22210 ;
  assign n22212 = ~n22191 & n22210 ;
  assign n22213 = ~n22211 & ~n22212 ;
  assign n22214 = ~n21857 & n22213 ;
  assign n22215 = n4249 & n7337 ;
  assign n22216 = ~n7334 & n22215 ;
  assign n22217 = n4249 & ~n7337 ;
  assign n22218 = ~n6605 & n22217 ;
  assign n22219 = ~n7333 & n22218 ;
  assign n22220 = \b[34]  & n4647 ;
  assign n22221 = n4644 & n22220 ;
  assign n22222 = ~\a[27]  & \b[35]  ;
  assign n22223 = n4241 & n22222 ;
  assign n22224 = ~n22221 & ~n22223 ;
  assign n22225 = \b[36]  & n4247 ;
  assign n22226 = \a[27]  & \b[35]  ;
  assign n22227 = n4238 & n22226 ;
  assign n22228 = \a[29]  & ~n22227 ;
  assign n22229 = ~n22225 & n22228 ;
  assign n22230 = n22224 & n22229 ;
  assign n22231 = ~n22219 & n22230 ;
  assign n22232 = ~n22216 & n22231 ;
  assign n22233 = ~n22225 & ~n22227 ;
  assign n22234 = n22224 & n22233 ;
  assign n22235 = ~n22219 & n22234 ;
  assign n22236 = ~n22216 & n22235 ;
  assign n22237 = ~\a[29]  & ~n22236 ;
  assign n22238 = ~n22232 & ~n22237 ;
  assign n22239 = ~n21497 & ~n22213 ;
  assign n22240 = ~n21856 & n22239 ;
  assign n22241 = ~n22238 & ~n22240 ;
  assign n22242 = ~n22214 & n22241 ;
  assign n22243 = ~n22213 & n22238 ;
  assign n22244 = n21857 & n22243 ;
  assign n22245 = n22213 & n22238 ;
  assign n22246 = ~n21857 & n22245 ;
  assign n22247 = ~n22244 & ~n22246 ;
  assign n22248 = ~n22242 & n22247 ;
  assign n22249 = n3402 & ~n8602 ;
  assign n22250 = ~n8600 & n22249 ;
  assign n22251 = \b[37]  & n3733 ;
  assign n22252 = n3730 & n22251 ;
  assign n22253 = \b[39]  & n3400 ;
  assign n22254 = \a[23]  & \b[38]  ;
  assign n22255 = n3731 & n22254 ;
  assign n22256 = ~\a[24]  & \b[38]  ;
  assign n22257 = n3394 & n22256 ;
  assign n22258 = ~n22255 & ~n22257 ;
  assign n22259 = ~n22253 & n22258 ;
  assign n22260 = ~n22252 & n22259 ;
  assign n22261 = ~n22250 & n22260 ;
  assign n22262 = ~\a[26]  & ~n22261 ;
  assign n22263 = \a[26]  & n22260 ;
  assign n22264 = ~n22250 & n22263 ;
  assign n22265 = ~n22262 & ~n22264 ;
  assign n22266 = ~n22248 & n22265 ;
  assign n22267 = ~n21855 & n22266 ;
  assign n22268 = n22248 & n22265 ;
  assign n22269 = n21855 & n22268 ;
  assign n22270 = ~n22267 & ~n22269 ;
  assign n22271 = ~n22248 & ~n22265 ;
  assign n22272 = n21855 & n22271 ;
  assign n22273 = n22248 & ~n22265 ;
  assign n22274 = ~n21855 & n22273 ;
  assign n22275 = ~n22272 & ~n22274 ;
  assign n22276 = n22270 & n22275 ;
  assign n22277 = ~n21852 & ~n22276 ;
  assign n22278 = ~n21828 & n22277 ;
  assign n22279 = ~n21852 & n22276 ;
  assign n22280 = n21828 & n22279 ;
  assign n22281 = ~n22278 & ~n22280 ;
  assign n22282 = n21852 & ~n22276 ;
  assign n22283 = n21828 & n22282 ;
  assign n22284 = n21852 & n22276 ;
  assign n22285 = ~n21828 & n22284 ;
  assign n22286 = ~n22283 & ~n22285 ;
  assign n22287 = n22281 & n22286 ;
  assign n22288 = ~n21827 & ~n22287 ;
  assign n22289 = n21810 & n22288 ;
  assign n22290 = ~n21827 & n22287 ;
  assign n22291 = ~n21810 & n22290 ;
  assign n22292 = ~n22289 & ~n22291 ;
  assign n22293 = n21827 & ~n22287 ;
  assign n22294 = ~n21810 & n22293 ;
  assign n22295 = n21827 & n22287 ;
  assign n22296 = n21810 & n22295 ;
  assign n22297 = ~n22294 & ~n22296 ;
  assign n22298 = n22292 & n22297 ;
  assign n22299 = ~n21807 & n22298 ;
  assign n22300 = n1467 & n12478 ;
  assign n22301 = ~n12475 & n22300 ;
  assign n22302 = n1467 & ~n12478 ;
  assign n22303 = ~n12433 & n22302 ;
  assign n22304 = ~n12474 & n22303 ;
  assign n22305 = \b[46]  & n1652 ;
  assign n22306 = n1649 & n22305 ;
  assign n22307 = ~\a[15]  & \b[47]  ;
  assign n22308 = n1459 & n22307 ;
  assign n22309 = ~n22306 & ~n22308 ;
  assign n22310 = \b[48]  & n1465 ;
  assign n22311 = \a[15]  & \b[47]  ;
  assign n22312 = n1456 & n22311 ;
  assign n22313 = \a[17]  & ~n22312 ;
  assign n22314 = ~n22310 & n22313 ;
  assign n22315 = n22309 & n22314 ;
  assign n22316 = ~n22304 & n22315 ;
  assign n22317 = ~n22301 & n22316 ;
  assign n22318 = ~n22310 & ~n22312 ;
  assign n22319 = n22309 & n22318 ;
  assign n22320 = ~n22304 & n22319 ;
  assign n22321 = ~n22301 & n22320 ;
  assign n22322 = ~\a[17]  & ~n22321 ;
  assign n22323 = ~n22317 & ~n22322 ;
  assign n22324 = n21575 & ~n22298 ;
  assign n22325 = ~n21806 & n22324 ;
  assign n22326 = ~n22323 & ~n22325 ;
  assign n22327 = ~n22299 & n22326 ;
  assign n22328 = ~n22298 & n22323 ;
  assign n22329 = n21807 & n22328 ;
  assign n22330 = n22298 & n22323 ;
  assign n22331 = ~n21807 & n22330 ;
  assign n22332 = ~n22329 & ~n22331 ;
  assign n22333 = ~n22327 & n22332 ;
  assign n22334 = ~n21805 & ~n22333 ;
  assign n22335 = n21788 & n22334 ;
  assign n22336 = ~n21805 & n22333 ;
  assign n22337 = ~n21788 & n22336 ;
  assign n22338 = ~n22335 & ~n22337 ;
  assign n22339 = n21805 & ~n22333 ;
  assign n22340 = ~n21788 & n22339 ;
  assign n22341 = n21805 & n22333 ;
  assign n22342 = n21788 & n22341 ;
  assign n22343 = ~n22340 & ~n22342 ;
  assign n22344 = n22338 & n22343 ;
  assign n22345 = ~n21785 & n22344 ;
  assign n22346 = ~n21619 & ~n22344 ;
  assign n22347 = ~n21784 & n22346 ;
  assign n22348 = n646 & ~n16398 ;
  assign n22349 = ~n15241 & n22348 ;
  assign n22350 = ~n16404 & n22349 ;
  assign n22351 = n646 & n16398 ;
  assign n22352 = n15241 & n22351 ;
  assign n22353 = n16400 & n22351 ;
  assign n22354 = ~n15239 & n22353 ;
  assign n22355 = ~n22352 & ~n22354 ;
  assign n22356 = ~n22350 & n22355 ;
  assign n22357 = \b[52]  & n796 ;
  assign n22358 = n793 & n22357 ;
  assign n22359 = ~\a[9]  & \b[53]  ;
  assign n22360 = n638 & n22359 ;
  assign n22361 = ~n22358 & ~n22360 ;
  assign n22362 = \b[54]  & n644 ;
  assign n22363 = \a[9]  & \b[53]  ;
  assign n22364 = n635 & n22363 ;
  assign n22365 = \a[11]  & ~n22364 ;
  assign n22366 = ~n22362 & n22365 ;
  assign n22367 = n22361 & n22366 ;
  assign n22368 = n22356 & n22367 ;
  assign n22369 = ~n22362 & ~n22364 ;
  assign n22370 = n22361 & n22369 ;
  assign n22371 = n22356 & n22370 ;
  assign n22372 = ~\a[11]  & ~n22371 ;
  assign n22373 = ~n22368 & ~n22372 ;
  assign n22374 = ~n22347 & ~n22373 ;
  assign n22375 = ~n22345 & n22374 ;
  assign n22376 = ~n22344 & n22373 ;
  assign n22377 = n21785 & n22376 ;
  assign n22378 = n22344 & n22373 ;
  assign n22379 = ~n21785 & n22378 ;
  assign n22380 = ~n22377 & ~n22379 ;
  assign n22381 = ~n22375 & n22380 ;
  assign n22382 = n252 & n20260 ;
  assign n22383 = ~n20257 & n22382 ;
  assign n22384 = n252 & ~n20260 ;
  assign n22385 = ~n19545 & n22384 ;
  assign n22386 = ~n20256 & n22385 ;
  assign n22387 = \b[58]  & n303 ;
  assign n22388 = n300 & n22387 ;
  assign n22389 = ~\a[3]  & \b[59]  ;
  assign n22390 = n244 & n22389 ;
  assign n22391 = ~n22388 & ~n22390 ;
  assign n22392 = \b[60]  & n250 ;
  assign n22393 = \a[3]  & \b[59]  ;
  assign n22394 = n241 & n22393 ;
  assign n22395 = \a[5]  & ~n22394 ;
  assign n22396 = ~n22392 & n22395 ;
  assign n22397 = n22391 & n22396 ;
  assign n22398 = ~n22386 & n22397 ;
  assign n22399 = ~n22383 & n22398 ;
  assign n22400 = ~n22392 & ~n22394 ;
  assign n22401 = n22391 & n22400 ;
  assign n22402 = ~n22386 & n22401 ;
  assign n22403 = ~n22383 & n22402 ;
  assign n22404 = ~\a[5]  & ~n22403 ;
  assign n22405 = ~n22399 & ~n22404 ;
  assign n22406 = n430 & ~n17690 ;
  assign n22407 = ~n17688 & n22406 ;
  assign n22408 = \b[57]  & n428 ;
  assign n22409 = \a[6]  & \b[56]  ;
  assign n22410 = n419 & n22409 ;
  assign n22411 = ~n22408 & ~n22410 ;
  assign n22412 = \b[55]  & n486 ;
  assign n22413 = n483 & n22412 ;
  assign n22414 = ~\a[6]  & \b[56]  ;
  assign n22415 = n422 & n22414 ;
  assign n22416 = ~n22413 & ~n22415 ;
  assign n22417 = n22411 & n22416 ;
  assign n22418 = ~n22407 & n22417 ;
  assign n22419 = ~\a[8]  & ~n22418 ;
  assign n22420 = \a[8]  & n22417 ;
  assign n22421 = ~n22407 & n22420 ;
  assign n22422 = ~n22419 & ~n22421 ;
  assign n22423 = ~n22405 & ~n22422 ;
  assign n22424 = ~n22381 & n22423 ;
  assign n22425 = ~n21783 & n22424 ;
  assign n22426 = ~n22405 & n22422 ;
  assign n22427 = ~n22381 & n22426 ;
  assign n22428 = n21783 & n22427 ;
  assign n22429 = ~n22425 & ~n22428 ;
  assign n22430 = n22381 & n22423 ;
  assign n22431 = n21783 & n22430 ;
  assign n22432 = n22381 & n22426 ;
  assign n22433 = ~n21783 & n22432 ;
  assign n22434 = ~n22431 & ~n22433 ;
  assign n22435 = n22429 & n22434 ;
  assign n22436 = ~n22404 & ~n22422 ;
  assign n22437 = ~n22381 & n22436 ;
  assign n22438 = n21783 & n22437 ;
  assign n22439 = ~n22404 & n22422 ;
  assign n22440 = ~n22381 & n22439 ;
  assign n22441 = ~n21783 & n22440 ;
  assign n22442 = ~n22438 & ~n22441 ;
  assign n22443 = n22381 & n22436 ;
  assign n22444 = ~n21783 & n22443 ;
  assign n22445 = n22381 & n22439 ;
  assign n22446 = n21783 & n22445 ;
  assign n22447 = ~n22444 & ~n22446 ;
  assign n22448 = n22442 & n22447 ;
  assign n22449 = ~n22399 & ~n22448 ;
  assign n22450 = n22435 & ~n22449 ;
  assign n22451 = n21780 & ~n22450 ;
  assign n22452 = ~n21780 & n22435 ;
  assign n22453 = ~n22449 & n22452 ;
  assign n22454 = ~n22451 & ~n22453 ;
  assign n22455 = ~n21695 & ~n21699 ;
  assign n22456 = \b[62]  & ~\b[63]  ;
  assign n22457 = ~\b[62]  & \b[63]  ;
  assign n22458 = ~n22456 & ~n22457 ;
  assign n22459 = ~n22455 & ~n22458 ;
  assign n22460 = ~n21695 & n22458 ;
  assign n22461 = ~n21699 & n22460 ;
  assign n22462 = n134 & ~n22461 ;
  assign n22463 = ~n22459 & n22462 ;
  assign n22464 = \a[0]  & \b[63]  ;
  assign n22465 = n133 & n22464 ;
  assign n22466 = \b[62]  & n141 ;
  assign n22467 = ~\a[1]  & \b[61]  ;
  assign n22468 = n10416 & n22467 ;
  assign n22469 = ~n22466 & ~n22468 ;
  assign n22470 = ~n22465 & n22469 ;
  assign n22471 = \a[2]  & n22470 ;
  assign n22472 = ~n22463 & n22471 ;
  assign n22473 = ~n22463 & n22470 ;
  assign n22474 = ~\a[2]  & ~n22473 ;
  assign n22475 = ~n22472 & ~n22474 ;
  assign n22476 = n21731 & ~n21760 ;
  assign n22477 = n22475 & ~n22476 ;
  assign n22478 = ~n22475 & n22476 ;
  assign n22479 = ~n22477 & ~n22478 ;
  assign n22480 = ~n22454 & ~n22479 ;
  assign n22481 = n22454 & n22479 ;
  assign n22482 = ~n22480 & ~n22481 ;
  assign n22483 = ~n21768 & n22482 ;
  assign n22484 = ~n21772 & n22483 ;
  assign n22485 = ~n21768 & ~n21772 ;
  assign n22486 = ~n22482 & ~n22485 ;
  assign n22487 = ~n22484 & ~n22486 ;
  assign n22488 = ~n22454 & n22478 ;
  assign n22489 = n22475 & n22476 ;
  assign n22490 = n22454 & n22489 ;
  assign n22491 = ~n22488 & ~n22490 ;
  assign n22492 = ~n21768 & n22491 ;
  assign n22493 = ~n21772 & n22492 ;
  assign n22494 = ~n22454 & n22477 ;
  assign n22495 = ~n22475 & ~n22476 ;
  assign n22496 = n22454 & n22495 ;
  assign n22497 = ~n22494 & ~n22496 ;
  assign n22498 = n21783 & n22381 ;
  assign n22499 = ~n22375 & ~n22498 ;
  assign n22500 = ~n21619 & n22338 ;
  assign n22501 = ~n21784 & n22500 ;
  assign n22502 = n22343 & ~n22501 ;
  assign n22503 = n646 & ~n16446 ;
  assign n22504 = ~n16444 & n22503 ;
  assign n22505 = \b[55]  & n644 ;
  assign n22506 = \a[9]  & \b[54]  ;
  assign n22507 = n635 & n22506 ;
  assign n22508 = ~n22505 & ~n22507 ;
  assign n22509 = \b[53]  & n796 ;
  assign n22510 = n793 & n22509 ;
  assign n22511 = ~\a[9]  & \b[54]  ;
  assign n22512 = n638 & n22511 ;
  assign n22513 = ~n22510 & ~n22512 ;
  assign n22514 = n22508 & n22513 ;
  assign n22515 = ~n22504 & n22514 ;
  assign n22516 = ~\a[11]  & ~n22515 ;
  assign n22517 = \a[11]  & n22514 ;
  assign n22518 = ~n22504 & n22517 ;
  assign n22519 = ~n22516 & ~n22518 ;
  assign n22520 = n21788 & n22333 ;
  assign n22521 = ~n22327 & ~n22520 ;
  assign n22522 = n21575 & n22292 ;
  assign n22523 = ~n21806 & n22522 ;
  assign n22524 = n22297 & ~n22523 ;
  assign n22525 = n1467 & ~n13524 ;
  assign n22526 = ~n13522 & n22525 ;
  assign n22527 = \b[49]  & n1465 ;
  assign n22528 = \a[15]  & \b[48]  ;
  assign n22529 = n1456 & n22528 ;
  assign n22530 = ~n22527 & ~n22529 ;
  assign n22531 = \b[47]  & n1652 ;
  assign n22532 = n1649 & n22531 ;
  assign n22533 = ~\a[15]  & \b[48]  ;
  assign n22534 = n1459 & n22533 ;
  assign n22535 = ~n22532 & ~n22534 ;
  assign n22536 = n22530 & n22535 ;
  assign n22537 = ~n22526 & n22536 ;
  assign n22538 = ~\a[17]  & ~n22537 ;
  assign n22539 = \a[17]  & n22536 ;
  assign n22540 = ~n22526 & n22539 ;
  assign n22541 = ~n22538 & ~n22540 ;
  assign n22542 = n21810 & n22287 ;
  assign n22543 = n22281 & ~n22542 ;
  assign n22544 = n1965 & n11906 ;
  assign n22545 = ~n11903 & n22544 ;
  assign n22546 = n1965 & ~n11906 ;
  assign n22547 = ~n11392 & n22546 ;
  assign n22548 = ~n11902 & n22547 ;
  assign n22549 = \b[44]  & n2218 ;
  assign n22550 = n2216 & n22549 ;
  assign n22551 = ~\a[18]  & \b[45]  ;
  assign n22552 = n1957 & n22551 ;
  assign n22553 = ~n22550 & ~n22552 ;
  assign n22554 = \b[46]  & n1963 ;
  assign n22555 = \a[18]  & \b[45]  ;
  assign n22556 = n2210 & n22555 ;
  assign n22557 = \a[20]  & ~n22556 ;
  assign n22558 = ~n22554 & n22557 ;
  assign n22559 = n22553 & n22558 ;
  assign n22560 = ~n22548 & n22559 ;
  assign n22561 = ~n22545 & n22560 ;
  assign n22562 = ~n22554 & ~n22556 ;
  assign n22563 = n22553 & n22562 ;
  assign n22564 = ~n22548 & n22563 ;
  assign n22565 = ~n22545 & n22564 ;
  assign n22566 = ~\a[20]  & ~n22565 ;
  assign n22567 = ~n22561 & ~n22566 ;
  assign n22568 = n2622 & ~n10409 ;
  assign n22569 = ~n10407 & n22568 ;
  assign n22570 = \b[43]  & n2620 ;
  assign n22571 = \a[21]  & \b[42]  ;
  assign n22572 = n20849 & n22571 ;
  assign n22573 = ~n22570 & ~n22572 ;
  assign n22574 = \b[41]  & n2912 ;
  assign n22575 = n2909 & n22574 ;
  assign n22576 = ~\a[21]  & \b[42]  ;
  assign n22577 = n2614 & n22576 ;
  assign n22578 = ~n22575 & ~n22577 ;
  assign n22579 = n22573 & n22578 ;
  assign n22580 = ~n22569 & n22579 ;
  assign n22581 = ~\a[23]  & ~n22580 ;
  assign n22582 = \a[23]  & n22579 ;
  assign n22583 = ~n22569 & n22582 ;
  assign n22584 = ~n22581 & ~n22583 ;
  assign n22585 = ~n21541 & n22275 ;
  assign n22586 = ~n21549 & n22585 ;
  assign n22587 = n22270 & ~n22586 ;
  assign n22588 = n21855 & n22248 ;
  assign n22589 = ~n22242 & ~n22588 ;
  assign n22590 = ~n21497 & ~n22211 ;
  assign n22591 = ~n22212 & ~n22590 ;
  assign n22592 = n21503 & ~n22212 ;
  assign n22593 = n21135 & n22592 ;
  assign n22594 = ~n22591 & ~n22593 ;
  assign n22595 = ~n22182 & ~n22189 ;
  assign n22596 = ~n21433 & n22142 ;
  assign n22597 = ~n21858 & n22596 ;
  assign n22598 = n22147 & ~n22597 ;
  assign n22599 = n21862 & n22118 ;
  assign n22600 = n22112 & ~n22599 ;
  assign n22601 = n21388 & ~n22081 ;
  assign n22602 = ~n21863 & n22601 ;
  assign n22603 = ~n22082 & ~n22602 ;
  assign n22604 = ~n22076 & ~n22078 ;
  assign n22605 = n21366 & n22037 ;
  assign n22606 = ~n21885 & n22605 ;
  assign n22607 = n22042 & ~n22606 ;
  assign n22608 = n21889 & n22015 ;
  assign n22609 = ~n22014 & ~n22608 ;
  assign n22610 = ~n21330 & n21998 ;
  assign n22611 = ~n21332 & n22610 ;
  assign n22612 = n22003 & ~n22611 ;
  assign n22613 = n21917 & n21969 ;
  assign n22614 = ~n21968 & ~n22613 ;
  assign n22615 = ~n21961 & ~n21964 ;
  assign n22616 = n222 & n20521 ;
  assign n22617 = \b[2]  & n21315 ;
  assign n22618 = n21312 & n22617 ;
  assign n22619 = \b[4]  & n20519 ;
  assign n22620 = \a[59]  & \b[3]  ;
  assign n22621 = n21313 & n22620 ;
  assign n22622 = ~\a[60]  & \b[3]  ;
  assign n22623 = n20513 & n22622 ;
  assign n22624 = ~n22621 & ~n22623 ;
  assign n22625 = ~n22619 & n22624 ;
  assign n22626 = ~n22618 & n22625 ;
  assign n22627 = ~n22616 & n22626 ;
  assign n22628 = ~\a[62]  & ~n22627 ;
  assign n22629 = \b[1]  & n21958 ;
  assign n22630 = \b[0]  & n21957 ;
  assign n22631 = ~n22629 & ~n22630 ;
  assign n22632 = \a[62]  & ~n22618 ;
  assign n22633 = n22625 & n22632 ;
  assign n22634 = ~n22616 & n22633 ;
  assign n22635 = n22631 & ~n22634 ;
  assign n22636 = ~n22628 & n22635 ;
  assign n22637 = \a[62]  & ~\a[63]  ;
  assign n22638 = \b[1]  & n22637 ;
  assign n22639 = ~n22630 & ~n22638 ;
  assign n22640 = ~n22618 & ~n22639 ;
  assign n22641 = n22625 & n22640 ;
  assign n22642 = ~n22616 & n22641 ;
  assign n22643 = ~\a[62]  & \a[63]  ;
  assign n22644 = \b[1]  & n22643 ;
  assign n22645 = ~n22627 & n22644 ;
  assign n22646 = ~n22642 & ~n22645 ;
  assign n22647 = ~n22636 & n22646 ;
  assign n22648 = n22615 & n22647 ;
  assign n22649 = ~n22615 & ~n22647 ;
  assign n22650 = ~n22648 & ~n22649 ;
  assign n22651 = ~n380 & n18516 ;
  assign n22652 = ~n322 & n18516 ;
  assign n22653 = ~n326 & n22652 ;
  assign n22654 = ~n22651 & ~n22653 ;
  assign n22655 = ~n383 & ~n22654 ;
  assign n22656 = \b[5]  & n19183 ;
  assign n22657 = n19180 & n22656 ;
  assign n22658 = \b[7]  & n18514 ;
  assign n22659 = \a[56]  & \b[6]  ;
  assign n22660 = n19181 & n22659 ;
  assign n22661 = ~\a[57]  & \b[6]  ;
  assign n22662 = n18508 & n22661 ;
  assign n22663 = ~n22660 & ~n22662 ;
  assign n22664 = ~n22658 & n22663 ;
  assign n22665 = ~n22657 & n22664 ;
  assign n22666 = ~\a[59]  & n22665 ;
  assign n22667 = ~n22655 & n22666 ;
  assign n22668 = \a[59]  & ~n22665 ;
  assign n22669 = \a[59]  & ~n383 ;
  assign n22670 = ~n22654 & n22669 ;
  assign n22671 = ~n22668 & ~n22670 ;
  assign n22672 = ~n22667 & n22671 ;
  assign n22673 = n22650 & ~n22672 ;
  assign n22674 = ~n22650 & n22672 ;
  assign n22675 = ~n22673 & ~n22674 ;
  assign n22676 = n685 & n16655 ;
  assign n22677 = ~n682 & n22676 ;
  assign n22678 = n11610 & n16655 ;
  assign n22679 = ~n681 & n22678 ;
  assign n22680 = \b[8]  & n17308 ;
  assign n22681 = n17305 & n22680 ;
  assign n22682 = ~\a[54]  & \b[9]  ;
  assign n22683 = n16647 & n22682 ;
  assign n22684 = ~n22681 & ~n22683 ;
  assign n22685 = \b[10]  & n16653 ;
  assign n22686 = \a[54]  & \b[9]  ;
  assign n22687 = n16644 & n22686 ;
  assign n22688 = \a[56]  & ~n22687 ;
  assign n22689 = ~n22685 & n22688 ;
  assign n22690 = n22684 & n22689 ;
  assign n22691 = ~n22679 & n22690 ;
  assign n22692 = ~n22677 & n22691 ;
  assign n22693 = ~n22685 & ~n22687 ;
  assign n22694 = n22684 & n22693 ;
  assign n22695 = ~n22679 & n22694 ;
  assign n22696 = ~n22677 & n22695 ;
  assign n22697 = ~\a[56]  & ~n22696 ;
  assign n22698 = ~n22692 & ~n22697 ;
  assign n22699 = ~n22675 & ~n22698 ;
  assign n22700 = ~n22614 & n22699 ;
  assign n22701 = n22675 & ~n22698 ;
  assign n22702 = n22614 & n22701 ;
  assign n22703 = ~n22700 & ~n22702 ;
  assign n22704 = ~n22675 & n22698 ;
  assign n22705 = n22614 & n22704 ;
  assign n22706 = n22675 & n22698 ;
  assign n22707 = ~n22614 & n22706 ;
  assign n22708 = ~n22705 & ~n22707 ;
  assign n22709 = n22703 & n22708 ;
  assign n22710 = ~n948 & n14793 ;
  assign n22711 = ~n908 & n14793 ;
  assign n22712 = ~n912 & n22711 ;
  assign n22713 = ~n22710 & ~n22712 ;
  assign n22714 = ~n951 & ~n22713 ;
  assign n22715 = \b[11]  & n15517 ;
  assign n22716 = n15514 & n22715 ;
  assign n22717 = ~\a[51]  & \b[12]  ;
  assign n22718 = n14785 & n22717 ;
  assign n22719 = ~n22716 & ~n22718 ;
  assign n22720 = \b[13]  & n14791 ;
  assign n22721 = \a[51]  & \b[12]  ;
  assign n22722 = n14782 & n22721 ;
  assign n22723 = \a[53]  & ~n22722 ;
  assign n22724 = ~n22720 & n22723 ;
  assign n22725 = n22719 & n22724 ;
  assign n22726 = ~n22714 & n22725 ;
  assign n22727 = ~n22720 & ~n22722 ;
  assign n22728 = n22719 & n22727 ;
  assign n22729 = ~\a[53]  & ~n22728 ;
  assign n22730 = ~\a[53]  & ~n951 ;
  assign n22731 = ~n22713 & n22730 ;
  assign n22732 = ~n22729 & ~n22731 ;
  assign n22733 = ~n22726 & n22732 ;
  assign n22734 = ~n22709 & n22733 ;
  assign n22735 = ~n22612 & n22734 ;
  assign n22736 = n22709 & n22733 ;
  assign n22737 = n22612 & n22736 ;
  assign n22738 = ~n22735 & ~n22737 ;
  assign n22739 = ~n22709 & ~n22733 ;
  assign n22740 = n22612 & n22739 ;
  assign n22741 = n22709 & ~n22733 ;
  assign n22742 = ~n22612 & n22741 ;
  assign n22743 = ~n22740 & ~n22742 ;
  assign n22744 = n22738 & n22743 ;
  assign n22745 = n1512 & n13125 ;
  assign n22746 = ~n1509 & n22745 ;
  assign n22747 = ~n1512 & n13125 ;
  assign n22748 = ~n1228 & n22747 ;
  assign n22749 = ~n1508 & n22748 ;
  assign n22750 = \b[14]  & n13794 ;
  assign n22751 = n13792 & n22750 ;
  assign n22752 = ~\a[48]  & \b[15]  ;
  assign n22753 = n13117 & n22752 ;
  assign n22754 = ~n22751 & ~n22753 ;
  assign n22755 = \b[16]  & n13123 ;
  assign n22756 = \a[48]  & \b[15]  ;
  assign n22757 = n13786 & n22756 ;
  assign n22758 = \a[50]  & ~n22757 ;
  assign n22759 = ~n22755 & n22758 ;
  assign n22760 = n22754 & n22759 ;
  assign n22761 = ~n22749 & n22760 ;
  assign n22762 = ~n22746 & n22761 ;
  assign n22763 = ~n22755 & ~n22757 ;
  assign n22764 = n22754 & n22763 ;
  assign n22765 = ~n22749 & n22764 ;
  assign n22766 = ~n22746 & n22765 ;
  assign n22767 = ~\a[50]  & ~n22766 ;
  assign n22768 = ~n22762 & ~n22767 ;
  assign n22769 = ~n22744 & ~n22768 ;
  assign n22770 = ~n22609 & n22769 ;
  assign n22771 = n22744 & ~n22768 ;
  assign n22772 = n22609 & n22771 ;
  assign n22773 = ~n22770 & ~n22772 ;
  assign n22774 = ~n22609 & ~n22744 ;
  assign n22775 = ~n22014 & n22744 ;
  assign n22776 = ~n22608 & n22775 ;
  assign n22777 = n22768 & ~n22776 ;
  assign n22778 = ~n22774 & n22777 ;
  assign n22779 = n22773 & ~n22778 ;
  assign n22780 = ~n2076 & n11572 ;
  assign n22781 = ~n1874 & n11572 ;
  assign n22782 = ~n1878 & n22781 ;
  assign n22783 = ~n22780 & ~n22782 ;
  assign n22784 = ~n2079 & ~n22783 ;
  assign n22785 = \b[17]  & n12159 ;
  assign n22786 = n12156 & n22785 ;
  assign n22787 = ~\a[45]  & \b[18]  ;
  assign n22788 = n11564 & n22787 ;
  assign n22789 = ~n22786 & ~n22788 ;
  assign n22790 = \b[19]  & n11570 ;
  assign n22791 = \a[45]  & \b[18]  ;
  assign n22792 = n11561 & n22791 ;
  assign n22793 = \a[47]  & ~n22792 ;
  assign n22794 = ~n22790 & n22793 ;
  assign n22795 = n22789 & n22794 ;
  assign n22796 = ~n22784 & n22795 ;
  assign n22797 = ~n22790 & ~n22792 ;
  assign n22798 = n22789 & n22797 ;
  assign n22799 = ~\a[47]  & ~n22798 ;
  assign n22800 = ~\a[47]  & ~n2079 ;
  assign n22801 = ~n22783 & n22800 ;
  assign n22802 = ~n22799 & ~n22801 ;
  assign n22803 = ~n22796 & n22802 ;
  assign n22804 = ~n22779 & n22803 ;
  assign n22805 = ~n22607 & n22804 ;
  assign n22806 = n22779 & n22803 ;
  assign n22807 = n22607 & n22806 ;
  assign n22808 = ~n22805 & ~n22807 ;
  assign n22809 = ~n22779 & ~n22803 ;
  assign n22810 = n22607 & n22809 ;
  assign n22811 = n22779 & ~n22803 ;
  assign n22812 = ~n22607 & n22811 ;
  assign n22813 = ~n22810 & ~n22812 ;
  assign n22814 = n22808 & n22813 ;
  assign n22815 = n2768 & n10082 ;
  assign n22816 = ~n2765 & n22815 ;
  assign n22817 = ~n2768 & n10082 ;
  assign n22818 = ~n2518 & n22817 ;
  assign n22819 = ~n2764 & n22818 ;
  assign n22820 = \b[20]  & n10681 ;
  assign n22821 = n10678 & n22820 ;
  assign n22822 = \b[22]  & n10080 ;
  assign n22823 = \a[42]  & \b[21]  ;
  assign n22824 = n10071 & n22823 ;
  assign n22825 = ~\a[42]  & \b[21]  ;
  assign n22826 = n10074 & n22825 ;
  assign n22827 = ~n22824 & ~n22826 ;
  assign n22828 = ~n22822 & n22827 ;
  assign n22829 = ~n22821 & n22828 ;
  assign n22830 = ~n22819 & n22829 ;
  assign n22831 = ~n22816 & n22830 ;
  assign n22832 = ~\a[44]  & ~n22831 ;
  assign n22833 = \a[44]  & n22829 ;
  assign n22834 = ~n22819 & n22833 ;
  assign n22835 = ~n22816 & n22834 ;
  assign n22836 = ~n22832 & ~n22835 ;
  assign n22837 = ~n22814 & ~n22836 ;
  assign n22838 = ~n22604 & n22837 ;
  assign n22839 = n22814 & ~n22836 ;
  assign n22840 = n22604 & n22839 ;
  assign n22841 = ~n22838 & ~n22840 ;
  assign n22842 = n22814 & n22836 ;
  assign n22843 = ~n22604 & n22842 ;
  assign n22844 = ~n22814 & n22836 ;
  assign n22845 = n22604 & n22844 ;
  assign n22846 = ~n22843 & ~n22845 ;
  assign n22847 = n22841 & n22846 ;
  assign n22848 = ~n3564 & n8759 ;
  assign n22849 = ~n3282 & n8759 ;
  assign n22850 = ~n3560 & n22849 ;
  assign n22851 = ~n22848 & ~n22850 ;
  assign n22852 = ~n3567 & ~n22851 ;
  assign n22853 = \b[23]  & n9301 ;
  assign n22854 = n9298 & n22853 ;
  assign n22855 = ~\a[39]  & \b[24]  ;
  assign n22856 = n8751 & n22855 ;
  assign n22857 = ~n22854 & ~n22856 ;
  assign n22858 = \b[25]  & n8757 ;
  assign n22859 = \a[39]  & \b[24]  ;
  assign n22860 = n8748 & n22859 ;
  assign n22861 = \a[41]  & ~n22860 ;
  assign n22862 = ~n22858 & n22861 ;
  assign n22863 = n22857 & n22862 ;
  assign n22864 = ~n22852 & n22863 ;
  assign n22865 = ~n22858 & ~n22860 ;
  assign n22866 = n22857 & n22865 ;
  assign n22867 = ~\a[41]  & ~n22866 ;
  assign n22868 = ~\a[41]  & ~n3567 ;
  assign n22869 = ~n22851 & n22868 ;
  assign n22870 = ~n22867 & ~n22869 ;
  assign n22871 = ~n22864 & n22870 ;
  assign n22872 = ~n22847 & ~n22871 ;
  assign n22873 = n22603 & n22872 ;
  assign n22874 = n22847 & ~n22871 ;
  assign n22875 = ~n22603 & n22874 ;
  assign n22876 = ~n22873 & ~n22875 ;
  assign n22877 = ~n22847 & n22871 ;
  assign n22878 = ~n22603 & n22877 ;
  assign n22879 = n22847 & n22871 ;
  assign n22880 = n22603 & n22879 ;
  assign n22881 = ~n22878 & ~n22880 ;
  assign n22882 = n22876 & n22881 ;
  assign n22883 = ~n22600 & n22882 ;
  assign n22884 = n22112 & ~n22882 ;
  assign n22885 = ~n22599 & n22884 ;
  assign n22886 = n4456 & n7534 ;
  assign n22887 = ~n18723 & n22886 ;
  assign n22888 = n7534 & n16805 ;
  assign n22889 = ~n4452 & n22888 ;
  assign n22890 = \b[26]  & n7973 ;
  assign n22891 = n7970 & n22890 ;
  assign n22892 = ~\a[36]  & \b[27]  ;
  assign n22893 = n7526 & n22892 ;
  assign n22894 = ~n22891 & ~n22893 ;
  assign n22895 = \b[28]  & n7532 ;
  assign n22896 = \a[36]  & \b[27]  ;
  assign n22897 = n17801 & n22896 ;
  assign n22898 = \a[38]  & ~n22897 ;
  assign n22899 = ~n22895 & n22898 ;
  assign n22900 = n22894 & n22899 ;
  assign n22901 = ~n22889 & n22900 ;
  assign n22902 = ~n22887 & n22901 ;
  assign n22903 = ~n22895 & ~n22897 ;
  assign n22904 = n22894 & n22903 ;
  assign n22905 = ~n22889 & n22904 ;
  assign n22906 = ~n22887 & n22905 ;
  assign n22907 = ~\a[38]  & ~n22906 ;
  assign n22908 = ~n22902 & ~n22907 ;
  assign n22909 = ~n22885 & ~n22908 ;
  assign n22910 = ~n22883 & n22909 ;
  assign n22911 = ~n22882 & n22908 ;
  assign n22912 = n22600 & n22911 ;
  assign n22913 = n22882 & n22908 ;
  assign n22914 = ~n22600 & n22913 ;
  assign n22915 = ~n22912 & ~n22914 ;
  assign n22916 = ~n22910 & n22915 ;
  assign n22917 = ~n5462 & n6309 ;
  assign n22918 = ~n5460 & n22917 ;
  assign n22919 = \b[31]  & n6307 ;
  assign n22920 = \a[33]  & \b[30]  ;
  assign n22921 = n6298 & n22920 ;
  assign n22922 = ~n22919 & ~n22921 ;
  assign n22923 = \b[29]  & n6778 ;
  assign n22924 = n6775 & n22923 ;
  assign n22925 = ~\a[33]  & \b[30]  ;
  assign n22926 = n6301 & n22925 ;
  assign n22927 = ~n22924 & ~n22926 ;
  assign n22928 = n22922 & n22927 ;
  assign n22929 = ~n22918 & n22928 ;
  assign n22930 = ~\a[35]  & ~n22929 ;
  assign n22931 = \a[35]  & n22928 ;
  assign n22932 = ~n22918 & n22931 ;
  assign n22933 = ~n22930 & ~n22932 ;
  assign n22934 = ~n22916 & n22933 ;
  assign n22935 = ~n22598 & n22934 ;
  assign n22936 = n22916 & n22933 ;
  assign n22937 = n22598 & n22936 ;
  assign n22938 = ~n22935 & ~n22937 ;
  assign n22939 = ~n22916 & ~n22933 ;
  assign n22940 = n22598 & n22939 ;
  assign n22941 = n22916 & ~n22933 ;
  assign n22942 = ~n22598 & n22941 ;
  assign n22943 = ~n22940 & ~n22942 ;
  assign n22944 = n22938 & n22943 ;
  assign n22945 = n5211 & n6565 ;
  assign n22946 = ~n6562 & n22945 ;
  assign n22947 = ~n5850 & ~n6565 ;
  assign n22948 = n5211 & n22947 ;
  assign n22949 = ~n6561 & n22948 ;
  assign n22950 = \b[32]  & n5595 ;
  assign n22951 = n5592 & n22950 ;
  assign n22952 = ~\a[30]  & \b[33]  ;
  assign n22953 = n5203 & n22952 ;
  assign n22954 = ~n22951 & ~n22953 ;
  assign n22955 = \b[34]  & n5209 ;
  assign n22956 = \a[30]  & \b[33]  ;
  assign n22957 = n5200 & n22956 ;
  assign n22958 = \a[32]  & ~n22957 ;
  assign n22959 = ~n22955 & n22958 ;
  assign n22960 = n22954 & n22959 ;
  assign n22961 = ~n22949 & n22960 ;
  assign n22962 = ~n22946 & n22961 ;
  assign n22963 = ~n22955 & ~n22957 ;
  assign n22964 = n22954 & n22963 ;
  assign n22965 = ~n22949 & n22964 ;
  assign n22966 = ~n22946 & n22965 ;
  assign n22967 = ~\a[32]  & ~n22966 ;
  assign n22968 = ~n22962 & ~n22967 ;
  assign n22969 = ~n22944 & ~n22968 ;
  assign n22970 = ~n22595 & n22969 ;
  assign n22971 = n22944 & ~n22968 ;
  assign n22972 = n22595 & n22971 ;
  assign n22973 = ~n22970 & ~n22972 ;
  assign n22974 = n22944 & n22968 ;
  assign n22975 = ~n22595 & n22974 ;
  assign n22976 = ~n22944 & n22968 ;
  assign n22977 = n22595 & n22976 ;
  assign n22978 = ~n22975 & ~n22977 ;
  assign n22979 = n22973 & n22978 ;
  assign n22980 = n4249 & ~n7761 ;
  assign n22981 = ~n7759 & n22980 ;
  assign n22982 = \b[37]  & n4247 ;
  assign n22983 = \a[27]  & \b[36]  ;
  assign n22984 = n4238 & n22983 ;
  assign n22985 = ~n22982 & ~n22984 ;
  assign n22986 = \b[35]  & n4647 ;
  assign n22987 = n4644 & n22986 ;
  assign n22988 = ~\a[27]  & \b[36]  ;
  assign n22989 = n4241 & n22988 ;
  assign n22990 = ~n22987 & ~n22989 ;
  assign n22991 = n22985 & n22990 ;
  assign n22992 = ~n22981 & n22991 ;
  assign n22993 = ~\a[29]  & ~n22992 ;
  assign n22994 = \a[29]  & n22991 ;
  assign n22995 = ~n22981 & n22994 ;
  assign n22996 = ~n22993 & ~n22995 ;
  assign n22997 = ~n22979 & ~n22996 ;
  assign n22998 = ~n22594 & n22997 ;
  assign n22999 = n22979 & ~n22996 ;
  assign n23000 = n22594 & n22999 ;
  assign n23001 = ~n22998 & ~n23000 ;
  assign n23002 = ~n22979 & n22996 ;
  assign n23003 = n22594 & n23002 ;
  assign n23004 = n22979 & n22996 ;
  assign n23005 = ~n22594 & n23004 ;
  assign n23006 = ~n23003 & ~n23005 ;
  assign n23007 = n23001 & n23006 ;
  assign n23008 = ~n22589 & n23007 ;
  assign n23009 = ~n22242 & ~n23007 ;
  assign n23010 = ~n22588 & n23009 ;
  assign n23011 = n3402 & n9044 ;
  assign n23012 = ~n9041 & n23011 ;
  assign n23013 = n3402 & ~n9044 ;
  assign n23014 = ~n8597 & n23013 ;
  assign n23015 = ~n9040 & n23014 ;
  assign n23016 = \b[38]  & n3733 ;
  assign n23017 = n3730 & n23016 ;
  assign n23018 = ~\a[24]  & \b[39]  ;
  assign n23019 = n3394 & n23018 ;
  assign n23020 = ~n23017 & ~n23019 ;
  assign n23021 = \b[40]  & n3400 ;
  assign n23022 = \a[24]  & \b[39]  ;
  assign n23023 = n3391 & n23022 ;
  assign n23024 = \a[26]  & ~n23023 ;
  assign n23025 = ~n23021 & n23024 ;
  assign n23026 = n23020 & n23025 ;
  assign n23027 = ~n23015 & n23026 ;
  assign n23028 = ~n23012 & n23027 ;
  assign n23029 = ~n23021 & ~n23023 ;
  assign n23030 = n23020 & n23029 ;
  assign n23031 = ~n23015 & n23030 ;
  assign n23032 = ~n23012 & n23031 ;
  assign n23033 = ~\a[26]  & ~n23032 ;
  assign n23034 = ~n23028 & ~n23033 ;
  assign n23035 = ~n23010 & ~n23034 ;
  assign n23036 = ~n23008 & n23035 ;
  assign n23037 = ~n23007 & n23034 ;
  assign n23038 = n22589 & n23037 ;
  assign n23039 = n23007 & n23034 ;
  assign n23040 = ~n22589 & n23039 ;
  assign n23041 = ~n23038 & ~n23040 ;
  assign n23042 = ~n23036 & n23041 ;
  assign n23043 = n22587 & n23042 ;
  assign n23044 = ~n22587 & ~n23042 ;
  assign n23045 = ~n23043 & ~n23044 ;
  assign n23046 = ~n22584 & n23045 ;
  assign n23047 = n22584 & ~n23045 ;
  assign n23048 = ~n23046 & ~n23047 ;
  assign n23049 = ~n22567 & ~n23048 ;
  assign n23050 = ~n22543 & n23049 ;
  assign n23051 = ~n22567 & n23048 ;
  assign n23052 = n22543 & n23051 ;
  assign n23053 = ~n23050 & ~n23052 ;
  assign n23054 = n22567 & ~n23048 ;
  assign n23055 = n22543 & n23054 ;
  assign n23056 = n22567 & n23048 ;
  assign n23057 = ~n22543 & n23056 ;
  assign n23058 = ~n23055 & ~n23057 ;
  assign n23059 = n23053 & n23058 ;
  assign n23060 = ~n22541 & ~n23059 ;
  assign n23061 = n22524 & n23060 ;
  assign n23062 = ~n22541 & n23059 ;
  assign n23063 = ~n22524 & n23062 ;
  assign n23064 = ~n23061 & ~n23063 ;
  assign n23065 = n22541 & ~n23059 ;
  assign n23066 = ~n22524 & n23065 ;
  assign n23067 = n22541 & n23059 ;
  assign n23068 = n22524 & n23067 ;
  assign n23069 = ~n23066 & ~n23068 ;
  assign n23070 = n23064 & n23069 ;
  assign n23071 = ~n22521 & n23070 ;
  assign n23072 = ~n847 & ~n14093 ;
  assign n23073 = ~n15201 & n23072 ;
  assign n23074 = ~n15197 & n23073 ;
  assign n23075 = ~n996 & n23074 ;
  assign n23076 = n999 & n15201 ;
  assign n23077 = ~n15198 & n23076 ;
  assign n23078 = ~n23075 & ~n23077 ;
  assign n23079 = \b[50]  & n1182 ;
  assign n23080 = n1179 & n23079 ;
  assign n23081 = \b[52]  & n997 ;
  assign n23082 = \a[11]  & \b[51]  ;
  assign n23083 = n1180 & n23082 ;
  assign n23084 = ~\a[12]  & \b[51]  ;
  assign n23085 = n7674 & n23084 ;
  assign n23086 = ~n23083 & ~n23085 ;
  assign n23087 = ~n23081 & n23086 ;
  assign n23088 = ~n23080 & n23087 ;
  assign n23089 = n23078 & n23088 ;
  assign n23090 = ~\a[14]  & ~n23089 ;
  assign n23091 = \a[14]  & n23088 ;
  assign n23092 = n23078 & n23091 ;
  assign n23093 = ~n23090 & ~n23092 ;
  assign n23094 = ~n22327 & ~n23070 ;
  assign n23095 = ~n22520 & n23094 ;
  assign n23096 = ~n23093 & ~n23095 ;
  assign n23097 = ~n23071 & n23096 ;
  assign n23098 = ~n23070 & n23093 ;
  assign n23099 = n22521 & n23098 ;
  assign n23100 = n23070 & n23093 ;
  assign n23101 = ~n22521 & n23100 ;
  assign n23102 = ~n23099 & ~n23101 ;
  assign n23103 = ~n23097 & n23102 ;
  assign n23104 = ~n22519 & ~n23103 ;
  assign n23105 = n22502 & n23104 ;
  assign n23106 = ~n22519 & n23103 ;
  assign n23107 = ~n22502 & n23106 ;
  assign n23108 = ~n23105 & ~n23107 ;
  assign n23109 = n22519 & ~n23103 ;
  assign n23110 = ~n22502 & n23109 ;
  assign n23111 = n22519 & n23103 ;
  assign n23112 = n22502 & n23111 ;
  assign n23113 = ~n23110 & ~n23112 ;
  assign n23114 = n23108 & n23113 ;
  assign n23115 = ~n22499 & n23114 ;
  assign n23116 = ~n22375 & ~n23114 ;
  assign n23117 = ~n22498 & n23116 ;
  assign n23118 = ~n359 & ~n17685 ;
  assign n23119 = ~n18940 & n23118 ;
  assign n23120 = ~n18936 & n23119 ;
  assign n23121 = ~n427 & n23120 ;
  assign n23122 = n430 & n18940 ;
  assign n23123 = ~n18937 & n23122 ;
  assign n23124 = ~n23121 & ~n23123 ;
  assign n23125 = \b[56]  & n486 ;
  assign n23126 = n483 & n23125 ;
  assign n23127 = ~\a[6]  & \b[57]  ;
  assign n23128 = n422 & n23127 ;
  assign n23129 = ~n23126 & ~n23128 ;
  assign n23130 = \b[58]  & n428 ;
  assign n23131 = \a[6]  & \b[57]  ;
  assign n23132 = n419 & n23131 ;
  assign n23133 = \a[8]  & ~n23132 ;
  assign n23134 = ~n23130 & n23133 ;
  assign n23135 = n23129 & n23134 ;
  assign n23136 = n23124 & n23135 ;
  assign n23137 = ~n23130 & ~n23132 ;
  assign n23138 = n23129 & n23137 ;
  assign n23139 = n23124 & n23138 ;
  assign n23140 = ~\a[8]  & ~n23139 ;
  assign n23141 = ~n23136 & ~n23140 ;
  assign n23142 = ~n23117 & ~n23141 ;
  assign n23143 = ~n23115 & n23142 ;
  assign n23144 = ~n23114 & n23141 ;
  assign n23145 = n22499 & n23144 ;
  assign n23146 = n23114 & n23141 ;
  assign n23147 = ~n22499 & n23146 ;
  assign n23148 = ~n23145 & ~n23147 ;
  assign n23149 = ~n23143 & n23148 ;
  assign n23150 = ~n22381 & n22422 ;
  assign n23151 = ~n21783 & n23150 ;
  assign n23152 = n22381 & n22422 ;
  assign n23153 = n21783 & n23152 ;
  assign n23154 = ~n23151 & ~n23153 ;
  assign n23155 = ~n22381 & ~n22422 ;
  assign n23156 = n21783 & n23155 ;
  assign n23157 = n22381 & ~n22422 ;
  assign n23158 = ~n21783 & n23157 ;
  assign n23159 = ~n23156 & ~n23158 ;
  assign n23160 = n22405 & n23159 ;
  assign n23161 = n23154 & ~n23160 ;
  assign n23162 = ~\a[1]  & \b[62]  ;
  assign n23163 = n10416 & n23162 ;
  assign n23164 = \b[63]  & n141 ;
  assign n23165 = ~n23163 & ~n23164 ;
  assign n23166 = ~\a[2]  & ~n23165 ;
  assign n23167 = \b[60]  & \b[62]  ;
  assign n23168 = ~n20965 & n23167 ;
  assign n23169 = ~\b[60]  & ~\b[62]  ;
  assign n23170 = ~n20259 & n23169 ;
  assign n23171 = ~n20964 & n23170 ;
  assign n23172 = n21696 & ~n23171 ;
  assign n23173 = ~n23168 & n23172 ;
  assign n23174 = n134 & ~n22458 ;
  assign n23175 = ~\a[2]  & n23174 ;
  assign n23176 = ~n23173 & n23175 ;
  assign n23177 = ~n23166 & ~n23176 ;
  assign n23178 = ~n23173 & n23174 ;
  assign n23179 = \a[2]  & n23165 ;
  assign n23180 = ~n23178 & n23179 ;
  assign n23181 = n23177 & ~n23180 ;
  assign n23182 = n252 & ~n20971 ;
  assign n23183 = ~n20969 & n23182 ;
  assign n23184 = \b[61]  & n250 ;
  assign n23185 = \a[3]  & \b[60]  ;
  assign n23186 = n241 & n23185 ;
  assign n23187 = ~\a[3]  & \b[60]  ;
  assign n23188 = n244 & n23187 ;
  assign n23189 = ~n23186 & ~n23188 ;
  assign n23190 = ~n23184 & n23189 ;
  assign n23191 = \b[59]  & n303 ;
  assign n23192 = n300 & n23191 ;
  assign n23193 = \a[5]  & ~n23192 ;
  assign n23194 = n23190 & n23193 ;
  assign n23195 = ~n23183 & n23194 ;
  assign n23196 = n23190 & ~n23192 ;
  assign n23197 = ~n23183 & n23196 ;
  assign n23198 = ~\a[5]  & ~n23197 ;
  assign n23199 = ~n23195 & ~n23198 ;
  assign n23200 = ~n23181 & ~n23199 ;
  assign n23201 = ~n23161 & n23200 ;
  assign n23202 = ~n23149 & n23201 ;
  assign n23203 = ~n23181 & n23199 ;
  assign n23204 = n23161 & n23203 ;
  assign n23205 = ~n23149 & n23204 ;
  assign n23206 = ~n23202 & ~n23205 ;
  assign n23207 = ~n23161 & n23203 ;
  assign n23208 = n23149 & n23207 ;
  assign n23209 = n23161 & n23200 ;
  assign n23210 = n23149 & n23209 ;
  assign n23211 = ~n23208 & ~n23210 ;
  assign n23212 = n23206 & n23211 ;
  assign n23213 = n23181 & n23199 ;
  assign n23214 = ~n23161 & n23213 ;
  assign n23215 = ~n23149 & n23214 ;
  assign n23216 = n23181 & ~n23199 ;
  assign n23217 = n23161 & n23216 ;
  assign n23218 = ~n23149 & n23217 ;
  assign n23219 = ~n23215 & ~n23218 ;
  assign n23220 = ~n23161 & n23216 ;
  assign n23221 = n23149 & n23220 ;
  assign n23222 = n23161 & n23213 ;
  assign n23223 = n23149 & n23222 ;
  assign n23224 = ~n23221 & ~n23223 ;
  assign n23225 = n23219 & n23224 ;
  assign n23226 = n23212 & n23225 ;
  assign n23227 = ~n22453 & n22475 ;
  assign n23228 = ~n22451 & ~n23227 ;
  assign n23229 = n23226 & n23228 ;
  assign n23230 = ~n23226 & ~n23228 ;
  assign n23231 = ~n23229 & ~n23230 ;
  assign n23232 = n22497 & n23231 ;
  assign n23233 = ~n22493 & n23232 ;
  assign n23234 = ~n22493 & n22497 ;
  assign n23235 = ~n23231 & ~n23234 ;
  assign n23236 = ~n23233 & ~n23235 ;
  assign n23237 = ~n23141 & ~n23199 ;
  assign n23238 = ~n23114 & n23237 ;
  assign n23239 = n22499 & n23238 ;
  assign n23240 = n23141 & ~n23199 ;
  assign n23241 = ~n23114 & n23240 ;
  assign n23242 = ~n22499 & n23241 ;
  assign n23243 = ~n23239 & ~n23242 ;
  assign n23244 = n23114 & n23237 ;
  assign n23245 = ~n22499 & n23244 ;
  assign n23246 = n23114 & n23240 ;
  assign n23247 = n22499 & n23246 ;
  assign n23248 = ~n23245 & ~n23247 ;
  assign n23249 = n23243 & n23248 ;
  assign n23250 = ~n23141 & n23199 ;
  assign n23251 = ~n23114 & n23250 ;
  assign n23252 = ~n22499 & n23251 ;
  assign n23253 = n23141 & n23199 ;
  assign n23254 = ~n23114 & n23253 ;
  assign n23255 = n22499 & n23254 ;
  assign n23256 = ~n23252 & ~n23255 ;
  assign n23257 = n23114 & n23250 ;
  assign n23258 = n22499 & n23257 ;
  assign n23259 = n23114 & n23253 ;
  assign n23260 = ~n22499 & n23259 ;
  assign n23261 = ~n23258 & ~n23260 ;
  assign n23262 = n23256 & n23261 ;
  assign n23263 = n23161 & n23262 ;
  assign n23264 = n23249 & n23263 ;
  assign n23265 = n23181 & ~n23264 ;
  assign n23266 = ~n23161 & ~n23199 ;
  assign n23267 = n23149 & n23266 ;
  assign n23268 = ~n23161 & n23199 ;
  assign n23269 = ~n23149 & n23268 ;
  assign n23270 = ~n23267 & ~n23269 ;
  assign n23271 = ~n23265 & n23270 ;
  assign n23272 = ~n23143 & n23199 ;
  assign n23273 = ~n133 & n22464 ;
  assign n23274 = ~n21694 & n23273 ;
  assign n23275 = ~n23171 & n23274 ;
  assign n23276 = ~\a[1]  & \b[63]  ;
  assign n23277 = ~\a[0]  & n23276 ;
  assign n23278 = \a[2]  & ~n23277 ;
  assign n23279 = ~n23275 & ~n23278 ;
  assign n23280 = \a[2]  & ~n21694 ;
  assign n23281 = n23273 & n23280 ;
  assign n23282 = ~n23171 & n23281 ;
  assign n23283 = ~n23279 & ~n23282 ;
  assign n23284 = n23148 & n23283 ;
  assign n23285 = ~n23272 & n23284 ;
  assign n23286 = n23148 & ~n23272 ;
  assign n23287 = ~n23283 & ~n23286 ;
  assign n23288 = ~n23285 & ~n23287 ;
  assign n23289 = ~n22375 & n23108 ;
  assign n23290 = ~n22498 & n23289 ;
  assign n23291 = n23113 & ~n23290 ;
  assign n23292 = n22502 & n23103 ;
  assign n23293 = ~n23097 & ~n23292 ;
  assign n23294 = ~n22327 & n23064 ;
  assign n23295 = ~n22520 & n23294 ;
  assign n23296 = n23069 & ~n23295 ;
  assign n23297 = n22524 & n23059 ;
  assign n23298 = n23053 & ~n23297 ;
  assign n23299 = n1467 & n14052 ;
  assign n23300 = ~n14049 & n23299 ;
  assign n23301 = n1467 & ~n14052 ;
  assign n23302 = ~n13519 & n23301 ;
  assign n23303 = ~n14048 & n23302 ;
  assign n23304 = \b[48]  & n1652 ;
  assign n23305 = n1649 & n23304 ;
  assign n23306 = ~\a[15]  & \b[49]  ;
  assign n23307 = n1459 & n23306 ;
  assign n23308 = ~n23305 & ~n23307 ;
  assign n23309 = \b[50]  & n1465 ;
  assign n23310 = \a[15]  & \b[49]  ;
  assign n23311 = n1456 & n23310 ;
  assign n23312 = \a[17]  & ~n23311 ;
  assign n23313 = ~n23309 & n23312 ;
  assign n23314 = n23308 & n23313 ;
  assign n23315 = ~n23303 & n23314 ;
  assign n23316 = ~n23300 & n23315 ;
  assign n23317 = ~n23309 & ~n23311 ;
  assign n23318 = n23308 & n23317 ;
  assign n23319 = ~n23303 & n23318 ;
  assign n23320 = ~n23300 & n23319 ;
  assign n23321 = ~\a[17]  & ~n23320 ;
  assign n23322 = ~n23316 & ~n23321 ;
  assign n23323 = n22281 & ~n23046 ;
  assign n23324 = ~n22542 & n23323 ;
  assign n23325 = ~n23047 & ~n23324 ;
  assign n23326 = n1965 & ~n12438 ;
  assign n23327 = ~n12436 & n23326 ;
  assign n23328 = \b[47]  & n1963 ;
  assign n23329 = \a[18]  & \b[46]  ;
  assign n23330 = n2210 & n23329 ;
  assign n23331 = ~n23328 & ~n23330 ;
  assign n23332 = \b[45]  & n2218 ;
  assign n23333 = n2216 & n23332 ;
  assign n23334 = ~\a[18]  & \b[46]  ;
  assign n23335 = n1957 & n23334 ;
  assign n23336 = ~n23333 & ~n23335 ;
  assign n23337 = n23331 & n23336 ;
  assign n23338 = ~n23327 & n23337 ;
  assign n23339 = ~\a[20]  & ~n23338 ;
  assign n23340 = \a[20]  & n23337 ;
  assign n23341 = ~n23327 & n23340 ;
  assign n23342 = ~n23339 & ~n23341 ;
  assign n23343 = ~n23036 & ~n23043 ;
  assign n23344 = n2622 & ~n10892 ;
  assign n23345 = ~n10890 & n23344 ;
  assign n23346 = \b[42]  & n2912 ;
  assign n23347 = n2909 & n23346 ;
  assign n23348 = ~\a[21]  & \b[43]  ;
  assign n23349 = n2614 & n23348 ;
  assign n23350 = ~n23347 & ~n23349 ;
  assign n23351 = \b[44]  & n2620 ;
  assign n23352 = \a[21]  & \b[43]  ;
  assign n23353 = n20849 & n23352 ;
  assign n23354 = \a[23]  & ~n23353 ;
  assign n23355 = ~n23351 & n23354 ;
  assign n23356 = n23350 & n23355 ;
  assign n23357 = ~n23345 & n23356 ;
  assign n23358 = ~n23351 & ~n23353 ;
  assign n23359 = n23350 & n23358 ;
  assign n23360 = ~n23345 & n23359 ;
  assign n23361 = ~\a[23]  & ~n23360 ;
  assign n23362 = ~n23357 & ~n23361 ;
  assign n23363 = ~n22242 & n23001 ;
  assign n23364 = ~n22588 & n23363 ;
  assign n23365 = n23006 & ~n23364 ;
  assign n23366 = ~n22594 & n22979 ;
  assign n23367 = n22973 & ~n23366 ;
  assign n23368 = n5211 & ~n6610 ;
  assign n23369 = ~n6608 & n23368 ;
  assign n23370 = \b[33]  & n5595 ;
  assign n23371 = n5592 & n23370 ;
  assign n23372 = ~\a[30]  & \b[34]  ;
  assign n23373 = n5203 & n23372 ;
  assign n23374 = ~n23371 & ~n23373 ;
  assign n23375 = \b[35]  & n5209 ;
  assign n23376 = \a[30]  & \b[34]  ;
  assign n23377 = n5200 & n23376 ;
  assign n23378 = \a[32]  & ~n23377 ;
  assign n23379 = ~n23375 & n23378 ;
  assign n23380 = n23374 & n23379 ;
  assign n23381 = ~n23369 & n23380 ;
  assign n23382 = ~n23375 & ~n23377 ;
  assign n23383 = n23374 & n23382 ;
  assign n23384 = ~n23369 & n23383 ;
  assign n23385 = ~\a[32]  & ~n23384 ;
  assign n23386 = ~n23381 & ~n23385 ;
  assign n23387 = ~n22182 & n22943 ;
  assign n23388 = ~n22189 & n23387 ;
  assign n23389 = n22938 & ~n23388 ;
  assign n23390 = n22598 & n22916 ;
  assign n23391 = ~n22910 & ~n23390 ;
  assign n23392 = n22112 & n22876 ;
  assign n23393 = ~n22599 & n23392 ;
  assign n23394 = n22881 & ~n23393 ;
  assign n23395 = n22603 & n22847 ;
  assign n23396 = n22841 & ~n23395 ;
  assign n23397 = ~n3022 & n10082 ;
  assign n23398 = ~n3020 & n23397 ;
  assign n23399 = \b[21]  & n10681 ;
  assign n23400 = n10678 & n23399 ;
  assign n23401 = \b[23]  & n10080 ;
  assign n23402 = \a[42]  & \b[22]  ;
  assign n23403 = n10071 & n23402 ;
  assign n23404 = ~\a[42]  & \b[22]  ;
  assign n23405 = n10074 & n23404 ;
  assign n23406 = ~n23403 & ~n23405 ;
  assign n23407 = ~n23401 & n23406 ;
  assign n23408 = ~n23400 & n23407 ;
  assign n23409 = ~\a[44]  & n23408 ;
  assign n23410 = ~n23398 & n23409 ;
  assign n23411 = ~n23398 & n23408 ;
  assign n23412 = \a[44]  & ~n23411 ;
  assign n23413 = ~n23410 & ~n23412 ;
  assign n23414 = ~n22076 & n22813 ;
  assign n23415 = ~n22078 & n23414 ;
  assign n23416 = n22808 & ~n23415 ;
  assign n23417 = n22607 & n22779 ;
  assign n23418 = n22773 & ~n23417 ;
  assign n23419 = ~n22014 & n22743 ;
  assign n23420 = ~n22608 & n23419 ;
  assign n23421 = n22738 & ~n23420 ;
  assign n23422 = ~n1694 & n13125 ;
  assign n23423 = ~n1692 & n23422 ;
  assign n23424 = \b[17]  & n13123 ;
  assign n23425 = \a[48]  & \b[16]  ;
  assign n23426 = n13786 & n23425 ;
  assign n23427 = ~n23424 & ~n23426 ;
  assign n23428 = \b[15]  & n13794 ;
  assign n23429 = n13792 & n23428 ;
  assign n23430 = ~\a[48]  & \b[16]  ;
  assign n23431 = n13117 & n23430 ;
  assign n23432 = ~n23429 & ~n23431 ;
  assign n23433 = n23427 & n23432 ;
  assign n23434 = ~n23423 & n23433 ;
  assign n23435 = ~\a[50]  & ~n23434 ;
  assign n23436 = \a[50]  & n23433 ;
  assign n23437 = ~n23423 & n23436 ;
  assign n23438 = ~n23435 & ~n23437 ;
  assign n23439 = n22612 & n22709 ;
  assign n23440 = n22703 & ~n23439 ;
  assign n23441 = ~n21968 & ~n22674 ;
  assign n23442 = ~n22613 & n23441 ;
  assign n23443 = ~n22673 & ~n23442 ;
  assign n23444 = ~n725 & n16655 ;
  assign n23445 = ~n684 & n16655 ;
  assign n23446 = ~n721 & n23445 ;
  assign n23447 = ~n23444 & ~n23446 ;
  assign n23448 = ~n728 & ~n23447 ;
  assign n23449 = \b[9]  & n17308 ;
  assign n23450 = n17305 & n23449 ;
  assign n23451 = ~\a[54]  & \b[10]  ;
  assign n23452 = n16647 & n23451 ;
  assign n23453 = ~n23450 & ~n23452 ;
  assign n23454 = \b[11]  & n16653 ;
  assign n23455 = \a[54]  & \b[10]  ;
  assign n23456 = n16644 & n23455 ;
  assign n23457 = \a[56]  & ~n23456 ;
  assign n23458 = ~n23454 & n23457 ;
  assign n23459 = n23453 & n23458 ;
  assign n23460 = ~n23448 & n23459 ;
  assign n23461 = ~n23454 & ~n23456 ;
  assign n23462 = n23453 & n23461 ;
  assign n23463 = ~\a[56]  & ~n23462 ;
  assign n23464 = ~\a[56]  & ~n728 ;
  assign n23465 = ~n23447 & n23464 ;
  assign n23466 = ~n23463 & ~n23465 ;
  assign n23467 = ~n23460 & n23466 ;
  assign n23468 = n22636 & n22646 ;
  assign n23469 = ~n21961 & n22646 ;
  assign n23470 = ~n21964 & n23469 ;
  assign n23471 = ~n23468 & ~n23470 ;
  assign n23472 = ~n273 & n20521 ;
  assign n23473 = ~n271 & n23472 ;
  assign n23474 = \b[3]  & n21315 ;
  assign n23475 = n21312 & n23474 ;
  assign n23476 = \b[5]  & n20519 ;
  assign n23477 = \a[59]  & \b[4]  ;
  assign n23478 = n21313 & n23477 ;
  assign n23479 = ~\a[60]  & \b[4]  ;
  assign n23480 = n20513 & n23479 ;
  assign n23481 = ~n23478 & ~n23480 ;
  assign n23482 = ~n23476 & n23481 ;
  assign n23483 = ~n23475 & n23482 ;
  assign n23484 = ~n23473 & n23483 ;
  assign n23485 = \b[2]  & n22643 ;
  assign n23486 = ~n23484 & n23485 ;
  assign n23487 = \b[1]  & n21957 ;
  assign n23488 = \b[2]  & n22637 ;
  assign n23489 = ~n23487 & ~n23488 ;
  assign n23490 = n23483 & ~n23489 ;
  assign n23491 = ~n23473 & n23490 ;
  assign n23492 = ~n23486 & ~n23491 ;
  assign n23493 = ~\a[62]  & ~n23484 ;
  assign n23494 = \b[2]  & n21958 ;
  assign n23495 = ~n23487 & ~n23494 ;
  assign n23496 = \a[62]  & n23483 ;
  assign n23497 = ~n23473 & n23496 ;
  assign n23498 = n23495 & ~n23497 ;
  assign n23499 = ~n23493 & n23498 ;
  assign n23500 = n23492 & ~n23499 ;
  assign n23501 = ~n23471 & ~n23500 ;
  assign n23502 = n23471 & n23500 ;
  assign n23503 = ~n23501 & ~n23502 ;
  assign n23504 = ~n505 & ~n17912 ;
  assign n23505 = ~n18513 & n23504 ;
  assign n23506 = n502 & n23505 ;
  assign n23507 = n505 & ~n17912 ;
  assign n23508 = ~n18513 & n23507 ;
  assign n23509 = ~n502 & n23508 ;
  assign n23510 = ~n23506 & ~n23509 ;
  assign n23511 = \b[6]  & n19183 ;
  assign n23512 = n19180 & n23511 ;
  assign n23513 = ~\a[57]  & \b[7]  ;
  assign n23514 = n18508 & n23513 ;
  assign n23515 = ~n23512 & ~n23514 ;
  assign n23516 = \b[8]  & n18514 ;
  assign n23517 = \a[57]  & \b[7]  ;
  assign n23518 = n18505 & n23517 ;
  assign n23519 = \a[59]  & ~n23518 ;
  assign n23520 = ~n23516 & n23519 ;
  assign n23521 = n23515 & n23520 ;
  assign n23522 = n23510 & n23521 ;
  assign n23523 = ~n23516 & ~n23518 ;
  assign n23524 = n23515 & n23523 ;
  assign n23525 = n23510 & n23524 ;
  assign n23526 = ~\a[59]  & ~n23525 ;
  assign n23527 = ~n23522 & ~n23526 ;
  assign n23528 = n23503 & ~n23527 ;
  assign n23529 = ~n23503 & n23527 ;
  assign n23530 = ~n23528 & ~n23529 ;
  assign n23531 = n23467 & ~n23530 ;
  assign n23532 = ~n23443 & n23531 ;
  assign n23533 = n23467 & n23530 ;
  assign n23534 = n23443 & n23533 ;
  assign n23535 = ~n23532 & ~n23534 ;
  assign n23536 = ~n23467 & ~n23530 ;
  assign n23537 = n23443 & n23536 ;
  assign n23538 = ~n23467 & n23530 ;
  assign n23539 = ~n23443 & n23538 ;
  assign n23540 = ~n23537 & ~n23539 ;
  assign n23541 = n23535 & n23540 ;
  assign n23542 = ~n23440 & n23541 ;
  assign n23543 = n22703 & ~n23541 ;
  assign n23544 = ~n23439 & n23543 ;
  assign n23545 = n1087 & n14793 ;
  assign n23546 = ~n1084 & n23545 ;
  assign n23547 = n14793 & n21340 ;
  assign n23548 = ~n1083 & n23547 ;
  assign n23549 = \b[12]  & n15517 ;
  assign n23550 = n15514 & n23549 ;
  assign n23551 = ~\a[51]  & \b[13]  ;
  assign n23552 = n14785 & n23551 ;
  assign n23553 = ~n23550 & ~n23552 ;
  assign n23554 = \b[14]  & n14791 ;
  assign n23555 = \a[51]  & \b[13]  ;
  assign n23556 = n14782 & n23555 ;
  assign n23557 = \a[53]  & ~n23556 ;
  assign n23558 = ~n23554 & n23557 ;
  assign n23559 = n23553 & n23558 ;
  assign n23560 = ~n23548 & n23559 ;
  assign n23561 = ~n23546 & n23560 ;
  assign n23562 = ~n23554 & ~n23556 ;
  assign n23563 = n23553 & n23562 ;
  assign n23564 = ~n23548 & n23563 ;
  assign n23565 = ~n23546 & n23564 ;
  assign n23566 = ~\a[53]  & ~n23565 ;
  assign n23567 = ~n23561 & ~n23566 ;
  assign n23568 = ~n23544 & ~n23567 ;
  assign n23569 = ~n23542 & n23568 ;
  assign n23570 = ~n23541 & n23567 ;
  assign n23571 = n23440 & n23570 ;
  assign n23572 = n23541 & n23567 ;
  assign n23573 = ~n23440 & n23572 ;
  assign n23574 = ~n23571 & ~n23573 ;
  assign n23575 = ~n23569 & n23574 ;
  assign n23576 = ~n23438 & ~n23575 ;
  assign n23577 = n23421 & n23576 ;
  assign n23578 = ~n23438 & n23575 ;
  assign n23579 = ~n23421 & n23578 ;
  assign n23580 = ~n23577 & ~n23579 ;
  assign n23581 = n23438 & ~n23575 ;
  assign n23582 = ~n23421 & n23581 ;
  assign n23583 = n23438 & n23575 ;
  assign n23584 = n23421 & n23583 ;
  assign n23585 = ~n23582 & ~n23584 ;
  assign n23586 = n23580 & n23585 ;
  assign n23587 = ~n23418 & n23586 ;
  assign n23588 = n22773 & ~n23586 ;
  assign n23589 = ~n23417 & n23588 ;
  assign n23590 = n2293 & n11572 ;
  assign n23591 = ~n19247 & n23590 ;
  assign n23592 = ~n2293 & n11572 ;
  assign n23593 = ~n2074 & n23592 ;
  assign n23594 = ~n2289 & n23593 ;
  assign n23595 = \b[18]  & n12159 ;
  assign n23596 = n12156 & n23595 ;
  assign n23597 = ~\a[45]  & \b[19]  ;
  assign n23598 = n11564 & n23597 ;
  assign n23599 = ~n23596 & ~n23598 ;
  assign n23600 = \b[20]  & n11570 ;
  assign n23601 = \a[45]  & \b[19]  ;
  assign n23602 = n11561 & n23601 ;
  assign n23603 = \a[47]  & ~n23602 ;
  assign n23604 = ~n23600 & n23603 ;
  assign n23605 = n23599 & n23604 ;
  assign n23606 = ~n23594 & n23605 ;
  assign n23607 = ~n23591 & n23606 ;
  assign n23608 = ~n23600 & ~n23602 ;
  assign n23609 = n23599 & n23608 ;
  assign n23610 = ~n23594 & n23609 ;
  assign n23611 = ~n23591 & n23610 ;
  assign n23612 = ~\a[47]  & ~n23611 ;
  assign n23613 = ~n23607 & ~n23612 ;
  assign n23614 = ~n23589 & ~n23613 ;
  assign n23615 = ~n23587 & n23614 ;
  assign n23616 = ~n23586 & n23613 ;
  assign n23617 = n23418 & n23616 ;
  assign n23618 = n23586 & n23613 ;
  assign n23619 = ~n23418 & n23618 ;
  assign n23620 = ~n23617 & ~n23619 ;
  assign n23621 = ~n23615 & n23620 ;
  assign n23622 = n23416 & n23621 ;
  assign n23623 = ~n23416 & ~n23621 ;
  assign n23624 = ~n23622 & ~n23623 ;
  assign n23625 = n23413 & n23624 ;
  assign n23626 = ~n23413 & ~n23624 ;
  assign n23627 = ~n23625 & ~n23626 ;
  assign n23628 = n3604 & n8759 ;
  assign n23629 = ~n19292 & n23628 ;
  assign n23630 = n8759 & n12021 ;
  assign n23631 = ~n3600 & n23630 ;
  assign n23632 = \b[24]  & n9301 ;
  assign n23633 = n9298 & n23632 ;
  assign n23634 = ~\a[39]  & \b[25]  ;
  assign n23635 = n8751 & n23634 ;
  assign n23636 = ~n23633 & ~n23635 ;
  assign n23637 = \b[26]  & n8757 ;
  assign n23638 = \a[39]  & \b[25]  ;
  assign n23639 = n8748 & n23638 ;
  assign n23640 = \a[41]  & ~n23639 ;
  assign n23641 = ~n23637 & n23640 ;
  assign n23642 = n23636 & n23641 ;
  assign n23643 = ~n23631 & n23642 ;
  assign n23644 = ~n23629 & n23643 ;
  assign n23645 = ~n23637 & ~n23639 ;
  assign n23646 = n23636 & n23645 ;
  assign n23647 = ~n23631 & n23646 ;
  assign n23648 = ~n23629 & n23647 ;
  assign n23649 = ~\a[41]  & ~n23648 ;
  assign n23650 = ~n23644 & ~n23649 ;
  assign n23651 = ~n23627 & ~n23650 ;
  assign n23652 = ~n23396 & n23651 ;
  assign n23653 = n23627 & ~n23650 ;
  assign n23654 = n23396 & n23653 ;
  assign n23655 = ~n23652 & ~n23654 ;
  assign n23656 = ~n23627 & n23650 ;
  assign n23657 = n23396 & n23656 ;
  assign n23658 = n23627 & n23650 ;
  assign n23659 = ~n23396 & n23658 ;
  assign n23660 = ~n23657 & ~n23659 ;
  assign n23661 = n23655 & n23660 ;
  assign n23662 = ~n4499 & n7534 ;
  assign n23663 = ~n4455 & n7534 ;
  assign n23664 = ~n4495 & n23663 ;
  assign n23665 = ~n23662 & ~n23664 ;
  assign n23666 = ~n4502 & ~n23665 ;
  assign n23667 = \b[27]  & n7973 ;
  assign n23668 = n7970 & n23667 ;
  assign n23669 = ~\a[36]  & \b[28]  ;
  assign n23670 = n7526 & n23669 ;
  assign n23671 = ~n23668 & ~n23670 ;
  assign n23672 = \b[29]  & n7532 ;
  assign n23673 = \a[36]  & \b[28]  ;
  assign n23674 = n17801 & n23673 ;
  assign n23675 = \a[38]  & ~n23674 ;
  assign n23676 = ~n23672 & n23675 ;
  assign n23677 = n23671 & n23676 ;
  assign n23678 = ~n23666 & n23677 ;
  assign n23679 = ~n23672 & ~n23674 ;
  assign n23680 = n23671 & n23679 ;
  assign n23681 = ~\a[38]  & ~n23680 ;
  assign n23682 = ~\a[38]  & ~n4502 ;
  assign n23683 = ~n23665 & n23682 ;
  assign n23684 = ~n23681 & ~n23683 ;
  assign n23685 = ~n23678 & n23684 ;
  assign n23686 = ~n23661 & ~n23685 ;
  assign n23687 = n23394 & n23686 ;
  assign n23688 = n23661 & ~n23685 ;
  assign n23689 = ~n23394 & n23688 ;
  assign n23690 = ~n23687 & ~n23689 ;
  assign n23691 = ~n23661 & n23685 ;
  assign n23692 = ~n23394 & n23691 ;
  assign n23693 = n23661 & n23685 ;
  assign n23694 = n23394 & n23693 ;
  assign n23695 = ~n23692 & ~n23694 ;
  assign n23696 = n23690 & n23695 ;
  assign n23697 = ~n23391 & n23696 ;
  assign n23698 = ~n22910 & ~n23696 ;
  assign n23699 = ~n23390 & n23698 ;
  assign n23700 = n5810 & n6309 ;
  assign n23701 = ~n5807 & n23700 ;
  assign n23702 = n6309 & n19029 ;
  assign n23703 = ~n5806 & n23702 ;
  assign n23704 = \b[30]  & n6778 ;
  assign n23705 = n6775 & n23704 ;
  assign n23706 = ~\a[33]  & \b[31]  ;
  assign n23707 = n6301 & n23706 ;
  assign n23708 = ~n23705 & ~n23707 ;
  assign n23709 = \b[32]  & n6307 ;
  assign n23710 = \a[33]  & \b[31]  ;
  assign n23711 = n6298 & n23710 ;
  assign n23712 = \a[35]  & ~n23711 ;
  assign n23713 = ~n23709 & n23712 ;
  assign n23714 = n23708 & n23713 ;
  assign n23715 = ~n23703 & n23714 ;
  assign n23716 = ~n23701 & n23715 ;
  assign n23717 = ~n23709 & ~n23711 ;
  assign n23718 = n23708 & n23717 ;
  assign n23719 = ~n23703 & n23718 ;
  assign n23720 = ~n23701 & n23719 ;
  assign n23721 = ~\a[35]  & ~n23720 ;
  assign n23722 = ~n23716 & ~n23721 ;
  assign n23723 = ~n23699 & ~n23722 ;
  assign n23724 = ~n23697 & n23723 ;
  assign n23725 = ~n23696 & n23722 ;
  assign n23726 = n23391 & n23725 ;
  assign n23727 = n23696 & n23722 ;
  assign n23728 = ~n23391 & n23727 ;
  assign n23729 = ~n23726 & ~n23728 ;
  assign n23730 = ~n23724 & n23729 ;
  assign n23731 = n23389 & n23730 ;
  assign n23732 = ~n23389 & ~n23730 ;
  assign n23733 = ~n23731 & ~n23732 ;
  assign n23734 = ~n23386 & n23733 ;
  assign n23735 = n23386 & ~n23733 ;
  assign n23736 = ~n23734 & ~n23735 ;
  assign n23737 = n4249 & n8175 ;
  assign n23738 = ~n8172 & n23737 ;
  assign n23739 = n4249 & ~n8175 ;
  assign n23740 = ~n7756 & n23739 ;
  assign n23741 = ~n8171 & n23740 ;
  assign n23742 = \b[36]  & n4647 ;
  assign n23743 = n4644 & n23742 ;
  assign n23744 = ~\a[27]  & \b[37]  ;
  assign n23745 = n4241 & n23744 ;
  assign n23746 = ~n23743 & ~n23745 ;
  assign n23747 = \b[38]  & n4247 ;
  assign n23748 = \a[27]  & \b[37]  ;
  assign n23749 = n4238 & n23748 ;
  assign n23750 = \a[29]  & ~n23749 ;
  assign n23751 = ~n23747 & n23750 ;
  assign n23752 = n23746 & n23751 ;
  assign n23753 = ~n23741 & n23752 ;
  assign n23754 = ~n23738 & n23753 ;
  assign n23755 = ~n23747 & ~n23749 ;
  assign n23756 = n23746 & n23755 ;
  assign n23757 = ~n23741 & n23756 ;
  assign n23758 = ~n23738 & n23757 ;
  assign n23759 = ~\a[29]  & ~n23758 ;
  assign n23760 = ~n23754 & ~n23759 ;
  assign n23761 = ~n23736 & ~n23760 ;
  assign n23762 = ~n23367 & n23761 ;
  assign n23763 = n23736 & ~n23760 ;
  assign n23764 = n23367 & n23763 ;
  assign n23765 = ~n23762 & ~n23764 ;
  assign n23766 = ~n23736 & n23760 ;
  assign n23767 = n23367 & n23766 ;
  assign n23768 = n23736 & n23760 ;
  assign n23769 = ~n23367 & n23768 ;
  assign n23770 = ~n23767 & ~n23769 ;
  assign n23771 = n23765 & n23770 ;
  assign n23772 = ~n23365 & ~n23771 ;
  assign n23773 = n23006 & n23771 ;
  assign n23774 = ~n23364 & n23773 ;
  assign n23775 = n3402 & ~n9482 ;
  assign n23776 = ~n9480 & n23775 ;
  assign n23777 = \b[41]  & n3400 ;
  assign n23778 = \a[24]  & \b[40]  ;
  assign n23779 = n3391 & n23778 ;
  assign n23780 = ~n23777 & ~n23779 ;
  assign n23781 = \b[39]  & n3733 ;
  assign n23782 = n3730 & n23781 ;
  assign n23783 = ~\a[24]  & \b[40]  ;
  assign n23784 = n3394 & n23783 ;
  assign n23785 = ~n23782 & ~n23784 ;
  assign n23786 = n23780 & n23785 ;
  assign n23787 = ~n23776 & n23786 ;
  assign n23788 = ~\a[26]  & ~n23787 ;
  assign n23789 = \a[26]  & n23786 ;
  assign n23790 = ~n23776 & n23789 ;
  assign n23791 = ~n23788 & ~n23790 ;
  assign n23792 = ~n23774 & ~n23791 ;
  assign n23793 = ~n23772 & n23792 ;
  assign n23794 = ~n23771 & n23791 ;
  assign n23795 = ~n23365 & n23794 ;
  assign n23796 = n23771 & n23791 ;
  assign n23797 = n23365 & n23796 ;
  assign n23798 = ~n23795 & ~n23797 ;
  assign n23799 = ~n23793 & n23798 ;
  assign n23800 = ~n23362 & ~n23799 ;
  assign n23801 = ~n23343 & n23800 ;
  assign n23802 = ~n23362 & n23799 ;
  assign n23803 = n23343 & n23802 ;
  assign n23804 = ~n23801 & ~n23803 ;
  assign n23805 = n23362 & ~n23799 ;
  assign n23806 = n23343 & n23805 ;
  assign n23807 = n23362 & n23799 ;
  assign n23808 = ~n23343 & n23807 ;
  assign n23809 = ~n23806 & ~n23808 ;
  assign n23810 = n23804 & n23809 ;
  assign n23811 = ~n23342 & ~n23810 ;
  assign n23812 = n23325 & n23811 ;
  assign n23813 = ~n23342 & n23810 ;
  assign n23814 = ~n23325 & n23813 ;
  assign n23815 = ~n23812 & ~n23814 ;
  assign n23816 = n23342 & ~n23810 ;
  assign n23817 = ~n23325 & n23816 ;
  assign n23818 = n23342 & n23810 ;
  assign n23819 = n23325 & n23818 ;
  assign n23820 = ~n23817 & ~n23819 ;
  assign n23821 = n23815 & n23820 ;
  assign n23822 = n23322 & ~n23821 ;
  assign n23823 = n23298 & n23822 ;
  assign n23824 = n23322 & n23821 ;
  assign n23825 = ~n23298 & n23824 ;
  assign n23826 = ~n23823 & ~n23825 ;
  assign n23827 = ~n23298 & n23821 ;
  assign n23828 = n23053 & ~n23821 ;
  assign n23829 = ~n23297 & n23828 ;
  assign n23830 = ~n23322 & ~n23829 ;
  assign n23831 = ~n23827 & n23830 ;
  assign n23832 = n23826 & ~n23831 ;
  assign n23833 = n999 & ~n15246 ;
  assign n23834 = ~n15244 & n23833 ;
  assign n23835 = \b[51]  & n1182 ;
  assign n23836 = n1179 & n23835 ;
  assign n23837 = \b[53]  & n997 ;
  assign n23838 = \a[11]  & \b[52]  ;
  assign n23839 = n1180 & n23838 ;
  assign n23840 = ~\a[12]  & \b[52]  ;
  assign n23841 = n7674 & n23840 ;
  assign n23842 = ~n23839 & ~n23841 ;
  assign n23843 = ~n23837 & n23842 ;
  assign n23844 = ~n23836 & n23843 ;
  assign n23845 = ~n23834 & n23844 ;
  assign n23846 = ~\a[14]  & ~n23845 ;
  assign n23847 = \a[14]  & n23844 ;
  assign n23848 = ~n23834 & n23847 ;
  assign n23849 = ~n23846 & ~n23848 ;
  assign n23850 = ~n23832 & ~n23849 ;
  assign n23851 = n23296 & n23850 ;
  assign n23852 = n23832 & ~n23849 ;
  assign n23853 = ~n23296 & n23852 ;
  assign n23854 = ~n23851 & ~n23853 ;
  assign n23855 = ~n23832 & n23849 ;
  assign n23856 = ~n23296 & n23855 ;
  assign n23857 = n23832 & n23849 ;
  assign n23858 = n23296 & n23857 ;
  assign n23859 = ~n23856 & ~n23858 ;
  assign n23860 = n23854 & n23859 ;
  assign n23861 = ~n551 & ~n16441 ;
  assign n23862 = ~n17647 & n23861 ;
  assign n23863 = ~n17643 & n23862 ;
  assign n23864 = ~n643 & n23863 ;
  assign n23865 = n646 & n17647 ;
  assign n23866 = ~n17644 & n23865 ;
  assign n23867 = ~n23864 & ~n23866 ;
  assign n23868 = \b[54]  & n796 ;
  assign n23869 = n793 & n23868 ;
  assign n23870 = ~\a[9]  & \b[55]  ;
  assign n23871 = n638 & n23870 ;
  assign n23872 = ~n23869 & ~n23871 ;
  assign n23873 = \b[56]  & n644 ;
  assign n23874 = \a[9]  & \b[55]  ;
  assign n23875 = n635 & n23874 ;
  assign n23876 = \a[11]  & ~n23875 ;
  assign n23877 = ~n23873 & n23876 ;
  assign n23878 = n23872 & n23877 ;
  assign n23879 = n23867 & n23878 ;
  assign n23880 = ~n23873 & ~n23875 ;
  assign n23881 = n23872 & n23880 ;
  assign n23882 = n23867 & n23881 ;
  assign n23883 = ~\a[11]  & ~n23882 ;
  assign n23884 = ~n23879 & ~n23883 ;
  assign n23885 = ~n23860 & n23884 ;
  assign n23886 = n23293 & n23885 ;
  assign n23887 = n23860 & n23884 ;
  assign n23888 = ~n23293 & n23887 ;
  assign n23889 = ~n23886 & ~n23888 ;
  assign n23890 = ~n23293 & n23860 ;
  assign n23891 = ~n23097 & ~n23860 ;
  assign n23892 = ~n23292 & n23891 ;
  assign n23893 = ~n23884 & ~n23892 ;
  assign n23894 = ~n23890 & n23893 ;
  assign n23895 = n23889 & ~n23894 ;
  assign n23896 = n430 & ~n19550 ;
  assign n23897 = ~n19548 & n23896 ;
  assign n23898 = \b[57]  & n486 ;
  assign n23899 = n483 & n23898 ;
  assign n23900 = ~\a[6]  & \b[58]  ;
  assign n23901 = n422 & n23900 ;
  assign n23902 = ~n23899 & ~n23901 ;
  assign n23903 = \b[59]  & n428 ;
  assign n23904 = \a[6]  & \b[58]  ;
  assign n23905 = n419 & n23904 ;
  assign n23906 = \a[8]  & ~n23905 ;
  assign n23907 = ~n23903 & n23906 ;
  assign n23908 = n23902 & n23907 ;
  assign n23909 = ~n23897 & n23908 ;
  assign n23910 = ~n23903 & ~n23905 ;
  assign n23911 = n23902 & n23910 ;
  assign n23912 = ~n23897 & n23911 ;
  assign n23913 = ~\a[8]  & ~n23912 ;
  assign n23914 = ~n23909 & ~n23913 ;
  assign n23915 = n252 & ~n21699 ;
  assign n23916 = ~n21697 & n23915 ;
  assign n23917 = \b[60]  & n303 ;
  assign n23918 = n300 & n23917 ;
  assign n23919 = ~\a[3]  & \b[61]  ;
  assign n23920 = n244 & n23919 ;
  assign n23921 = ~n23918 & ~n23920 ;
  assign n23922 = \b[62]  & n250 ;
  assign n23923 = \a[3]  & \b[61]  ;
  assign n23924 = n241 & n23923 ;
  assign n23925 = \a[5]  & ~n23924 ;
  assign n23926 = ~n23922 & n23925 ;
  assign n23927 = n23921 & n23926 ;
  assign n23928 = ~n23916 & n23927 ;
  assign n23929 = ~n23922 & ~n23924 ;
  assign n23930 = n23921 & n23929 ;
  assign n23931 = ~n23916 & n23930 ;
  assign n23932 = ~\a[5]  & ~n23931 ;
  assign n23933 = ~n23928 & ~n23932 ;
  assign n23934 = n23914 & ~n23933 ;
  assign n23935 = ~n23895 & n23934 ;
  assign n23936 = ~n23291 & n23935 ;
  assign n23937 = ~n23914 & ~n23933 ;
  assign n23938 = n23895 & n23937 ;
  assign n23939 = ~n23291 & n23938 ;
  assign n23940 = ~n23936 & ~n23939 ;
  assign n23941 = ~n23895 & n23937 ;
  assign n23942 = n23291 & n23941 ;
  assign n23943 = n23895 & n23934 ;
  assign n23944 = n23291 & n23943 ;
  assign n23945 = ~n23942 & ~n23944 ;
  assign n23946 = n23940 & n23945 ;
  assign n23947 = n23895 & ~n23914 ;
  assign n23948 = ~n23291 & n23947 ;
  assign n23949 = ~n23895 & n23914 ;
  assign n23950 = ~n23291 & n23949 ;
  assign n23951 = ~n23948 & ~n23950 ;
  assign n23952 = ~n23884 & ~n23914 ;
  assign n23953 = ~n23860 & n23952 ;
  assign n23954 = n23293 & n23953 ;
  assign n23955 = n23884 & ~n23914 ;
  assign n23956 = ~n23860 & n23955 ;
  assign n23957 = ~n23293 & n23956 ;
  assign n23958 = ~n23954 & ~n23957 ;
  assign n23959 = n23860 & n23952 ;
  assign n23960 = ~n23293 & n23959 ;
  assign n23961 = n23860 & n23955 ;
  assign n23962 = n23293 & n23961 ;
  assign n23963 = ~n23960 & ~n23962 ;
  assign n23964 = n23958 & n23963 ;
  assign n23965 = ~n23884 & n23914 ;
  assign n23966 = ~n23860 & n23965 ;
  assign n23967 = ~n23293 & n23966 ;
  assign n23968 = n23884 & n23914 ;
  assign n23969 = ~n23860 & n23968 ;
  assign n23970 = n23293 & n23969 ;
  assign n23971 = ~n23967 & ~n23970 ;
  assign n23972 = n23860 & n23965 ;
  assign n23973 = n23293 & n23972 ;
  assign n23974 = n23860 & n23968 ;
  assign n23975 = ~n23293 & n23974 ;
  assign n23976 = ~n23973 & ~n23975 ;
  assign n23977 = n23971 & n23976 ;
  assign n23978 = n23964 & n23977 ;
  assign n23979 = n23291 & n23978 ;
  assign n23980 = n23933 & ~n23979 ;
  assign n23981 = n23951 & n23980 ;
  assign n23982 = n23946 & ~n23981 ;
  assign n23983 = n23288 & ~n23982 ;
  assign n23984 = ~n23288 & n23982 ;
  assign n23985 = ~n23983 & ~n23984 ;
  assign n23986 = ~n23271 & ~n23985 ;
  assign n23987 = n23271 & n23985 ;
  assign n23988 = ~n23986 & ~n23987 ;
  assign n23989 = n23229 & n23988 ;
  assign n23990 = n23233 & n23988 ;
  assign n23991 = ~n23989 & ~n23990 ;
  assign n23992 = ~n23229 & ~n23988 ;
  assign n23993 = ~n23233 & n23992 ;
  assign n23994 = n23991 & ~n23993 ;
  assign n23995 = n430 & n20260 ;
  assign n23996 = ~n20257 & n23995 ;
  assign n23997 = n430 & ~n20260 ;
  assign n23998 = ~n19545 & n23997 ;
  assign n23999 = ~n20256 & n23998 ;
  assign n24000 = \b[58]  & n486 ;
  assign n24001 = n483 & n24000 ;
  assign n24002 = ~\a[6]  & \b[59]  ;
  assign n24003 = n422 & n24002 ;
  assign n24004 = ~n24001 & ~n24003 ;
  assign n24005 = \b[60]  & n428 ;
  assign n24006 = \a[6]  & \b[59]  ;
  assign n24007 = n419 & n24006 ;
  assign n24008 = \a[8]  & ~n24007 ;
  assign n24009 = ~n24005 & n24008 ;
  assign n24010 = n24004 & n24009 ;
  assign n24011 = ~n23999 & n24010 ;
  assign n24012 = ~n23996 & n24011 ;
  assign n24013 = ~n24005 & ~n24007 ;
  assign n24014 = n24004 & n24013 ;
  assign n24015 = ~n23999 & n24014 ;
  assign n24016 = ~n23996 & n24015 ;
  assign n24017 = ~\a[8]  & ~n24016 ;
  assign n24018 = ~n24012 & ~n24017 ;
  assign n24019 = \a[8]  & ~n23912 ;
  assign n24020 = ~\a[8]  & n23912 ;
  assign n24021 = ~n24019 & ~n24020 ;
  assign n24022 = n23889 & n24021 ;
  assign n24023 = ~n23894 & ~n24022 ;
  assign n24024 = ~n24018 & ~n24023 ;
  assign n24025 = ~n23894 & n24018 ;
  assign n24026 = ~n24022 & n24025 ;
  assign n24027 = ~n23097 & n23854 ;
  assign n24028 = ~n23292 & n24027 ;
  assign n24029 = n23296 & n23832 ;
  assign n24030 = ~n23831 & ~n24029 ;
  assign n24031 = n23053 & n23815 ;
  assign n24032 = ~n23297 & n24031 ;
  assign n24033 = n23820 & ~n24032 ;
  assign n24034 = n23325 & n23810 ;
  assign n24035 = n23804 & ~n24034 ;
  assign n24036 = n1965 & n12478 ;
  assign n24037 = ~n12475 & n24036 ;
  assign n24038 = n1965 & ~n12478 ;
  assign n24039 = ~n12433 & n24038 ;
  assign n24040 = ~n12474 & n24039 ;
  assign n24041 = \b[46]  & n2218 ;
  assign n24042 = n2216 & n24041 ;
  assign n24043 = ~\a[18]  & \b[47]  ;
  assign n24044 = n1957 & n24043 ;
  assign n24045 = ~n24042 & ~n24044 ;
  assign n24046 = \b[48]  & n1963 ;
  assign n24047 = \a[18]  & \b[47]  ;
  assign n24048 = n2210 & n24047 ;
  assign n24049 = \a[20]  & ~n24048 ;
  assign n24050 = ~n24046 & n24049 ;
  assign n24051 = n24045 & n24050 ;
  assign n24052 = ~n24040 & n24051 ;
  assign n24053 = ~n24037 & n24052 ;
  assign n24054 = ~n24046 & ~n24048 ;
  assign n24055 = n24045 & n24054 ;
  assign n24056 = ~n24040 & n24055 ;
  assign n24057 = ~n24037 & n24056 ;
  assign n24058 = ~\a[20]  & ~n24057 ;
  assign n24059 = ~n24053 & ~n24058 ;
  assign n24060 = ~n23036 & ~n23793 ;
  assign n24061 = ~n23043 & n24060 ;
  assign n24062 = n23798 & ~n24061 ;
  assign n24063 = n2622 & ~n11397 ;
  assign n24064 = ~n11395 & n24063 ;
  assign n24065 = \b[43]  & n2912 ;
  assign n24066 = n2909 & n24065 ;
  assign n24067 = ~\a[21]  & \b[44]  ;
  assign n24068 = n2614 & n24067 ;
  assign n24069 = ~n24066 & ~n24068 ;
  assign n24070 = \b[45]  & n2620 ;
  assign n24071 = \a[21]  & \b[44]  ;
  assign n24072 = n20849 & n24071 ;
  assign n24073 = \a[23]  & ~n24072 ;
  assign n24074 = ~n24070 & n24073 ;
  assign n24075 = n24069 & n24074 ;
  assign n24076 = ~n24064 & n24075 ;
  assign n24077 = ~n24070 & ~n24072 ;
  assign n24078 = n24069 & n24077 ;
  assign n24079 = ~n24064 & n24078 ;
  assign n24080 = ~\a[23]  & ~n24079 ;
  assign n24081 = ~n24076 & ~n24080 ;
  assign n24082 = ~n24062 & n24081 ;
  assign n24083 = n23798 & ~n24081 ;
  assign n24084 = ~n24061 & n24083 ;
  assign n24085 = n23765 & ~n23774 ;
  assign n24086 = n3402 & n9930 ;
  assign n24087 = ~n9927 & n24086 ;
  assign n24088 = n3402 & ~n9930 ;
  assign n24089 = ~n9477 & n24088 ;
  assign n24090 = ~n9926 & n24089 ;
  assign n24091 = \b[40]  & n3733 ;
  assign n24092 = n3730 & n24091 ;
  assign n24093 = ~\a[24]  & \b[41]  ;
  assign n24094 = n3394 & n24093 ;
  assign n24095 = ~n24092 & ~n24094 ;
  assign n24096 = \b[42]  & n3400 ;
  assign n24097 = \a[24]  & \b[41]  ;
  assign n24098 = n3391 & n24097 ;
  assign n24099 = \a[26]  & ~n24098 ;
  assign n24100 = ~n24096 & n24099 ;
  assign n24101 = n24095 & n24100 ;
  assign n24102 = ~n24090 & n24101 ;
  assign n24103 = ~n24087 & n24102 ;
  assign n24104 = ~n24096 & ~n24098 ;
  assign n24105 = n24095 & n24104 ;
  assign n24106 = ~n24090 & n24105 ;
  assign n24107 = ~n24087 & n24106 ;
  assign n24108 = ~\a[26]  & ~n24107 ;
  assign n24109 = ~n24103 & ~n24108 ;
  assign n24110 = n22973 & ~n23734 ;
  assign n24111 = ~n23366 & n24110 ;
  assign n24112 = ~n23735 & ~n24111 ;
  assign n24113 = n4249 & ~n8602 ;
  assign n24114 = ~n8600 & n24113 ;
  assign n24115 = \b[37]  & n4647 ;
  assign n24116 = n4644 & n24115 ;
  assign n24117 = ~\a[27]  & \b[38]  ;
  assign n24118 = n4241 & n24117 ;
  assign n24119 = ~n24116 & ~n24118 ;
  assign n24120 = \b[39]  & n4247 ;
  assign n24121 = \a[27]  & \b[38]  ;
  assign n24122 = n4238 & n24121 ;
  assign n24123 = \a[29]  & ~n24122 ;
  assign n24124 = ~n24120 & n24123 ;
  assign n24125 = n24119 & n24124 ;
  assign n24126 = ~n24114 & n24125 ;
  assign n24127 = ~n24120 & ~n24122 ;
  assign n24128 = n24119 & n24127 ;
  assign n24129 = ~n24114 & n24128 ;
  assign n24130 = ~\a[29]  & ~n24129 ;
  assign n24131 = ~n24126 & ~n24130 ;
  assign n24132 = ~n24112 & n24131 ;
  assign n24133 = ~n23735 & ~n24131 ;
  assign n24134 = ~n24111 & n24133 ;
  assign n24135 = ~n23724 & ~n23731 ;
  assign n24136 = n5211 & n7337 ;
  assign n24137 = ~n7334 & n24136 ;
  assign n24138 = ~n6605 & ~n7337 ;
  assign n24139 = n5211 & n24138 ;
  assign n24140 = ~n7333 & n24139 ;
  assign n24141 = \b[34]  & n5595 ;
  assign n24142 = n5592 & n24141 ;
  assign n24143 = ~\a[30]  & \b[35]  ;
  assign n24144 = n5203 & n24143 ;
  assign n24145 = ~n24142 & ~n24144 ;
  assign n24146 = \b[36]  & n5209 ;
  assign n24147 = \a[30]  & \b[35]  ;
  assign n24148 = n5200 & n24147 ;
  assign n24149 = \a[32]  & ~n24148 ;
  assign n24150 = ~n24146 & n24149 ;
  assign n24151 = n24145 & n24150 ;
  assign n24152 = ~n24140 & n24151 ;
  assign n24153 = ~n24137 & n24152 ;
  assign n24154 = ~n24146 & ~n24148 ;
  assign n24155 = n24145 & n24154 ;
  assign n24156 = ~n24140 & n24155 ;
  assign n24157 = ~n24137 & n24156 ;
  assign n24158 = ~\a[32]  & ~n24157 ;
  assign n24159 = ~n24153 & ~n24158 ;
  assign n24160 = ~n22910 & n23690 ;
  assign n24161 = ~n23390 & n24160 ;
  assign n24162 = n23695 & ~n24161 ;
  assign n24163 = n23394 & n23661 ;
  assign n24164 = n23655 & ~n24163 ;
  assign n24165 = n22841 & ~n23625 ;
  assign n24166 = ~n23395 & n24165 ;
  assign n24167 = ~n23626 & ~n24166 ;
  assign n24168 = ~n23615 & ~n23622 ;
  assign n24169 = n22773 & n23580 ;
  assign n24170 = ~n23417 & n24169 ;
  assign n24171 = n23585 & ~n24170 ;
  assign n24172 = n23421 & n23575 ;
  assign n24173 = ~n23569 & ~n24172 ;
  assign n24174 = n22703 & n23540 ;
  assign n24175 = ~n23439 & n24174 ;
  assign n24176 = n23535 & ~n24175 ;
  assign n24177 = n23443 & n23530 ;
  assign n24178 = ~n23528 & ~n24177 ;
  assign n24179 = ~n909 & ~n16016 ;
  assign n24180 = ~n16652 & n24179 ;
  assign n24181 = n906 & n24180 ;
  assign n24182 = n909 & ~n16016 ;
  assign n24183 = ~n16652 & n24182 ;
  assign n24184 = ~n906 & n24183 ;
  assign n24185 = ~n24181 & ~n24184 ;
  assign n24186 = \b[10]  & n17308 ;
  assign n24187 = n17305 & n24186 ;
  assign n24188 = ~\a[54]  & \b[11]  ;
  assign n24189 = n16647 & n24188 ;
  assign n24190 = ~n24187 & ~n24189 ;
  assign n24191 = \b[12]  & n16653 ;
  assign n24192 = \a[54]  & \b[11]  ;
  assign n24193 = n16644 & n24192 ;
  assign n24194 = \a[56]  & ~n24193 ;
  assign n24195 = ~n24191 & n24194 ;
  assign n24196 = n24190 & n24195 ;
  assign n24197 = n24185 & n24196 ;
  assign n24198 = ~n24191 & ~n24193 ;
  assign n24199 = n24190 & n24198 ;
  assign n24200 = n24185 & n24199 ;
  assign n24201 = ~\a[56]  & ~n24200 ;
  assign n24202 = ~n24197 & ~n24201 ;
  assign n24203 = n23492 & ~n23502 ;
  assign n24204 = ~n323 & ~n19861 ;
  assign n24205 = ~n20518 & n24204 ;
  assign n24206 = n320 & n24205 ;
  assign n24207 = n323 & ~n19861 ;
  assign n24208 = ~n20518 & n24207 ;
  assign n24209 = ~n320 & n24208 ;
  assign n24210 = ~n24206 & ~n24209 ;
  assign n24211 = \b[4]  & n21315 ;
  assign n24212 = n21312 & n24211 ;
  assign n24213 = \b[6]  & n20519 ;
  assign n24214 = \a[59]  & \b[5]  ;
  assign n24215 = n21313 & n24214 ;
  assign n24216 = ~\a[60]  & \b[5]  ;
  assign n24217 = n20513 & n24216 ;
  assign n24218 = ~n24215 & ~n24217 ;
  assign n24219 = ~n24213 & n24218 ;
  assign n24220 = ~n24212 & n24219 ;
  assign n24221 = n24210 & n24220 ;
  assign n24222 = \b[3]  & n21958 ;
  assign n24223 = \b[2]  & n21957 ;
  assign n24224 = ~\a[2]  & ~n24223 ;
  assign n24225 = ~n24222 & n24224 ;
  assign n24226 = \a[2]  & \b[3]  ;
  assign n24227 = n21958 & n24226 ;
  assign n24228 = \a[2]  & \b[2]  ;
  assign n24229 = n21957 & n24228 ;
  assign n24230 = ~\a[62]  & ~n24229 ;
  assign n24231 = ~n24227 & n24230 ;
  assign n24232 = ~n24225 & n24231 ;
  assign n24233 = ~n24221 & n24232 ;
  assign n24234 = \a[62]  & ~n24229 ;
  assign n24235 = ~n24227 & n24234 ;
  assign n24236 = ~n24225 & n24235 ;
  assign n24237 = n24220 & n24236 ;
  assign n24238 = n24210 & n24237 ;
  assign n24239 = ~n24233 & ~n24238 ;
  assign n24240 = ~\a[62]  & ~n24221 ;
  assign n24241 = ~n24227 & ~n24229 ;
  assign n24242 = ~n24225 & n24241 ;
  assign n24243 = \a[62]  & n24220 ;
  assign n24244 = n24210 & n24243 ;
  assign n24245 = ~n24242 & ~n24244 ;
  assign n24246 = ~n24240 & n24245 ;
  assign n24247 = n24239 & ~n24246 ;
  assign n24248 = ~n24203 & n24247 ;
  assign n24249 = n23492 & ~n24247 ;
  assign n24250 = ~n23502 & n24249 ;
  assign n24251 = ~n589 & n18516 ;
  assign n24252 = ~n587 & n24251 ;
  assign n24253 = \b[9]  & n18514 ;
  assign n24254 = \a[57]  & \b[8]  ;
  assign n24255 = n18505 & n24254 ;
  assign n24256 = ~n24253 & ~n24255 ;
  assign n24257 = \b[7]  & n19183 ;
  assign n24258 = n19180 & n24257 ;
  assign n24259 = ~\a[57]  & \b[8]  ;
  assign n24260 = n18508 & n24259 ;
  assign n24261 = ~n24258 & ~n24260 ;
  assign n24262 = n24256 & n24261 ;
  assign n24263 = ~n24252 & n24262 ;
  assign n24264 = ~\a[59]  & ~n24263 ;
  assign n24265 = \a[59]  & n24262 ;
  assign n24266 = ~n24252 & n24265 ;
  assign n24267 = ~n24264 & ~n24266 ;
  assign n24268 = ~n24250 & n24267 ;
  assign n24269 = ~n24248 & n24268 ;
  assign n24270 = ~n24248 & ~n24250 ;
  assign n24271 = ~n24267 & ~n24270 ;
  assign n24272 = ~n24269 & ~n24271 ;
  assign n24273 = n24202 & ~n24272 ;
  assign n24274 = n24178 & n24273 ;
  assign n24275 = n24202 & n24272 ;
  assign n24276 = ~n24178 & n24275 ;
  assign n24277 = ~n24274 & ~n24276 ;
  assign n24278 = ~n24202 & ~n24272 ;
  assign n24279 = ~n24178 & n24278 ;
  assign n24280 = ~n24202 & n24272 ;
  assign n24281 = n24178 & n24280 ;
  assign n24282 = ~n24279 & ~n24281 ;
  assign n24283 = n24277 & n24282 ;
  assign n24284 = ~n1233 & n14793 ;
  assign n24285 = ~n1231 & n24284 ;
  assign n24286 = \b[15]  & n14791 ;
  assign n24287 = \a[51]  & \b[14]  ;
  assign n24288 = n14782 & n24287 ;
  assign n24289 = ~n24286 & ~n24288 ;
  assign n24290 = \b[13]  & n15517 ;
  assign n24291 = n15514 & n24290 ;
  assign n24292 = ~\a[51]  & \b[14]  ;
  assign n24293 = n14785 & n24292 ;
  assign n24294 = ~n24291 & ~n24293 ;
  assign n24295 = n24289 & n24294 ;
  assign n24296 = ~n24285 & n24295 ;
  assign n24297 = ~\a[53]  & ~n24296 ;
  assign n24298 = \a[53]  & n24295 ;
  assign n24299 = ~n24285 & n24298 ;
  assign n24300 = ~n24297 & ~n24299 ;
  assign n24301 = ~n24283 & ~n24300 ;
  assign n24302 = ~n24176 & n24301 ;
  assign n24303 = n24283 & ~n24300 ;
  assign n24304 = n24176 & n24303 ;
  assign n24305 = ~n24302 & ~n24304 ;
  assign n24306 = ~n24283 & n24300 ;
  assign n24307 = n24176 & n24306 ;
  assign n24308 = n24283 & n24300 ;
  assign n24309 = ~n24176 & n24308 ;
  assign n24310 = ~n24307 & ~n24309 ;
  assign n24311 = n24305 & n24310 ;
  assign n24312 = n1875 & n13125 ;
  assign n24313 = ~n1872 & n24312 ;
  assign n24314 = ~n1875 & n13125 ;
  assign n24315 = ~n1689 & n24314 ;
  assign n24316 = ~n1871 & n24315 ;
  assign n24317 = \b[16]  & n13794 ;
  assign n24318 = n13792 & n24317 ;
  assign n24319 = ~\a[48]  & \b[17]  ;
  assign n24320 = n13117 & n24319 ;
  assign n24321 = ~n24318 & ~n24320 ;
  assign n24322 = \b[18]  & n13123 ;
  assign n24323 = \a[48]  & \b[17]  ;
  assign n24324 = n13786 & n24323 ;
  assign n24325 = \a[50]  & ~n24324 ;
  assign n24326 = ~n24322 & n24325 ;
  assign n24327 = n24321 & n24326 ;
  assign n24328 = ~n24316 & n24327 ;
  assign n24329 = ~n24313 & n24328 ;
  assign n24330 = ~n24322 & ~n24324 ;
  assign n24331 = n24321 & n24330 ;
  assign n24332 = ~n24316 & n24331 ;
  assign n24333 = ~n24313 & n24332 ;
  assign n24334 = ~\a[50]  & ~n24333 ;
  assign n24335 = ~n24329 & ~n24334 ;
  assign n24336 = ~n24311 & n24335 ;
  assign n24337 = n24173 & n24336 ;
  assign n24338 = n24311 & n24335 ;
  assign n24339 = ~n24173 & n24338 ;
  assign n24340 = ~n24337 & ~n24339 ;
  assign n24341 = ~n24173 & n24311 ;
  assign n24342 = ~n23569 & ~n24311 ;
  assign n24343 = ~n24172 & n24342 ;
  assign n24344 = ~n24335 & ~n24343 ;
  assign n24345 = ~n24341 & n24344 ;
  assign n24346 = n24340 & ~n24345 ;
  assign n24347 = ~n2523 & n11572 ;
  assign n24348 = ~n2521 & n24347 ;
  assign n24349 = \b[21]  & n11570 ;
  assign n24350 = \a[45]  & \b[20]  ;
  assign n24351 = n11561 & n24350 ;
  assign n24352 = ~n24349 & ~n24351 ;
  assign n24353 = \b[19]  & n12159 ;
  assign n24354 = n12156 & n24353 ;
  assign n24355 = ~\a[45]  & \b[20]  ;
  assign n24356 = n11564 & n24355 ;
  assign n24357 = ~n24354 & ~n24356 ;
  assign n24358 = n24352 & n24357 ;
  assign n24359 = ~n24348 & n24358 ;
  assign n24360 = ~\a[47]  & ~n24359 ;
  assign n24361 = \a[47]  & n24358 ;
  assign n24362 = ~n24348 & n24361 ;
  assign n24363 = ~n24360 & ~n24362 ;
  assign n24364 = ~n24346 & n24363 ;
  assign n24365 = ~n24171 & n24364 ;
  assign n24366 = n24346 & n24363 ;
  assign n24367 = n24171 & n24366 ;
  assign n24368 = ~n24365 & ~n24367 ;
  assign n24369 = ~n24346 & ~n24363 ;
  assign n24370 = n24171 & n24369 ;
  assign n24371 = n24346 & ~n24363 ;
  assign n24372 = ~n24171 & n24371 ;
  assign n24373 = ~n24370 & ~n24372 ;
  assign n24374 = n24368 & n24373 ;
  assign n24375 = n3283 & n10082 ;
  assign n24376 = ~n3280 & n24375 ;
  assign n24377 = ~n3283 & n10082 ;
  assign n24378 = ~n3017 & n24377 ;
  assign n24379 = ~n3279 & n24378 ;
  assign n24380 = \b[22]  & n10681 ;
  assign n24381 = n10678 & n24380 ;
  assign n24382 = ~\a[42]  & \b[23]  ;
  assign n24383 = n10074 & n24382 ;
  assign n24384 = ~n24381 & ~n24383 ;
  assign n24385 = \b[24]  & n10080 ;
  assign n24386 = \a[42]  & \b[23]  ;
  assign n24387 = n10071 & n24386 ;
  assign n24388 = \a[44]  & ~n24387 ;
  assign n24389 = ~n24385 & n24388 ;
  assign n24390 = n24384 & n24389 ;
  assign n24391 = ~n24379 & n24390 ;
  assign n24392 = ~n24376 & n24391 ;
  assign n24393 = ~n24385 & ~n24387 ;
  assign n24394 = n24384 & n24393 ;
  assign n24395 = ~n24379 & n24394 ;
  assign n24396 = ~n24376 & n24395 ;
  assign n24397 = ~\a[44]  & ~n24396 ;
  assign n24398 = ~n24392 & ~n24397 ;
  assign n24399 = n24374 & n24398 ;
  assign n24400 = ~n24168 & n24399 ;
  assign n24401 = ~n24374 & n24398 ;
  assign n24402 = n24168 & n24401 ;
  assign n24403 = ~n24400 & ~n24402 ;
  assign n24404 = ~n24374 & ~n24398 ;
  assign n24405 = ~n24168 & n24404 ;
  assign n24406 = n24374 & ~n24398 ;
  assign n24407 = n24168 & n24406 ;
  assign n24408 = ~n24405 & ~n24407 ;
  assign n24409 = n24403 & n24408 ;
  assign n24410 = ~n4145 & n8759 ;
  assign n24411 = ~n3603 & n8759 ;
  assign n24412 = ~n4141 & n24411 ;
  assign n24413 = ~n24410 & ~n24412 ;
  assign n24414 = ~n4148 & ~n24413 ;
  assign n24415 = \b[25]  & n9301 ;
  assign n24416 = n9298 & n24415 ;
  assign n24417 = ~\a[39]  & \b[26]  ;
  assign n24418 = n8751 & n24417 ;
  assign n24419 = ~n24416 & ~n24418 ;
  assign n24420 = \b[27]  & n8757 ;
  assign n24421 = \a[39]  & \b[26]  ;
  assign n24422 = n8748 & n24421 ;
  assign n24423 = \a[41]  & ~n24422 ;
  assign n24424 = ~n24420 & n24423 ;
  assign n24425 = n24419 & n24424 ;
  assign n24426 = ~n24414 & n24425 ;
  assign n24427 = ~n24420 & ~n24422 ;
  assign n24428 = n24419 & n24427 ;
  assign n24429 = ~\a[41]  & ~n24428 ;
  assign n24430 = ~\a[41]  & ~n4148 ;
  assign n24431 = ~n24413 & n24430 ;
  assign n24432 = ~n24429 & ~n24431 ;
  assign n24433 = ~n24426 & n24432 ;
  assign n24434 = ~n24409 & ~n24433 ;
  assign n24435 = n24167 & n24434 ;
  assign n24436 = n24409 & ~n24433 ;
  assign n24437 = ~n24167 & n24436 ;
  assign n24438 = ~n24435 & ~n24437 ;
  assign n24439 = ~n24409 & n24433 ;
  assign n24440 = ~n24167 & n24439 ;
  assign n24441 = n24409 & n24433 ;
  assign n24442 = n24167 & n24441 ;
  assign n24443 = ~n24440 & ~n24442 ;
  assign n24444 = n24438 & n24443 ;
  assign n24445 = ~n5105 & ~n7098 ;
  assign n24446 = ~n7531 & n24445 ;
  assign n24447 = n5102 & n24446 ;
  assign n24448 = n5105 & ~n7098 ;
  assign n24449 = ~n7531 & n24448 ;
  assign n24450 = ~n5102 & n24449 ;
  assign n24451 = ~n24447 & ~n24450 ;
  assign n24452 = \b[28]  & n7973 ;
  assign n24453 = n7970 & n24452 ;
  assign n24454 = ~\a[36]  & \b[29]  ;
  assign n24455 = n7526 & n24454 ;
  assign n24456 = ~n24453 & ~n24455 ;
  assign n24457 = \b[30]  & n7532 ;
  assign n24458 = \a[36]  & \b[29]  ;
  assign n24459 = n17801 & n24458 ;
  assign n24460 = \a[38]  & ~n24459 ;
  assign n24461 = ~n24457 & n24460 ;
  assign n24462 = n24456 & n24461 ;
  assign n24463 = n24451 & n24462 ;
  assign n24464 = ~n24457 & ~n24459 ;
  assign n24465 = n24456 & n24464 ;
  assign n24466 = n24451 & n24465 ;
  assign n24467 = ~\a[38]  & ~n24466 ;
  assign n24468 = ~n24463 & ~n24467 ;
  assign n24469 = ~n24444 & n24468 ;
  assign n24470 = n24164 & n24469 ;
  assign n24471 = n24444 & n24468 ;
  assign n24472 = ~n24164 & n24471 ;
  assign n24473 = ~n24470 & ~n24472 ;
  assign n24474 = ~n24164 & n24444 ;
  assign n24475 = n23655 & ~n24444 ;
  assign n24476 = ~n24163 & n24475 ;
  assign n24477 = ~n24468 & ~n24476 ;
  assign n24478 = ~n24474 & n24477 ;
  assign n24479 = n24473 & ~n24478 ;
  assign n24480 = ~n5852 & n6309 ;
  assign n24481 = ~n5809 & n6309 ;
  assign n24482 = ~n5848 & n24481 ;
  assign n24483 = ~n24480 & ~n24482 ;
  assign n24484 = ~n5855 & ~n24483 ;
  assign n24485 = \b[31]  & n6778 ;
  assign n24486 = n6775 & n24485 ;
  assign n24487 = ~\a[33]  & \b[32]  ;
  assign n24488 = n6301 & n24487 ;
  assign n24489 = ~n24486 & ~n24488 ;
  assign n24490 = \b[33]  & n6307 ;
  assign n24491 = \a[33]  & \b[32]  ;
  assign n24492 = n6298 & n24491 ;
  assign n24493 = \a[35]  & ~n24492 ;
  assign n24494 = ~n24490 & n24493 ;
  assign n24495 = n24489 & n24494 ;
  assign n24496 = ~n24484 & n24495 ;
  assign n24497 = ~n24490 & ~n24492 ;
  assign n24498 = n24489 & n24497 ;
  assign n24499 = ~\a[35]  & ~n24498 ;
  assign n24500 = ~\a[35]  & ~n5855 ;
  assign n24501 = ~n24483 & n24500 ;
  assign n24502 = ~n24499 & ~n24501 ;
  assign n24503 = ~n24496 & n24502 ;
  assign n24504 = ~n24479 & n24503 ;
  assign n24505 = ~n24162 & n24504 ;
  assign n24506 = n24479 & n24503 ;
  assign n24507 = n24162 & n24506 ;
  assign n24508 = ~n24505 & ~n24507 ;
  assign n24509 = n24479 & ~n24503 ;
  assign n24510 = ~n24162 & n24509 ;
  assign n24511 = ~n24479 & ~n24503 ;
  assign n24512 = n24162 & n24511 ;
  assign n24513 = ~n24510 & ~n24512 ;
  assign n24514 = n24508 & n24513 ;
  assign n24515 = ~n24159 & n24514 ;
  assign n24516 = n24135 & n24515 ;
  assign n24517 = n24159 & n24514 ;
  assign n24518 = ~n24135 & n24517 ;
  assign n24519 = ~n24516 & ~n24518 ;
  assign n24520 = ~n24159 & ~n24514 ;
  assign n24521 = ~n24135 & n24520 ;
  assign n24522 = n24159 & ~n24514 ;
  assign n24523 = n24135 & n24522 ;
  assign n24524 = ~n24521 & ~n24523 ;
  assign n24525 = n24519 & n24524 ;
  assign n24526 = ~n24134 & n24525 ;
  assign n24527 = ~n24132 & n24526 ;
  assign n24528 = ~n24131 & ~n24159 ;
  assign n24529 = ~n24514 & n24528 ;
  assign n24530 = ~n24135 & n24529 ;
  assign n24531 = ~n24131 & n24159 ;
  assign n24532 = n24514 & n24531 ;
  assign n24533 = ~n24135 & n24532 ;
  assign n24534 = ~n24530 & ~n24533 ;
  assign n24535 = ~n24514 & n24531 ;
  assign n24536 = n24135 & n24535 ;
  assign n24537 = n24514 & n24528 ;
  assign n24538 = n24135 & n24537 ;
  assign n24539 = ~n24536 & ~n24538 ;
  assign n24540 = n24534 & n24539 ;
  assign n24541 = n24112 & ~n24540 ;
  assign n24542 = n24131 & ~n24525 ;
  assign n24543 = ~n24112 & n24542 ;
  assign n24544 = ~n24541 & ~n24543 ;
  assign n24545 = ~n24527 & n24544 ;
  assign n24546 = ~n24109 & ~n24545 ;
  assign n24547 = ~n24085 & n24546 ;
  assign n24548 = n24109 & n24545 ;
  assign n24549 = ~n24085 & n24548 ;
  assign n24550 = n23765 & ~n24109 ;
  assign n24551 = n24545 & n24550 ;
  assign n24552 = ~n23774 & n24551 ;
  assign n24553 = n23765 & n24109 ;
  assign n24554 = ~n24545 & n24553 ;
  assign n24555 = ~n23774 & n24554 ;
  assign n24556 = ~n24552 & ~n24555 ;
  assign n24557 = ~n24549 & n24556 ;
  assign n24558 = ~n24547 & n24557 ;
  assign n24559 = ~n24084 & n24558 ;
  assign n24560 = ~n24082 & n24559 ;
  assign n24561 = n24084 & ~n24558 ;
  assign n24562 = n24081 & ~n24558 ;
  assign n24563 = ~n24062 & n24562 ;
  assign n24564 = ~n24561 & ~n24563 ;
  assign n24565 = ~n24560 & n24564 ;
  assign n24566 = ~n24059 & ~n24565 ;
  assign n24567 = ~n24035 & n24566 ;
  assign n24568 = n24059 & n24565 ;
  assign n24569 = ~n24035 & n24568 ;
  assign n24570 = n23804 & ~n24059 ;
  assign n24571 = n24565 & n24570 ;
  assign n24572 = ~n24034 & n24571 ;
  assign n24573 = n23804 & n24059 ;
  assign n24574 = ~n24565 & n24573 ;
  assign n24575 = ~n24034 & n24574 ;
  assign n24576 = ~n24572 & ~n24575 ;
  assign n24577 = ~n24569 & n24576 ;
  assign n24578 = ~n24567 & n24577 ;
  assign n24579 = n999 & ~n16398 ;
  assign n24580 = ~n15241 & n24579 ;
  assign n24581 = ~n16404 & n24580 ;
  assign n24582 = n999 & n16398 ;
  assign n24583 = n15241 & n24582 ;
  assign n24584 = n16400 & n24582 ;
  assign n24585 = ~n15239 & n24584 ;
  assign n24586 = ~n24583 & ~n24585 ;
  assign n24587 = ~n24581 & n24586 ;
  assign n24588 = \b[52]  & n1182 ;
  assign n24589 = n1179 & n24588 ;
  assign n24590 = \b[54]  & n997 ;
  assign n24591 = \a[11]  & \b[53]  ;
  assign n24592 = n1180 & n24591 ;
  assign n24593 = ~\a[12]  & \b[53]  ;
  assign n24594 = n7674 & n24593 ;
  assign n24595 = ~n24592 & ~n24594 ;
  assign n24596 = ~n24590 & n24595 ;
  assign n24597 = ~n24589 & n24596 ;
  assign n24598 = n24587 & n24597 ;
  assign n24599 = ~\a[14]  & ~n24598 ;
  assign n24600 = \a[14]  & n24597 ;
  assign n24601 = n24587 & n24600 ;
  assign n24602 = ~n24599 & ~n24601 ;
  assign n24603 = n1467 & ~n14098 ;
  assign n24604 = ~n14096 & n24603 ;
  assign n24605 = \b[49]  & n1652 ;
  assign n24606 = n1649 & n24605 ;
  assign n24607 = ~\a[15]  & \b[50]  ;
  assign n24608 = n1459 & n24607 ;
  assign n24609 = ~n24606 & ~n24608 ;
  assign n24610 = \b[51]  & n1465 ;
  assign n24611 = \a[15]  & \b[50]  ;
  assign n24612 = n1456 & n24611 ;
  assign n24613 = \a[17]  & ~n24612 ;
  assign n24614 = ~n24610 & n24613 ;
  assign n24615 = n24609 & n24614 ;
  assign n24616 = ~n24604 & n24615 ;
  assign n24617 = ~n24610 & ~n24612 ;
  assign n24618 = n24609 & n24617 ;
  assign n24619 = ~n24604 & n24618 ;
  assign n24620 = ~\a[17]  & ~n24619 ;
  assign n24621 = ~n24616 & ~n24620 ;
  assign n24622 = n24602 & n24621 ;
  assign n24623 = ~n24578 & n24622 ;
  assign n24624 = ~n24033 & n24623 ;
  assign n24625 = n24602 & ~n24621 ;
  assign n24626 = n24578 & n24625 ;
  assign n24627 = ~n24033 & n24626 ;
  assign n24628 = ~n24624 & ~n24627 ;
  assign n24629 = ~n24578 & n24625 ;
  assign n24630 = n24033 & n24629 ;
  assign n24631 = n24578 & n24622 ;
  assign n24632 = n24033 & n24631 ;
  assign n24633 = ~n24630 & ~n24632 ;
  assign n24634 = n24628 & n24633 ;
  assign n24635 = ~n24602 & ~n24621 ;
  assign n24636 = ~n24578 & n24635 ;
  assign n24637 = ~n24033 & n24636 ;
  assign n24638 = ~n24602 & n24621 ;
  assign n24639 = n24578 & n24638 ;
  assign n24640 = ~n24033 & n24639 ;
  assign n24641 = ~n24637 & ~n24640 ;
  assign n24642 = ~n24578 & n24638 ;
  assign n24643 = n24033 & n24642 ;
  assign n24644 = n24578 & n24635 ;
  assign n24645 = n24033 & n24644 ;
  assign n24646 = ~n24643 & ~n24645 ;
  assign n24647 = n24641 & n24646 ;
  assign n24648 = n24634 & n24647 ;
  assign n24649 = ~n24030 & ~n24648 ;
  assign n24650 = n24030 & n24648 ;
  assign n24651 = ~n24649 & ~n24650 ;
  assign n24652 = n646 & ~n17690 ;
  assign n24653 = ~n17688 & n24652 ;
  assign n24654 = \b[55]  & n796 ;
  assign n24655 = n793 & n24654 ;
  assign n24656 = ~\a[9]  & \b[56]  ;
  assign n24657 = n638 & n24656 ;
  assign n24658 = ~n24655 & ~n24657 ;
  assign n24659 = \b[57]  & n644 ;
  assign n24660 = \a[9]  & \b[56]  ;
  assign n24661 = n635 & n24660 ;
  assign n24662 = \a[11]  & ~n24661 ;
  assign n24663 = ~n24659 & n24662 ;
  assign n24664 = n24658 & n24663 ;
  assign n24665 = ~n24653 & n24664 ;
  assign n24666 = ~n24659 & ~n24661 ;
  assign n24667 = n24658 & n24666 ;
  assign n24668 = ~n24653 & n24667 ;
  assign n24669 = ~\a[11]  & ~n24668 ;
  assign n24670 = ~n24665 & ~n24669 ;
  assign n24671 = n23859 & ~n24670 ;
  assign n24672 = ~n24651 & n24671 ;
  assign n24673 = ~n24028 & n24672 ;
  assign n24674 = n23859 & ~n24028 ;
  assign n24675 = ~n24651 & n24670 ;
  assign n24676 = ~n24674 & n24675 ;
  assign n24677 = ~n24673 & ~n24676 ;
  assign n24678 = ~n24028 & n24671 ;
  assign n24679 = n24651 & ~n24670 ;
  assign n24680 = n23859 & n24651 ;
  assign n24681 = ~n24028 & n24680 ;
  assign n24682 = ~n24679 & ~n24681 ;
  assign n24683 = ~n24678 & ~n24682 ;
  assign n24684 = n24677 & ~n24683 ;
  assign n24685 = ~n24026 & n24684 ;
  assign n24686 = ~n24024 & n24685 ;
  assign n24687 = ~n24024 & ~n24026 ;
  assign n24688 = ~n24684 & ~n24687 ;
  assign n24689 = ~n24686 & ~n24688 ;
  assign n24690 = n252 & ~n22461 ;
  assign n24691 = ~n22459 & n24690 ;
  assign n24692 = \b[63]  & n250 ;
  assign n24693 = \a[3]  & \b[62]  ;
  assign n24694 = n241 & n24693 ;
  assign n24695 = ~n24692 & ~n24694 ;
  assign n24696 = \b[61]  & n303 ;
  assign n24697 = n300 & n24696 ;
  assign n24698 = ~\a[3]  & \b[62]  ;
  assign n24699 = n244 & n24698 ;
  assign n24700 = ~n24697 & ~n24699 ;
  assign n24701 = n24695 & n24700 ;
  assign n24702 = ~n24691 & n24701 ;
  assign n24703 = ~\a[5]  & ~n24702 ;
  assign n24704 = \a[5]  & n24701 ;
  assign n24705 = ~n24691 & n24704 ;
  assign n24706 = ~n24703 & ~n24705 ;
  assign n24707 = n23951 & ~n23980 ;
  assign n24708 = n24706 & ~n24707 ;
  assign n24709 = ~n24706 & n24707 ;
  assign n24710 = ~n24708 & ~n24709 ;
  assign n24711 = ~n24689 & n24710 ;
  assign n24712 = n24689 & n24708 ;
  assign n24713 = n24689 & n24709 ;
  assign n24714 = ~n24712 & ~n24713 ;
  assign n24715 = ~n24711 & n24714 ;
  assign n24716 = ~n23285 & n23982 ;
  assign n24717 = ~n23287 & ~n24716 ;
  assign n24718 = ~n24715 & ~n24717 ;
  assign n24719 = n24715 & n24717 ;
  assign n24720 = ~n24718 & ~n24719 ;
  assign n24721 = ~n23987 & n24720 ;
  assign n24722 = ~n23989 & n24721 ;
  assign n24723 = ~n23990 & n24722 ;
  assign n24724 = ~n23987 & ~n23989 ;
  assign n24725 = ~n23990 & n24724 ;
  assign n24726 = ~n24720 & ~n24725 ;
  assign n24727 = ~n24723 & ~n24726 ;
  assign n24728 = ~n23987 & ~n24719 ;
  assign n24729 = ~n23989 & n24728 ;
  assign n24730 = ~n23990 & n24729 ;
  assign n24731 = ~n24689 & ~n24708 ;
  assign n24732 = ~n24709 & ~n24731 ;
  assign n24733 = n23820 & ~n24621 ;
  assign n24734 = ~n24032 & n24733 ;
  assign n24735 = ~n24033 & n24621 ;
  assign n24736 = n24578 & ~n24734 ;
  assign n24737 = ~n24735 & n24736 ;
  assign n24738 = ~n24734 & ~n24737 ;
  assign n24739 = n999 & ~n16446 ;
  assign n24740 = ~n16444 & n24739 ;
  assign n24741 = \b[53]  & n1182 ;
  assign n24742 = n1179 & n24741 ;
  assign n24743 = \b[55]  & n997 ;
  assign n24744 = \a[11]  & \b[54]  ;
  assign n24745 = n1180 & n24744 ;
  assign n24746 = ~\a[12]  & \b[54]  ;
  assign n24747 = n7674 & n24746 ;
  assign n24748 = ~n24745 & ~n24747 ;
  assign n24749 = ~n24743 & n24748 ;
  assign n24750 = ~n24742 & n24749 ;
  assign n24751 = ~n24740 & n24750 ;
  assign n24752 = \a[14]  & ~n24751 ;
  assign n24753 = ~\a[14]  & n24751 ;
  assign n24754 = ~n24752 & ~n24753 ;
  assign n24755 = ~n24738 & n24754 ;
  assign n24756 = ~\a[14]  & ~n24751 ;
  assign n24757 = \a[14]  & n24750 ;
  assign n24758 = ~n24740 & n24757 ;
  assign n24759 = ~n24756 & ~n24758 ;
  assign n24760 = ~n24734 & n24759 ;
  assign n24761 = ~n24737 & n24760 ;
  assign n24762 = ~n23804 & ~n24059 ;
  assign n24763 = n23810 & ~n24059 ;
  assign n24764 = n23325 & n24763 ;
  assign n24765 = ~n24762 & ~n24764 ;
  assign n24766 = ~n24572 & n24765 ;
  assign n24767 = ~n24569 & n24766 ;
  assign n24768 = n1467 & n15201 ;
  assign n24769 = ~n15198 & n24768 ;
  assign n24770 = n1467 & ~n15201 ;
  assign n24771 = ~n14093 & n24770 ;
  assign n24772 = ~n15197 & n24771 ;
  assign n24773 = \b[52]  & n1465 ;
  assign n24774 = \a[15]  & \b[51]  ;
  assign n24775 = n1456 & n24774 ;
  assign n24776 = ~n24773 & ~n24775 ;
  assign n24777 = \b[50]  & n1652 ;
  assign n24778 = n1649 & n24777 ;
  assign n24779 = ~\a[15]  & \b[51]  ;
  assign n24780 = n1459 & n24779 ;
  assign n24781 = ~n24778 & ~n24780 ;
  assign n24782 = n24776 & n24781 ;
  assign n24783 = ~n24772 & n24782 ;
  assign n24784 = ~n24769 & n24783 ;
  assign n24785 = \a[17]  & ~n24784 ;
  assign n24786 = ~\a[17]  & n24784 ;
  assign n24787 = ~n24785 & ~n24786 ;
  assign n24788 = ~n24767 & n24787 ;
  assign n24789 = ~\a[17]  & ~n24784 ;
  assign n24790 = \a[17]  & n24782 ;
  assign n24791 = ~n24772 & n24790 ;
  assign n24792 = ~n24769 & n24791 ;
  assign n24793 = ~n24789 & ~n24792 ;
  assign n24794 = n24767 & n24793 ;
  assign n24795 = ~n24788 & ~n24794 ;
  assign n24796 = n1965 & ~n13524 ;
  assign n24797 = ~n13522 & n24796 ;
  assign n24798 = \b[49]  & n1963 ;
  assign n24799 = \a[18]  & \b[48]  ;
  assign n24800 = n2210 & n24799 ;
  assign n24801 = ~n24798 & ~n24800 ;
  assign n24802 = \b[47]  & n2218 ;
  assign n24803 = n2216 & n24802 ;
  assign n24804 = ~\a[18]  & \b[48]  ;
  assign n24805 = n1957 & n24804 ;
  assign n24806 = ~n24803 & ~n24805 ;
  assign n24807 = n24801 & n24806 ;
  assign n24808 = ~n24797 & n24807 ;
  assign n24809 = ~\a[20]  & ~n24808 ;
  assign n24810 = \a[20]  & n24807 ;
  assign n24811 = ~n24797 & n24810 ;
  assign n24812 = ~n24809 & ~n24811 ;
  assign n24813 = ~n24084 & n24812 ;
  assign n24814 = ~n24560 & n24813 ;
  assign n24815 = ~n24084 & ~n24560 ;
  assign n24816 = \a[20]  & ~n24808 ;
  assign n24817 = ~\a[20]  & n24808 ;
  assign n24818 = ~n24816 & ~n24817 ;
  assign n24819 = ~n24815 & n24818 ;
  assign n24820 = ~n24814 & ~n24819 ;
  assign n24821 = ~n24549 & ~n24552 ;
  assign n24822 = ~n24085 & ~n24109 ;
  assign n24823 = n24821 & ~n24822 ;
  assign n24824 = n2622 & n11906 ;
  assign n24825 = ~n11903 & n24824 ;
  assign n24826 = n2622 & ~n11906 ;
  assign n24827 = ~n11392 & n24826 ;
  assign n24828 = ~n11902 & n24827 ;
  assign n24829 = \b[46]  & n2620 ;
  assign n24830 = \a[21]  & \b[45]  ;
  assign n24831 = n20849 & n24830 ;
  assign n24832 = ~n24829 & ~n24831 ;
  assign n24833 = \b[44]  & n2912 ;
  assign n24834 = n2909 & n24833 ;
  assign n24835 = ~\a[21]  & \b[45]  ;
  assign n24836 = n2614 & n24835 ;
  assign n24837 = ~n24834 & ~n24836 ;
  assign n24838 = n24832 & n24837 ;
  assign n24839 = ~n24828 & n24838 ;
  assign n24840 = ~n24825 & n24839 ;
  assign n24841 = \a[23]  & ~n24840 ;
  assign n24842 = ~\a[23]  & n24840 ;
  assign n24843 = ~n24841 & ~n24842 ;
  assign n24844 = ~n24823 & n24843 ;
  assign n24845 = ~n24134 & ~n24527 ;
  assign n24846 = n3402 & ~n10409 ;
  assign n24847 = ~n10407 & n24846 ;
  assign n24848 = \b[43]  & n3400 ;
  assign n24849 = \a[24]  & \b[42]  ;
  assign n24850 = n3391 & n24849 ;
  assign n24851 = ~n24848 & ~n24850 ;
  assign n24852 = \b[41]  & n3733 ;
  assign n24853 = n3730 & n24852 ;
  assign n24854 = ~\a[24]  & \b[42]  ;
  assign n24855 = n3394 & n24854 ;
  assign n24856 = ~n24853 & ~n24855 ;
  assign n24857 = n24851 & n24856 ;
  assign n24858 = ~n24847 & n24857 ;
  assign n24859 = \a[26]  & ~n24858 ;
  assign n24860 = ~\a[26]  & n24858 ;
  assign n24861 = ~n24859 & ~n24860 ;
  assign n24862 = ~n24845 & n24861 ;
  assign n24863 = ~\a[26]  & ~n24858 ;
  assign n24864 = \a[26]  & n24857 ;
  assign n24865 = ~n24847 & n24864 ;
  assign n24866 = ~n24863 & ~n24865 ;
  assign n24867 = ~n24134 & n24866 ;
  assign n24868 = ~n24527 & n24867 ;
  assign n24869 = n23724 & ~n24159 ;
  assign n24870 = n23729 & ~n24159 ;
  assign n24871 = n23389 & n24870 ;
  assign n24872 = ~n24869 & ~n24871 ;
  assign n24873 = n24519 & n24872 ;
  assign n24874 = n4249 & n9044 ;
  assign n24875 = ~n9041 & n24874 ;
  assign n24876 = n4249 & ~n9044 ;
  assign n24877 = ~n8597 & n24876 ;
  assign n24878 = ~n9040 & n24877 ;
  assign n24879 = \b[40]  & n4247 ;
  assign n24880 = \a[27]  & \b[39]  ;
  assign n24881 = n4238 & n24880 ;
  assign n24882 = ~n24879 & ~n24881 ;
  assign n24883 = \b[38]  & n4647 ;
  assign n24884 = n4644 & n24883 ;
  assign n24885 = ~\a[27]  & \b[39]  ;
  assign n24886 = n4241 & n24885 ;
  assign n24887 = ~n24884 & ~n24886 ;
  assign n24888 = n24882 & n24887 ;
  assign n24889 = ~n24878 & n24888 ;
  assign n24890 = ~n24875 & n24889 ;
  assign n24891 = \a[29]  & ~n24890 ;
  assign n24892 = ~\a[29]  & n24890 ;
  assign n24893 = ~n24891 & ~n24892 ;
  assign n24894 = ~n24873 & n24893 ;
  assign n24895 = n24162 & n24479 ;
  assign n24896 = ~n24162 & ~n24479 ;
  assign n24897 = ~n24503 & ~n24896 ;
  assign n24898 = ~n24895 & ~n24897 ;
  assign n24899 = n5211 & ~n7761 ;
  assign n24900 = ~n7759 & n24899 ;
  assign n24901 = \b[37]  & n5209 ;
  assign n24902 = \a[30]  & \b[36]  ;
  assign n24903 = n5200 & n24902 ;
  assign n24904 = ~n24901 & ~n24903 ;
  assign n24905 = \b[35]  & n5595 ;
  assign n24906 = n5592 & n24905 ;
  assign n24907 = ~\a[30]  & \b[36]  ;
  assign n24908 = n5203 & n24907 ;
  assign n24909 = ~n24906 & ~n24908 ;
  assign n24910 = n24904 & n24909 ;
  assign n24911 = ~n24900 & n24910 ;
  assign n24912 = \a[32]  & ~n24911 ;
  assign n24913 = ~\a[32]  & n24911 ;
  assign n24914 = ~n24912 & ~n24913 ;
  assign n24915 = ~n24898 & n24914 ;
  assign n24916 = ~\a[32]  & ~n24911 ;
  assign n24917 = \a[32]  & n24910 ;
  assign n24918 = ~n24900 & n24917 ;
  assign n24919 = ~n24916 & ~n24918 ;
  assign n24920 = ~n24895 & n24919 ;
  assign n24921 = ~n24897 & n24920 ;
  assign n24922 = ~n24915 & ~n24921 ;
  assign n24923 = n23655 & n24468 ;
  assign n24924 = ~n24163 & n24923 ;
  assign n24925 = ~n24469 & ~n24924 ;
  assign n24926 = ~n24476 & n24925 ;
  assign n24927 = ~n5952 & ~n6565 ;
  assign n24928 = ~n6306 & n24927 ;
  assign n24929 = n6562 & n24928 ;
  assign n24930 = ~n5952 & n6565 ;
  assign n24931 = ~n6306 & n24930 ;
  assign n24932 = ~n6562 & n24931 ;
  assign n24933 = ~n24929 & ~n24932 ;
  assign n24934 = \b[32]  & n6778 ;
  assign n24935 = n6775 & n24934 ;
  assign n24936 = ~\a[33]  & \b[33]  ;
  assign n24937 = n6301 & n24936 ;
  assign n24938 = ~n24935 & ~n24937 ;
  assign n24939 = \b[34]  & n6307 ;
  assign n24940 = \a[33]  & \b[33]  ;
  assign n24941 = n6298 & n24940 ;
  assign n24942 = \a[35]  & ~n24941 ;
  assign n24943 = ~n24939 & n24942 ;
  assign n24944 = n24938 & n24943 ;
  assign n24945 = n24933 & n24944 ;
  assign n24946 = ~n24939 & ~n24941 ;
  assign n24947 = n24938 & n24946 ;
  assign n24948 = n24933 & n24947 ;
  assign n24949 = ~\a[35]  & ~n24948 ;
  assign n24950 = ~n24945 & ~n24949 ;
  assign n24951 = ~n24168 & n24374 ;
  assign n24952 = n24168 & ~n24374 ;
  assign n24953 = ~n24398 & ~n24952 ;
  assign n24954 = ~n24951 & ~n24953 ;
  assign n24955 = n24171 & n24346 ;
  assign n24956 = n24373 & ~n24955 ;
  assign n24957 = ~n23569 & n24335 ;
  assign n24958 = ~n24172 & n24957 ;
  assign n24959 = ~n24336 & ~n24958 ;
  assign n24960 = ~n24343 & n24959 ;
  assign n24961 = ~n24238 & n24241 ;
  assign n24962 = ~n24233 & n24961 ;
  assign n24963 = \b[5]  & n21315 ;
  assign n24964 = n21312 & n24963 ;
  assign n24965 = \b[7]  & n20519 ;
  assign n24966 = \a[59]  & \b[6]  ;
  assign n24967 = n21313 & n24966 ;
  assign n24968 = ~\a[60]  & \b[6]  ;
  assign n24969 = n20513 & n24968 ;
  assign n24970 = ~n24967 & ~n24969 ;
  assign n24971 = ~n24965 & n24970 ;
  assign n24972 = ~n24964 & n24971 ;
  assign n24973 = \b[4]  & n21958 ;
  assign n24974 = \b[3]  & n21957 ;
  assign n24975 = ~\a[2]  & ~n24974 ;
  assign n24976 = ~n24973 & n24975 ;
  assign n24977 = \a[2]  & \b[4]  ;
  assign n24978 = n21958 & n24977 ;
  assign n24979 = n21957 & n24226 ;
  assign n24980 = ~\a[62]  & ~n24979 ;
  assign n24981 = ~n24978 & n24980 ;
  assign n24982 = ~n24976 & n24981 ;
  assign n24983 = ~n24972 & n24982 ;
  assign n24984 = ~n380 & n20521 ;
  assign n24985 = ~n322 & n20521 ;
  assign n24986 = ~n326 & n24985 ;
  assign n24987 = ~n24984 & ~n24986 ;
  assign n24988 = ~n383 & n24982 ;
  assign n24989 = ~n24987 & n24988 ;
  assign n24990 = ~n24983 & ~n24989 ;
  assign n24991 = ~n383 & ~n24987 ;
  assign n24992 = \a[62]  & ~n24979 ;
  assign n24993 = ~n24978 & n24992 ;
  assign n24994 = ~n24976 & n24993 ;
  assign n24995 = n24972 & n24994 ;
  assign n24996 = ~n24991 & n24995 ;
  assign n24997 = n24990 & ~n24996 ;
  assign n24998 = ~\a[62]  & ~n24972 ;
  assign n24999 = ~\a[62]  & ~n383 ;
  assign n25000 = ~n24987 & n24999 ;
  assign n25001 = ~n24998 & ~n25000 ;
  assign n25002 = ~n24978 & ~n24979 ;
  assign n25003 = ~n24976 & n25002 ;
  assign n25004 = \a[62]  & n24972 ;
  assign n25005 = ~n24991 & n25004 ;
  assign n25006 = ~n25003 & ~n25005 ;
  assign n25007 = n25001 & n25006 ;
  assign n25008 = n24997 & ~n25007 ;
  assign n25009 = n24962 & ~n25008 ;
  assign n25010 = ~n24962 & n24997 ;
  assign n25011 = ~n25007 & n25010 ;
  assign n25012 = ~n25009 & ~n25011 ;
  assign n25013 = n685 & n18516 ;
  assign n25014 = ~n682 & n25013 ;
  assign n25015 = ~n685 & n18516 ;
  assign n25016 = ~n584 & n25015 ;
  assign n25017 = ~n681 & n25016 ;
  assign n25018 = \b[8]  & n19183 ;
  assign n25019 = n19180 & n25018 ;
  assign n25020 = ~\a[57]  & \b[9]  ;
  assign n25021 = n18508 & n25020 ;
  assign n25022 = ~n25019 & ~n25021 ;
  assign n25023 = \b[10]  & n18514 ;
  assign n25024 = \a[57]  & \b[9]  ;
  assign n25025 = n18505 & n25024 ;
  assign n25026 = \a[59]  & ~n25025 ;
  assign n25027 = ~n25023 & n25026 ;
  assign n25028 = n25022 & n25027 ;
  assign n25029 = ~n25017 & n25028 ;
  assign n25030 = ~n25014 & n25029 ;
  assign n25031 = ~n25023 & ~n25025 ;
  assign n25032 = n25022 & n25031 ;
  assign n25033 = ~n25017 & n25032 ;
  assign n25034 = ~n25014 & n25033 ;
  assign n25035 = ~\a[59]  & ~n25034 ;
  assign n25036 = ~n25030 & ~n25035 ;
  assign n25037 = n25012 & ~n25036 ;
  assign n25038 = ~n25012 & n25036 ;
  assign n25039 = ~n25037 & ~n25038 ;
  assign n25040 = ~n24248 & n24267 ;
  assign n25041 = ~n24250 & ~n25040 ;
  assign n25042 = ~n25039 & ~n25041 ;
  assign n25043 = n25039 & n25041 ;
  assign n25044 = ~n25042 & ~n25043 ;
  assign n25045 = ~n948 & n16655 ;
  assign n25046 = ~n908 & n16655 ;
  assign n25047 = ~n912 & n25046 ;
  assign n25048 = ~n25045 & ~n25047 ;
  assign n25049 = ~n951 & ~n25048 ;
  assign n25050 = \b[11]  & n17308 ;
  assign n25051 = n17305 & n25050 ;
  assign n25052 = ~\a[54]  & \b[12]  ;
  assign n25053 = n16647 & n25052 ;
  assign n25054 = ~n25051 & ~n25053 ;
  assign n25055 = \b[13]  & n16653 ;
  assign n25056 = \a[54]  & \b[12]  ;
  assign n25057 = n16644 & n25056 ;
  assign n25058 = \a[56]  & ~n25057 ;
  assign n25059 = ~n25055 & n25058 ;
  assign n25060 = n25054 & n25059 ;
  assign n25061 = ~n25049 & n25060 ;
  assign n25062 = ~n25055 & ~n25057 ;
  assign n25063 = n25054 & n25062 ;
  assign n25064 = ~\a[56]  & ~n25063 ;
  assign n25065 = ~\a[56]  & ~n951 ;
  assign n25066 = ~n25048 & n25065 ;
  assign n25067 = ~n25064 & ~n25066 ;
  assign n25068 = ~n25061 & n25067 ;
  assign n25069 = ~n25044 & n25068 ;
  assign n25070 = n25044 & ~n25068 ;
  assign n25071 = ~n25069 & ~n25070 ;
  assign n25072 = n24178 & n24272 ;
  assign n25073 = ~n23528 & n24202 ;
  assign n25074 = ~n24177 & n25073 ;
  assign n25075 = ~n24275 & ~n25074 ;
  assign n25076 = ~n25072 & n25075 ;
  assign n25077 = n25071 & n25076 ;
  assign n25078 = ~n25071 & ~n25076 ;
  assign n25079 = ~n25077 & ~n25078 ;
  assign n25080 = n1512 & n14793 ;
  assign n25081 = ~n1509 & n25080 ;
  assign n25082 = ~n1512 & n14793 ;
  assign n25083 = ~n1228 & n25082 ;
  assign n25084 = ~n1508 & n25083 ;
  assign n25085 = \b[14]  & n15517 ;
  assign n25086 = n15514 & n25085 ;
  assign n25087 = ~\a[51]  & \b[15]  ;
  assign n25088 = n14785 & n25087 ;
  assign n25089 = ~n25086 & ~n25088 ;
  assign n25090 = \b[16]  & n14791 ;
  assign n25091 = \a[51]  & \b[15]  ;
  assign n25092 = n14782 & n25091 ;
  assign n25093 = \a[53]  & ~n25092 ;
  assign n25094 = ~n25090 & n25093 ;
  assign n25095 = n25089 & n25094 ;
  assign n25096 = ~n25084 & n25095 ;
  assign n25097 = ~n25081 & n25096 ;
  assign n25098 = ~n25090 & ~n25092 ;
  assign n25099 = n25089 & n25098 ;
  assign n25100 = ~n25084 & n25099 ;
  assign n25101 = ~n25081 & n25100 ;
  assign n25102 = ~\a[53]  & ~n25101 ;
  assign n25103 = ~n25097 & ~n25102 ;
  assign n25104 = ~n25079 & n25103 ;
  assign n25105 = n25079 & ~n25103 ;
  assign n25106 = ~n25104 & ~n25105 ;
  assign n25107 = n24176 & ~n24283 ;
  assign n25108 = n23535 & ~n24300 ;
  assign n25109 = ~n24175 & n25108 ;
  assign n25110 = ~n24301 & ~n25109 ;
  assign n25111 = ~n25107 & n25110 ;
  assign n25112 = ~n25106 & n25111 ;
  assign n25113 = n25106 & ~n25111 ;
  assign n25114 = ~n25112 & ~n25113 ;
  assign n25115 = ~n2079 & n13125 ;
  assign n25116 = ~n2077 & n25115 ;
  assign n25117 = \b[17]  & n13794 ;
  assign n25118 = n13792 & n25117 ;
  assign n25119 = ~\a[48]  & \b[18]  ;
  assign n25120 = n13117 & n25119 ;
  assign n25121 = ~n25118 & ~n25120 ;
  assign n25122 = \b[19]  & n13123 ;
  assign n25123 = \a[48]  & \b[18]  ;
  assign n25124 = n13786 & n25123 ;
  assign n25125 = \a[50]  & ~n25124 ;
  assign n25126 = ~n25122 & n25125 ;
  assign n25127 = n25121 & n25126 ;
  assign n25128 = ~n25116 & n25127 ;
  assign n25129 = ~n25122 & ~n25124 ;
  assign n25130 = n25121 & n25129 ;
  assign n25131 = ~n25116 & n25130 ;
  assign n25132 = ~\a[50]  & ~n25131 ;
  assign n25133 = ~n25128 & ~n25132 ;
  assign n25134 = n25114 & ~n25133 ;
  assign n25135 = ~n25114 & n25133 ;
  assign n25136 = ~n25134 & ~n25135 ;
  assign n25137 = n2768 & n11572 ;
  assign n25138 = ~n2765 & n25137 ;
  assign n25139 = ~n2768 & n11572 ;
  assign n25140 = ~n2518 & n25139 ;
  assign n25141 = ~n2764 & n25140 ;
  assign n25142 = \b[20]  & n12159 ;
  assign n25143 = n12156 & n25142 ;
  assign n25144 = ~\a[45]  & \b[21]  ;
  assign n25145 = n11564 & n25144 ;
  assign n25146 = ~n25143 & ~n25145 ;
  assign n25147 = \b[22]  & n11570 ;
  assign n25148 = \a[45]  & \b[21]  ;
  assign n25149 = n11561 & n25148 ;
  assign n25150 = \a[47]  & ~n25149 ;
  assign n25151 = ~n25147 & n25150 ;
  assign n25152 = n25146 & n25151 ;
  assign n25153 = ~n25141 & n25152 ;
  assign n25154 = ~n25138 & n25153 ;
  assign n25155 = ~n25147 & ~n25149 ;
  assign n25156 = n25146 & n25155 ;
  assign n25157 = ~n25141 & n25156 ;
  assign n25158 = ~n25138 & n25157 ;
  assign n25159 = ~\a[47]  & ~n25158 ;
  assign n25160 = ~n25154 & ~n25159 ;
  assign n25161 = ~n25136 & n25160 ;
  assign n25162 = ~n24960 & n25161 ;
  assign n25163 = n25136 & n25160 ;
  assign n25164 = n24960 & n25163 ;
  assign n25165 = ~n25162 & ~n25164 ;
  assign n25166 = n25136 & ~n25160 ;
  assign n25167 = ~n24960 & n25166 ;
  assign n25168 = ~n25136 & ~n25160 ;
  assign n25169 = n24960 & n25168 ;
  assign n25170 = ~n25167 & ~n25169 ;
  assign n25171 = n25165 & n25170 ;
  assign n25172 = ~n24956 & n25171 ;
  assign n25173 = ~n3567 & n10082 ;
  assign n25174 = ~n3565 & n25173 ;
  assign n25175 = \b[23]  & n10681 ;
  assign n25176 = n10678 & n25175 ;
  assign n25177 = ~\a[42]  & \b[24]  ;
  assign n25178 = n10074 & n25177 ;
  assign n25179 = ~n25176 & ~n25178 ;
  assign n25180 = \b[25]  & n10080 ;
  assign n25181 = \a[42]  & \b[24]  ;
  assign n25182 = n10071 & n25181 ;
  assign n25183 = \a[44]  & ~n25182 ;
  assign n25184 = ~n25180 & n25183 ;
  assign n25185 = n25179 & n25184 ;
  assign n25186 = ~n25174 & n25185 ;
  assign n25187 = ~n25180 & ~n25182 ;
  assign n25188 = n25179 & n25187 ;
  assign n25189 = ~n25174 & n25188 ;
  assign n25190 = ~\a[44]  & ~n25189 ;
  assign n25191 = ~n25186 & ~n25190 ;
  assign n25192 = ~n24955 & ~n25171 ;
  assign n25193 = n24373 & n25192 ;
  assign n25194 = ~n25191 & ~n25193 ;
  assign n25195 = ~n25172 & n25194 ;
  assign n25196 = ~n25171 & n25191 ;
  assign n25197 = n24956 & n25196 ;
  assign n25198 = n25171 & n25191 ;
  assign n25199 = ~n24956 & n25198 ;
  assign n25200 = ~n25197 & ~n25199 ;
  assign n25201 = ~n25195 & n25200 ;
  assign n25202 = n4456 & n8759 ;
  assign n25203 = ~n18723 & n25202 ;
  assign n25204 = n8759 & n16805 ;
  assign n25205 = ~n4452 & n25204 ;
  assign n25206 = \b[26]  & n9301 ;
  assign n25207 = n9298 & n25206 ;
  assign n25208 = ~\a[39]  & \b[27]  ;
  assign n25209 = n8751 & n25208 ;
  assign n25210 = ~n25207 & ~n25209 ;
  assign n25211 = \b[28]  & n8757 ;
  assign n25212 = \a[39]  & \b[27]  ;
  assign n25213 = n8748 & n25212 ;
  assign n25214 = \a[41]  & ~n25213 ;
  assign n25215 = ~n25211 & n25214 ;
  assign n25216 = n25210 & n25215 ;
  assign n25217 = ~n25205 & n25216 ;
  assign n25218 = ~n25203 & n25217 ;
  assign n25219 = ~n25211 & ~n25213 ;
  assign n25220 = n25210 & n25219 ;
  assign n25221 = ~n25205 & n25220 ;
  assign n25222 = ~n25203 & n25221 ;
  assign n25223 = ~\a[41]  & ~n25222 ;
  assign n25224 = ~n25218 & ~n25223 ;
  assign n25225 = n25201 & n25224 ;
  assign n25226 = ~n24954 & n25225 ;
  assign n25227 = ~n25201 & n25224 ;
  assign n25228 = n24954 & n25227 ;
  assign n25229 = ~n25226 & ~n25228 ;
  assign n25230 = ~n25201 & ~n25224 ;
  assign n25231 = ~n24954 & n25230 ;
  assign n25232 = n25201 & ~n25224 ;
  assign n25233 = n24954 & n25232 ;
  assign n25234 = ~n25231 & ~n25233 ;
  assign n25235 = n25229 & n25234 ;
  assign n25236 = n24167 & n24409 ;
  assign n25237 = ~n23626 & ~n24433 ;
  assign n25238 = ~n24166 & n25237 ;
  assign n25239 = ~n24436 & ~n25238 ;
  assign n25240 = ~n25236 & n25239 ;
  assign n25241 = ~n25235 & n25240 ;
  assign n25242 = n25235 & ~n25240 ;
  assign n25243 = ~n25241 & ~n25242 ;
  assign n25244 = ~n5459 & n7534 ;
  assign n25245 = ~n5104 & n7534 ;
  assign n25246 = ~n5455 & n25245 ;
  assign n25247 = ~n25244 & ~n25246 ;
  assign n25248 = ~n5462 & ~n25247 ;
  assign n25249 = \b[29]  & n7973 ;
  assign n25250 = n7970 & n25249 ;
  assign n25251 = ~\a[36]  & \b[30]  ;
  assign n25252 = n7526 & n25251 ;
  assign n25253 = ~n25250 & ~n25252 ;
  assign n25254 = \b[31]  & n7532 ;
  assign n25255 = \a[36]  & \b[30]  ;
  assign n25256 = n17801 & n25255 ;
  assign n25257 = \a[38]  & ~n25256 ;
  assign n25258 = ~n25254 & n25257 ;
  assign n25259 = n25253 & n25258 ;
  assign n25260 = ~n25248 & n25259 ;
  assign n25261 = ~n25254 & ~n25256 ;
  assign n25262 = n25253 & n25261 ;
  assign n25263 = ~\a[38]  & ~n25262 ;
  assign n25264 = ~\a[38]  & ~n5462 ;
  assign n25265 = ~n25247 & n25264 ;
  assign n25266 = ~n25263 & ~n25265 ;
  assign n25267 = ~n25260 & n25266 ;
  assign n25268 = ~n25243 & n25267 ;
  assign n25269 = n25243 & ~n25267 ;
  assign n25270 = ~n25268 & ~n25269 ;
  assign n25271 = n24950 & ~n25270 ;
  assign n25272 = n24926 & n25271 ;
  assign n25273 = n24950 & n25270 ;
  assign n25274 = ~n24926 & n25273 ;
  assign n25275 = ~n25272 & ~n25274 ;
  assign n25276 = ~n24950 & ~n25270 ;
  assign n25277 = ~n24926 & n25276 ;
  assign n25278 = ~n24950 & n25270 ;
  assign n25279 = n24926 & n25278 ;
  assign n25280 = ~n25277 & ~n25279 ;
  assign n25281 = n25275 & n25280 ;
  assign n25282 = ~n24922 & n25281 ;
  assign n25283 = ~n24921 & ~n25281 ;
  assign n25284 = ~n24915 & n25283 ;
  assign n25285 = ~n25282 & ~n25284 ;
  assign n25286 = ~\a[29]  & ~n24890 ;
  assign n25287 = \a[29]  & n24888 ;
  assign n25288 = ~n24878 & n25287 ;
  assign n25289 = ~n24875 & n25288 ;
  assign n25290 = ~n25286 & ~n25289 ;
  assign n25291 = n24872 & n25290 ;
  assign n25292 = n24519 & n25291 ;
  assign n25293 = n25285 & ~n25292 ;
  assign n25294 = ~n24894 & n25293 ;
  assign n25295 = ~n24894 & ~n25292 ;
  assign n25296 = ~n25285 & ~n25295 ;
  assign n25297 = ~n25294 & ~n25296 ;
  assign n25298 = ~n24868 & n25297 ;
  assign n25299 = ~n24862 & n25298 ;
  assign n25300 = ~n24862 & ~n24868 ;
  assign n25301 = ~n25297 & ~n25300 ;
  assign n25302 = ~n25299 & ~n25301 ;
  assign n25303 = ~\a[23]  & ~n24840 ;
  assign n25304 = \a[23]  & n24838 ;
  assign n25305 = ~n24828 & n25304 ;
  assign n25306 = ~n24825 & n25305 ;
  assign n25307 = ~n25303 & ~n25306 ;
  assign n25308 = ~n24822 & n25307 ;
  assign n25309 = n24821 & n25308 ;
  assign n25310 = n25302 & ~n25309 ;
  assign n25311 = ~n24844 & n25310 ;
  assign n25312 = ~n24844 & ~n25309 ;
  assign n25313 = ~n25302 & ~n25312 ;
  assign n25314 = ~n25311 & ~n25313 ;
  assign n25315 = ~n24820 & n25314 ;
  assign n25316 = ~n24814 & ~n25314 ;
  assign n25317 = ~n24819 & n25316 ;
  assign n25318 = ~n25315 & ~n25317 ;
  assign n25319 = n24795 & n25318 ;
  assign n25320 = ~n24795 & ~n25318 ;
  assign n25321 = ~n25319 & ~n25320 ;
  assign n25322 = ~n24761 & ~n25321 ;
  assign n25323 = ~n24755 & n25322 ;
  assign n25324 = ~n24755 & ~n24761 ;
  assign n25325 = n25321 & ~n25324 ;
  assign n25326 = ~n25323 & ~n25325 ;
  assign n25327 = n23831 & ~n24602 ;
  assign n25328 = n23832 & ~n24602 ;
  assign n25329 = n23296 & n25328 ;
  assign n25330 = ~n25327 & ~n25329 ;
  assign n25331 = ~n23831 & n24602 ;
  assign n25332 = ~n24029 & n25331 ;
  assign n25333 = n25330 & n25332 ;
  assign n25334 = ~n24578 & n24734 ;
  assign n25335 = ~n24578 & n24621 ;
  assign n25336 = ~n24033 & n25335 ;
  assign n25337 = ~n25334 & ~n25336 ;
  assign n25338 = ~n24737 & n25337 ;
  assign n25339 = n25330 & ~n25338 ;
  assign n25340 = ~n25333 & ~n25339 ;
  assign n25341 = ~n551 & ~n17685 ;
  assign n25342 = ~n18940 & n25341 ;
  assign n25343 = ~n18936 & n25342 ;
  assign n25344 = ~n643 & n25343 ;
  assign n25345 = n646 & n18940 ;
  assign n25346 = ~n18937 & n25345 ;
  assign n25347 = ~n25344 & ~n25346 ;
  assign n25348 = \b[58]  & n644 ;
  assign n25349 = \a[9]  & \b[57]  ;
  assign n25350 = n635 & n25349 ;
  assign n25351 = ~n25348 & ~n25350 ;
  assign n25352 = \b[56]  & n796 ;
  assign n25353 = n793 & n25352 ;
  assign n25354 = ~\a[9]  & \b[57]  ;
  assign n25355 = n638 & n25354 ;
  assign n25356 = ~n25353 & ~n25355 ;
  assign n25357 = n25351 & n25356 ;
  assign n25358 = n25347 & n25357 ;
  assign n25359 = \a[11]  & ~n25358 ;
  assign n25360 = ~\a[11]  & n25358 ;
  assign n25361 = ~n25359 & ~n25360 ;
  assign n25362 = n25340 & n25361 ;
  assign n25363 = ~\a[11]  & ~n25358 ;
  assign n25364 = \a[11]  & n25357 ;
  assign n25365 = n25347 & n25364 ;
  assign n25366 = ~n25363 & ~n25365 ;
  assign n25367 = ~n25340 & n25366 ;
  assign n25368 = ~n25362 & ~n25367 ;
  assign n25369 = n25326 & n25368 ;
  assign n25370 = ~n25326 & ~n25368 ;
  assign n25371 = ~n25369 & ~n25370 ;
  assign n25372 = n24670 & ~n24674 ;
  assign n25373 = n24651 & ~n24678 ;
  assign n25374 = ~n25372 & ~n25373 ;
  assign n25375 = n430 & ~n20971 ;
  assign n25376 = ~n20969 & n25375 ;
  assign n25377 = \b[61]  & n428 ;
  assign n25378 = \a[6]  & \b[60]  ;
  assign n25379 = n419 & n25378 ;
  assign n25380 = ~n25377 & ~n25379 ;
  assign n25381 = \b[59]  & n486 ;
  assign n25382 = n483 & n25381 ;
  assign n25383 = ~\a[6]  & \b[60]  ;
  assign n25384 = n422 & n25383 ;
  assign n25385 = ~n25382 & ~n25384 ;
  assign n25386 = n25380 & n25385 ;
  assign n25387 = ~n25376 & n25386 ;
  assign n25388 = \a[8]  & ~n25387 ;
  assign n25389 = ~\a[8]  & n25387 ;
  assign n25390 = ~n25388 & ~n25389 ;
  assign n25391 = n25374 & n25390 ;
  assign n25392 = ~\a[8]  & ~n25387 ;
  assign n25393 = \a[8]  & n25386 ;
  assign n25394 = ~n25376 & n25393 ;
  assign n25395 = ~n25392 & ~n25394 ;
  assign n25396 = ~n25374 & n25395 ;
  assign n25397 = ~n25391 & ~n25396 ;
  assign n25398 = n25371 & n25397 ;
  assign n25399 = ~n25371 & ~n25397 ;
  assign n25400 = ~n25398 & ~n25399 ;
  assign n25401 = ~n24024 & n24684 ;
  assign n25402 = \b[62]  & n303 ;
  assign n25403 = n300 & n25402 ;
  assign n25404 = ~\a[3]  & \b[63]  ;
  assign n25405 = n244 & n25404 ;
  assign n25406 = \a[3]  & \b[63]  ;
  assign n25407 = n241 & n25406 ;
  assign n25408 = ~n25405 & ~n25407 ;
  assign n25409 = ~n25403 & n25408 ;
  assign n25410 = ~\a[5]  & ~n25409 ;
  assign n25411 = n252 & ~n22458 ;
  assign n25412 = ~\a[5]  & n25411 ;
  assign n25413 = ~n23173 & n25412 ;
  assign n25414 = ~n25410 & ~n25413 ;
  assign n25415 = ~n23173 & n25411 ;
  assign n25416 = \a[5]  & n25409 ;
  assign n25417 = ~n25415 & n25416 ;
  assign n25418 = n25414 & ~n25417 ;
  assign n25419 = ~n24026 & ~n25418 ;
  assign n25420 = ~n25401 & n25419 ;
  assign n25421 = n24026 & n25418 ;
  assign n25422 = n24684 & n25418 ;
  assign n25423 = ~n24024 & n25422 ;
  assign n25424 = ~n25421 & ~n25423 ;
  assign n25425 = ~n25420 & n25424 ;
  assign n25426 = n25400 & n25425 ;
  assign n25427 = ~n25400 & ~n25425 ;
  assign n25428 = ~n25426 & ~n25427 ;
  assign n25429 = ~n24732 & n25428 ;
  assign n25430 = n24732 & ~n25428 ;
  assign n25431 = ~n25429 & ~n25430 ;
  assign n25432 = ~n24718 & n25431 ;
  assign n25433 = ~n24730 & n25432 ;
  assign n25434 = ~n24718 & ~n24730 ;
  assign n25435 = ~n25431 & ~n25434 ;
  assign n25436 = ~n25433 & ~n25435 ;
  assign n25437 = ~n25429 & ~n25433 ;
  assign n25438 = ~n25400 & ~n25420 ;
  assign n25439 = n25424 & ~n25438 ;
  assign n25440 = n25326 & ~n25367 ;
  assign n25441 = ~n25362 & ~n25440 ;
  assign n25442 = n430 & ~n21699 ;
  assign n25443 = ~n21697 & n25442 ;
  assign n25444 = \b[62]  & n428 ;
  assign n25445 = \a[6]  & \b[61]  ;
  assign n25446 = n419 & n25445 ;
  assign n25447 = ~n25444 & ~n25446 ;
  assign n25448 = \b[60]  & n486 ;
  assign n25449 = n483 & n25448 ;
  assign n25450 = ~\a[6]  & \b[61]  ;
  assign n25451 = n422 & n25450 ;
  assign n25452 = ~n25449 & ~n25451 ;
  assign n25453 = n25447 & n25452 ;
  assign n25454 = ~n25443 & n25453 ;
  assign n25455 = \a[8]  & ~n25454 ;
  assign n25456 = ~\a[8]  & n25454 ;
  assign n25457 = ~n25455 & ~n25456 ;
  assign n25458 = ~n25441 & n25457 ;
  assign n25459 = ~n24755 & n24761 ;
  assign n25460 = ~n24755 & n25321 ;
  assign n25461 = n646 & ~n19550 ;
  assign n25462 = ~n19548 & n25461 ;
  assign n25463 = \b[59]  & n644 ;
  assign n25464 = \a[9]  & \b[58]  ;
  assign n25465 = n635 & n25464 ;
  assign n25466 = ~n25463 & ~n25465 ;
  assign n25467 = \b[57]  & n796 ;
  assign n25468 = n793 & n25467 ;
  assign n25469 = ~\a[9]  & \b[58]  ;
  assign n25470 = n638 & n25469 ;
  assign n25471 = ~n25468 & ~n25470 ;
  assign n25472 = n25466 & n25471 ;
  assign n25473 = ~n25462 & n25472 ;
  assign n25474 = ~\a[11]  & ~n25473 ;
  assign n25475 = \a[11]  & n25472 ;
  assign n25476 = ~n25462 & n25475 ;
  assign n25477 = ~n25474 & ~n25476 ;
  assign n25478 = ~n25460 & ~n25477 ;
  assign n25479 = ~n25459 & n25478 ;
  assign n25480 = ~n24755 & ~n25322 ;
  assign n25481 = n25477 & n25480 ;
  assign n25482 = ~n24788 & n25318 ;
  assign n25483 = ~n24788 & n24794 ;
  assign n25484 = ~n25482 & ~n25483 ;
  assign n25485 = n999 & n17647 ;
  assign n25486 = ~n17644 & n25485 ;
  assign n25487 = n999 & ~n17647 ;
  assign n25488 = ~n16441 & n25487 ;
  assign n25489 = ~n17643 & n25488 ;
  assign n25490 = \b[54]  & n1182 ;
  assign n25491 = n1179 & n25490 ;
  assign n25492 = \b[56]  & n997 ;
  assign n25493 = \a[11]  & \b[55]  ;
  assign n25494 = n1180 & n25493 ;
  assign n25495 = ~\a[12]  & \b[55]  ;
  assign n25496 = n7674 & n25495 ;
  assign n25497 = ~n25494 & ~n25496 ;
  assign n25498 = ~n25492 & n25497 ;
  assign n25499 = ~n25491 & n25498 ;
  assign n25500 = ~n25489 & n25499 ;
  assign n25501 = ~n25486 & n25500 ;
  assign n25502 = \a[14]  & ~n25501 ;
  assign n25503 = ~\a[14]  & n25501 ;
  assign n25504 = ~n25502 & ~n25503 ;
  assign n25505 = n25484 & n25504 ;
  assign n25506 = ~\a[14]  & ~n25501 ;
  assign n25507 = \a[14]  & n25499 ;
  assign n25508 = ~n25489 & n25507 ;
  assign n25509 = ~n25486 & n25508 ;
  assign n25510 = ~n25506 & ~n25509 ;
  assign n25511 = ~n25484 & n25510 ;
  assign n25512 = ~n25505 & ~n25511 ;
  assign n25513 = n1467 & ~n15246 ;
  assign n25514 = ~n15244 & n25513 ;
  assign n25515 = \b[53]  & n1465 ;
  assign n25516 = \a[15]  & \b[52]  ;
  assign n25517 = n1456 & n25516 ;
  assign n25518 = ~n25515 & ~n25517 ;
  assign n25519 = \b[51]  & n1652 ;
  assign n25520 = n1649 & n25519 ;
  assign n25521 = ~\a[15]  & \b[52]  ;
  assign n25522 = n1459 & n25521 ;
  assign n25523 = ~n25520 & ~n25522 ;
  assign n25524 = n25518 & n25523 ;
  assign n25525 = ~n25514 & n25524 ;
  assign n25526 = ~\a[17]  & ~n25525 ;
  assign n25527 = \a[17]  & n25524 ;
  assign n25528 = ~n25514 & n25527 ;
  assign n25529 = n24814 & ~n25528 ;
  assign n25530 = ~n25314 & ~n25528 ;
  assign n25531 = ~n24819 & n25530 ;
  assign n25532 = ~n25529 & ~n25531 ;
  assign n25533 = ~n25526 & ~n25532 ;
  assign n25534 = ~n24819 & ~n25314 ;
  assign n25535 = \a[17]  & ~n25525 ;
  assign n25536 = ~\a[17]  & n25525 ;
  assign n25537 = ~n25535 & ~n25536 ;
  assign n25538 = ~n24814 & n25537 ;
  assign n25539 = ~n25534 & n25538 ;
  assign n25540 = ~n24862 & n24868 ;
  assign n25541 = ~n24862 & ~n25297 ;
  assign n25542 = n2622 & ~n12438 ;
  assign n25543 = ~n12436 & n25542 ;
  assign n25544 = \b[47]  & n2620 ;
  assign n25545 = \a[21]  & \b[46]  ;
  assign n25546 = n20849 & n25545 ;
  assign n25547 = ~n25544 & ~n25546 ;
  assign n25548 = \b[45]  & n2912 ;
  assign n25549 = n2909 & n25548 ;
  assign n25550 = ~\a[21]  & \b[46]  ;
  assign n25551 = n2614 & n25550 ;
  assign n25552 = ~n25549 & ~n25551 ;
  assign n25553 = n25547 & n25552 ;
  assign n25554 = ~n25543 & n25553 ;
  assign n25555 = ~\a[23]  & ~n25554 ;
  assign n25556 = \a[23]  & n25553 ;
  assign n25557 = ~n25543 & n25556 ;
  assign n25558 = ~n25555 & ~n25557 ;
  assign n25559 = ~n25541 & ~n25558 ;
  assign n25560 = ~n25540 & n25559 ;
  assign n25561 = ~n24862 & ~n25298 ;
  assign n25562 = n25558 & n25561 ;
  assign n25563 = ~n24894 & ~n25293 ;
  assign n25564 = n3402 & ~n10892 ;
  assign n25565 = ~n10890 & n25564 ;
  assign n25566 = \b[44]  & n3400 ;
  assign n25567 = \a[24]  & \b[43]  ;
  assign n25568 = n3391 & n25567 ;
  assign n25569 = ~n25566 & ~n25568 ;
  assign n25570 = \b[42]  & n3733 ;
  assign n25571 = n3730 & n25570 ;
  assign n25572 = ~\a[24]  & \b[43]  ;
  assign n25573 = n3394 & n25572 ;
  assign n25574 = ~n25571 & ~n25573 ;
  assign n25575 = n25569 & n25574 ;
  assign n25576 = ~n25565 & n25575 ;
  assign n25577 = \a[26]  & ~n25576 ;
  assign n25578 = ~\a[26]  & n25576 ;
  assign n25579 = ~n25577 & ~n25578 ;
  assign n25580 = ~n25563 & n25579 ;
  assign n25581 = ~\a[26]  & ~n25576 ;
  assign n25582 = \a[26]  & n25575 ;
  assign n25583 = ~n25565 & n25582 ;
  assign n25584 = ~n25581 & ~n25583 ;
  assign n25585 = n25563 & n25584 ;
  assign n25586 = ~n25580 & ~n25585 ;
  assign n25587 = ~n24915 & ~n25283 ;
  assign n25588 = n4249 & ~n9482 ;
  assign n25589 = ~n9480 & n25588 ;
  assign n25590 = \b[41]  & n4247 ;
  assign n25591 = \a[27]  & \b[40]  ;
  assign n25592 = n4238 & n25591 ;
  assign n25593 = ~n25590 & ~n25592 ;
  assign n25594 = \b[39]  & n4647 ;
  assign n25595 = n4644 & n25594 ;
  assign n25596 = ~\a[27]  & \b[40]  ;
  assign n25597 = n4241 & n25596 ;
  assign n25598 = ~n25595 & ~n25597 ;
  assign n25599 = n25593 & n25598 ;
  assign n25600 = ~n25589 & n25599 ;
  assign n25601 = ~\a[29]  & ~n25600 ;
  assign n25602 = \a[29]  & n25599 ;
  assign n25603 = ~n25589 & n25602 ;
  assign n25604 = ~n25601 & ~n25603 ;
  assign n25605 = n25587 & n25604 ;
  assign n25606 = ~n24915 & n25281 ;
  assign n25607 = ~n24895 & n24913 ;
  assign n25608 = ~n24897 & n25607 ;
  assign n25609 = ~n24895 & n24912 ;
  assign n25610 = ~n24897 & n25609 ;
  assign n25611 = ~n25608 & ~n25610 ;
  assign n25612 = ~n25604 & n25611 ;
  assign n25613 = ~n25606 & n25612 ;
  assign n25614 = ~n25605 & ~n25613 ;
  assign n25615 = n24926 & n25270 ;
  assign n25616 = ~n24476 & ~n24950 ;
  assign n25617 = n24925 & n25616 ;
  assign n25618 = ~n25278 & ~n25617 ;
  assign n25619 = ~n25615 & n25618 ;
  assign n25620 = n5211 & n8175 ;
  assign n25621 = ~n8172 & n25620 ;
  assign n25622 = ~n7756 & ~n8175 ;
  assign n25623 = n5211 & n25622 ;
  assign n25624 = ~n8171 & n25623 ;
  assign n25625 = \b[38]  & n5209 ;
  assign n25626 = \a[30]  & \b[37]  ;
  assign n25627 = n5200 & n25626 ;
  assign n25628 = ~n25625 & ~n25627 ;
  assign n25629 = \b[36]  & n5595 ;
  assign n25630 = n5592 & n25629 ;
  assign n25631 = ~\a[30]  & \b[37]  ;
  assign n25632 = n5203 & n25631 ;
  assign n25633 = ~n25630 & ~n25632 ;
  assign n25634 = n25628 & n25633 ;
  assign n25635 = ~n25624 & n25634 ;
  assign n25636 = ~n25621 & n25635 ;
  assign n25637 = \a[32]  & ~n25636 ;
  assign n25638 = ~\a[32]  & n25636 ;
  assign n25639 = ~n25637 & ~n25638 ;
  assign n25640 = ~n25619 & n25639 ;
  assign n25641 = ~\a[32]  & ~n25636 ;
  assign n25642 = \a[32]  & n25634 ;
  assign n25643 = ~n25624 & n25642 ;
  assign n25644 = ~n25621 & n25643 ;
  assign n25645 = ~n25641 & ~n25644 ;
  assign n25646 = n25619 & n25645 ;
  assign n25647 = ~n25640 & ~n25646 ;
  assign n25648 = ~n24954 & n25201 ;
  assign n25649 = n24954 & ~n25201 ;
  assign n25650 = ~n25224 & ~n25649 ;
  assign n25651 = ~n25648 & ~n25650 ;
  assign n25652 = ~n24955 & n25191 ;
  assign n25653 = n24373 & n25652 ;
  assign n25654 = ~n25196 & ~n25653 ;
  assign n25655 = ~n25193 & n25654 ;
  assign n25656 = ~n24960 & ~n25136 ;
  assign n25657 = n24960 & n25136 ;
  assign n25658 = n25160 & ~n25657 ;
  assign n25659 = ~n25656 & ~n25658 ;
  assign n25660 = ~n1694 & n14793 ;
  assign n25661 = ~n1692 & n25660 ;
  assign n25662 = \b[15]  & n15517 ;
  assign n25663 = n15514 & n25662 ;
  assign n25664 = ~\a[51]  & \b[16]  ;
  assign n25665 = n14785 & n25664 ;
  assign n25666 = ~n25663 & ~n25665 ;
  assign n25667 = \b[17]  & n14791 ;
  assign n25668 = \a[51]  & \b[16]  ;
  assign n25669 = n14782 & n25668 ;
  assign n25670 = \a[53]  & ~n25669 ;
  assign n25671 = ~n25667 & n25670 ;
  assign n25672 = n25666 & n25671 ;
  assign n25673 = ~n25661 & n25672 ;
  assign n25674 = ~n25667 & ~n25669 ;
  assign n25675 = n25666 & n25674 ;
  assign n25676 = ~n25661 & n25675 ;
  assign n25677 = ~\a[53]  & ~n25676 ;
  assign n25678 = ~n25673 & ~n25677 ;
  assign n25679 = ~n25043 & n25068 ;
  assign n25680 = ~n25042 & ~n25679 ;
  assign n25681 = n24997 & n25002 ;
  assign n25682 = ~n505 & ~n19861 ;
  assign n25683 = ~n20518 & n25682 ;
  assign n25684 = n502 & n25683 ;
  assign n25685 = n505 & ~n19861 ;
  assign n25686 = ~n20518 & n25685 ;
  assign n25687 = ~n502 & n25686 ;
  assign n25688 = ~n25684 & ~n25687 ;
  assign n25689 = \b[6]  & n21315 ;
  assign n25690 = n21312 & n25689 ;
  assign n25691 = \b[8]  & n20519 ;
  assign n25692 = \a[59]  & \b[7]  ;
  assign n25693 = n21313 & n25692 ;
  assign n25694 = ~\a[60]  & \b[7]  ;
  assign n25695 = n20513 & n25694 ;
  assign n25696 = ~n25693 & ~n25695 ;
  assign n25697 = ~n25691 & n25696 ;
  assign n25698 = ~n25690 & n25697 ;
  assign n25699 = n25688 & n25698 ;
  assign n25700 = \b[5]  & n21958 ;
  assign n25701 = \b[4]  & n21957 ;
  assign n25702 = ~\a[2]  & ~n25701 ;
  assign n25703 = ~n25700 & n25702 ;
  assign n25704 = \a[2]  & \b[5]  ;
  assign n25705 = n21958 & n25704 ;
  assign n25706 = n21957 & n24977 ;
  assign n25707 = ~\a[62]  & ~n25706 ;
  assign n25708 = ~n25705 & n25707 ;
  assign n25709 = ~n25703 & n25708 ;
  assign n25710 = ~n25699 & n25709 ;
  assign n25711 = \a[62]  & ~n25706 ;
  assign n25712 = ~n25705 & n25711 ;
  assign n25713 = ~n25703 & n25712 ;
  assign n25714 = n25698 & n25713 ;
  assign n25715 = n25688 & n25714 ;
  assign n25716 = ~n25710 & ~n25715 ;
  assign n25717 = ~\a[62]  & ~n25699 ;
  assign n25718 = ~n25705 & ~n25706 ;
  assign n25719 = ~n25703 & n25718 ;
  assign n25720 = \a[62]  & n25698 ;
  assign n25721 = n25688 & n25720 ;
  assign n25722 = ~n25719 & ~n25721 ;
  assign n25723 = ~n25717 & n25722 ;
  assign n25724 = n25716 & ~n25723 ;
  assign n25725 = n25681 & ~n25724 ;
  assign n25726 = ~n25681 & n25724 ;
  assign n25727 = ~n25725 & ~n25726 ;
  assign n25728 = ~n728 & n18516 ;
  assign n25729 = ~n726 & n25728 ;
  assign n25730 = \b[9]  & n19183 ;
  assign n25731 = n19180 & n25730 ;
  assign n25732 = ~\a[57]  & \b[10]  ;
  assign n25733 = n18508 & n25732 ;
  assign n25734 = ~n25731 & ~n25733 ;
  assign n25735 = \b[11]  & n18514 ;
  assign n25736 = \a[57]  & \b[10]  ;
  assign n25737 = n18505 & n25736 ;
  assign n25738 = \a[59]  & ~n25737 ;
  assign n25739 = ~n25735 & n25738 ;
  assign n25740 = n25734 & n25739 ;
  assign n25741 = ~n25729 & n25740 ;
  assign n25742 = ~n25735 & ~n25737 ;
  assign n25743 = n25734 & n25742 ;
  assign n25744 = ~n25729 & n25743 ;
  assign n25745 = ~\a[59]  & ~n25744 ;
  assign n25746 = ~n25741 & ~n25745 ;
  assign n25747 = n25727 & ~n25746 ;
  assign n25748 = ~n25727 & n25746 ;
  assign n25749 = ~n25011 & n25036 ;
  assign n25750 = ~n25009 & ~n25749 ;
  assign n25751 = ~n25748 & n25750 ;
  assign n25752 = ~n25747 & n25751 ;
  assign n25753 = ~n25746 & ~n25750 ;
  assign n25754 = n25727 & n25753 ;
  assign n25755 = ~n25727 & ~n25750 ;
  assign n25756 = n25746 & n25755 ;
  assign n25757 = ~n25754 & ~n25756 ;
  assign n25758 = ~n25752 & n25757 ;
  assign n25759 = n1087 & n16655 ;
  assign n25760 = ~n1084 & n25759 ;
  assign n25761 = n16655 & n21340 ;
  assign n25762 = ~n1083 & n25761 ;
  assign n25763 = \b[12]  & n17308 ;
  assign n25764 = n17305 & n25763 ;
  assign n25765 = ~\a[54]  & \b[13]  ;
  assign n25766 = n16647 & n25765 ;
  assign n25767 = ~n25764 & ~n25766 ;
  assign n25768 = \b[14]  & n16653 ;
  assign n25769 = \a[54]  & \b[13]  ;
  assign n25770 = n16644 & n25769 ;
  assign n25771 = \a[56]  & ~n25770 ;
  assign n25772 = ~n25768 & n25771 ;
  assign n25773 = n25767 & n25772 ;
  assign n25774 = ~n25762 & n25773 ;
  assign n25775 = ~n25760 & n25774 ;
  assign n25776 = ~n25768 & ~n25770 ;
  assign n25777 = n25767 & n25776 ;
  assign n25778 = ~n25762 & n25777 ;
  assign n25779 = ~n25760 & n25778 ;
  assign n25780 = ~\a[56]  & ~n25779 ;
  assign n25781 = ~n25775 & ~n25780 ;
  assign n25782 = ~n25758 & ~n25781 ;
  assign n25783 = n25758 & n25781 ;
  assign n25784 = ~n25782 & ~n25783 ;
  assign n25785 = n25680 & ~n25784 ;
  assign n25786 = ~n25680 & n25784 ;
  assign n25787 = ~n25785 & ~n25786 ;
  assign n25788 = n25678 & n25787 ;
  assign n25789 = ~n25678 & ~n25787 ;
  assign n25790 = ~n25788 & ~n25789 ;
  assign n25791 = ~n25078 & ~n25103 ;
  assign n25792 = ~n25077 & ~n25791 ;
  assign n25793 = n2293 & n13125 ;
  assign n25794 = ~n19247 & n25793 ;
  assign n25795 = ~n2293 & n13125 ;
  assign n25796 = ~n2074 & n25795 ;
  assign n25797 = ~n2289 & n25796 ;
  assign n25798 = \b[18]  & n13794 ;
  assign n25799 = n13792 & n25798 ;
  assign n25800 = ~\a[48]  & \b[19]  ;
  assign n25801 = n13117 & n25800 ;
  assign n25802 = ~n25799 & ~n25801 ;
  assign n25803 = \b[20]  & n13123 ;
  assign n25804 = \a[48]  & \b[19]  ;
  assign n25805 = n13786 & n25804 ;
  assign n25806 = \a[50]  & ~n25805 ;
  assign n25807 = ~n25803 & n25806 ;
  assign n25808 = n25802 & n25807 ;
  assign n25809 = ~n25797 & n25808 ;
  assign n25810 = ~n25794 & n25809 ;
  assign n25811 = ~n25803 & ~n25805 ;
  assign n25812 = n25802 & n25811 ;
  assign n25813 = ~n25797 & n25812 ;
  assign n25814 = ~n25794 & n25813 ;
  assign n25815 = ~\a[50]  & ~n25814 ;
  assign n25816 = ~n25810 & ~n25815 ;
  assign n25817 = ~n25792 & n25816 ;
  assign n25818 = ~n25790 & n25817 ;
  assign n25819 = n25792 & n25816 ;
  assign n25820 = n25790 & n25819 ;
  assign n25821 = ~n25818 & ~n25820 ;
  assign n25822 = n25792 & ~n25816 ;
  assign n25823 = ~n25790 & n25822 ;
  assign n25824 = ~n25792 & ~n25816 ;
  assign n25825 = n25790 & n25824 ;
  assign n25826 = ~n25823 & ~n25825 ;
  assign n25827 = n25821 & n25826 ;
  assign n25828 = ~n25113 & n25133 ;
  assign n25829 = ~n25112 & ~n25828 ;
  assign n25830 = ~n3022 & n11572 ;
  assign n25831 = ~n3020 & n25830 ;
  assign n25832 = \b[21]  & n12159 ;
  assign n25833 = n12156 & n25832 ;
  assign n25834 = ~\a[45]  & \b[22]  ;
  assign n25835 = n11564 & n25834 ;
  assign n25836 = ~n25833 & ~n25835 ;
  assign n25837 = \b[23]  & n11570 ;
  assign n25838 = \a[45]  & \b[22]  ;
  assign n25839 = n11561 & n25838 ;
  assign n25840 = \a[47]  & ~n25839 ;
  assign n25841 = ~n25837 & n25840 ;
  assign n25842 = n25836 & n25841 ;
  assign n25843 = ~n25831 & n25842 ;
  assign n25844 = ~n25837 & ~n25839 ;
  assign n25845 = n25836 & n25844 ;
  assign n25846 = ~n25831 & n25845 ;
  assign n25847 = ~\a[47]  & ~n25846 ;
  assign n25848 = ~n25843 & ~n25847 ;
  assign n25849 = ~n25829 & ~n25848 ;
  assign n25850 = n25827 & n25849 ;
  assign n25851 = n25829 & ~n25848 ;
  assign n25852 = ~n25827 & n25851 ;
  assign n25853 = ~n25850 & ~n25852 ;
  assign n25854 = ~n25829 & n25848 ;
  assign n25855 = ~n25827 & n25854 ;
  assign n25856 = n25829 & n25848 ;
  assign n25857 = n25827 & n25856 ;
  assign n25858 = ~n25855 & ~n25857 ;
  assign n25859 = n25853 & n25858 ;
  assign n25860 = n3604 & n10082 ;
  assign n25861 = ~n19292 & n25860 ;
  assign n25862 = ~n3604 & n10082 ;
  assign n25863 = ~n3562 & n25862 ;
  assign n25864 = ~n3600 & n25863 ;
  assign n25865 = \b[24]  & n10681 ;
  assign n25866 = n10678 & n25865 ;
  assign n25867 = ~\a[42]  & \b[25]  ;
  assign n25868 = n10074 & n25867 ;
  assign n25869 = ~n25866 & ~n25868 ;
  assign n25870 = \b[26]  & n10080 ;
  assign n25871 = \a[42]  & \b[25]  ;
  assign n25872 = n10071 & n25871 ;
  assign n25873 = \a[44]  & ~n25872 ;
  assign n25874 = ~n25870 & n25873 ;
  assign n25875 = n25869 & n25874 ;
  assign n25876 = ~n25864 & n25875 ;
  assign n25877 = ~n25861 & n25876 ;
  assign n25878 = ~n25870 & ~n25872 ;
  assign n25879 = n25869 & n25878 ;
  assign n25880 = ~n25864 & n25879 ;
  assign n25881 = ~n25861 & n25880 ;
  assign n25882 = ~\a[44]  & ~n25881 ;
  assign n25883 = ~n25877 & ~n25882 ;
  assign n25884 = ~n25859 & n25883 ;
  assign n25885 = ~n25659 & n25884 ;
  assign n25886 = n25859 & n25883 ;
  assign n25887 = n25659 & n25886 ;
  assign n25888 = ~n25885 & ~n25887 ;
  assign n25889 = n25859 & ~n25883 ;
  assign n25890 = ~n25659 & n25889 ;
  assign n25891 = ~n25859 & ~n25883 ;
  assign n25892 = n25659 & n25891 ;
  assign n25893 = ~n25890 & ~n25892 ;
  assign n25894 = n25888 & n25893 ;
  assign n25895 = ~n4499 & n8759 ;
  assign n25896 = ~n4455 & n8759 ;
  assign n25897 = ~n4495 & n25896 ;
  assign n25898 = ~n25895 & ~n25897 ;
  assign n25899 = ~n4502 & ~n25898 ;
  assign n25900 = \b[27]  & n9301 ;
  assign n25901 = n9298 & n25900 ;
  assign n25902 = ~\a[39]  & \b[28]  ;
  assign n25903 = n8751 & n25902 ;
  assign n25904 = ~n25901 & ~n25903 ;
  assign n25905 = \b[29]  & n8757 ;
  assign n25906 = \a[39]  & \b[28]  ;
  assign n25907 = n8748 & n25906 ;
  assign n25908 = \a[41]  & ~n25907 ;
  assign n25909 = ~n25905 & n25908 ;
  assign n25910 = n25904 & n25909 ;
  assign n25911 = ~n25899 & n25910 ;
  assign n25912 = ~n25905 & ~n25907 ;
  assign n25913 = n25904 & n25912 ;
  assign n25914 = ~\a[41]  & ~n25913 ;
  assign n25915 = ~\a[41]  & ~n4502 ;
  assign n25916 = ~n25898 & n25915 ;
  assign n25917 = ~n25914 & ~n25916 ;
  assign n25918 = ~n25911 & n25917 ;
  assign n25919 = ~n25894 & ~n25918 ;
  assign n25920 = n25655 & n25919 ;
  assign n25921 = n25894 & ~n25918 ;
  assign n25922 = ~n25655 & n25921 ;
  assign n25923 = ~n25920 & ~n25922 ;
  assign n25924 = ~n25894 & n25918 ;
  assign n25925 = ~n25655 & n25924 ;
  assign n25926 = n25894 & n25918 ;
  assign n25927 = n25655 & n25926 ;
  assign n25928 = ~n25925 & ~n25927 ;
  assign n25929 = n25923 & n25928 ;
  assign n25930 = n5810 & n7534 ;
  assign n25931 = ~n5807 & n25930 ;
  assign n25932 = n7534 & n19029 ;
  assign n25933 = ~n5806 & n25932 ;
  assign n25934 = \b[30]  & n7973 ;
  assign n25935 = n7970 & n25934 ;
  assign n25936 = ~\a[36]  & \b[31]  ;
  assign n25937 = n7526 & n25936 ;
  assign n25938 = ~n25935 & ~n25937 ;
  assign n25939 = \b[32]  & n7532 ;
  assign n25940 = \a[36]  & \b[31]  ;
  assign n25941 = n17801 & n25940 ;
  assign n25942 = \a[38]  & ~n25941 ;
  assign n25943 = ~n25939 & n25942 ;
  assign n25944 = n25938 & n25943 ;
  assign n25945 = ~n25933 & n25944 ;
  assign n25946 = ~n25931 & n25945 ;
  assign n25947 = ~n25939 & ~n25941 ;
  assign n25948 = n25938 & n25947 ;
  assign n25949 = ~n25933 & n25948 ;
  assign n25950 = ~n25931 & n25949 ;
  assign n25951 = ~\a[38]  & ~n25950 ;
  assign n25952 = ~n25946 & ~n25951 ;
  assign n25953 = ~n25929 & n25952 ;
  assign n25954 = n25651 & n25953 ;
  assign n25955 = n25929 & n25952 ;
  assign n25956 = ~n25651 & n25955 ;
  assign n25957 = ~n25954 & ~n25956 ;
  assign n25958 = ~n25651 & n25929 ;
  assign n25959 = ~n25648 & ~n25929 ;
  assign n25960 = ~n25650 & n25959 ;
  assign n25961 = ~n25952 & ~n25960 ;
  assign n25962 = ~n25958 & n25961 ;
  assign n25963 = n25957 & ~n25962 ;
  assign n25964 = ~n25242 & n25267 ;
  assign n25965 = ~n25241 & ~n25964 ;
  assign n25966 = n25963 & n25965 ;
  assign n25967 = ~n25963 & ~n25965 ;
  assign n25968 = ~n25966 & ~n25967 ;
  assign n25969 = n6309 & ~n6610 ;
  assign n25970 = ~n6608 & n25969 ;
  assign n25971 = \b[33]  & n6778 ;
  assign n25972 = n6775 & n25971 ;
  assign n25973 = ~\a[33]  & \b[34]  ;
  assign n25974 = n6301 & n25973 ;
  assign n25975 = ~n25972 & ~n25974 ;
  assign n25976 = \b[35]  & n6307 ;
  assign n25977 = \a[33]  & \b[34]  ;
  assign n25978 = n6298 & n25977 ;
  assign n25979 = \a[35]  & ~n25978 ;
  assign n25980 = ~n25976 & n25979 ;
  assign n25981 = n25975 & n25980 ;
  assign n25982 = ~n25970 & n25981 ;
  assign n25983 = ~n25976 & ~n25978 ;
  assign n25984 = n25975 & n25983 ;
  assign n25985 = ~n25970 & n25984 ;
  assign n25986 = ~\a[35]  & ~n25985 ;
  assign n25987 = ~n25982 & ~n25986 ;
  assign n25988 = ~n25968 & n25987 ;
  assign n25989 = n25968 & ~n25987 ;
  assign n25990 = ~n25988 & ~n25989 ;
  assign n25991 = n25647 & n25990 ;
  assign n25992 = ~n25647 & ~n25990 ;
  assign n25993 = ~n25991 & ~n25992 ;
  assign n25994 = n25614 & n25993 ;
  assign n25995 = ~n25614 & ~n25993 ;
  assign n25996 = ~n25994 & ~n25995 ;
  assign n25997 = n25586 & n25996 ;
  assign n25998 = ~n25586 & ~n25996 ;
  assign n25999 = ~n25997 & ~n25998 ;
  assign n26000 = ~n25562 & n25999 ;
  assign n26001 = ~n25560 & n26000 ;
  assign n26002 = ~n25560 & ~n25562 ;
  assign n26003 = ~n25999 & ~n26002 ;
  assign n26004 = ~n26001 & ~n26003 ;
  assign n26005 = ~n24844 & ~n25310 ;
  assign n26006 = n1965 & n14052 ;
  assign n26007 = ~n14049 & n26006 ;
  assign n26008 = n1965 & ~n14052 ;
  assign n26009 = ~n13519 & n26008 ;
  assign n26010 = ~n14048 & n26009 ;
  assign n26011 = \b[50]  & n1963 ;
  assign n26012 = \a[18]  & \b[49]  ;
  assign n26013 = n2210 & n26012 ;
  assign n26014 = ~n26011 & ~n26013 ;
  assign n26015 = \b[48]  & n2218 ;
  assign n26016 = n2216 & n26015 ;
  assign n26017 = ~\a[18]  & \b[49]  ;
  assign n26018 = n1957 & n26017 ;
  assign n26019 = ~n26016 & ~n26018 ;
  assign n26020 = n26014 & n26019 ;
  assign n26021 = ~n26010 & n26020 ;
  assign n26022 = ~n26007 & n26021 ;
  assign n26023 = \a[20]  & ~n26022 ;
  assign n26024 = ~\a[20]  & n26022 ;
  assign n26025 = ~n26023 & ~n26024 ;
  assign n26026 = ~n26005 & n26025 ;
  assign n26027 = ~\a[20]  & ~n26022 ;
  assign n26028 = \a[20]  & n26020 ;
  assign n26029 = ~n26010 & n26028 ;
  assign n26030 = ~n26007 & n26029 ;
  assign n26031 = ~n26027 & ~n26030 ;
  assign n26032 = n26005 & n26031 ;
  assign n26033 = ~n26026 & ~n26032 ;
  assign n26034 = n26004 & n26033 ;
  assign n26035 = ~n26004 & ~n26033 ;
  assign n26036 = ~n26034 & ~n26035 ;
  assign n26037 = ~n25539 & n26036 ;
  assign n26038 = ~n25533 & n26037 ;
  assign n26039 = ~n25533 & ~n25539 ;
  assign n26040 = ~n26036 & ~n26039 ;
  assign n26041 = ~n26038 & ~n26040 ;
  assign n26042 = n25512 & n26041 ;
  assign n26043 = ~n25512 & ~n26041 ;
  assign n26044 = ~n26042 & ~n26043 ;
  assign n26045 = ~n25481 & n26044 ;
  assign n26046 = ~n25479 & n26045 ;
  assign n26047 = ~n25479 & ~n25481 ;
  assign n26048 = ~n26044 & ~n26047 ;
  assign n26049 = ~n26046 & ~n26048 ;
  assign n26050 = ~\a[8]  & ~n25454 ;
  assign n26051 = \a[8]  & n25453 ;
  assign n26052 = ~n25443 & n26051 ;
  assign n26053 = ~n26050 & ~n26052 ;
  assign n26054 = ~n25362 & n26053 ;
  assign n26055 = ~n25440 & n26054 ;
  assign n26056 = n26049 & ~n26055 ;
  assign n26057 = ~n25458 & n26056 ;
  assign n26058 = ~n25458 & ~n26055 ;
  assign n26059 = ~n26049 & ~n26058 ;
  assign n26060 = ~n26057 & ~n26059 ;
  assign n26061 = \b[63]  & n252 ;
  assign n26062 = ~n21694 & n26061 ;
  assign n26063 = ~n23171 & n26062 ;
  assign n26064 = \a[2]  & \a[4]  ;
  assign n26065 = \a[3]  & ~\a[5]  ;
  assign n26066 = n26064 & n26065 ;
  assign n26067 = ~\a[2]  & ~\a[4]  ;
  assign n26068 = ~\a[3]  & \a[5]  ;
  assign n26069 = n26067 & n26068 ;
  assign n26070 = ~n26066 & ~n26069 ;
  assign n26071 = \b[63]  & ~n26070 ;
  assign n26072 = \a[5]  & ~n26071 ;
  assign n26073 = ~n26063 & n26072 ;
  assign n26074 = ~n26063 & ~n26071 ;
  assign n26075 = ~\a[5]  & ~n26074 ;
  assign n26076 = ~n26073 & ~n26075 ;
  assign n26077 = n25391 & ~n26076 ;
  assign n26078 = n25371 & ~n26076 ;
  assign n26079 = ~n25396 & n26078 ;
  assign n26080 = ~n26077 & ~n26079 ;
  assign n26081 = n25371 & ~n25396 ;
  assign n26082 = ~n25391 & n26076 ;
  assign n26083 = ~n26081 & n26082 ;
  assign n26084 = n26080 & ~n26083 ;
  assign n26085 = n26060 & n26084 ;
  assign n26086 = ~n26060 & ~n26084 ;
  assign n26087 = ~n26085 & ~n26086 ;
  assign n26088 = n25439 & n26087 ;
  assign n26089 = ~n25439 & ~n26087 ;
  assign n26090 = ~n26088 & ~n26089 ;
  assign n26091 = ~n25437 & n26090 ;
  assign n26092 = ~n25429 & ~n26090 ;
  assign n26093 = ~n25433 & n26092 ;
  assign n26094 = ~n26091 & ~n26093 ;
  assign n26095 = ~n25429 & ~n26088 ;
  assign n26096 = ~n25433 & n26095 ;
  assign n26097 = ~n26060 & n26080 ;
  assign n26098 = n26080 & n26083 ;
  assign n26099 = ~n26097 & ~n26098 ;
  assign n26100 = ~n25458 & ~n26056 ;
  assign n26101 = n430 & ~n22461 ;
  assign n26102 = ~n22459 & n26101 ;
  assign n26103 = \b[63]  & n428 ;
  assign n26104 = \a[6]  & \b[62]  ;
  assign n26105 = n419 & n26104 ;
  assign n26106 = ~n26103 & ~n26105 ;
  assign n26107 = \b[61]  & n486 ;
  assign n26108 = n483 & n26107 ;
  assign n26109 = ~\a[6]  & \b[62]  ;
  assign n26110 = n422 & n26109 ;
  assign n26111 = ~n26108 & ~n26110 ;
  assign n26112 = n26106 & n26111 ;
  assign n26113 = ~n26102 & n26112 ;
  assign n26114 = ~\a[8]  & ~n26113 ;
  assign n26115 = \a[8]  & n26112 ;
  assign n26116 = ~n26102 & n26115 ;
  assign n26117 = ~n26114 & ~n26116 ;
  assign n26118 = ~n25479 & ~n26045 ;
  assign n26119 = ~n25505 & ~n26041 ;
  assign n26120 = ~n25505 & n25511 ;
  assign n26121 = ~n26119 & ~n26120 ;
  assign n26122 = ~n25539 & ~n26036 ;
  assign n26123 = ~n25533 & ~n26122 ;
  assign n26124 = n1965 & ~n14098 ;
  assign n26125 = ~n14096 & n26124 ;
  assign n26126 = \b[51]  & n1963 ;
  assign n26127 = \a[18]  & \b[50]  ;
  assign n26128 = n2210 & n26127 ;
  assign n26129 = ~n26126 & ~n26128 ;
  assign n26130 = \b[49]  & n2218 ;
  assign n26131 = n2216 & n26130 ;
  assign n26132 = ~\a[18]  & \b[50]  ;
  assign n26133 = n1957 & n26132 ;
  assign n26134 = ~n26131 & ~n26133 ;
  assign n26135 = n26129 & n26134 ;
  assign n26136 = ~n26125 & n26135 ;
  assign n26137 = ~\a[20]  & ~n26136 ;
  assign n26138 = \a[20]  & n26135 ;
  assign n26139 = ~n26125 & n26138 ;
  assign n26140 = ~n26137 & ~n26139 ;
  assign n26141 = n26026 & ~n26140 ;
  assign n26142 = n26004 & ~n26140 ;
  assign n26143 = ~n26032 & n26142 ;
  assign n26144 = ~n26141 & ~n26143 ;
  assign n26145 = n26004 & ~n26032 ;
  assign n26146 = ~n26026 & n26140 ;
  assign n26147 = ~n26145 & n26146 ;
  assign n26148 = n26144 & ~n26147 ;
  assign n26149 = n1467 & ~n16398 ;
  assign n26150 = ~n15241 & n26149 ;
  assign n26151 = ~n16404 & n26150 ;
  assign n26152 = n1467 & n16398 ;
  assign n26153 = n15241 & n26152 ;
  assign n26154 = n16400 & n26152 ;
  assign n26155 = ~n15239 & n26154 ;
  assign n26156 = ~n26153 & ~n26155 ;
  assign n26157 = ~n26151 & n26156 ;
  assign n26158 = \b[52]  & n1652 ;
  assign n26159 = n1649 & n26158 ;
  assign n26160 = ~\a[15]  & \b[53]  ;
  assign n26161 = n1459 & n26160 ;
  assign n26162 = ~n26159 & ~n26161 ;
  assign n26163 = \b[54]  & n1465 ;
  assign n26164 = \a[15]  & \b[53]  ;
  assign n26165 = n1456 & n26164 ;
  assign n26166 = \a[17]  & ~n26165 ;
  assign n26167 = ~n26163 & n26166 ;
  assign n26168 = n26162 & n26167 ;
  assign n26169 = n26157 & n26168 ;
  assign n26170 = ~n26163 & ~n26165 ;
  assign n26171 = n26162 & n26170 ;
  assign n26172 = n26157 & n26171 ;
  assign n26173 = ~\a[17]  & ~n26172 ;
  assign n26174 = ~n26169 & ~n26173 ;
  assign n26175 = ~n25560 & ~n26000 ;
  assign n26176 = ~n25580 & ~n25996 ;
  assign n26177 = ~n25580 & n25585 ;
  assign n26178 = ~n26176 & ~n26177 ;
  assign n26179 = ~n25613 & ~n25993 ;
  assign n26180 = ~n25605 & ~n26179 ;
  assign n26181 = n5211 & ~n8602 ;
  assign n26182 = ~n8600 & n26181 ;
  assign n26183 = \b[37]  & n5595 ;
  assign n26184 = n5592 & n26183 ;
  assign n26185 = ~\a[30]  & \b[38]  ;
  assign n26186 = n5203 & n26185 ;
  assign n26187 = ~n26184 & ~n26186 ;
  assign n26188 = \b[39]  & n5209 ;
  assign n26189 = \a[30]  & \b[38]  ;
  assign n26190 = n5200 & n26189 ;
  assign n26191 = \a[32]  & ~n26190 ;
  assign n26192 = ~n26188 & n26191 ;
  assign n26193 = n26187 & n26192 ;
  assign n26194 = ~n26182 & n26193 ;
  assign n26195 = ~n26188 & ~n26190 ;
  assign n26196 = n26187 & n26195 ;
  assign n26197 = ~n26182 & n26196 ;
  assign n26198 = ~\a[32]  & ~n26197 ;
  assign n26199 = ~n26194 & ~n26198 ;
  assign n26200 = n25646 & n26199 ;
  assign n26201 = ~n25990 & n26199 ;
  assign n26202 = ~n25640 & n26201 ;
  assign n26203 = ~n26200 & ~n26202 ;
  assign n26204 = ~n25640 & ~n25990 ;
  assign n26205 = ~n25646 & ~n26199 ;
  assign n26206 = ~n26204 & n26205 ;
  assign n26207 = n26203 & ~n26206 ;
  assign n26208 = n4249 & n9930 ;
  assign n26209 = ~n9927 & n26208 ;
  assign n26210 = n4249 & ~n9930 ;
  assign n26211 = ~n9477 & n26210 ;
  assign n26212 = ~n9926 & n26211 ;
  assign n26213 = \b[40]  & n4647 ;
  assign n26214 = n4644 & n26213 ;
  assign n26215 = ~\a[27]  & \b[41]  ;
  assign n26216 = n4241 & n26215 ;
  assign n26217 = ~n26214 & ~n26216 ;
  assign n26218 = \b[42]  & n4247 ;
  assign n26219 = \a[27]  & \b[41]  ;
  assign n26220 = n4238 & n26219 ;
  assign n26221 = \a[29]  & ~n26220 ;
  assign n26222 = ~n26218 & n26221 ;
  assign n26223 = n26217 & n26222 ;
  assign n26224 = ~n26212 & n26223 ;
  assign n26225 = ~n26209 & n26224 ;
  assign n26226 = ~n26218 & ~n26220 ;
  assign n26227 = n26217 & n26226 ;
  assign n26228 = ~n26212 & n26227 ;
  assign n26229 = ~n26209 & n26228 ;
  assign n26230 = ~\a[29]  & ~n26229 ;
  assign n26231 = ~n26225 & ~n26230 ;
  assign n26232 = ~n25958 & ~n25962 ;
  assign n26233 = ~n1230 & n16655 ;
  assign n26234 = ~n1086 & n16655 ;
  assign n26235 = ~n1226 & n26234 ;
  assign n26236 = ~n26233 & ~n26235 ;
  assign n26237 = ~n1233 & ~n26236 ;
  assign n26238 = \b[13]  & n17308 ;
  assign n26239 = n17305 & n26238 ;
  assign n26240 = ~\a[54]  & \b[14]  ;
  assign n26241 = n16647 & n26240 ;
  assign n26242 = ~n26239 & ~n26241 ;
  assign n26243 = \b[15]  & n16653 ;
  assign n26244 = \a[54]  & \b[14]  ;
  assign n26245 = n16644 & n26244 ;
  assign n26246 = \a[56]  & ~n26245 ;
  assign n26247 = ~n26243 & n26246 ;
  assign n26248 = n26242 & n26247 ;
  assign n26249 = ~n26237 & n26248 ;
  assign n26250 = ~n26243 & ~n26245 ;
  assign n26251 = n26242 & n26250 ;
  assign n26252 = ~\a[56]  & ~n26251 ;
  assign n26253 = ~\a[56]  & ~n1233 ;
  assign n26254 = ~n26236 & n26253 ;
  assign n26255 = ~n26252 & ~n26254 ;
  assign n26256 = ~n26249 & n26255 ;
  assign n26257 = ~n25726 & n25746 ;
  assign n26258 = ~n25725 & ~n26257 ;
  assign n26259 = ~n909 & ~n17912 ;
  assign n26260 = ~n18513 & n26259 ;
  assign n26261 = n906 & n26260 ;
  assign n26262 = n909 & ~n17912 ;
  assign n26263 = ~n18513 & n26262 ;
  assign n26264 = ~n906 & n26263 ;
  assign n26265 = ~n26261 & ~n26264 ;
  assign n26266 = \b[10]  & n19183 ;
  assign n26267 = n19180 & n26266 ;
  assign n26268 = ~\a[57]  & \b[11]  ;
  assign n26269 = n18508 & n26268 ;
  assign n26270 = ~n26267 & ~n26269 ;
  assign n26271 = \b[12]  & n18514 ;
  assign n26272 = \a[57]  & \b[11]  ;
  assign n26273 = n18505 & n26272 ;
  assign n26274 = \a[59]  & ~n26273 ;
  assign n26275 = ~n26271 & n26274 ;
  assign n26276 = n26270 & n26275 ;
  assign n26277 = n26265 & n26276 ;
  assign n26278 = ~n26271 & ~n26273 ;
  assign n26279 = n26270 & n26278 ;
  assign n26280 = n26265 & n26279 ;
  assign n26281 = ~\a[59]  & ~n26280 ;
  assign n26282 = ~n26277 & ~n26281 ;
  assign n26283 = ~\a[2]  & ~\a[5]  ;
  assign n26284 = \a[2]  & \a[5]  ;
  assign n26285 = ~n26283 & ~n26284 ;
  assign n26286 = \b[6]  & n21958 ;
  assign n26287 = \b[5]  & n21957 ;
  assign n26288 = ~n26286 & ~n26287 ;
  assign n26289 = ~n26285 & ~n26288 ;
  assign n26290 = n26285 & ~n26287 ;
  assign n26291 = ~n26286 & n26290 ;
  assign n26292 = ~n26289 & ~n26291 ;
  assign n26293 = n25718 & n26292 ;
  assign n26294 = ~n25715 & n26293 ;
  assign n26295 = ~n25710 & n26294 ;
  assign n26296 = ~n25715 & n25718 ;
  assign n26297 = ~n25710 & n26296 ;
  assign n26298 = ~n26292 & ~n26297 ;
  assign n26299 = ~n26295 & ~n26298 ;
  assign n26300 = ~n586 & n20521 ;
  assign n26301 = ~n504 & n20521 ;
  assign n26302 = ~n508 & n26301 ;
  assign n26303 = ~n26300 & ~n26302 ;
  assign n26304 = ~n589 & ~n26303 ;
  assign n26305 = \b[7]  & n21315 ;
  assign n26306 = n21312 & n26305 ;
  assign n26307 = ~\a[60]  & \b[8]  ;
  assign n26308 = n20513 & n26307 ;
  assign n26309 = ~n26306 & ~n26308 ;
  assign n26310 = \b[9]  & n20519 ;
  assign n26311 = \a[60]  & \b[8]  ;
  assign n26312 = n20510 & n26311 ;
  assign n26313 = \a[62]  & ~n26312 ;
  assign n26314 = ~n26310 & n26313 ;
  assign n26315 = n26309 & n26314 ;
  assign n26316 = ~n26304 & n26315 ;
  assign n26317 = ~n26310 & ~n26312 ;
  assign n26318 = n26309 & n26317 ;
  assign n26319 = ~\a[62]  & ~n26318 ;
  assign n26320 = ~\a[62]  & ~n589 ;
  assign n26321 = ~n26303 & n26320 ;
  assign n26322 = ~n26319 & ~n26321 ;
  assign n26323 = ~n26316 & n26322 ;
  assign n26324 = ~n26299 & n26323 ;
  assign n26325 = ~n26295 & ~n26323 ;
  assign n26326 = ~n26298 & n26325 ;
  assign n26327 = ~n26324 & ~n26326 ;
  assign n26328 = ~n26282 & n26327 ;
  assign n26329 = n26282 & ~n26327 ;
  assign n26330 = ~n26328 & ~n26329 ;
  assign n26331 = n26258 & n26330 ;
  assign n26332 = ~n26258 & ~n26330 ;
  assign n26333 = ~n26331 & ~n26332 ;
  assign n26334 = ~n25752 & n25781 ;
  assign n26335 = n25757 & ~n26334 ;
  assign n26336 = ~n26333 & ~n26335 ;
  assign n26337 = n26256 & n26336 ;
  assign n26338 = n26333 & ~n26335 ;
  assign n26339 = ~n26256 & n26338 ;
  assign n26340 = ~n26337 & ~n26339 ;
  assign n26341 = n25757 & ~n26256 ;
  assign n26342 = ~n26334 & n26341 ;
  assign n26343 = ~n26333 & n26342 ;
  assign n26344 = n25757 & n26256 ;
  assign n26345 = ~n26334 & n26344 ;
  assign n26346 = n26333 & n26345 ;
  assign n26347 = ~n26343 & ~n26346 ;
  assign n26348 = n1875 & n14793 ;
  assign n26349 = ~n1872 & n26348 ;
  assign n26350 = ~n1875 & n14793 ;
  assign n26351 = ~n1689 & n26350 ;
  assign n26352 = ~n1871 & n26351 ;
  assign n26353 = \b[16]  & n15517 ;
  assign n26354 = n15514 & n26353 ;
  assign n26355 = ~\a[51]  & \b[17]  ;
  assign n26356 = n14785 & n26355 ;
  assign n26357 = ~n26354 & ~n26356 ;
  assign n26358 = \b[18]  & n14791 ;
  assign n26359 = \a[51]  & \b[17]  ;
  assign n26360 = n14782 & n26359 ;
  assign n26361 = \a[53]  & ~n26360 ;
  assign n26362 = ~n26358 & n26361 ;
  assign n26363 = n26357 & n26362 ;
  assign n26364 = ~n26352 & n26363 ;
  assign n26365 = ~n26349 & n26364 ;
  assign n26366 = ~n26358 & ~n26360 ;
  assign n26367 = n26357 & n26366 ;
  assign n26368 = ~n26352 & n26367 ;
  assign n26369 = ~n26349 & n26368 ;
  assign n26370 = ~\a[53]  & ~n26369 ;
  assign n26371 = ~n26365 & ~n26370 ;
  assign n26372 = n26347 & ~n26371 ;
  assign n26373 = n26340 & n26372 ;
  assign n26374 = n26340 & n26347 ;
  assign n26375 = n26371 & ~n26374 ;
  assign n26376 = ~n26373 & ~n26375 ;
  assign n26377 = n25678 & ~n25785 ;
  assign n26378 = ~n25786 & ~n26377 ;
  assign n26379 = ~n26376 & ~n26378 ;
  assign n26380 = ~n26373 & n26378 ;
  assign n26381 = ~n26375 & n26380 ;
  assign n26382 = ~n2523 & n13125 ;
  assign n26383 = ~n2521 & n26382 ;
  assign n26384 = \b[21]  & n13123 ;
  assign n26385 = \a[48]  & \b[20]  ;
  assign n26386 = n13786 & n26385 ;
  assign n26387 = ~n26384 & ~n26386 ;
  assign n26388 = \b[19]  & n13794 ;
  assign n26389 = n13792 & n26388 ;
  assign n26390 = ~\a[48]  & \b[20]  ;
  assign n26391 = n13117 & n26390 ;
  assign n26392 = ~n26389 & ~n26391 ;
  assign n26393 = n26387 & n26392 ;
  assign n26394 = ~n26383 & n26393 ;
  assign n26395 = ~\a[50]  & ~n26394 ;
  assign n26396 = \a[50]  & n26393 ;
  assign n26397 = ~n26383 & n26396 ;
  assign n26398 = ~n26395 & ~n26397 ;
  assign n26399 = ~n26381 & ~n26398 ;
  assign n26400 = ~n26379 & n26399 ;
  assign n26401 = ~n26378 & n26398 ;
  assign n26402 = ~n26376 & n26401 ;
  assign n26403 = n26378 & n26398 ;
  assign n26404 = n26376 & n26403 ;
  assign n26405 = ~n26402 & ~n26404 ;
  assign n26406 = ~n26400 & n26405 ;
  assign n26407 = n3283 & n11572 ;
  assign n26408 = ~n3280 & n26407 ;
  assign n26409 = ~n3283 & n11572 ;
  assign n26410 = ~n3017 & n26409 ;
  assign n26411 = ~n3279 & n26410 ;
  assign n26412 = \b[22]  & n12159 ;
  assign n26413 = n12156 & n26412 ;
  assign n26414 = ~\a[45]  & \b[23]  ;
  assign n26415 = n11564 & n26414 ;
  assign n26416 = ~n26413 & ~n26415 ;
  assign n26417 = \b[24]  & n11570 ;
  assign n26418 = \a[45]  & \b[23]  ;
  assign n26419 = n11561 & n26418 ;
  assign n26420 = \a[47]  & ~n26419 ;
  assign n26421 = ~n26417 & n26420 ;
  assign n26422 = n26416 & n26421 ;
  assign n26423 = ~n26411 & n26422 ;
  assign n26424 = ~n26408 & n26423 ;
  assign n26425 = ~n26417 & ~n26419 ;
  assign n26426 = n26416 & n26425 ;
  assign n26427 = ~n26411 & n26426 ;
  assign n26428 = ~n26408 & n26427 ;
  assign n26429 = ~\a[47]  & ~n26428 ;
  assign n26430 = ~n26424 & ~n26429 ;
  assign n26431 = ~n25790 & ~n25792 ;
  assign n26432 = n25826 & ~n26431 ;
  assign n26433 = ~n26430 & ~n26432 ;
  assign n26434 = ~n26406 & n26433 ;
  assign n26435 = ~n26430 & n26432 ;
  assign n26436 = n26406 & n26435 ;
  assign n26437 = ~n26434 & ~n26436 ;
  assign n26438 = n26430 & n26432 ;
  assign n26439 = ~n26406 & n26438 ;
  assign n26440 = n26430 & ~n26432 ;
  assign n26441 = n26406 & n26440 ;
  assign n26442 = ~n26439 & ~n26441 ;
  assign n26443 = n26437 & n26442 ;
  assign n26444 = ~n25827 & ~n25829 ;
  assign n26445 = n25827 & n25829 ;
  assign n26446 = n25848 & ~n26445 ;
  assign n26447 = ~n26444 & ~n26446 ;
  assign n26448 = ~n4148 & n10082 ;
  assign n26449 = ~n4146 & n26448 ;
  assign n26450 = \b[27]  & n10080 ;
  assign n26451 = \a[42]  & \b[26]  ;
  assign n26452 = n10071 & n26451 ;
  assign n26453 = ~n26450 & ~n26452 ;
  assign n26454 = \b[25]  & n10681 ;
  assign n26455 = n10678 & n26454 ;
  assign n26456 = ~\a[42]  & \b[26]  ;
  assign n26457 = n10074 & n26456 ;
  assign n26458 = ~n26455 & ~n26457 ;
  assign n26459 = n26453 & n26458 ;
  assign n26460 = ~n26449 & n26459 ;
  assign n26461 = ~\a[44]  & ~n26460 ;
  assign n26462 = \a[44]  & n26459 ;
  assign n26463 = ~n26449 & n26462 ;
  assign n26464 = ~n26461 & ~n26463 ;
  assign n26465 = ~n26447 & ~n26464 ;
  assign n26466 = n26443 & n26465 ;
  assign n26467 = n26447 & ~n26464 ;
  assign n26468 = ~n26443 & n26467 ;
  assign n26469 = ~n26466 & ~n26468 ;
  assign n26470 = ~n26447 & n26464 ;
  assign n26471 = ~n26443 & n26470 ;
  assign n26472 = n26447 & n26464 ;
  assign n26473 = n26443 & n26472 ;
  assign n26474 = ~n26471 & ~n26473 ;
  assign n26475 = n26469 & n26474 ;
  assign n26476 = ~n25659 & ~n25859 ;
  assign n26477 = n25659 & n25859 ;
  assign n26478 = n25883 & ~n26477 ;
  assign n26479 = ~n26476 & ~n26478 ;
  assign n26480 = ~n26475 & ~n26479 ;
  assign n26481 = n26475 & n26479 ;
  assign n26482 = ~n26480 & ~n26481 ;
  assign n26483 = ~n5105 & ~n8272 ;
  assign n26484 = ~n8756 & n26483 ;
  assign n26485 = n5102 & n26484 ;
  assign n26486 = n5105 & ~n8272 ;
  assign n26487 = ~n8756 & n26486 ;
  assign n26488 = ~n5102 & n26487 ;
  assign n26489 = ~n26485 & ~n26488 ;
  assign n26490 = \b[28]  & n9301 ;
  assign n26491 = n9298 & n26490 ;
  assign n26492 = ~\a[39]  & \b[29]  ;
  assign n26493 = n8751 & n26492 ;
  assign n26494 = ~n26491 & ~n26493 ;
  assign n26495 = \b[30]  & n8757 ;
  assign n26496 = \a[39]  & \b[29]  ;
  assign n26497 = n8748 & n26496 ;
  assign n26498 = \a[41]  & ~n26497 ;
  assign n26499 = ~n26495 & n26498 ;
  assign n26500 = n26494 & n26499 ;
  assign n26501 = n26489 & n26500 ;
  assign n26502 = ~n26495 & ~n26497 ;
  assign n26503 = n26494 & n26502 ;
  assign n26504 = n26489 & n26503 ;
  assign n26505 = ~\a[41]  & ~n26504 ;
  assign n26506 = ~n26501 & ~n26505 ;
  assign n26507 = ~n26482 & n26506 ;
  assign n26508 = n26482 & ~n26506 ;
  assign n26509 = ~n26507 & ~n26508 ;
  assign n26510 = ~n5852 & n7534 ;
  assign n26511 = ~n5809 & n7534 ;
  assign n26512 = ~n5848 & n26511 ;
  assign n26513 = ~n26510 & ~n26512 ;
  assign n26514 = ~n5855 & ~n26513 ;
  assign n26515 = \b[31]  & n7973 ;
  assign n26516 = n7970 & n26515 ;
  assign n26517 = ~\a[36]  & \b[32]  ;
  assign n26518 = n7526 & n26517 ;
  assign n26519 = ~n26516 & ~n26518 ;
  assign n26520 = \b[33]  & n7532 ;
  assign n26521 = \a[36]  & \b[32]  ;
  assign n26522 = n17801 & n26521 ;
  assign n26523 = \a[38]  & ~n26522 ;
  assign n26524 = ~n26520 & n26523 ;
  assign n26525 = n26519 & n26524 ;
  assign n26526 = ~n26514 & n26525 ;
  assign n26527 = ~n26520 & ~n26522 ;
  assign n26528 = n26519 & n26527 ;
  assign n26529 = ~\a[38]  & ~n26528 ;
  assign n26530 = ~\a[38]  & ~n5855 ;
  assign n26531 = ~n26513 & n26530 ;
  assign n26532 = ~n26529 & ~n26531 ;
  assign n26533 = ~n26526 & n26532 ;
  assign n26534 = n25655 & n25894 ;
  assign n26535 = ~n25193 & ~n25918 ;
  assign n26536 = n25654 & n26535 ;
  assign n26537 = ~n25921 & ~n26536 ;
  assign n26538 = ~n26534 & n26537 ;
  assign n26539 = ~n26533 & n26538 ;
  assign n26540 = n26509 & n26539 ;
  assign n26541 = ~n26533 & ~n26538 ;
  assign n26542 = ~n26509 & n26541 ;
  assign n26543 = ~n26540 & ~n26542 ;
  assign n26544 = n26533 & n26538 ;
  assign n26545 = ~n26509 & n26544 ;
  assign n26546 = n26533 & ~n26538 ;
  assign n26547 = n26509 & n26546 ;
  assign n26548 = ~n26545 & ~n26547 ;
  assign n26549 = n26543 & n26548 ;
  assign n26550 = ~n26232 & n26549 ;
  assign n26551 = n6309 & n7337 ;
  assign n26552 = ~n7334 & n26551 ;
  assign n26553 = n6309 & n24138 ;
  assign n26554 = ~n7333 & n26553 ;
  assign n26555 = \b[34]  & n6778 ;
  assign n26556 = n6775 & n26555 ;
  assign n26557 = ~\a[33]  & \b[35]  ;
  assign n26558 = n6301 & n26557 ;
  assign n26559 = ~n26556 & ~n26558 ;
  assign n26560 = \b[36]  & n6307 ;
  assign n26561 = \a[33]  & \b[35]  ;
  assign n26562 = n6298 & n26561 ;
  assign n26563 = \a[35]  & ~n26562 ;
  assign n26564 = ~n26560 & n26563 ;
  assign n26565 = n26559 & n26564 ;
  assign n26566 = ~n26554 & n26565 ;
  assign n26567 = ~n26552 & n26566 ;
  assign n26568 = ~n26560 & ~n26562 ;
  assign n26569 = n26559 & n26568 ;
  assign n26570 = ~n26554 & n26569 ;
  assign n26571 = ~n26552 & n26570 ;
  assign n26572 = ~\a[35]  & ~n26571 ;
  assign n26573 = ~n26567 & ~n26572 ;
  assign n26574 = ~n25958 & ~n26549 ;
  assign n26575 = ~n25962 & n26574 ;
  assign n26576 = ~n26573 & ~n26575 ;
  assign n26577 = ~n26550 & n26576 ;
  assign n26578 = ~n26549 & n26573 ;
  assign n26579 = n26232 & n26578 ;
  assign n26580 = n26549 & n26573 ;
  assign n26581 = ~n26232 & n26580 ;
  assign n26582 = ~n26579 & ~n26581 ;
  assign n26583 = ~n26577 & n26582 ;
  assign n26584 = ~n25966 & n25987 ;
  assign n26585 = ~n25967 & ~n26584 ;
  assign n26586 = ~n26583 & ~n26585 ;
  assign n26587 = n26583 & n26585 ;
  assign n26588 = ~n26586 & ~n26587 ;
  assign n26589 = ~n26231 & n26588 ;
  assign n26590 = ~n26207 & n26589 ;
  assign n26591 = ~n26231 & ~n26588 ;
  assign n26592 = n26207 & n26591 ;
  assign n26593 = ~n26590 & ~n26592 ;
  assign n26594 = ~n26180 & ~n26593 ;
  assign n26595 = n26231 & n26588 ;
  assign n26596 = ~n26207 & n26595 ;
  assign n26597 = n26231 & ~n26588 ;
  assign n26598 = n26207 & n26597 ;
  assign n26599 = ~n26596 & ~n26598 ;
  assign n26600 = ~n25605 & ~n26599 ;
  assign n26601 = ~n26179 & n26600 ;
  assign n26602 = ~n26594 & ~n26601 ;
  assign n26603 = n26207 & n26588 ;
  assign n26604 = ~n26207 & ~n26588 ;
  assign n26605 = ~n26603 & ~n26604 ;
  assign n26606 = n26231 & ~n26605 ;
  assign n26607 = ~n26180 & n26606 ;
  assign n26608 = ~n26207 & n26591 ;
  assign n26609 = n26207 & n26589 ;
  assign n26610 = ~n26608 & ~n26609 ;
  assign n26611 = ~n25605 & ~n26610 ;
  assign n26612 = ~n26179 & n26611 ;
  assign n26613 = ~n26607 & ~n26612 ;
  assign n26614 = n26602 & n26613 ;
  assign n26615 = n2622 & n12478 ;
  assign n26616 = ~n12475 & n26615 ;
  assign n26617 = n2622 & ~n12478 ;
  assign n26618 = ~n12433 & n26617 ;
  assign n26619 = ~n12474 & n26618 ;
  assign n26620 = \b[46]  & n2912 ;
  assign n26621 = n2909 & n26620 ;
  assign n26622 = ~\a[21]  & \b[47]  ;
  assign n26623 = n2614 & n26622 ;
  assign n26624 = ~n26621 & ~n26623 ;
  assign n26625 = \b[48]  & n2620 ;
  assign n26626 = \a[21]  & \b[47]  ;
  assign n26627 = n20849 & n26626 ;
  assign n26628 = \a[23]  & ~n26627 ;
  assign n26629 = ~n26625 & n26628 ;
  assign n26630 = n26624 & n26629 ;
  assign n26631 = ~n26619 & n26630 ;
  assign n26632 = ~n26616 & n26631 ;
  assign n26633 = ~n26625 & ~n26627 ;
  assign n26634 = n26624 & n26633 ;
  assign n26635 = ~n26619 & n26634 ;
  assign n26636 = ~n26616 & n26635 ;
  assign n26637 = ~\a[23]  & ~n26636 ;
  assign n26638 = ~n26632 & ~n26637 ;
  assign n26639 = n3402 & ~n11397 ;
  assign n26640 = ~n11395 & n26639 ;
  assign n26641 = \b[45]  & n3400 ;
  assign n26642 = \a[24]  & \b[44]  ;
  assign n26643 = n3391 & n26642 ;
  assign n26644 = ~n26641 & ~n26643 ;
  assign n26645 = \b[43]  & n3733 ;
  assign n26646 = n3730 & n26645 ;
  assign n26647 = ~\a[24]  & \b[44]  ;
  assign n26648 = n3394 & n26647 ;
  assign n26649 = ~n26646 & ~n26648 ;
  assign n26650 = n26644 & n26649 ;
  assign n26651 = ~n26640 & n26650 ;
  assign n26652 = ~\a[26]  & ~n26651 ;
  assign n26653 = \a[26]  & n26650 ;
  assign n26654 = ~n26640 & n26653 ;
  assign n26655 = ~n26652 & ~n26654 ;
  assign n26656 = ~n26638 & ~n26655 ;
  assign n26657 = ~n26614 & n26656 ;
  assign n26658 = ~n26178 & n26657 ;
  assign n26659 = ~n26638 & n26655 ;
  assign n26660 = n26614 & n26659 ;
  assign n26661 = ~n26178 & n26660 ;
  assign n26662 = ~n26658 & ~n26661 ;
  assign n26663 = n26614 & n26656 ;
  assign n26664 = n26178 & n26663 ;
  assign n26665 = ~n26614 & n26659 ;
  assign n26666 = n26178 & n26665 ;
  assign n26667 = ~n26664 & ~n26666 ;
  assign n26668 = n26662 & n26667 ;
  assign n26669 = ~n26175 & ~n26668 ;
  assign n26670 = n26638 & ~n26655 ;
  assign n26671 = ~n26614 & n26670 ;
  assign n26672 = ~n26178 & n26671 ;
  assign n26673 = n26638 & n26655 ;
  assign n26674 = n26614 & n26673 ;
  assign n26675 = ~n26178 & n26674 ;
  assign n26676 = ~n26672 & ~n26675 ;
  assign n26677 = n26614 & n26670 ;
  assign n26678 = n26178 & n26677 ;
  assign n26679 = ~n26614 & n26673 ;
  assign n26680 = n26178 & n26679 ;
  assign n26681 = ~n26678 & ~n26680 ;
  assign n26682 = n26676 & n26681 ;
  assign n26683 = n26175 & ~n26682 ;
  assign n26684 = ~n26669 & ~n26683 ;
  assign n26685 = ~n26178 & n26655 ;
  assign n26686 = n25996 & ~n26655 ;
  assign n26687 = ~n25585 & n26686 ;
  assign n26688 = n25580 & ~n26655 ;
  assign n26689 = ~n26687 & ~n26688 ;
  assign n26690 = n26614 & n26689 ;
  assign n26691 = ~n26685 & n26690 ;
  assign n26692 = ~n26614 & ~n26655 ;
  assign n26693 = n26178 & n26692 ;
  assign n26694 = ~n26614 & n26655 ;
  assign n26695 = ~n26178 & n26694 ;
  assign n26696 = ~n26693 & ~n26695 ;
  assign n26697 = ~n26691 & n26696 ;
  assign n26698 = n26638 & ~n26697 ;
  assign n26699 = ~n26175 & n26698 ;
  assign n26700 = ~n26178 & n26663 ;
  assign n26701 = ~n26178 & n26665 ;
  assign n26702 = ~n26700 & ~n26701 ;
  assign n26703 = n26178 & n26657 ;
  assign n26704 = n26178 & n26660 ;
  assign n26705 = ~n26703 & ~n26704 ;
  assign n26706 = n26702 & n26705 ;
  assign n26707 = n26175 & ~n26706 ;
  assign n26708 = ~n26699 & ~n26707 ;
  assign n26709 = n26684 & n26708 ;
  assign n26710 = ~n26174 & ~n26709 ;
  assign n26711 = ~n26148 & n26710 ;
  assign n26712 = ~n26174 & n26709 ;
  assign n26713 = n26148 & n26712 ;
  assign n26714 = ~n26711 & ~n26713 ;
  assign n26715 = ~n26123 & ~n26714 ;
  assign n26716 = n26174 & ~n26709 ;
  assign n26717 = ~n26148 & n26716 ;
  assign n26718 = n26174 & n26709 ;
  assign n26719 = n26148 & n26718 ;
  assign n26720 = ~n26717 & ~n26719 ;
  assign n26721 = n26123 & ~n26720 ;
  assign n26722 = ~n26715 & ~n26721 ;
  assign n26723 = n26148 & ~n26709 ;
  assign n26724 = ~n26148 & n26709 ;
  assign n26725 = ~n26723 & ~n26724 ;
  assign n26726 = n26174 & ~n26725 ;
  assign n26727 = ~n26123 & n26726 ;
  assign n26728 = n26148 & n26710 ;
  assign n26729 = ~n26148 & n26712 ;
  assign n26730 = ~n26728 & ~n26729 ;
  assign n26731 = n26123 & ~n26730 ;
  assign n26732 = ~n26727 & ~n26731 ;
  assign n26733 = n26722 & n26732 ;
  assign n26734 = n646 & n20260 ;
  assign n26735 = ~n20257 & n26734 ;
  assign n26736 = n646 & ~n20260 ;
  assign n26737 = ~n19545 & n26736 ;
  assign n26738 = ~n20256 & n26737 ;
  assign n26739 = \b[58]  & n796 ;
  assign n26740 = n793 & n26739 ;
  assign n26741 = ~\a[9]  & \b[59]  ;
  assign n26742 = n638 & n26741 ;
  assign n26743 = ~n26740 & ~n26742 ;
  assign n26744 = \b[60]  & n644 ;
  assign n26745 = \a[9]  & \b[59]  ;
  assign n26746 = n635 & n26745 ;
  assign n26747 = \a[11]  & ~n26746 ;
  assign n26748 = ~n26744 & n26747 ;
  assign n26749 = n26743 & n26748 ;
  assign n26750 = ~n26738 & n26749 ;
  assign n26751 = ~n26735 & n26750 ;
  assign n26752 = ~n26744 & ~n26746 ;
  assign n26753 = n26743 & n26752 ;
  assign n26754 = ~n26738 & n26753 ;
  assign n26755 = ~n26735 & n26754 ;
  assign n26756 = ~\a[11]  & ~n26755 ;
  assign n26757 = ~n26751 & ~n26756 ;
  assign n26758 = n999 & ~n17690 ;
  assign n26759 = ~n17688 & n26758 ;
  assign n26760 = \b[55]  & n1182 ;
  assign n26761 = n1179 & n26760 ;
  assign n26762 = \b[57]  & n997 ;
  assign n26763 = \a[11]  & \b[56]  ;
  assign n26764 = n1180 & n26763 ;
  assign n26765 = ~\a[12]  & \b[56]  ;
  assign n26766 = n7674 & n26765 ;
  assign n26767 = ~n26764 & ~n26766 ;
  assign n26768 = ~n26762 & n26767 ;
  assign n26769 = ~n26761 & n26768 ;
  assign n26770 = ~n26759 & n26769 ;
  assign n26771 = ~\a[14]  & ~n26770 ;
  assign n26772 = \a[14]  & n26769 ;
  assign n26773 = ~n26759 & n26772 ;
  assign n26774 = ~n26771 & ~n26773 ;
  assign n26775 = ~n26757 & ~n26774 ;
  assign n26776 = ~n26733 & n26775 ;
  assign n26777 = ~n26121 & n26776 ;
  assign n26778 = ~n26757 & n26774 ;
  assign n26779 = n26733 & n26778 ;
  assign n26780 = ~n26121 & n26779 ;
  assign n26781 = ~n26777 & ~n26780 ;
  assign n26782 = ~n26733 & n26778 ;
  assign n26783 = n26121 & n26782 ;
  assign n26784 = n26733 & n26775 ;
  assign n26785 = n26121 & n26784 ;
  assign n26786 = ~n26783 & ~n26785 ;
  assign n26787 = n26781 & n26786 ;
  assign n26788 = ~n26118 & ~n26787 ;
  assign n26789 = n26757 & ~n26774 ;
  assign n26790 = ~n26733 & n26789 ;
  assign n26791 = ~n26121 & n26790 ;
  assign n26792 = n26757 & n26774 ;
  assign n26793 = n26733 & n26792 ;
  assign n26794 = ~n26121 & n26793 ;
  assign n26795 = ~n26791 & ~n26794 ;
  assign n26796 = ~n26733 & n26792 ;
  assign n26797 = n26121 & n26796 ;
  assign n26798 = n26733 & n26789 ;
  assign n26799 = n26121 & n26798 ;
  assign n26800 = ~n26797 & ~n26799 ;
  assign n26801 = n26795 & n26800 ;
  assign n26802 = n26118 & ~n26801 ;
  assign n26803 = ~n26788 & ~n26802 ;
  assign n26804 = ~n26121 & n26774 ;
  assign n26805 = n26041 & ~n26774 ;
  assign n26806 = ~n25511 & n26805 ;
  assign n26807 = n25505 & ~n26774 ;
  assign n26808 = ~n26806 & ~n26807 ;
  assign n26809 = n26733 & n26808 ;
  assign n26810 = ~n26804 & n26809 ;
  assign n26811 = ~n26733 & n26774 ;
  assign n26812 = ~n26121 & n26811 ;
  assign n26813 = ~n26733 & ~n26774 ;
  assign n26814 = n26121 & n26813 ;
  assign n26815 = ~n26812 & ~n26814 ;
  assign n26816 = ~n26810 & n26815 ;
  assign n26817 = n26757 & ~n26816 ;
  assign n26818 = ~n26118 & n26817 ;
  assign n26819 = ~n26121 & n26782 ;
  assign n26820 = ~n26121 & n26784 ;
  assign n26821 = ~n26819 & ~n26820 ;
  assign n26822 = n26121 & n26776 ;
  assign n26823 = n26121 & n26779 ;
  assign n26824 = ~n26822 & ~n26823 ;
  assign n26825 = n26821 & n26824 ;
  assign n26826 = n26118 & ~n26825 ;
  assign n26827 = ~n26818 & ~n26826 ;
  assign n26828 = n26803 & n26827 ;
  assign n26829 = ~n26117 & ~n26828 ;
  assign n26830 = n26100 & n26829 ;
  assign n26831 = n26117 & ~n26828 ;
  assign n26832 = ~n26100 & n26831 ;
  assign n26833 = ~n26830 & ~n26832 ;
  assign n26834 = ~n26117 & n26828 ;
  assign n26835 = ~n26100 & n26834 ;
  assign n26836 = n26117 & n26828 ;
  assign n26837 = n26100 & n26836 ;
  assign n26838 = ~n26835 & ~n26837 ;
  assign n26839 = n26833 & n26838 ;
  assign n26840 = n26099 & n26839 ;
  assign n26841 = ~n26099 & ~n26839 ;
  assign n26842 = ~n26840 & ~n26841 ;
  assign n26843 = ~n26089 & n26842 ;
  assign n26844 = ~n26096 & n26843 ;
  assign n26845 = ~n26089 & ~n26096 ;
  assign n26846 = ~n26842 & ~n26845 ;
  assign n26847 = ~n26844 & ~n26846 ;
  assign n26848 = ~n26840 & ~n26844 ;
  assign n26849 = n26100 & n26117 ;
  assign n26850 = ~n26100 & ~n26117 ;
  assign n26851 = n26828 & ~n26850 ;
  assign n26852 = ~n26849 & ~n26851 ;
  assign n26853 = ~n26118 & ~n26757 ;
  assign n26854 = ~n26816 & ~n26853 ;
  assign n26855 = \b[62]  & n486 ;
  assign n26856 = n483 & n26855 ;
  assign n26857 = ~\a[6]  & \b[63]  ;
  assign n26858 = n422 & n26857 ;
  assign n26859 = \a[6]  & \b[63]  ;
  assign n26860 = n419 & n26859 ;
  assign n26861 = ~n26858 & ~n26860 ;
  assign n26862 = ~n26856 & n26861 ;
  assign n26863 = ~\a[8]  & ~n26862 ;
  assign n26864 = n430 & ~n22458 ;
  assign n26865 = ~\a[8]  & n26864 ;
  assign n26866 = ~n23173 & n26865 ;
  assign n26867 = ~n26863 & ~n26866 ;
  assign n26868 = ~n23173 & n26864 ;
  assign n26869 = \a[8]  & n26862 ;
  assign n26870 = ~n26868 & n26869 ;
  assign n26871 = n26867 & ~n26870 ;
  assign n26872 = n26118 & n26757 ;
  assign n26873 = ~n26871 & ~n26872 ;
  assign n26874 = ~n26854 & n26873 ;
  assign n26875 = n26871 & n26872 ;
  assign n26876 = ~n26816 & n26871 ;
  assign n26877 = ~n26853 & n26876 ;
  assign n26878 = ~n26875 & ~n26877 ;
  assign n26879 = ~n26874 & n26878 ;
  assign n26880 = ~n26733 & n26808 ;
  assign n26881 = ~n26804 & ~n26880 ;
  assign n26882 = n646 & ~n20971 ;
  assign n26883 = ~n20969 & n26882 ;
  assign n26884 = \b[61]  & n644 ;
  assign n26885 = \a[9]  & \b[60]  ;
  assign n26886 = n635 & n26885 ;
  assign n26887 = ~n26884 & ~n26886 ;
  assign n26888 = \b[59]  & n796 ;
  assign n26889 = n793 & n26888 ;
  assign n26890 = ~\a[9]  & \b[60]  ;
  assign n26891 = n638 & n26890 ;
  assign n26892 = ~n26889 & ~n26891 ;
  assign n26893 = n26887 & n26892 ;
  assign n26894 = ~n26883 & n26893 ;
  assign n26895 = ~\a[11]  & ~n26894 ;
  assign n26896 = \a[11]  & n26893 ;
  assign n26897 = ~n26883 & n26896 ;
  assign n26898 = ~n26895 & ~n26897 ;
  assign n26899 = ~n26881 & n26898 ;
  assign n26900 = \a[11]  & ~n26894 ;
  assign n26901 = ~\a[11]  & n26894 ;
  assign n26902 = ~n26900 & ~n26901 ;
  assign n26903 = n26881 & n26902 ;
  assign n26904 = ~n26899 & ~n26903 ;
  assign n26905 = n26123 & ~n26174 ;
  assign n26906 = ~n847 & ~n17685 ;
  assign n26907 = ~n18940 & n26906 ;
  assign n26908 = ~n18936 & n26907 ;
  assign n26909 = ~n996 & n26908 ;
  assign n26910 = n999 & n18940 ;
  assign n26911 = ~n18937 & n26910 ;
  assign n26912 = ~n26909 & ~n26911 ;
  assign n26913 = \b[58]  & n997 ;
  assign n26914 = \a[11]  & \b[57]  ;
  assign n26915 = n1180 & n26914 ;
  assign n26916 = ~\a[12]  & \b[57]  ;
  assign n26917 = n7674 & n26916 ;
  assign n26918 = ~n26915 & ~n26917 ;
  assign n26919 = ~n26913 & n26918 ;
  assign n26920 = \b[56]  & n1182 ;
  assign n26921 = n1179 & n26920 ;
  assign n26922 = \a[14]  & ~n26921 ;
  assign n26923 = n26919 & n26922 ;
  assign n26924 = n26912 & n26923 ;
  assign n26925 = n26919 & ~n26921 ;
  assign n26926 = n26912 & n26925 ;
  assign n26927 = ~\a[14]  & ~n26926 ;
  assign n26928 = ~n26924 & ~n26927 ;
  assign n26929 = ~n26905 & n26928 ;
  assign n26930 = n26722 & n26929 ;
  assign n26931 = ~n26174 & ~n26928 ;
  assign n26932 = n26123 & n26931 ;
  assign n26933 = n26725 & n26931 ;
  assign n26934 = n26725 & ~n26928 ;
  assign n26935 = n26123 & n26934 ;
  assign n26936 = ~n26933 & ~n26935 ;
  assign n26937 = ~n26932 & n26936 ;
  assign n26938 = n1467 & ~n16446 ;
  assign n26939 = ~n16444 & n26938 ;
  assign n26940 = \b[55]  & n1465 ;
  assign n26941 = \a[15]  & \b[54]  ;
  assign n26942 = n1456 & n26941 ;
  assign n26943 = ~n26940 & ~n26942 ;
  assign n26944 = \b[53]  & n1652 ;
  assign n26945 = n1649 & n26944 ;
  assign n26946 = ~\a[15]  & \b[54]  ;
  assign n26947 = n1459 & n26946 ;
  assign n26948 = ~n26945 & ~n26947 ;
  assign n26949 = n26943 & n26948 ;
  assign n26950 = ~n26939 & n26949 ;
  assign n26951 = ~\a[17]  & ~n26950 ;
  assign n26952 = \a[17]  & n26949 ;
  assign n26953 = ~n26939 & n26952 ;
  assign n26954 = n26147 & ~n26953 ;
  assign n26955 = n26709 & ~n26953 ;
  assign n26956 = n26144 & n26955 ;
  assign n26957 = ~n26954 & ~n26956 ;
  assign n26958 = ~n26951 & ~n26957 ;
  assign n26959 = n26144 & n26709 ;
  assign n26960 = ~n26951 & ~n26953 ;
  assign n26961 = ~n26147 & ~n26960 ;
  assign n26962 = ~n26959 & n26961 ;
  assign n26963 = ~n26175 & ~n26638 ;
  assign n26964 = ~n26697 & ~n26963 ;
  assign n26965 = n1965 & n15201 ;
  assign n26966 = ~n15198 & n26965 ;
  assign n26967 = n1965 & ~n15201 ;
  assign n26968 = ~n14093 & n26967 ;
  assign n26969 = ~n15197 & n26968 ;
  assign n26970 = \b[50]  & n2218 ;
  assign n26971 = n2216 & n26970 ;
  assign n26972 = ~\a[18]  & \b[51]  ;
  assign n26973 = n1957 & n26972 ;
  assign n26974 = ~n26971 & ~n26973 ;
  assign n26975 = \b[52]  & n1963 ;
  assign n26976 = \a[18]  & \b[51]  ;
  assign n26977 = n2210 & n26976 ;
  assign n26978 = \a[20]  & ~n26977 ;
  assign n26979 = ~n26975 & n26978 ;
  assign n26980 = n26974 & n26979 ;
  assign n26981 = ~n26969 & n26980 ;
  assign n26982 = ~n26966 & n26981 ;
  assign n26983 = ~n26975 & ~n26977 ;
  assign n26984 = n26974 & n26983 ;
  assign n26985 = ~n26969 & n26984 ;
  assign n26986 = ~n26966 & n26985 ;
  assign n26987 = ~\a[20]  & ~n26986 ;
  assign n26988 = ~n26982 & ~n26987 ;
  assign n26989 = n26175 & n26638 ;
  assign n26990 = ~n26988 & ~n26989 ;
  assign n26991 = ~n26964 & n26990 ;
  assign n26992 = n26988 & n26989 ;
  assign n26993 = ~n26697 & n26988 ;
  assign n26994 = ~n26963 & n26993 ;
  assign n26995 = ~n26992 & ~n26994 ;
  assign n26996 = ~n25605 & ~n26231 ;
  assign n26997 = ~n26179 & n26996 ;
  assign n26998 = ~n26601 & ~n26997 ;
  assign n26999 = ~n26594 & n26998 ;
  assign n27000 = n3402 & n11906 ;
  assign n27001 = ~n11903 & n27000 ;
  assign n27002 = n3402 & ~n11906 ;
  assign n27003 = ~n11392 & n27002 ;
  assign n27004 = ~n11902 & n27003 ;
  assign n27005 = \b[44]  & n3733 ;
  assign n27006 = n3730 & n27005 ;
  assign n27007 = ~\a[24]  & \b[45]  ;
  assign n27008 = n3394 & n27007 ;
  assign n27009 = ~n27006 & ~n27008 ;
  assign n27010 = \b[46]  & n3400 ;
  assign n27011 = \a[24]  & \b[45]  ;
  assign n27012 = n3391 & n27011 ;
  assign n27013 = \a[26]  & ~n27012 ;
  assign n27014 = ~n27010 & n27013 ;
  assign n27015 = n27009 & n27014 ;
  assign n27016 = ~n27004 & n27015 ;
  assign n27017 = ~n27001 & n27016 ;
  assign n27018 = ~n27010 & ~n27012 ;
  assign n27019 = n27009 & n27018 ;
  assign n27020 = ~n27004 & n27019 ;
  assign n27021 = ~n27001 & n27020 ;
  assign n27022 = ~\a[26]  & ~n27021 ;
  assign n27023 = ~n27017 & ~n27022 ;
  assign n27024 = ~n26203 & ~n26206 ;
  assign n27025 = ~n26206 & ~n26588 ;
  assign n27026 = ~n27024 & ~n27025 ;
  assign n27027 = n4249 & ~n10409 ;
  assign n27028 = ~n10407 & n27027 ;
  assign n27029 = \b[43]  & n4247 ;
  assign n27030 = \a[27]  & \b[42]  ;
  assign n27031 = n4238 & n27030 ;
  assign n27032 = ~n27029 & ~n27031 ;
  assign n27033 = \b[41]  & n4647 ;
  assign n27034 = n4644 & n27033 ;
  assign n27035 = ~\a[27]  & \b[42]  ;
  assign n27036 = n4241 & n27035 ;
  assign n27037 = ~n27034 & ~n27036 ;
  assign n27038 = n27032 & n27037 ;
  assign n27039 = ~n27028 & n27038 ;
  assign n27040 = \a[29]  & ~n27039 ;
  assign n27041 = ~\a[29]  & n27039 ;
  assign n27042 = ~n27040 & ~n27041 ;
  assign n27043 = n27026 & n27042 ;
  assign n27044 = ~\a[29]  & ~n27039 ;
  assign n27045 = \a[29]  & n27038 ;
  assign n27046 = ~n27028 & n27045 ;
  assign n27047 = ~n27044 & ~n27046 ;
  assign n27048 = ~n27026 & n27047 ;
  assign n27049 = ~n27043 & ~n27048 ;
  assign n27050 = ~n26577 & ~n26585 ;
  assign n27051 = n26582 & ~n27050 ;
  assign n27052 = n5211 & n9044 ;
  assign n27053 = ~n9041 & n27052 ;
  assign n27054 = ~n8597 & ~n9044 ;
  assign n27055 = n5211 & n27054 ;
  assign n27056 = ~n9040 & n27055 ;
  assign n27057 = \b[40]  & n5209 ;
  assign n27058 = \a[30]  & \b[39]  ;
  assign n27059 = n5200 & n27058 ;
  assign n27060 = ~n27057 & ~n27059 ;
  assign n27061 = \b[38]  & n5595 ;
  assign n27062 = n5592 & n27061 ;
  assign n27063 = ~\a[30]  & \b[39]  ;
  assign n27064 = n5203 & n27063 ;
  assign n27065 = ~n27062 & ~n27064 ;
  assign n27066 = n27060 & n27065 ;
  assign n27067 = ~n27056 & n27066 ;
  assign n27068 = ~n27053 & n27067 ;
  assign n27069 = ~\a[32]  & ~n27068 ;
  assign n27070 = \a[32]  & ~n27059 ;
  assign n27071 = ~n27057 & n27070 ;
  assign n27072 = n27065 & n27071 ;
  assign n27073 = ~n27056 & n27072 ;
  assign n27074 = ~n27053 & n27073 ;
  assign n27075 = ~n27069 & ~n27074 ;
  assign n27076 = ~n27051 & n27075 ;
  assign n27077 = \a[32]  & ~n27068 ;
  assign n27078 = ~\a[32]  & n27068 ;
  assign n27079 = ~n27077 & ~n27078 ;
  assign n27080 = n26582 & n27079 ;
  assign n27081 = ~n27050 & n27080 ;
  assign n27082 = ~n25958 & n26543 ;
  assign n27083 = ~n25962 & n27082 ;
  assign n27084 = n26548 & ~n27083 ;
  assign n27085 = n6309 & ~n7761 ;
  assign n27086 = ~n7759 & n27085 ;
  assign n27087 = \b[35]  & n6778 ;
  assign n27088 = n6775 & n27087 ;
  assign n27089 = ~\a[33]  & \b[36]  ;
  assign n27090 = n6301 & n27089 ;
  assign n27091 = ~n27088 & ~n27090 ;
  assign n27092 = \b[37]  & n6307 ;
  assign n27093 = \a[33]  & \b[36]  ;
  assign n27094 = n6298 & n27093 ;
  assign n27095 = \a[35]  & ~n27094 ;
  assign n27096 = ~n27092 & n27095 ;
  assign n27097 = n27091 & n27096 ;
  assign n27098 = ~n27086 & n27097 ;
  assign n27099 = ~n27092 & ~n27094 ;
  assign n27100 = n27091 & n27099 ;
  assign n27101 = ~n27086 & n27100 ;
  assign n27102 = ~\a[35]  & ~n27101 ;
  assign n27103 = ~n27098 & ~n27102 ;
  assign n27104 = n26469 & ~n26479 ;
  assign n27105 = n26474 & ~n27104 ;
  assign n27106 = ~n26400 & n26432 ;
  assign n27107 = n26405 & ~n27106 ;
  assign n27108 = ~n26256 & n26333 ;
  assign n27109 = n26347 & ~n27108 ;
  assign n27110 = ~n26258 & ~n26328 ;
  assign n27111 = ~n26329 & ~n27110 ;
  assign n27112 = ~n26298 & n26323 ;
  assign n27113 = ~n26295 & ~n27112 ;
  assign n27114 = n685 & n20521 ;
  assign n27115 = ~n682 & n27114 ;
  assign n27116 = n11610 & n20521 ;
  assign n27117 = ~n681 & n27116 ;
  assign n27118 = \b[10]  & n20519 ;
  assign n27119 = \a[60]  & \b[9]  ;
  assign n27120 = n20510 & n27119 ;
  assign n27121 = ~n27118 & ~n27120 ;
  assign n27122 = \b[8]  & n21315 ;
  assign n27123 = n21312 & n27122 ;
  assign n27124 = ~\a[60]  & \b[9]  ;
  assign n27125 = n20513 & n27124 ;
  assign n27126 = ~n27123 & ~n27125 ;
  assign n27127 = n27121 & n27126 ;
  assign n27128 = ~n27117 & n27127 ;
  assign n27129 = ~n27115 & n27128 ;
  assign n27130 = ~n26283 & ~n26287 ;
  assign n27131 = ~n26286 & n27130 ;
  assign n27132 = ~n26284 & ~n27131 ;
  assign n27133 = \b[7]  & n21958 ;
  assign n27134 = \b[6]  & n21957 ;
  assign n27135 = ~n27133 & ~n27134 ;
  assign n27136 = ~\a[62]  & ~n27135 ;
  assign n27137 = n27132 & n27136 ;
  assign n27138 = ~\a[62]  & n27135 ;
  assign n27139 = ~n27132 & n27138 ;
  assign n27140 = ~n27137 & ~n27139 ;
  assign n27141 = ~n27129 & ~n27140 ;
  assign n27142 = \a[62]  & ~n27135 ;
  assign n27143 = n27132 & n27142 ;
  assign n27144 = \a[62]  & n27135 ;
  assign n27145 = ~n27132 & n27144 ;
  assign n27146 = ~n27143 & ~n27145 ;
  assign n27147 = n27127 & ~n27146 ;
  assign n27148 = ~n27117 & n27147 ;
  assign n27149 = ~n27115 & n27148 ;
  assign n27150 = ~n27141 & ~n27149 ;
  assign n27151 = ~\a[62]  & ~n27129 ;
  assign n27152 = n27132 & n27135 ;
  assign n27153 = ~n27132 & ~n27135 ;
  assign n27154 = ~n27152 & ~n27153 ;
  assign n27155 = \a[62]  & n27127 ;
  assign n27156 = ~n27117 & n27155 ;
  assign n27157 = ~n27115 & n27156 ;
  assign n27158 = ~n27154 & ~n27157 ;
  assign n27159 = ~n27151 & n27158 ;
  assign n27160 = n27150 & ~n27159 ;
  assign n27161 = n27113 & n27160 ;
  assign n27162 = ~n27113 & ~n27160 ;
  assign n27163 = ~n27161 & ~n27162 ;
  assign n27164 = ~n948 & n18516 ;
  assign n27165 = ~n908 & n18516 ;
  assign n27166 = ~n912 & n27165 ;
  assign n27167 = ~n27164 & ~n27166 ;
  assign n27168 = ~n951 & ~n27167 ;
  assign n27169 = \b[11]  & n19183 ;
  assign n27170 = n19180 & n27169 ;
  assign n27171 = ~\a[57]  & \b[12]  ;
  assign n27172 = n18508 & n27171 ;
  assign n27173 = ~n27170 & ~n27172 ;
  assign n27174 = \b[13]  & n18514 ;
  assign n27175 = \a[57]  & \b[12]  ;
  assign n27176 = n18505 & n27175 ;
  assign n27177 = \a[59]  & ~n27176 ;
  assign n27178 = ~n27174 & n27177 ;
  assign n27179 = n27173 & n27178 ;
  assign n27180 = ~n27168 & n27179 ;
  assign n27181 = ~n27174 & ~n27176 ;
  assign n27182 = n27173 & n27181 ;
  assign n27183 = ~\a[59]  & ~n27182 ;
  assign n27184 = ~\a[59]  & ~n951 ;
  assign n27185 = ~n27167 & n27184 ;
  assign n27186 = ~n27183 & ~n27185 ;
  assign n27187 = ~n27180 & n27186 ;
  assign n27188 = n27163 & ~n27187 ;
  assign n27189 = ~n27163 & n27187 ;
  assign n27190 = ~n27188 & ~n27189 ;
  assign n27191 = ~n27111 & ~n27190 ;
  assign n27192 = n27111 & n27190 ;
  assign n27193 = ~n27191 & ~n27192 ;
  assign n27194 = n1512 & n16655 ;
  assign n27195 = ~n1509 & n27194 ;
  assign n27196 = n10165 & n16655 ;
  assign n27197 = ~n1508 & n27196 ;
  assign n27198 = \b[14]  & n17308 ;
  assign n27199 = n17305 & n27198 ;
  assign n27200 = ~\a[54]  & \b[15]  ;
  assign n27201 = n16647 & n27200 ;
  assign n27202 = ~n27199 & ~n27201 ;
  assign n27203 = \b[16]  & n16653 ;
  assign n27204 = \a[54]  & \b[15]  ;
  assign n27205 = n16644 & n27204 ;
  assign n27206 = \a[56]  & ~n27205 ;
  assign n27207 = ~n27203 & n27206 ;
  assign n27208 = n27202 & n27207 ;
  assign n27209 = ~n27197 & n27208 ;
  assign n27210 = ~n27195 & n27209 ;
  assign n27211 = ~n27203 & ~n27205 ;
  assign n27212 = n27202 & n27211 ;
  assign n27213 = ~n27197 & n27212 ;
  assign n27214 = ~n27195 & n27213 ;
  assign n27215 = ~\a[56]  & ~n27214 ;
  assign n27216 = ~n27210 & ~n27215 ;
  assign n27217 = ~n27193 & n27216 ;
  assign n27218 = n27193 & ~n27216 ;
  assign n27219 = ~n27217 & ~n27218 ;
  assign n27220 = n27109 & ~n27219 ;
  assign n27221 = ~n27109 & n27219 ;
  assign n27222 = ~n27220 & ~n27221 ;
  assign n27223 = ~n2079 & n14793 ;
  assign n27224 = ~n2077 & n27223 ;
  assign n27225 = \b[17]  & n15517 ;
  assign n27226 = n15514 & n27225 ;
  assign n27227 = ~\a[51]  & \b[18]  ;
  assign n27228 = n14785 & n27227 ;
  assign n27229 = ~n27226 & ~n27228 ;
  assign n27230 = \b[19]  & n14791 ;
  assign n27231 = \a[51]  & \b[18]  ;
  assign n27232 = n14782 & n27231 ;
  assign n27233 = \a[53]  & ~n27232 ;
  assign n27234 = ~n27230 & n27233 ;
  assign n27235 = n27229 & n27234 ;
  assign n27236 = ~n27224 & n27235 ;
  assign n27237 = ~n27230 & ~n27232 ;
  assign n27238 = n27229 & n27237 ;
  assign n27239 = ~n27224 & n27238 ;
  assign n27240 = ~\a[53]  & ~n27239 ;
  assign n27241 = ~n27236 & ~n27240 ;
  assign n27242 = n27222 & ~n27241 ;
  assign n27243 = ~n27222 & n27241 ;
  assign n27244 = ~n27242 & ~n27243 ;
  assign n27245 = ~n26373 & ~n26378 ;
  assign n27246 = ~n26375 & ~n27245 ;
  assign n27247 = n2768 & n13125 ;
  assign n27248 = ~n2765 & n27247 ;
  assign n27249 = ~n2768 & n13125 ;
  assign n27250 = ~n2518 & n27249 ;
  assign n27251 = ~n2764 & n27250 ;
  assign n27252 = \b[20]  & n13794 ;
  assign n27253 = n13792 & n27252 ;
  assign n27254 = ~\a[48]  & \b[21]  ;
  assign n27255 = n13117 & n27254 ;
  assign n27256 = ~n27253 & ~n27255 ;
  assign n27257 = \b[22]  & n13123 ;
  assign n27258 = \a[48]  & \b[21]  ;
  assign n27259 = n13786 & n27258 ;
  assign n27260 = \a[50]  & ~n27259 ;
  assign n27261 = ~n27257 & n27260 ;
  assign n27262 = n27256 & n27261 ;
  assign n27263 = ~n27251 & n27262 ;
  assign n27264 = ~n27248 & n27263 ;
  assign n27265 = ~n27257 & ~n27259 ;
  assign n27266 = n27256 & n27265 ;
  assign n27267 = ~n27251 & n27266 ;
  assign n27268 = ~n27248 & n27267 ;
  assign n27269 = ~\a[50]  & ~n27268 ;
  assign n27270 = ~n27264 & ~n27269 ;
  assign n27271 = ~n27246 & n27270 ;
  assign n27272 = ~n27244 & n27271 ;
  assign n27273 = n27246 & n27270 ;
  assign n27274 = n27244 & n27273 ;
  assign n27275 = ~n27272 & ~n27274 ;
  assign n27276 = n27246 & ~n27270 ;
  assign n27277 = ~n27244 & n27276 ;
  assign n27278 = ~n27246 & ~n27270 ;
  assign n27279 = n27244 & n27278 ;
  assign n27280 = ~n27277 & ~n27279 ;
  assign n27281 = n27275 & n27280 ;
  assign n27282 = ~n27107 & ~n27281 ;
  assign n27283 = n27107 & n27281 ;
  assign n27284 = ~n27282 & ~n27283 ;
  assign n27285 = ~n3567 & n11572 ;
  assign n27286 = ~n3565 & n27285 ;
  assign n27287 = \b[23]  & n12159 ;
  assign n27288 = n12156 & n27287 ;
  assign n27289 = ~\a[45]  & \b[24]  ;
  assign n27290 = n11564 & n27289 ;
  assign n27291 = ~n27288 & ~n27290 ;
  assign n27292 = \b[25]  & n11570 ;
  assign n27293 = \a[45]  & \b[24]  ;
  assign n27294 = n11561 & n27293 ;
  assign n27295 = \a[47]  & ~n27294 ;
  assign n27296 = ~n27292 & n27295 ;
  assign n27297 = n27291 & n27296 ;
  assign n27298 = ~n27286 & n27297 ;
  assign n27299 = ~n27292 & ~n27294 ;
  assign n27300 = n27291 & n27299 ;
  assign n27301 = ~n27286 & n27300 ;
  assign n27302 = ~\a[47]  & ~n27301 ;
  assign n27303 = ~n27298 & ~n27302 ;
  assign n27304 = n27284 & ~n27303 ;
  assign n27305 = ~n27284 & n27303 ;
  assign n27306 = ~n27304 & ~n27305 ;
  assign n27307 = n26437 & ~n26447 ;
  assign n27308 = n26442 & ~n27307 ;
  assign n27309 = n4456 & n10082 ;
  assign n27310 = ~n18723 & n27309 ;
  assign n27311 = ~n4456 & n10082 ;
  assign n27312 = ~n4143 & n27311 ;
  assign n27313 = ~n4452 & n27312 ;
  assign n27314 = \b[26]  & n10681 ;
  assign n27315 = n10678 & n27314 ;
  assign n27316 = ~\a[42]  & \b[27]  ;
  assign n27317 = n10074 & n27316 ;
  assign n27318 = ~n27315 & ~n27317 ;
  assign n27319 = \b[28]  & n10080 ;
  assign n27320 = \a[42]  & \b[27]  ;
  assign n27321 = n10071 & n27320 ;
  assign n27322 = \a[44]  & ~n27321 ;
  assign n27323 = ~n27319 & n27322 ;
  assign n27324 = n27318 & n27323 ;
  assign n27325 = ~n27313 & n27324 ;
  assign n27326 = ~n27310 & n27325 ;
  assign n27327 = ~n27319 & ~n27321 ;
  assign n27328 = n27318 & n27327 ;
  assign n27329 = ~n27313 & n27328 ;
  assign n27330 = ~n27310 & n27329 ;
  assign n27331 = ~\a[44]  & ~n27330 ;
  assign n27332 = ~n27326 & ~n27331 ;
  assign n27333 = ~n27308 & n27332 ;
  assign n27334 = ~n27306 & n27333 ;
  assign n27335 = n27308 & n27332 ;
  assign n27336 = n27306 & n27335 ;
  assign n27337 = ~n27334 & ~n27336 ;
  assign n27338 = n27308 & ~n27332 ;
  assign n27339 = ~n27306 & n27338 ;
  assign n27340 = ~n27308 & ~n27332 ;
  assign n27341 = n27306 & n27340 ;
  assign n27342 = ~n27339 & ~n27341 ;
  assign n27343 = n27337 & n27342 ;
  assign n27344 = ~n27105 & ~n27343 ;
  assign n27345 = n27105 & n27343 ;
  assign n27346 = ~n27344 & ~n27345 ;
  assign n27347 = ~n5459 & n8759 ;
  assign n27348 = ~n5104 & n8759 ;
  assign n27349 = ~n5455 & n27348 ;
  assign n27350 = ~n27347 & ~n27349 ;
  assign n27351 = ~n5462 & ~n27350 ;
  assign n27352 = \b[29]  & n9301 ;
  assign n27353 = n9298 & n27352 ;
  assign n27354 = ~\a[39]  & \b[30]  ;
  assign n27355 = n8751 & n27354 ;
  assign n27356 = ~n27353 & ~n27355 ;
  assign n27357 = \b[31]  & n8757 ;
  assign n27358 = \a[39]  & \b[30]  ;
  assign n27359 = n8748 & n27358 ;
  assign n27360 = \a[41]  & ~n27359 ;
  assign n27361 = ~n27357 & n27360 ;
  assign n27362 = n27356 & n27361 ;
  assign n27363 = ~n27351 & n27362 ;
  assign n27364 = ~n27357 & ~n27359 ;
  assign n27365 = n27356 & n27364 ;
  assign n27366 = ~\a[41]  & ~n27365 ;
  assign n27367 = ~\a[41]  & ~n5462 ;
  assign n27368 = ~n27350 & n27367 ;
  assign n27369 = ~n27366 & ~n27368 ;
  assign n27370 = ~n27363 & n27369 ;
  assign n27371 = ~n27346 & n27370 ;
  assign n27372 = n27346 & ~n27370 ;
  assign n27373 = ~n27371 & ~n27372 ;
  assign n27374 = ~n6565 & ~n7098 ;
  assign n27375 = ~n7531 & n27374 ;
  assign n27376 = n6562 & n27375 ;
  assign n27377 = n6565 & ~n7098 ;
  assign n27378 = ~n7531 & n27377 ;
  assign n27379 = ~n6562 & n27378 ;
  assign n27380 = ~n27376 & ~n27379 ;
  assign n27381 = \b[32]  & n7973 ;
  assign n27382 = n7970 & n27381 ;
  assign n27383 = ~\a[36]  & \b[33]  ;
  assign n27384 = n7526 & n27383 ;
  assign n27385 = ~n27382 & ~n27384 ;
  assign n27386 = \b[34]  & n7532 ;
  assign n27387 = \a[36]  & \b[33]  ;
  assign n27388 = n17801 & n27387 ;
  assign n27389 = \a[38]  & ~n27388 ;
  assign n27390 = ~n27386 & n27389 ;
  assign n27391 = n27385 & n27390 ;
  assign n27392 = n27380 & n27391 ;
  assign n27393 = ~n27386 & ~n27388 ;
  assign n27394 = n27385 & n27393 ;
  assign n27395 = n27380 & n27394 ;
  assign n27396 = ~\a[38]  & ~n27395 ;
  assign n27397 = ~n27392 & ~n27396 ;
  assign n27398 = ~n26508 & n26538 ;
  assign n27399 = ~n26507 & ~n27398 ;
  assign n27400 = ~n27397 & ~n27399 ;
  assign n27401 = n27373 & n27400 ;
  assign n27402 = ~n27397 & n27399 ;
  assign n27403 = ~n27373 & n27402 ;
  assign n27404 = ~n27401 & ~n27403 ;
  assign n27405 = n27397 & ~n27399 ;
  assign n27406 = ~n27373 & n27405 ;
  assign n27407 = n27397 & n27399 ;
  assign n27408 = n27373 & n27407 ;
  assign n27409 = ~n27406 & ~n27408 ;
  assign n27410 = n27404 & n27409 ;
  assign n27411 = n27103 & ~n27410 ;
  assign n27412 = n27084 & n27411 ;
  assign n27413 = n27103 & n27410 ;
  assign n27414 = ~n27084 & n27413 ;
  assign n27415 = ~n27412 & ~n27414 ;
  assign n27416 = ~n27103 & ~n27410 ;
  assign n27417 = ~n27084 & n27416 ;
  assign n27418 = ~n27103 & n27410 ;
  assign n27419 = n27084 & n27418 ;
  assign n27420 = ~n27417 & ~n27419 ;
  assign n27421 = n27415 & n27420 ;
  assign n27422 = ~n27081 & ~n27421 ;
  assign n27423 = ~n27076 & n27422 ;
  assign n27424 = n27081 & n27421 ;
  assign n27425 = n27075 & n27421 ;
  assign n27426 = ~n27051 & n27425 ;
  assign n27427 = ~n27424 & ~n27426 ;
  assign n27428 = ~n27423 & n27427 ;
  assign n27429 = n27049 & n27428 ;
  assign n27430 = ~n27049 & ~n27428 ;
  assign n27431 = ~n27429 & ~n27430 ;
  assign n27432 = n27023 & n27431 ;
  assign n27433 = ~n26999 & n27432 ;
  assign n27434 = ~n27023 & n27431 ;
  assign n27435 = n26999 & n27434 ;
  assign n27436 = ~n27433 & ~n27435 ;
  assign n27437 = n27023 & ~n27431 ;
  assign n27438 = n26999 & n27437 ;
  assign n27439 = ~n27023 & ~n27431 ;
  assign n27440 = ~n26999 & n27439 ;
  assign n27441 = ~n27438 & ~n27440 ;
  assign n27442 = n27436 & n27441 ;
  assign n27443 = ~n26614 & n26689 ;
  assign n27444 = ~n26685 & ~n27443 ;
  assign n27445 = n2622 & ~n13524 ;
  assign n27446 = ~n13522 & n27445 ;
  assign n27447 = \b[49]  & n2620 ;
  assign n27448 = \a[21]  & \b[48]  ;
  assign n27449 = n20849 & n27448 ;
  assign n27450 = ~n27447 & ~n27449 ;
  assign n27451 = \b[47]  & n2912 ;
  assign n27452 = n2909 & n27451 ;
  assign n27453 = ~\a[21]  & \b[48]  ;
  assign n27454 = n2614 & n27453 ;
  assign n27455 = ~n27452 & ~n27454 ;
  assign n27456 = n27450 & n27455 ;
  assign n27457 = ~n27446 & n27456 ;
  assign n27458 = \a[23]  & ~n27457 ;
  assign n27459 = ~\a[23]  & n27457 ;
  assign n27460 = ~n27458 & ~n27459 ;
  assign n27461 = n27444 & n27460 ;
  assign n27462 = ~\a[23]  & ~n27457 ;
  assign n27463 = \a[23]  & n27456 ;
  assign n27464 = ~n27446 & n27463 ;
  assign n27465 = ~n27462 & ~n27464 ;
  assign n27466 = ~n27444 & n27465 ;
  assign n27467 = ~n27461 & ~n27466 ;
  assign n27468 = n27442 & n27467 ;
  assign n27469 = ~n27442 & ~n27467 ;
  assign n27470 = ~n27468 & ~n27469 ;
  assign n27471 = n26995 & n27470 ;
  assign n27472 = ~n26991 & n27471 ;
  assign n27473 = ~n26995 & ~n27470 ;
  assign n27474 = ~n26964 & ~n26989 ;
  assign n27475 = ~n26988 & ~n27470 ;
  assign n27476 = n27474 & n27475 ;
  assign n27477 = ~n27473 & ~n27476 ;
  assign n27478 = ~n27472 & n27477 ;
  assign n27479 = ~n26962 & n27478 ;
  assign n27480 = ~n26958 & n27479 ;
  assign n27481 = n26962 & ~n27478 ;
  assign n27482 = ~n26951 & ~n27478 ;
  assign n27483 = ~n26957 & n27482 ;
  assign n27484 = ~n27481 & ~n27483 ;
  assign n27485 = ~n27480 & n27484 ;
  assign n27486 = n26937 & n27485 ;
  assign n27487 = ~n26930 & n27486 ;
  assign n27488 = ~n26937 & ~n27485 ;
  assign n27489 = ~n26905 & ~n27485 ;
  assign n27490 = n26722 & n27489 ;
  assign n27491 = n26928 & n27490 ;
  assign n27492 = ~n27488 & ~n27491 ;
  assign n27493 = ~n27487 & n27492 ;
  assign n27494 = n26904 & n27493 ;
  assign n27495 = ~n26904 & ~n27493 ;
  assign n27496 = ~n27494 & ~n27495 ;
  assign n27497 = n26879 & n27496 ;
  assign n27498 = ~n26879 & ~n27496 ;
  assign n27499 = ~n27497 & ~n27498 ;
  assign n27500 = n26852 & n27499 ;
  assign n27501 = ~n26852 & ~n27499 ;
  assign n27502 = ~n27500 & ~n27501 ;
  assign n27503 = ~n26848 & n27502 ;
  assign n27504 = ~n26840 & ~n27502 ;
  assign n27505 = ~n26844 & n27504 ;
  assign n27506 = ~n27503 & ~n27505 ;
  assign n27507 = ~n26840 & ~n27500 ;
  assign n27508 = ~n26844 & n27507 ;
  assign n27509 = ~n26903 & ~n27493 ;
  assign n27510 = n26899 & ~n26903 ;
  assign n27511 = ~n27509 & ~n27510 ;
  assign n27512 = \b[63]  & n430 ;
  assign n27513 = ~n21694 & n27512 ;
  assign n27514 = ~n23171 & n27513 ;
  assign n27515 = \a[5]  & \a[7]  ;
  assign n27516 = \a[6]  & ~\a[8]  ;
  assign n27517 = n27515 & n27516 ;
  assign n27518 = ~\a[5]  & ~\a[7]  ;
  assign n27519 = ~\a[6]  & \a[8]  ;
  assign n27520 = n27518 & n27519 ;
  assign n27521 = ~n27517 & ~n27520 ;
  assign n27522 = \b[63]  & ~n27521 ;
  assign n27523 = \a[8]  & ~n27522 ;
  assign n27524 = ~n27514 & n27523 ;
  assign n27525 = ~n27514 & ~n27522 ;
  assign n27526 = ~\a[8]  & ~n27525 ;
  assign n27527 = ~n27524 & ~n27526 ;
  assign n27528 = ~n27511 & n27527 ;
  assign n27529 = ~n26962 & ~n27478 ;
  assign n27530 = n26959 & n26960 ;
  assign n27531 = n26147 & n26960 ;
  assign n27532 = ~n27530 & ~n27531 ;
  assign n27533 = ~n27529 & n27532 ;
  assign n27534 = n999 & ~n19550 ;
  assign n27535 = ~n19548 & n27534 ;
  assign n27536 = \b[57]  & n1182 ;
  assign n27537 = n1179 & n27536 ;
  assign n27538 = \b[59]  & n997 ;
  assign n27539 = \a[11]  & \b[58]  ;
  assign n27540 = n1180 & n27539 ;
  assign n27541 = ~\a[12]  & \b[58]  ;
  assign n27542 = n7674 & n27541 ;
  assign n27543 = ~n27540 & ~n27542 ;
  assign n27544 = ~n27538 & n27543 ;
  assign n27545 = ~n27537 & n27544 ;
  assign n27546 = ~n27535 & n27545 ;
  assign n27547 = \a[14]  & ~n27546 ;
  assign n27548 = ~\a[14]  & n27546 ;
  assign n27549 = ~n27547 & ~n27548 ;
  assign n27550 = n27533 & n27549 ;
  assign n27551 = ~\a[14]  & ~n27546 ;
  assign n27552 = \a[14]  & n27545 ;
  assign n27553 = ~n27535 & n27552 ;
  assign n27554 = ~n27551 & ~n27553 ;
  assign n27555 = ~n27533 & n27554 ;
  assign n27556 = ~n27550 & ~n27555 ;
  assign n27557 = n1467 & n17647 ;
  assign n27558 = ~n17644 & n27557 ;
  assign n27559 = n1467 & ~n17647 ;
  assign n27560 = ~n16441 & n27559 ;
  assign n27561 = ~n17643 & n27560 ;
  assign n27562 = \b[56]  & n1465 ;
  assign n27563 = \a[15]  & \b[55]  ;
  assign n27564 = n1456 & n27563 ;
  assign n27565 = ~n27562 & ~n27564 ;
  assign n27566 = \b[54]  & n1652 ;
  assign n27567 = n1649 & n27566 ;
  assign n27568 = ~\a[15]  & \b[55]  ;
  assign n27569 = n1459 & n27568 ;
  assign n27570 = ~n27567 & ~n27569 ;
  assign n27571 = n27565 & n27570 ;
  assign n27572 = ~n27561 & n27571 ;
  assign n27573 = ~n27558 & n27572 ;
  assign n27574 = ~\a[17]  & ~n27573 ;
  assign n27575 = \a[17]  & n27571 ;
  assign n27576 = ~n27561 & n27575 ;
  assign n27577 = ~n27558 & n27576 ;
  assign n27578 = ~n26995 & ~n27577 ;
  assign n27579 = ~n27470 & ~n27577 ;
  assign n27580 = ~n26991 & n27579 ;
  assign n27581 = ~n27578 & ~n27580 ;
  assign n27582 = ~n27574 & ~n27581 ;
  assign n27583 = ~n26991 & ~n27470 ;
  assign n27584 = ~n27574 & ~n27577 ;
  assign n27585 = n26995 & ~n27584 ;
  assign n27586 = ~n27583 & n27585 ;
  assign n27587 = ~n26999 & ~n27023 ;
  assign n27588 = n2622 & n14052 ;
  assign n27589 = ~n14049 & n27588 ;
  assign n27590 = n2622 & ~n14052 ;
  assign n27591 = ~n13519 & n27590 ;
  assign n27592 = ~n14048 & n27591 ;
  assign n27593 = \b[50]  & n2620 ;
  assign n27594 = \a[21]  & \b[49]  ;
  assign n27595 = n20849 & n27594 ;
  assign n27596 = ~n27593 & ~n27595 ;
  assign n27597 = \b[48]  & n2912 ;
  assign n27598 = n2909 & n27597 ;
  assign n27599 = ~\a[21]  & \b[49]  ;
  assign n27600 = n2614 & n27599 ;
  assign n27601 = ~n27598 & ~n27600 ;
  assign n27602 = n27596 & n27601 ;
  assign n27603 = ~n27592 & n27602 ;
  assign n27604 = ~n27589 & n27603 ;
  assign n27605 = ~\a[23]  & ~n27604 ;
  assign n27606 = \a[23]  & ~n27595 ;
  assign n27607 = ~n27593 & n27606 ;
  assign n27608 = n27601 & n27607 ;
  assign n27609 = ~n27592 & n27608 ;
  assign n27610 = ~n27589 & n27609 ;
  assign n27611 = ~n27605 & ~n27610 ;
  assign n27612 = ~n27587 & n27611 ;
  assign n27613 = n27436 & n27612 ;
  assign n27614 = n27436 & ~n27587 ;
  assign n27615 = \a[23]  & ~n27604 ;
  assign n27616 = ~\a[23]  & n27604 ;
  assign n27617 = ~n27615 & ~n27616 ;
  assign n27618 = ~n27614 & n27617 ;
  assign n27619 = ~n27613 & ~n27618 ;
  assign n27620 = ~n27043 & ~n27428 ;
  assign n27621 = ~n27043 & n27048 ;
  assign n27622 = ~n27620 & ~n27621 ;
  assign n27623 = n3402 & ~n12438 ;
  assign n27624 = ~n12436 & n27623 ;
  assign n27625 = \b[47]  & n3400 ;
  assign n27626 = \a[23]  & ~\a[25]  ;
  assign n27627 = \a[24]  & \b[46]  ;
  assign n27628 = n27626 & n27627 ;
  assign n27629 = ~n27625 & ~n27628 ;
  assign n27630 = \b[45]  & n3733 ;
  assign n27631 = n3730 & n27630 ;
  assign n27632 = ~\a[24]  & \b[46]  ;
  assign n27633 = n3394 & n27632 ;
  assign n27634 = ~n27631 & ~n27633 ;
  assign n27635 = n27629 & n27634 ;
  assign n27636 = ~n27624 & n27635 ;
  assign n27637 = \a[26]  & ~n27636 ;
  assign n27638 = ~\a[26]  & n27636 ;
  assign n27639 = ~n27637 & ~n27638 ;
  assign n27640 = n27622 & n27639 ;
  assign n27641 = ~\a[26]  & ~n27636 ;
  assign n27642 = \a[26]  & n27635 ;
  assign n27643 = ~n27624 & n27642 ;
  assign n27644 = ~n27641 & ~n27643 ;
  assign n27645 = ~n27622 & n27644 ;
  assign n27646 = ~n27640 & ~n27645 ;
  assign n27647 = n27084 & n27410 ;
  assign n27648 = n26548 & ~n27103 ;
  assign n27649 = ~n27083 & n27648 ;
  assign n27650 = ~n27418 & ~n27649 ;
  assign n27651 = ~n27647 & n27650 ;
  assign n27652 = n5211 & ~n9482 ;
  assign n27653 = ~n9480 & n27652 ;
  assign n27654 = \b[41]  & n5209 ;
  assign n27655 = \a[30]  & \b[40]  ;
  assign n27656 = n5200 & n27655 ;
  assign n27657 = ~n27654 & ~n27656 ;
  assign n27658 = \b[39]  & n5595 ;
  assign n27659 = n5592 & n27658 ;
  assign n27660 = ~\a[30]  & \b[40]  ;
  assign n27661 = n5203 & n27660 ;
  assign n27662 = ~n27659 & ~n27661 ;
  assign n27663 = n27657 & n27662 ;
  assign n27664 = ~n27653 & n27663 ;
  assign n27665 = ~\a[32]  & ~n27664 ;
  assign n27666 = \a[32]  & ~n27656 ;
  assign n27667 = ~n27654 & n27666 ;
  assign n27668 = n27662 & n27667 ;
  assign n27669 = ~n27653 & n27668 ;
  assign n27670 = ~n27665 & ~n27669 ;
  assign n27671 = n27651 & n27670 ;
  assign n27672 = \a[32]  & ~n27664 ;
  assign n27673 = ~\a[32]  & n27664 ;
  assign n27674 = ~n27672 & ~n27673 ;
  assign n27675 = ~n27651 & n27674 ;
  assign n27676 = ~n27671 & ~n27675 ;
  assign n27677 = n27373 & n27399 ;
  assign n27678 = n27404 & ~n27677 ;
  assign n27679 = ~n3022 & n13125 ;
  assign n27680 = ~n3020 & n27679 ;
  assign n27681 = \b[21]  & n13794 ;
  assign n27682 = n13792 & n27681 ;
  assign n27683 = ~\a[48]  & \b[22]  ;
  assign n27684 = n13117 & n27683 ;
  assign n27685 = ~n27682 & ~n27684 ;
  assign n27686 = \b[23]  & n13123 ;
  assign n27687 = \a[48]  & \b[22]  ;
  assign n27688 = n13786 & n27687 ;
  assign n27689 = \a[50]  & ~n27688 ;
  assign n27690 = ~n27686 & n27689 ;
  assign n27691 = n27685 & n27690 ;
  assign n27692 = ~n27680 & n27691 ;
  assign n27693 = ~n27686 & ~n27688 ;
  assign n27694 = n27685 & n27693 ;
  assign n27695 = ~n27680 & n27694 ;
  assign n27696 = ~\a[50]  & ~n27695 ;
  assign n27697 = ~n27692 & ~n27696 ;
  assign n27698 = n1087 & n18516 ;
  assign n27699 = ~n1084 & n27698 ;
  assign n27700 = n18516 & n21340 ;
  assign n27701 = ~n1083 & n27700 ;
  assign n27702 = \b[12]  & n19183 ;
  assign n27703 = n19180 & n27702 ;
  assign n27704 = ~\a[57]  & \b[13]  ;
  assign n27705 = n18508 & n27704 ;
  assign n27706 = ~n27703 & ~n27705 ;
  assign n27707 = \b[14]  & n18514 ;
  assign n27708 = \a[57]  & \b[13]  ;
  assign n27709 = n18505 & n27708 ;
  assign n27710 = \a[59]  & ~n27709 ;
  assign n27711 = ~n27707 & n27710 ;
  assign n27712 = n27706 & n27711 ;
  assign n27713 = ~n27701 & n27712 ;
  assign n27714 = ~n27699 & n27713 ;
  assign n27715 = ~n27707 & ~n27709 ;
  assign n27716 = n27706 & n27715 ;
  assign n27717 = ~n27701 & n27716 ;
  assign n27718 = ~n27699 & n27717 ;
  assign n27719 = ~\a[59]  & ~n27718 ;
  assign n27720 = ~n27714 & ~n27719 ;
  assign n27721 = ~n725 & n20521 ;
  assign n27722 = ~n684 & n20521 ;
  assign n27723 = ~n721 & n27722 ;
  assign n27724 = ~n27721 & ~n27723 ;
  assign n27725 = ~n728 & ~n27724 ;
  assign n27726 = \b[9]  & n21315 ;
  assign n27727 = n21312 & n27726 ;
  assign n27728 = ~\a[60]  & \b[10]  ;
  assign n27729 = n20513 & n27728 ;
  assign n27730 = ~n27727 & ~n27729 ;
  assign n27731 = \b[11]  & n20519 ;
  assign n27732 = \a[60]  & \b[10]  ;
  assign n27733 = n20510 & n27732 ;
  assign n27734 = \a[62]  & ~n27733 ;
  assign n27735 = ~n27731 & n27734 ;
  assign n27736 = n27730 & n27735 ;
  assign n27737 = ~n27725 & n27736 ;
  assign n27738 = ~n27731 & ~n27733 ;
  assign n27739 = n27730 & n27738 ;
  assign n27740 = ~\a[62]  & ~n27739 ;
  assign n27741 = ~\a[62]  & ~n728 ;
  assign n27742 = ~n27724 & n27741 ;
  assign n27743 = ~n27740 & ~n27742 ;
  assign n27744 = ~n27737 & n27743 ;
  assign n27745 = ~n27149 & ~n27152 ;
  assign n27746 = ~n27141 & n27745 ;
  assign n27747 = \b[8]  & n21958 ;
  assign n27748 = \b[7]  & n21957 ;
  assign n27749 = ~n27747 & ~n27748 ;
  assign n27750 = n27135 & ~n27749 ;
  assign n27751 = ~n27135 & n27749 ;
  assign n27752 = ~n27750 & ~n27751 ;
  assign n27753 = n27746 & n27752 ;
  assign n27754 = ~n27746 & ~n27752 ;
  assign n27755 = ~n27753 & ~n27754 ;
  assign n27756 = ~n27744 & ~n27755 ;
  assign n27757 = n27744 & n27755 ;
  assign n27758 = ~n27756 & ~n27757 ;
  assign n27759 = n27720 & n27758 ;
  assign n27760 = ~n27720 & ~n27758 ;
  assign n27761 = ~n27759 & ~n27760 ;
  assign n27762 = ~n27161 & n27187 ;
  assign n27763 = ~n27162 & ~n27762 ;
  assign n27764 = n27761 & ~n27763 ;
  assign n27765 = ~n27761 & n27763 ;
  assign n27766 = ~n27764 & ~n27765 ;
  assign n27767 = ~n1691 & n16655 ;
  assign n27768 = ~n1511 & n16655 ;
  assign n27769 = ~n1515 & n27768 ;
  assign n27770 = ~n27767 & ~n27769 ;
  assign n27771 = ~n1694 & ~n27770 ;
  assign n27772 = \b[15]  & n17308 ;
  assign n27773 = n17305 & n27772 ;
  assign n27774 = ~\a[54]  & \b[16]  ;
  assign n27775 = n16647 & n27774 ;
  assign n27776 = ~n27773 & ~n27775 ;
  assign n27777 = \b[17]  & n16653 ;
  assign n27778 = \a[54]  & \b[16]  ;
  assign n27779 = n16644 & n27778 ;
  assign n27780 = \a[56]  & ~n27779 ;
  assign n27781 = ~n27777 & n27780 ;
  assign n27782 = n27776 & n27781 ;
  assign n27783 = ~n27771 & n27782 ;
  assign n27784 = ~n27777 & ~n27779 ;
  assign n27785 = n27776 & n27784 ;
  assign n27786 = ~\a[56]  & ~n27785 ;
  assign n27787 = ~\a[56]  & ~n1694 ;
  assign n27788 = ~n27770 & n27787 ;
  assign n27789 = ~n27786 & ~n27788 ;
  assign n27790 = ~n27783 & n27789 ;
  assign n27791 = n27766 & ~n27790 ;
  assign n27792 = ~n27766 & n27790 ;
  assign n27793 = ~n27791 & ~n27792 ;
  assign n27794 = ~n27192 & n27216 ;
  assign n27795 = ~n27191 & ~n27794 ;
  assign n27796 = ~n27793 & ~n27795 ;
  assign n27797 = n27793 & n27795 ;
  assign n27798 = ~n27796 & ~n27797 ;
  assign n27799 = n2293 & n14793 ;
  assign n27800 = ~n19247 & n27799 ;
  assign n27801 = ~n2293 & n14793 ;
  assign n27802 = ~n2074 & n27801 ;
  assign n27803 = ~n2289 & n27802 ;
  assign n27804 = \b[18]  & n15517 ;
  assign n27805 = n15514 & n27804 ;
  assign n27806 = ~\a[51]  & \b[19]  ;
  assign n27807 = n14785 & n27806 ;
  assign n27808 = ~n27805 & ~n27807 ;
  assign n27809 = \b[20]  & n14791 ;
  assign n27810 = \a[51]  & \b[19]  ;
  assign n27811 = n14782 & n27810 ;
  assign n27812 = \a[53]  & ~n27811 ;
  assign n27813 = ~n27809 & n27812 ;
  assign n27814 = n27808 & n27813 ;
  assign n27815 = ~n27803 & n27814 ;
  assign n27816 = ~n27800 & n27815 ;
  assign n27817 = ~n27809 & ~n27811 ;
  assign n27818 = n27808 & n27817 ;
  assign n27819 = ~n27803 & n27818 ;
  assign n27820 = ~n27800 & n27819 ;
  assign n27821 = ~\a[53]  & ~n27820 ;
  assign n27822 = ~n27816 & ~n27821 ;
  assign n27823 = ~n27798 & n27822 ;
  assign n27824 = n27798 & ~n27822 ;
  assign n27825 = ~n27823 & ~n27824 ;
  assign n27826 = ~n27221 & n27241 ;
  assign n27827 = ~n27220 & ~n27826 ;
  assign n27828 = n27825 & n27827 ;
  assign n27829 = ~n27825 & ~n27827 ;
  assign n27830 = ~n27828 & ~n27829 ;
  assign n27831 = n27697 & n27830 ;
  assign n27832 = ~n27697 & ~n27830 ;
  assign n27833 = ~n27831 & ~n27832 ;
  assign n27834 = ~n27244 & ~n27246 ;
  assign n27835 = n27244 & n27246 ;
  assign n27836 = n27270 & ~n27835 ;
  assign n27837 = ~n27834 & ~n27836 ;
  assign n27838 = n3604 & n11572 ;
  assign n27839 = ~n19292 & n27838 ;
  assign n27840 = ~n3604 & n11572 ;
  assign n27841 = ~n3562 & n27840 ;
  assign n27842 = ~n3600 & n27841 ;
  assign n27843 = \b[24]  & n12159 ;
  assign n27844 = n12156 & n27843 ;
  assign n27845 = ~\a[45]  & \b[25]  ;
  assign n27846 = n11564 & n27845 ;
  assign n27847 = ~n27844 & ~n27846 ;
  assign n27848 = \b[26]  & n11570 ;
  assign n27849 = \a[45]  & \b[25]  ;
  assign n27850 = n11561 & n27849 ;
  assign n27851 = \a[47]  & ~n27850 ;
  assign n27852 = ~n27848 & n27851 ;
  assign n27853 = n27847 & n27852 ;
  assign n27854 = ~n27842 & n27853 ;
  assign n27855 = ~n27839 & n27854 ;
  assign n27856 = ~n27848 & ~n27850 ;
  assign n27857 = n27847 & n27856 ;
  assign n27858 = ~n27842 & n27857 ;
  assign n27859 = ~n27839 & n27858 ;
  assign n27860 = ~\a[47]  & ~n27859 ;
  assign n27861 = ~n27855 & ~n27860 ;
  assign n27862 = ~n27837 & ~n27861 ;
  assign n27863 = ~n27833 & n27862 ;
  assign n27864 = n27837 & ~n27861 ;
  assign n27865 = n27833 & n27864 ;
  assign n27866 = ~n27863 & ~n27865 ;
  assign n27867 = ~n27837 & n27861 ;
  assign n27868 = n27833 & n27867 ;
  assign n27869 = n27837 & n27861 ;
  assign n27870 = ~n27833 & n27869 ;
  assign n27871 = ~n27868 & ~n27870 ;
  assign n27872 = n27866 & n27871 ;
  assign n27873 = ~n27283 & n27303 ;
  assign n27874 = ~n27282 & ~n27873 ;
  assign n27875 = ~n4502 & n10082 ;
  assign n27876 = ~n4500 & n27875 ;
  assign n27877 = \b[29]  & n10080 ;
  assign n27878 = \a[41]  & \b[28]  ;
  assign n27879 = n10679 & n27878 ;
  assign n27880 = ~\a[42]  & \b[28]  ;
  assign n27881 = n10074 & n27880 ;
  assign n27882 = ~n27879 & ~n27881 ;
  assign n27883 = ~n27877 & n27882 ;
  assign n27884 = \b[27]  & n10681 ;
  assign n27885 = n10678 & n27884 ;
  assign n27886 = \a[44]  & ~n27885 ;
  assign n27887 = n27883 & n27886 ;
  assign n27888 = ~n27876 & n27887 ;
  assign n27889 = n27883 & ~n27885 ;
  assign n27890 = ~n27876 & n27889 ;
  assign n27891 = ~\a[44]  & ~n27890 ;
  assign n27892 = ~n27888 & ~n27891 ;
  assign n27893 = ~n27874 & n27892 ;
  assign n27894 = ~n27872 & n27893 ;
  assign n27895 = n27874 & n27892 ;
  assign n27896 = n27872 & n27895 ;
  assign n27897 = ~n27894 & ~n27896 ;
  assign n27898 = ~n27874 & ~n27892 ;
  assign n27899 = n27872 & n27898 ;
  assign n27900 = n27874 & ~n27892 ;
  assign n27901 = ~n27872 & n27900 ;
  assign n27902 = ~n27899 & ~n27901 ;
  assign n27903 = n27897 & n27902 ;
  assign n27904 = ~n27306 & ~n27308 ;
  assign n27905 = n27306 & n27308 ;
  assign n27906 = n27332 & ~n27905 ;
  assign n27907 = ~n27904 & ~n27906 ;
  assign n27908 = ~n27903 & ~n27907 ;
  assign n27909 = n27903 & n27907 ;
  assign n27910 = ~n27908 & ~n27909 ;
  assign n27911 = n5810 & n8759 ;
  assign n27912 = ~n5807 & n27911 ;
  assign n27913 = ~n5810 & n8759 ;
  assign n27914 = ~n5457 & n27913 ;
  assign n27915 = ~n5806 & n27914 ;
  assign n27916 = \b[30]  & n9301 ;
  assign n27917 = n9298 & n27916 ;
  assign n27918 = ~\a[39]  & \b[31]  ;
  assign n27919 = n8751 & n27918 ;
  assign n27920 = ~n27917 & ~n27919 ;
  assign n27921 = \b[32]  & n8757 ;
  assign n27922 = \a[39]  & \b[31]  ;
  assign n27923 = n8748 & n27922 ;
  assign n27924 = \a[41]  & ~n27923 ;
  assign n27925 = ~n27921 & n27924 ;
  assign n27926 = n27920 & n27925 ;
  assign n27927 = ~n27915 & n27926 ;
  assign n27928 = ~n27912 & n27927 ;
  assign n27929 = ~n27921 & ~n27923 ;
  assign n27930 = n27920 & n27929 ;
  assign n27931 = ~n27915 & n27930 ;
  assign n27932 = ~n27912 & n27931 ;
  assign n27933 = ~\a[41]  & ~n27932 ;
  assign n27934 = ~n27928 & ~n27933 ;
  assign n27935 = ~n27910 & n27934 ;
  assign n27936 = n27910 & ~n27934 ;
  assign n27937 = ~n27935 & ~n27936 ;
  assign n27938 = ~n27345 & n27370 ;
  assign n27939 = ~n27344 & ~n27938 ;
  assign n27940 = ~n6610 & n7534 ;
  assign n27941 = ~n6608 & n27940 ;
  assign n27942 = \b[33]  & n7973 ;
  assign n27943 = n7970 & n27942 ;
  assign n27944 = ~\a[36]  & \b[34]  ;
  assign n27945 = n7526 & n27944 ;
  assign n27946 = ~n27943 & ~n27945 ;
  assign n27947 = \b[35]  & n7532 ;
  assign n27948 = \a[36]  & \b[34]  ;
  assign n27949 = n17801 & n27948 ;
  assign n27950 = \a[38]  & ~n27949 ;
  assign n27951 = ~n27947 & n27950 ;
  assign n27952 = n27946 & n27951 ;
  assign n27953 = ~n27941 & n27952 ;
  assign n27954 = ~n27947 & ~n27949 ;
  assign n27955 = n27946 & n27954 ;
  assign n27956 = ~n27941 & n27955 ;
  assign n27957 = ~\a[38]  & ~n27956 ;
  assign n27958 = ~n27953 & ~n27957 ;
  assign n27959 = ~n27939 & n27958 ;
  assign n27960 = ~n27937 & n27959 ;
  assign n27961 = n27939 & n27958 ;
  assign n27962 = n27937 & n27961 ;
  assign n27963 = ~n27960 & ~n27962 ;
  assign n27964 = ~n27939 & ~n27958 ;
  assign n27965 = n27937 & n27964 ;
  assign n27966 = n27939 & ~n27958 ;
  assign n27967 = ~n27937 & n27966 ;
  assign n27968 = ~n27965 & ~n27967 ;
  assign n27969 = n27963 & n27968 ;
  assign n27970 = n27678 & ~n27969 ;
  assign n27971 = ~n27678 & n27969 ;
  assign n27972 = ~n27970 & ~n27971 ;
  assign n27973 = n6309 & n8175 ;
  assign n27974 = ~n8172 & n27973 ;
  assign n27975 = n6309 & ~n8175 ;
  assign n27976 = ~n7756 & n27975 ;
  assign n27977 = ~n8171 & n27976 ;
  assign n27978 = \b[36]  & n6778 ;
  assign n27979 = n6775 & n27978 ;
  assign n27980 = ~\a[33]  & \b[37]  ;
  assign n27981 = n6301 & n27980 ;
  assign n27982 = ~n27979 & ~n27981 ;
  assign n27983 = \b[38]  & n6307 ;
  assign n27984 = \a[33]  & \b[37]  ;
  assign n27985 = n6298 & n27984 ;
  assign n27986 = \a[35]  & ~n27985 ;
  assign n27987 = ~n27983 & n27986 ;
  assign n27988 = n27982 & n27987 ;
  assign n27989 = ~n27977 & n27988 ;
  assign n27990 = ~n27974 & n27989 ;
  assign n27991 = ~n27983 & ~n27985 ;
  assign n27992 = n27982 & n27991 ;
  assign n27993 = ~n27977 & n27992 ;
  assign n27994 = ~n27974 & n27993 ;
  assign n27995 = ~\a[35]  & ~n27994 ;
  assign n27996 = ~n27990 & ~n27995 ;
  assign n27997 = n27972 & ~n27996 ;
  assign n27998 = ~n27972 & n27996 ;
  assign n27999 = ~n27997 & ~n27998 ;
  assign n28000 = n27676 & n27999 ;
  assign n28001 = ~n27676 & ~n27999 ;
  assign n28002 = ~n28000 & ~n28001 ;
  assign n28003 = ~n27081 & n27421 ;
  assign n28004 = ~n27076 & ~n28003 ;
  assign n28005 = ~n10886 & ~n10889 ;
  assign n28006 = ~n10404 & n10889 ;
  assign n28007 = ~n10885 & n28006 ;
  assign n28008 = n4249 & ~n28007 ;
  assign n28009 = ~n28005 & n28008 ;
  assign n28010 = \b[44]  & n4247 ;
  assign n28011 = \a[27]  & \b[43]  ;
  assign n28012 = n4238 & n28011 ;
  assign n28013 = ~n28010 & ~n28012 ;
  assign n28014 = \b[42]  & n4647 ;
  assign n28015 = n4644 & n28014 ;
  assign n28016 = ~\a[27]  & \b[43]  ;
  assign n28017 = n4241 & n28016 ;
  assign n28018 = ~n28015 & ~n28017 ;
  assign n28019 = n28013 & n28018 ;
  assign n28020 = ~n28009 & n28019 ;
  assign n28021 = \a[29]  & ~n28020 ;
  assign n28022 = ~\a[29]  & n28020 ;
  assign n28023 = ~n28021 & ~n28022 ;
  assign n28024 = n28004 & n28023 ;
  assign n28025 = ~\a[29]  & ~n28020 ;
  assign n28026 = \a[29]  & n28019 ;
  assign n28027 = ~n28009 & n28026 ;
  assign n28028 = ~n28025 & ~n28027 ;
  assign n28029 = ~n28004 & n28028 ;
  assign n28030 = ~n28024 & ~n28029 ;
  assign n28031 = n28002 & n28030 ;
  assign n28032 = ~n28002 & ~n28030 ;
  assign n28033 = ~n28031 & ~n28032 ;
  assign n28034 = n27646 & n28033 ;
  assign n28035 = ~n27646 & ~n28033 ;
  assign n28036 = ~n28034 & ~n28035 ;
  assign n28037 = ~n27619 & ~n28036 ;
  assign n28038 = ~n27613 & n28036 ;
  assign n28039 = ~n27618 & n28038 ;
  assign n28040 = ~n28037 & ~n28039 ;
  assign n28041 = ~n27461 & n27466 ;
  assign n28042 = ~n27442 & ~n27461 ;
  assign n28043 = ~n28041 & ~n28042 ;
  assign n28044 = n1965 & ~n15246 ;
  assign n28045 = ~n15244 & n28044 ;
  assign n28046 = \b[53]  & n1963 ;
  assign n28047 = \a[17]  & ~\a[19]  ;
  assign n28048 = \a[18]  & \b[52]  ;
  assign n28049 = n28047 & n28048 ;
  assign n28050 = ~n28046 & ~n28049 ;
  assign n28051 = \b[51]  & n2218 ;
  assign n28052 = n2216 & n28051 ;
  assign n28053 = ~\a[18]  & \b[52]  ;
  assign n28054 = n1957 & n28053 ;
  assign n28055 = ~n28052 & ~n28054 ;
  assign n28056 = n28050 & n28055 ;
  assign n28057 = ~n28045 & n28056 ;
  assign n28058 = \a[20]  & ~n28057 ;
  assign n28059 = ~\a[20]  & n28057 ;
  assign n28060 = ~n28058 & ~n28059 ;
  assign n28061 = n28043 & n28060 ;
  assign n28062 = ~\a[20]  & ~n28057 ;
  assign n28063 = \a[20]  & n28056 ;
  assign n28064 = ~n28045 & n28063 ;
  assign n28065 = ~n28062 & ~n28064 ;
  assign n28066 = ~n28043 & n28065 ;
  assign n28067 = ~n28061 & ~n28066 ;
  assign n28068 = n28040 & n28067 ;
  assign n28069 = ~n28040 & ~n28067 ;
  assign n28070 = ~n28068 & ~n28069 ;
  assign n28071 = ~n27586 & n28070 ;
  assign n28072 = ~n27582 & n28071 ;
  assign n28073 = ~n27582 & ~n27586 ;
  assign n28074 = ~n28070 & ~n28073 ;
  assign n28075 = ~n28072 & ~n28074 ;
  assign n28076 = n27556 & n28075 ;
  assign n28077 = ~n27556 & ~n28075 ;
  assign n28078 = ~n28076 & ~n28077 ;
  assign n28079 = n26937 & ~n27485 ;
  assign n28080 = n26930 & n26937 ;
  assign n28081 = ~n28079 & ~n28080 ;
  assign n28082 = n646 & n21696 ;
  assign n28083 = ~n21693 & n28082 ;
  assign n28084 = n646 & ~n21696 ;
  assign n28085 = ~n20966 & n28084 ;
  assign n28086 = ~n21692 & n28085 ;
  assign n28087 = \b[60]  & n796 ;
  assign n28088 = n793 & n28087 ;
  assign n28089 = \b[62]  & n644 ;
  assign n28090 = \a[8]  & \b[61]  ;
  assign n28091 = n794 & n28090 ;
  assign n28092 = ~\a[9]  & \b[61]  ;
  assign n28093 = n638 & n28092 ;
  assign n28094 = ~n28091 & ~n28093 ;
  assign n28095 = ~n28089 & n28094 ;
  assign n28096 = ~n28088 & n28095 ;
  assign n28097 = ~n28086 & n28096 ;
  assign n28098 = ~n28083 & n28097 ;
  assign n28099 = \a[11]  & ~n28098 ;
  assign n28100 = ~\a[11]  & n28098 ;
  assign n28101 = ~n28099 & ~n28100 ;
  assign n28102 = n28081 & n28101 ;
  assign n28103 = ~\a[11]  & ~n28098 ;
  assign n28104 = \a[11]  & n28096 ;
  assign n28105 = ~n28086 & n28104 ;
  assign n28106 = ~n28083 & n28105 ;
  assign n28107 = ~n28103 & ~n28106 ;
  assign n28108 = ~n28081 & n28107 ;
  assign n28109 = ~n28102 & ~n28108 ;
  assign n28110 = n28078 & n28109 ;
  assign n28111 = ~n28078 & ~n28109 ;
  assign n28112 = ~n28110 & ~n28111 ;
  assign n28113 = n27493 & ~n27527 ;
  assign n28114 = ~n26899 & n28113 ;
  assign n28115 = n26903 & ~n27527 ;
  assign n28116 = ~n28114 & ~n28115 ;
  assign n28117 = n28112 & n28116 ;
  assign n28118 = ~n27528 & n28117 ;
  assign n28119 = ~n27527 & ~n28112 ;
  assign n28120 = n27511 & n28119 ;
  assign n28121 = n27527 & ~n28112 ;
  assign n28122 = ~n27511 & n28121 ;
  assign n28123 = ~n28120 & ~n28122 ;
  assign n28124 = ~n28118 & n28123 ;
  assign n28125 = ~n26874 & ~n27496 ;
  assign n28126 = n26878 & ~n28125 ;
  assign n28127 = n28124 & n28126 ;
  assign n28128 = ~n28124 & ~n28126 ;
  assign n28129 = ~n28127 & ~n28128 ;
  assign n28130 = ~n27501 & n28129 ;
  assign n28131 = ~n27508 & n28130 ;
  assign n28132 = ~n27501 & ~n27508 ;
  assign n28133 = ~n28129 & ~n28132 ;
  assign n28134 = ~n28131 & ~n28133 ;
  assign n28135 = ~n28127 & ~n28131 ;
  assign n28136 = n28116 & ~n28118 ;
  assign n28137 = ~n28102 & n28108 ;
  assign n28138 = ~n28078 & ~n28102 ;
  assign n28139 = ~n28137 & ~n28138 ;
  assign n28140 = n646 & ~n22461 ;
  assign n28141 = ~n22459 & n28140 ;
  assign n28142 = \b[63]  & n644 ;
  assign n28143 = \a[8]  & ~\a[10]  ;
  assign n28144 = \a[9]  & \b[62]  ;
  assign n28145 = n28143 & n28144 ;
  assign n28146 = ~n28142 & ~n28145 ;
  assign n28147 = \b[61]  & n796 ;
  assign n28148 = n793 & n28147 ;
  assign n28149 = ~\a[9]  & \b[62]  ;
  assign n28150 = n638 & n28149 ;
  assign n28151 = ~n28148 & ~n28150 ;
  assign n28152 = n28146 & n28151 ;
  assign n28153 = ~n28141 & n28152 ;
  assign n28154 = ~\a[11]  & ~n28153 ;
  assign n28155 = \a[11]  & n28152 ;
  assign n28156 = ~n28141 & n28155 ;
  assign n28157 = ~n28154 & ~n28156 ;
  assign n28158 = ~n28139 & n28157 ;
  assign n28159 = ~n27550 & ~n28075 ;
  assign n28160 = ~n27550 & n27555 ;
  assign n28161 = ~n28159 & ~n28160 ;
  assign n28162 = n1467 & ~n17690 ;
  assign n28163 = ~n17688 & n28162 ;
  assign n28164 = \b[57]  & n1465 ;
  assign n28165 = \a[15]  & \b[56]  ;
  assign n28166 = n1456 & n28165 ;
  assign n28167 = ~n28164 & ~n28166 ;
  assign n28168 = \b[55]  & n1652 ;
  assign n28169 = n1649 & n28168 ;
  assign n28170 = ~\a[15]  & \b[56]  ;
  assign n28171 = n1459 & n28170 ;
  assign n28172 = ~n28169 & ~n28171 ;
  assign n28173 = n28167 & n28172 ;
  assign n28174 = ~n28163 & n28173 ;
  assign n28175 = ~\a[17]  & ~n28174 ;
  assign n28176 = \a[17]  & n28173 ;
  assign n28177 = ~n28163 & n28176 ;
  assign n28178 = ~n28175 & ~n28177 ;
  assign n28179 = ~n27586 & ~n28070 ;
  assign n28180 = ~n27582 & ~n28179 ;
  assign n28181 = n28178 & ~n28180 ;
  assign n28182 = ~n28178 & n28180 ;
  assign n28183 = ~n28181 & ~n28182 ;
  assign n28184 = n999 & n20260 ;
  assign n28185 = ~n20257 & n28184 ;
  assign n28186 = n999 & ~n20260 ;
  assign n28187 = ~n19545 & n28186 ;
  assign n28188 = ~n20256 & n28187 ;
  assign n28189 = \b[58]  & n1182 ;
  assign n28190 = n1179 & n28189 ;
  assign n28191 = ~\a[12]  & \b[59]  ;
  assign n28192 = n7674 & n28191 ;
  assign n28193 = ~n28190 & ~n28192 ;
  assign n28194 = \b[60]  & n997 ;
  assign n28195 = \a[11]  & ~\a[13]  ;
  assign n28196 = \a[12]  & \b[59]  ;
  assign n28197 = n28195 & n28196 ;
  assign n28198 = \a[14]  & ~n28197 ;
  assign n28199 = ~n28194 & n28198 ;
  assign n28200 = n28193 & n28199 ;
  assign n28201 = ~n28188 & n28200 ;
  assign n28202 = ~n28185 & n28201 ;
  assign n28203 = ~n28194 & ~n28197 ;
  assign n28204 = n28193 & n28203 ;
  assign n28205 = ~n28188 & n28204 ;
  assign n28206 = ~n28185 & n28205 ;
  assign n28207 = ~\a[14]  & ~n28206 ;
  assign n28208 = ~n28202 & ~n28207 ;
  assign n28209 = ~n27023 & n27605 ;
  assign n28210 = ~n26999 & n28209 ;
  assign n28211 = n27431 & n27605 ;
  assign n28212 = ~n26999 & n28211 ;
  assign n28213 = n27431 & n28209 ;
  assign n28214 = ~n28212 & ~n28213 ;
  assign n28215 = ~n28210 & n28214 ;
  assign n28216 = \a[23]  & n27587 ;
  assign n28217 = n26999 & n27023 ;
  assign n28218 = \a[23]  & n27431 ;
  assign n28219 = ~n28217 & n28218 ;
  assign n28220 = ~n28216 & ~n28219 ;
  assign n28221 = n27604 & ~n28220 ;
  assign n28222 = ~n28038 & ~n28221 ;
  assign n28223 = n28215 & n28222 ;
  assign n28224 = n2622 & ~n14098 ;
  assign n28225 = ~n14096 & n28224 ;
  assign n28226 = \b[49]  & n2912 ;
  assign n28227 = n2909 & n28226 ;
  assign n28228 = \b[51]  & n2620 ;
  assign n28229 = \a[20]  & \b[50]  ;
  assign n28230 = n2910 & n28229 ;
  assign n28231 = ~\a[21]  & \b[50]  ;
  assign n28232 = n2614 & n28231 ;
  assign n28233 = ~n28230 & ~n28232 ;
  assign n28234 = ~n28228 & n28233 ;
  assign n28235 = ~n28227 & n28234 ;
  assign n28236 = ~n28225 & n28235 ;
  assign n28237 = ~\a[23]  & ~n28236 ;
  assign n28238 = \a[23]  & n28235 ;
  assign n28239 = ~n28225 & n28238 ;
  assign n28240 = ~n28237 & ~n28239 ;
  assign n28241 = ~n27640 & ~n28033 ;
  assign n28242 = ~n27640 & n27645 ;
  assign n28243 = ~n28241 & ~n28242 ;
  assign n28244 = n4249 & ~n11397 ;
  assign n28245 = ~n11395 & n28244 ;
  assign n28246 = \b[43]  & n4647 ;
  assign n28247 = n4644 & n28246 ;
  assign n28248 = ~\a[27]  & \b[44]  ;
  assign n28249 = n4241 & n28248 ;
  assign n28250 = ~n28247 & ~n28249 ;
  assign n28251 = \b[45]  & n4247 ;
  assign n28252 = \a[27]  & \b[44]  ;
  assign n28253 = n4238 & n28252 ;
  assign n28254 = \a[29]  & ~n28253 ;
  assign n28255 = ~n28251 & n28254 ;
  assign n28256 = n28250 & n28255 ;
  assign n28257 = ~n28245 & n28256 ;
  assign n28258 = ~n28251 & ~n28253 ;
  assign n28259 = n28250 & n28258 ;
  assign n28260 = ~n28245 & n28259 ;
  assign n28261 = ~\a[29]  & ~n28260 ;
  assign n28262 = ~n28257 & ~n28261 ;
  assign n28263 = n28002 & ~n28262 ;
  assign n28264 = ~n28029 & n28263 ;
  assign n28265 = n28024 & ~n28262 ;
  assign n28266 = ~n28264 & ~n28265 ;
  assign n28267 = ~n28024 & n28029 ;
  assign n28268 = ~n28002 & ~n28024 ;
  assign n28269 = ~n28267 & ~n28268 ;
  assign n28270 = n28262 & ~n28269 ;
  assign n28271 = n28266 & ~n28270 ;
  assign n28272 = n5211 & n9930 ;
  assign n28273 = ~n9927 & n28272 ;
  assign n28274 = n5211 & ~n9930 ;
  assign n28275 = ~n9477 & n28274 ;
  assign n28276 = ~n9926 & n28275 ;
  assign n28277 = \b[40]  & n5595 ;
  assign n28278 = n5592 & n28277 ;
  assign n28279 = ~\a[30]  & \b[41]  ;
  assign n28280 = n5203 & n28279 ;
  assign n28281 = ~n28278 & ~n28280 ;
  assign n28282 = \b[42]  & n5209 ;
  assign n28283 = \a[30]  & \b[41]  ;
  assign n28284 = n5200 & n28283 ;
  assign n28285 = \a[32]  & ~n28284 ;
  assign n28286 = ~n28282 & n28285 ;
  assign n28287 = n28281 & n28286 ;
  assign n28288 = ~n28276 & n28287 ;
  assign n28289 = ~n28273 & n28288 ;
  assign n28290 = ~n28282 & ~n28284 ;
  assign n28291 = n28281 & n28290 ;
  assign n28292 = ~n28276 & n28291 ;
  assign n28293 = ~n28273 & n28292 ;
  assign n28294 = ~\a[32]  & ~n28293 ;
  assign n28295 = ~n28289 & ~n28294 ;
  assign n28296 = ~n27675 & ~n27999 ;
  assign n28297 = n27671 & ~n27675 ;
  assign n28298 = ~n28296 & ~n28297 ;
  assign n28299 = ~n27971 & n27996 ;
  assign n28300 = n27970 & ~n27971 ;
  assign n28301 = ~n28299 & ~n28300 ;
  assign n28302 = ~n3283 & ~n12606 ;
  assign n28303 = ~n13122 & n28302 ;
  assign n28304 = n3280 & n28303 ;
  assign n28305 = n3283 & ~n12606 ;
  assign n28306 = ~n13122 & n28305 ;
  assign n28307 = ~n3280 & n28306 ;
  assign n28308 = ~n28304 & ~n28307 ;
  assign n28309 = \b[22]  & n13794 ;
  assign n28310 = n13792 & n28309 ;
  assign n28311 = \b[24]  & n13123 ;
  assign n28312 = \a[48]  & \b[23]  ;
  assign n28313 = n13786 & n28312 ;
  assign n28314 = ~\a[48]  & \b[23]  ;
  assign n28315 = n13117 & n28314 ;
  assign n28316 = ~n28313 & ~n28315 ;
  assign n28317 = ~n28311 & n28316 ;
  assign n28318 = ~n28310 & n28317 ;
  assign n28319 = n28308 & n28318 ;
  assign n28320 = ~\a[50]  & ~n28319 ;
  assign n28321 = \a[50]  & n28318 ;
  assign n28322 = n28308 & n28321 ;
  assign n28323 = ~n28320 & ~n28322 ;
  assign n28324 = ~n27797 & n27822 ;
  assign n28325 = n27796 & ~n27797 ;
  assign n28326 = ~n28324 & ~n28325 ;
  assign n28327 = n27720 & ~n27756 ;
  assign n28328 = ~n27757 & ~n28327 ;
  assign n28329 = ~n1230 & n18516 ;
  assign n28330 = ~n1086 & n18516 ;
  assign n28331 = ~n1226 & n28330 ;
  assign n28332 = ~n28329 & ~n28331 ;
  assign n28333 = ~n1233 & ~n28332 ;
  assign n28334 = \b[15]  & n18514 ;
  assign n28335 = \a[56]  & \b[14]  ;
  assign n28336 = n19181 & n28335 ;
  assign n28337 = ~\a[57]  & \b[14]  ;
  assign n28338 = n18508 & n28337 ;
  assign n28339 = ~n28336 & ~n28338 ;
  assign n28340 = ~n28334 & n28339 ;
  assign n28341 = \b[13]  & n19183 ;
  assign n28342 = n19180 & n28341 ;
  assign n28343 = \a[59]  & ~n28342 ;
  assign n28344 = n28340 & n28343 ;
  assign n28345 = ~n28333 & n28344 ;
  assign n28346 = n28340 & ~n28342 ;
  assign n28347 = ~\a[59]  & ~n28346 ;
  assign n28348 = ~\a[59]  & ~n1233 ;
  assign n28349 = ~n28332 & n28348 ;
  assign n28350 = ~n28347 & ~n28349 ;
  assign n28351 = ~n28345 & n28350 ;
  assign n28352 = ~n909 & ~n19861 ;
  assign n28353 = ~n20518 & n28352 ;
  assign n28354 = n906 & n28353 ;
  assign n28355 = n909 & ~n19861 ;
  assign n28356 = ~n20518 & n28355 ;
  assign n28357 = ~n906 & n28356 ;
  assign n28358 = ~n28354 & ~n28357 ;
  assign n28359 = \b[10]  & n21315 ;
  assign n28360 = n21312 & n28359 ;
  assign n28361 = \b[12]  & n20519 ;
  assign n28362 = \a[59]  & \b[11]  ;
  assign n28363 = n21313 & n28362 ;
  assign n28364 = ~\a[60]  & \b[11]  ;
  assign n28365 = n20513 & n28364 ;
  assign n28366 = ~n28363 & ~n28365 ;
  assign n28367 = ~n28361 & n28366 ;
  assign n28368 = ~n28360 & n28367 ;
  assign n28369 = n28358 & n28368 ;
  assign n28370 = ~\a[62]  & ~n28369 ;
  assign n28371 = \a[62]  & n28368 ;
  assign n28372 = n28358 & n28371 ;
  assign n28373 = ~n28370 & ~n28372 ;
  assign n28374 = ~n27152 & ~n27751 ;
  assign n28375 = ~n27149 & n28374 ;
  assign n28376 = ~n27141 & n28375 ;
  assign n28377 = ~\a[8]  & n27748 ;
  assign n28378 = ~\a[8]  & \b[8]  ;
  assign n28379 = n21958 & n28378 ;
  assign n28380 = ~n28377 & ~n28379 ;
  assign n28381 = \a[8]  & ~n27748 ;
  assign n28382 = ~n27747 & n28381 ;
  assign n28383 = n28380 & ~n28382 ;
  assign n28384 = \b[9]  & n21958 ;
  assign n28385 = \b[8]  & n21957 ;
  assign n28386 = ~n28384 & ~n28385 ;
  assign n28387 = ~n28383 & ~n28386 ;
  assign n28388 = n28383 & n28386 ;
  assign n28389 = ~n28387 & ~n28388 ;
  assign n28390 = ~n27750 & ~n28389 ;
  assign n28391 = ~n28376 & n28390 ;
  assign n28392 = ~n27750 & ~n28376 ;
  assign n28393 = n28389 & ~n28392 ;
  assign n28394 = ~n28391 & ~n28393 ;
  assign n28395 = n28373 & ~n28394 ;
  assign n28396 = ~n28373 & n28394 ;
  assign n28397 = ~n28395 & ~n28396 ;
  assign n28398 = n28351 & ~n28397 ;
  assign n28399 = ~n28351 & n28397 ;
  assign n28400 = ~n28398 & ~n28399 ;
  assign n28401 = n28328 & n28400 ;
  assign n28402 = ~n28328 & n28398 ;
  assign n28403 = ~n28328 & n28399 ;
  assign n28404 = ~n28402 & ~n28403 ;
  assign n28405 = ~n28401 & n28404 ;
  assign n28406 = n1875 & n16655 ;
  assign n28407 = ~n1872 & n28406 ;
  assign n28408 = n5000 & n16655 ;
  assign n28409 = ~n1871 & n28408 ;
  assign n28410 = \b[16]  & n17308 ;
  assign n28411 = n17305 & n28410 ;
  assign n28412 = \b[18]  & n16653 ;
  assign n28413 = \a[53]  & \b[17]  ;
  assign n28414 = n17306 & n28413 ;
  assign n28415 = ~\a[54]  & \b[17]  ;
  assign n28416 = n16647 & n28415 ;
  assign n28417 = ~n28414 & ~n28416 ;
  assign n28418 = ~n28412 & n28417 ;
  assign n28419 = ~n28411 & n28418 ;
  assign n28420 = ~n28409 & n28419 ;
  assign n28421 = ~n28407 & n28420 ;
  assign n28422 = ~\a[56]  & ~n28421 ;
  assign n28423 = \a[56]  & n28419 ;
  assign n28424 = ~n28409 & n28423 ;
  assign n28425 = ~n28407 & n28424 ;
  assign n28426 = ~n28422 & ~n28425 ;
  assign n28427 = n28405 & ~n28426 ;
  assign n28428 = ~n28405 & n28426 ;
  assign n28429 = ~n28427 & ~n28428 ;
  assign n28430 = ~n27765 & n27790 ;
  assign n28431 = ~n27764 & ~n28430 ;
  assign n28432 = ~n28429 & ~n28431 ;
  assign n28433 = n28429 & n28431 ;
  assign n28434 = ~n28432 & ~n28433 ;
  assign n28435 = ~n2520 & n14793 ;
  assign n28436 = ~n2292 & n14793 ;
  assign n28437 = ~n2516 & n28436 ;
  assign n28438 = ~n28435 & ~n28437 ;
  assign n28439 = ~n2523 & ~n28438 ;
  assign n28440 = \b[19]  & n15517 ;
  assign n28441 = n15514 & n28440 ;
  assign n28442 = \b[21]  & n14791 ;
  assign n28443 = \a[50]  & \b[20]  ;
  assign n28444 = n15515 & n28443 ;
  assign n28445 = ~\a[51]  & \b[20]  ;
  assign n28446 = n14785 & n28445 ;
  assign n28447 = ~n28444 & ~n28446 ;
  assign n28448 = ~n28442 & n28447 ;
  assign n28449 = ~n28441 & n28448 ;
  assign n28450 = ~\a[53]  & n28449 ;
  assign n28451 = ~n28439 & n28450 ;
  assign n28452 = \a[53]  & ~n28449 ;
  assign n28453 = \a[53]  & ~n2523 ;
  assign n28454 = ~n28438 & n28453 ;
  assign n28455 = ~n28452 & ~n28454 ;
  assign n28456 = ~n28451 & n28455 ;
  assign n28457 = n28434 & n28456 ;
  assign n28458 = ~n28434 & ~n28456 ;
  assign n28459 = ~n28457 & ~n28458 ;
  assign n28460 = n28326 & n28459 ;
  assign n28461 = ~n28326 & ~n28459 ;
  assign n28462 = ~n28460 & ~n28461 ;
  assign n28463 = ~n28323 & n28462 ;
  assign n28464 = n28323 & ~n28462 ;
  assign n28465 = ~n28463 & ~n28464 ;
  assign n28466 = ~n4145 & n11572 ;
  assign n28467 = ~n3603 & n11572 ;
  assign n28468 = ~n4141 & n28467 ;
  assign n28469 = ~n28466 & ~n28468 ;
  assign n28470 = ~n4148 & ~n28469 ;
  assign n28471 = \b[25]  & n12159 ;
  assign n28472 = n12156 & n28471 ;
  assign n28473 = ~\a[45]  & \b[26]  ;
  assign n28474 = n11564 & n28473 ;
  assign n28475 = ~n28472 & ~n28474 ;
  assign n28476 = \b[27]  & n11570 ;
  assign n28477 = \a[45]  & \b[26]  ;
  assign n28478 = n11561 & n28477 ;
  assign n28479 = \a[47]  & ~n28478 ;
  assign n28480 = ~n28476 & n28479 ;
  assign n28481 = n28475 & n28480 ;
  assign n28482 = ~n28470 & n28481 ;
  assign n28483 = ~n28476 & ~n28478 ;
  assign n28484 = n28475 & n28483 ;
  assign n28485 = ~\a[47]  & ~n28484 ;
  assign n28486 = ~\a[47]  & ~n4148 ;
  assign n28487 = ~n28469 & n28486 ;
  assign n28488 = ~n28485 & ~n28487 ;
  assign n28489 = ~n28482 & n28488 ;
  assign n28490 = n27697 & ~n27828 ;
  assign n28491 = ~n27829 & ~n28490 ;
  assign n28492 = ~n28489 & n28491 ;
  assign n28493 = ~n28465 & n28492 ;
  assign n28494 = ~n28489 & ~n28491 ;
  assign n28495 = n28465 & n28494 ;
  assign n28496 = ~n28493 & ~n28495 ;
  assign n28497 = n28489 & ~n28491 ;
  assign n28498 = ~n28465 & n28497 ;
  assign n28499 = n28489 & n28491 ;
  assign n28500 = n28465 & n28499 ;
  assign n28501 = ~n28498 & ~n28500 ;
  assign n28502 = n28496 & n28501 ;
  assign n28503 = n27833 & ~n27837 ;
  assign n28504 = ~n27833 & n27837 ;
  assign n28505 = n27861 & ~n28504 ;
  assign n28506 = ~n28503 & ~n28505 ;
  assign n28507 = ~n5105 & ~n9646 ;
  assign n28508 = ~n10079 & n28507 ;
  assign n28509 = n5102 & n28508 ;
  assign n28510 = n5105 & ~n9646 ;
  assign n28511 = ~n10079 & n28510 ;
  assign n28512 = ~n5102 & n28511 ;
  assign n28513 = ~n28509 & ~n28512 ;
  assign n28514 = \b[28]  & n10681 ;
  assign n28515 = n10678 & n28514 ;
  assign n28516 = \b[30]  & n10080 ;
  assign n28517 = \a[41]  & \b[29]  ;
  assign n28518 = n10679 & n28517 ;
  assign n28519 = ~\a[42]  & \b[29]  ;
  assign n28520 = n10074 & n28519 ;
  assign n28521 = ~n28518 & ~n28520 ;
  assign n28522 = ~n28516 & n28521 ;
  assign n28523 = ~n28515 & n28522 ;
  assign n28524 = n28513 & n28523 ;
  assign n28525 = ~\a[44]  & ~n28524 ;
  assign n28526 = \a[44]  & n28523 ;
  assign n28527 = n28513 & n28526 ;
  assign n28528 = ~n28525 & ~n28527 ;
  assign n28529 = ~n28506 & n28528 ;
  assign n28530 = ~n28502 & n28529 ;
  assign n28531 = n28506 & n28528 ;
  assign n28532 = n28502 & n28531 ;
  assign n28533 = ~n28530 & ~n28532 ;
  assign n28534 = ~n28506 & ~n28528 ;
  assign n28535 = n28502 & n28534 ;
  assign n28536 = n28506 & ~n28528 ;
  assign n28537 = ~n28502 & n28536 ;
  assign n28538 = ~n28535 & ~n28537 ;
  assign n28539 = n28533 & n28538 ;
  assign n28540 = ~n5855 & n8759 ;
  assign n28541 = ~n5853 & n28540 ;
  assign n28542 = \b[31]  & n9301 ;
  assign n28543 = n9298 & n28542 ;
  assign n28544 = ~\a[39]  & \b[32]  ;
  assign n28545 = n8751 & n28544 ;
  assign n28546 = ~n28543 & ~n28545 ;
  assign n28547 = \b[33]  & n8757 ;
  assign n28548 = \a[39]  & \b[32]  ;
  assign n28549 = n8748 & n28548 ;
  assign n28550 = \a[41]  & ~n28549 ;
  assign n28551 = ~n28547 & n28550 ;
  assign n28552 = n28546 & n28551 ;
  assign n28553 = ~n28541 & n28552 ;
  assign n28554 = ~n28547 & ~n28549 ;
  assign n28555 = n28546 & n28554 ;
  assign n28556 = ~n28541 & n28555 ;
  assign n28557 = ~\a[41]  & ~n28556 ;
  assign n28558 = ~n28553 & ~n28557 ;
  assign n28559 = ~n27872 & ~n27874 ;
  assign n28560 = n27872 & n27874 ;
  assign n28561 = n27892 & ~n28560 ;
  assign n28562 = ~n28559 & ~n28561 ;
  assign n28563 = ~n28558 & ~n28562 ;
  assign n28564 = n28539 & n28563 ;
  assign n28565 = ~n28558 & n28562 ;
  assign n28566 = ~n28539 & n28565 ;
  assign n28567 = ~n28564 & ~n28566 ;
  assign n28568 = n28558 & ~n28562 ;
  assign n28569 = ~n28539 & n28568 ;
  assign n28570 = n28558 & n28562 ;
  assign n28571 = n28539 & n28570 ;
  assign n28572 = ~n28569 & ~n28571 ;
  assign n28573 = n28567 & n28572 ;
  assign n28574 = n7337 & n7534 ;
  assign n28575 = ~n7334 & n28574 ;
  assign n28576 = ~n7337 & n7534 ;
  assign n28577 = ~n6605 & n28576 ;
  assign n28578 = ~n7333 & n28577 ;
  assign n28579 = \b[34]  & n7973 ;
  assign n28580 = n7970 & n28579 ;
  assign n28581 = ~\a[36]  & \b[35]  ;
  assign n28582 = n7526 & n28581 ;
  assign n28583 = ~n28580 & ~n28582 ;
  assign n28584 = \b[36]  & n7532 ;
  assign n28585 = \a[36]  & \b[35]  ;
  assign n28586 = n17801 & n28585 ;
  assign n28587 = \a[38]  & ~n28586 ;
  assign n28588 = ~n28584 & n28587 ;
  assign n28589 = n28583 & n28588 ;
  assign n28590 = ~n28578 & n28589 ;
  assign n28591 = ~n28575 & n28590 ;
  assign n28592 = ~n28584 & ~n28586 ;
  assign n28593 = n28583 & n28592 ;
  assign n28594 = ~n28578 & n28593 ;
  assign n28595 = ~n28575 & n28594 ;
  assign n28596 = ~\a[38]  & ~n28595 ;
  assign n28597 = ~n28591 & ~n28596 ;
  assign n28598 = ~n27909 & n27934 ;
  assign n28599 = n27908 & ~n27909 ;
  assign n28600 = ~n28598 & ~n28599 ;
  assign n28601 = ~n28597 & n28600 ;
  assign n28602 = ~n28573 & n28601 ;
  assign n28603 = ~n28597 & ~n28600 ;
  assign n28604 = n28573 & n28603 ;
  assign n28605 = ~n28602 & ~n28604 ;
  assign n28606 = n28597 & ~n28600 ;
  assign n28607 = ~n28573 & n28606 ;
  assign n28608 = n28597 & n28600 ;
  assign n28609 = n28573 & n28608 ;
  assign n28610 = ~n28607 & ~n28609 ;
  assign n28611 = n28605 & n28610 ;
  assign n28612 = ~n27937 & ~n27939 ;
  assign n28613 = n27937 & n27939 ;
  assign n28614 = n27958 & ~n28613 ;
  assign n28615 = ~n28612 & ~n28614 ;
  assign n28616 = ~n28611 & ~n28615 ;
  assign n28617 = n28611 & n28615 ;
  assign n28618 = ~n28616 & ~n28617 ;
  assign n28619 = n6309 & ~n8602 ;
  assign n28620 = ~n8600 & n28619 ;
  assign n28621 = \b[37]  & n6778 ;
  assign n28622 = n6775 & n28621 ;
  assign n28623 = ~\a[33]  & \b[38]  ;
  assign n28624 = n6301 & n28623 ;
  assign n28625 = ~n28622 & ~n28624 ;
  assign n28626 = \b[39]  & n6307 ;
  assign n28627 = \a[33]  & \b[38]  ;
  assign n28628 = n6298 & n28627 ;
  assign n28629 = \a[35]  & ~n28628 ;
  assign n28630 = ~n28626 & n28629 ;
  assign n28631 = n28625 & n28630 ;
  assign n28632 = ~n28620 & n28631 ;
  assign n28633 = ~n28626 & ~n28628 ;
  assign n28634 = n28625 & n28633 ;
  assign n28635 = ~n28620 & n28634 ;
  assign n28636 = ~\a[35]  & ~n28635 ;
  assign n28637 = ~n28632 & ~n28636 ;
  assign n28638 = n28618 & ~n28637 ;
  assign n28639 = ~n28618 & n28637 ;
  assign n28640 = ~n28638 & ~n28639 ;
  assign n28641 = n28301 & n28640 ;
  assign n28642 = ~n28301 & ~n28640 ;
  assign n28643 = ~n28641 & ~n28642 ;
  assign n28644 = ~n28298 & ~n28643 ;
  assign n28645 = n28295 & n28644 ;
  assign n28646 = ~n28295 & n28301 ;
  assign n28647 = ~n28640 & n28646 ;
  assign n28648 = ~n28295 & ~n28301 ;
  assign n28649 = n28640 & n28648 ;
  assign n28650 = ~n28647 & ~n28649 ;
  assign n28651 = ~n28298 & ~n28650 ;
  assign n28652 = n28295 & n28301 ;
  assign n28653 = ~n28640 & n28652 ;
  assign n28654 = n28295 & ~n28301 ;
  assign n28655 = n28640 & n28654 ;
  assign n28656 = ~n28653 & ~n28655 ;
  assign n28657 = n28298 & ~n28656 ;
  assign n28658 = ~n28651 & ~n28657 ;
  assign n28659 = ~n28640 & n28648 ;
  assign n28660 = n28640 & n28646 ;
  assign n28661 = ~n28659 & ~n28660 ;
  assign n28662 = n28298 & ~n28661 ;
  assign n28663 = n28658 & ~n28662 ;
  assign n28664 = ~n28645 & n28663 ;
  assign n28665 = ~n28271 & ~n28664 ;
  assign n28666 = n3402 & n12478 ;
  assign n28667 = ~n12475 & n28666 ;
  assign n28668 = ~n12433 & ~n12478 ;
  assign n28669 = n3402 & n28668 ;
  assign n28670 = ~n12474 & n28669 ;
  assign n28671 = \b[46]  & n3733 ;
  assign n28672 = n3730 & n28671 ;
  assign n28673 = ~\a[24]  & \b[47]  ;
  assign n28674 = n3394 & n28673 ;
  assign n28675 = ~n28672 & ~n28674 ;
  assign n28676 = \b[48]  & n3400 ;
  assign n28677 = \a[24]  & \b[47]  ;
  assign n28678 = n27626 & n28677 ;
  assign n28679 = \a[26]  & ~n28678 ;
  assign n28680 = ~n28676 & n28679 ;
  assign n28681 = n28675 & n28680 ;
  assign n28682 = ~n28670 & n28681 ;
  assign n28683 = ~n28667 & n28682 ;
  assign n28684 = ~n28676 & ~n28678 ;
  assign n28685 = n28675 & n28684 ;
  assign n28686 = ~n28670 & n28685 ;
  assign n28687 = ~n28667 & n28686 ;
  assign n28688 = ~\a[26]  & ~n28687 ;
  assign n28689 = ~n28683 & ~n28688 ;
  assign n28690 = n28266 & n28664 ;
  assign n28691 = ~n28270 & n28690 ;
  assign n28692 = n28689 & ~n28691 ;
  assign n28693 = ~n28665 & n28692 ;
  assign n28694 = n28243 & n28693 ;
  assign n28695 = ~n28689 & ~n28691 ;
  assign n28696 = ~n28665 & n28695 ;
  assign n28697 = ~n28243 & n28696 ;
  assign n28698 = ~n28694 & ~n28697 ;
  assign n28699 = ~n28664 & n28689 ;
  assign n28700 = ~n28271 & n28699 ;
  assign n28701 = n28664 & n28689 ;
  assign n28702 = n28271 & n28701 ;
  assign n28703 = ~n28700 & ~n28702 ;
  assign n28704 = ~n28243 & ~n28703 ;
  assign n28705 = ~n28664 & ~n28689 ;
  assign n28706 = ~n28271 & n28705 ;
  assign n28707 = n28664 & ~n28689 ;
  assign n28708 = n28271 & n28707 ;
  assign n28709 = ~n28706 & ~n28708 ;
  assign n28710 = n28243 & ~n28709 ;
  assign n28711 = ~n28704 & ~n28710 ;
  assign n28712 = n28698 & n28711 ;
  assign n28713 = ~n28240 & n28712 ;
  assign n28714 = ~n28223 & n28713 ;
  assign n28715 = n28240 & n28712 ;
  assign n28716 = n28223 & n28715 ;
  assign n28717 = ~n28714 & ~n28716 ;
  assign n28718 = ~n28223 & ~n28240 ;
  assign n28719 = n28215 & n28240 ;
  assign n28720 = n28222 & n28719 ;
  assign n28721 = ~n28712 & ~n28720 ;
  assign n28722 = ~n28718 & n28721 ;
  assign n28723 = n28717 & ~n28722 ;
  assign n28724 = n28040 & ~n28066 ;
  assign n28725 = n1965 & ~n16398 ;
  assign n28726 = ~n15241 & n28725 ;
  assign n28727 = ~n16404 & n28726 ;
  assign n28728 = n1965 & n16398 ;
  assign n28729 = n15241 & n28728 ;
  assign n28730 = n16400 & n28728 ;
  assign n28731 = ~n15239 & n28730 ;
  assign n28732 = ~n28729 & ~n28731 ;
  assign n28733 = ~n28727 & n28732 ;
  assign n28734 = \b[52]  & n2218 ;
  assign n28735 = n2216 & n28734 ;
  assign n28736 = ~\a[18]  & \b[53]  ;
  assign n28737 = n1957 & n28736 ;
  assign n28738 = ~n28735 & ~n28737 ;
  assign n28739 = \b[54]  & n1963 ;
  assign n28740 = \a[18]  & \b[53]  ;
  assign n28741 = n28047 & n28740 ;
  assign n28742 = \a[20]  & ~n28741 ;
  assign n28743 = ~n28739 & n28742 ;
  assign n28744 = n28738 & n28743 ;
  assign n28745 = n28733 & n28744 ;
  assign n28746 = ~n28739 & ~n28741 ;
  assign n28747 = n28738 & n28746 ;
  assign n28748 = n28733 & n28747 ;
  assign n28749 = ~\a[20]  & ~n28748 ;
  assign n28750 = ~n28745 & ~n28749 ;
  assign n28751 = ~n28061 & n28750 ;
  assign n28752 = ~n28724 & n28751 ;
  assign n28753 = n28061 & ~n28750 ;
  assign n28754 = n28040 & ~n28750 ;
  assign n28755 = ~n28066 & n28754 ;
  assign n28756 = ~n28753 & ~n28755 ;
  assign n28757 = ~n28752 & n28756 ;
  assign n28758 = ~n28723 & ~n28757 ;
  assign n28759 = n28723 & n28757 ;
  assign n28760 = ~n28758 & ~n28759 ;
  assign n28761 = ~n28208 & ~n28760 ;
  assign n28762 = ~n28183 & n28761 ;
  assign n28763 = ~n28208 & n28760 ;
  assign n28764 = n28183 & n28763 ;
  assign n28765 = ~n28762 & ~n28764 ;
  assign n28766 = ~n28161 & ~n28765 ;
  assign n28767 = n28208 & ~n28760 ;
  assign n28768 = ~n28183 & n28767 ;
  assign n28769 = n28208 & n28760 ;
  assign n28770 = n28183 & n28769 ;
  assign n28771 = ~n28768 & ~n28770 ;
  assign n28772 = n28161 & ~n28771 ;
  assign n28773 = ~n28766 & ~n28772 ;
  assign n28774 = n28183 & ~n28760 ;
  assign n28775 = ~n28183 & n28760 ;
  assign n28776 = ~n28774 & ~n28775 ;
  assign n28777 = n28208 & ~n28776 ;
  assign n28778 = ~n28161 & n28777 ;
  assign n28779 = n28183 & n28761 ;
  assign n28780 = ~n28183 & n28763 ;
  assign n28781 = ~n28779 & ~n28780 ;
  assign n28782 = n28161 & ~n28781 ;
  assign n28783 = ~n28778 & ~n28782 ;
  assign n28784 = n28773 & n28783 ;
  assign n28785 = n28078 & ~n28157 ;
  assign n28786 = ~n28108 & n28785 ;
  assign n28787 = n28102 & ~n28157 ;
  assign n28788 = ~n28786 & ~n28787 ;
  assign n28789 = n28784 & n28788 ;
  assign n28790 = ~n28158 & n28789 ;
  assign n28791 = ~n28157 & ~n28784 ;
  assign n28792 = n28139 & n28791 ;
  assign n28793 = n28157 & ~n28784 ;
  assign n28794 = ~n28139 & n28793 ;
  assign n28795 = ~n28792 & ~n28794 ;
  assign n28796 = ~n28790 & n28795 ;
  assign n28797 = ~n28136 & n28796 ;
  assign n28798 = n28116 & ~n28796 ;
  assign n28799 = ~n28118 & n28798 ;
  assign n28800 = ~n28797 & ~n28799 ;
  assign n28801 = ~n28135 & n28800 ;
  assign n28802 = ~n28127 & ~n28800 ;
  assign n28803 = ~n28131 & n28802 ;
  assign n28804 = ~n28801 & ~n28803 ;
  assign n28805 = ~n28127 & ~n28797 ;
  assign n28806 = ~n28131 & n28805 ;
  assign n28807 = ~n28784 & n28788 ;
  assign n28808 = ~n28158 & ~n28807 ;
  assign n28809 = n999 & ~n20971 ;
  assign n28810 = ~n20969 & n28809 ;
  assign n28811 = \b[61]  & n997 ;
  assign n28812 = \a[12]  & \b[60]  ;
  assign n28813 = n28195 & n28812 ;
  assign n28814 = ~n28811 & ~n28813 ;
  assign n28815 = \b[59]  & n1182 ;
  assign n28816 = n1179 & n28815 ;
  assign n28817 = ~\a[12]  & \b[60]  ;
  assign n28818 = n7674 & n28817 ;
  assign n28819 = ~n28816 & ~n28818 ;
  assign n28820 = n28814 & n28819 ;
  assign n28821 = ~n28810 & n28820 ;
  assign n28822 = ~\a[14]  & ~n28821 ;
  assign n28823 = \a[14]  & n28820 ;
  assign n28824 = ~n28810 & n28823 ;
  assign n28825 = n28181 & ~n28824 ;
  assign n28826 = n28760 & ~n28824 ;
  assign n28827 = ~n28182 & n28826 ;
  assign n28828 = ~n28825 & ~n28827 ;
  assign n28829 = ~n28822 & ~n28828 ;
  assign n28830 = ~n28182 & n28760 ;
  assign n28831 = \a[14]  & ~n28821 ;
  assign n28832 = ~\a[14]  & n28821 ;
  assign n28833 = ~n28831 & ~n28832 ;
  assign n28834 = ~n28181 & n28833 ;
  assign n28835 = ~n28830 & n28834 ;
  assign n28836 = n1965 & ~n16446 ;
  assign n28837 = ~n16444 & n28836 ;
  assign n28838 = \b[55]  & n1963 ;
  assign n28839 = \a[18]  & \b[54]  ;
  assign n28840 = n28047 & n28839 ;
  assign n28841 = ~n28838 & ~n28840 ;
  assign n28842 = \b[53]  & n2218 ;
  assign n28843 = n2216 & n28842 ;
  assign n28844 = ~\a[18]  & \b[54]  ;
  assign n28845 = n1957 & n28844 ;
  assign n28846 = ~n28843 & ~n28845 ;
  assign n28847 = n28841 & n28846 ;
  assign n28848 = ~n28837 & n28847 ;
  assign n28849 = ~\a[20]  & ~n28848 ;
  assign n28850 = \a[20]  & ~n28840 ;
  assign n28851 = ~n28838 & n28850 ;
  assign n28852 = n28846 & n28851 ;
  assign n28853 = ~n28837 & n28852 ;
  assign n28854 = ~n28849 & ~n28853 ;
  assign n28855 = n28240 & n28854 ;
  assign n28856 = n28223 & n28855 ;
  assign n28857 = ~n28712 & n28854 ;
  assign n28858 = n28223 & n28857 ;
  assign n28859 = ~n28712 & n28855 ;
  assign n28860 = ~n28858 & ~n28859 ;
  assign n28861 = ~n28856 & n28860 ;
  assign n28862 = ~n28712 & ~n28718 ;
  assign n28863 = \a[20]  & ~n28848 ;
  assign n28864 = ~\a[20]  & n28848 ;
  assign n28865 = ~n28863 & ~n28864 ;
  assign n28866 = ~n28720 & n28865 ;
  assign n28867 = ~n28862 & n28866 ;
  assign n28868 = n28861 & ~n28867 ;
  assign n28869 = n2622 & n15201 ;
  assign n28870 = ~n15198 & n28869 ;
  assign n28871 = ~n14093 & ~n15201 ;
  assign n28872 = n2622 & n28871 ;
  assign n28873 = ~n15197 & n28872 ;
  assign n28874 = \b[52]  & n2620 ;
  assign n28875 = \a[20]  & \b[51]  ;
  assign n28876 = n2910 & n28875 ;
  assign n28877 = ~\a[21]  & \b[51]  ;
  assign n28878 = n2614 & n28877 ;
  assign n28879 = ~n28876 & ~n28878 ;
  assign n28880 = ~n28874 & n28879 ;
  assign n28881 = \b[50]  & n2912 ;
  assign n28882 = n2909 & n28881 ;
  assign n28883 = \a[23]  & ~n28882 ;
  assign n28884 = n28880 & n28883 ;
  assign n28885 = ~n28873 & n28884 ;
  assign n28886 = ~n28870 & n28885 ;
  assign n28887 = n28880 & ~n28882 ;
  assign n28888 = ~n28873 & n28887 ;
  assign n28889 = ~n28870 & n28888 ;
  assign n28890 = ~\a[23]  & ~n28889 ;
  assign n28891 = ~n28886 & ~n28890 ;
  assign n28892 = n28033 & ~n28689 ;
  assign n28893 = ~n27645 & n28892 ;
  assign n28894 = n27640 & ~n28689 ;
  assign n28895 = ~n28893 & ~n28894 ;
  assign n28896 = n28891 & n28895 ;
  assign n28897 = n28698 & n28896 ;
  assign n28898 = n4249 & n11906 ;
  assign n28899 = ~n11903 & n28898 ;
  assign n28900 = n4249 & ~n11906 ;
  assign n28901 = ~n11392 & n28900 ;
  assign n28902 = ~n11902 & n28901 ;
  assign n28903 = \b[44]  & n4647 ;
  assign n28904 = n4644 & n28903 ;
  assign n28905 = ~\a[27]  & \b[45]  ;
  assign n28906 = n4241 & n28905 ;
  assign n28907 = ~n28904 & ~n28906 ;
  assign n28908 = \b[46]  & n4247 ;
  assign n28909 = \a[27]  & \b[45]  ;
  assign n28910 = n4238 & n28909 ;
  assign n28911 = \a[29]  & ~n28910 ;
  assign n28912 = ~n28908 & n28911 ;
  assign n28913 = n28907 & n28912 ;
  assign n28914 = ~n28902 & n28913 ;
  assign n28915 = ~n28899 & n28914 ;
  assign n28916 = ~n28908 & ~n28910 ;
  assign n28917 = n28907 & n28916 ;
  assign n28918 = ~n28902 & n28917 ;
  assign n28919 = ~n28899 & n28918 ;
  assign n28920 = ~\a[29]  & ~n28919 ;
  assign n28921 = ~n28915 & ~n28920 ;
  assign n28922 = n28643 & ~n28921 ;
  assign n28923 = n28298 & n28922 ;
  assign n28924 = ~n28295 & ~n28921 ;
  assign n28925 = n28643 & n28924 ;
  assign n28926 = n28298 & n28924 ;
  assign n28927 = ~n28925 & ~n28926 ;
  assign n28928 = ~n28923 & n28927 ;
  assign n28929 = ~n28295 & n28298 ;
  assign n28930 = n28921 & ~n28929 ;
  assign n28931 = n28658 & n28930 ;
  assign n28932 = ~n28301 & ~n28638 ;
  assign n28933 = ~n28639 & ~n28932 ;
  assign n28934 = n5211 & ~n10409 ;
  assign n28935 = ~n10407 & n28934 ;
  assign n28936 = \b[43]  & n5209 ;
  assign n28937 = \a[30]  & \b[42]  ;
  assign n28938 = n5200 & n28937 ;
  assign n28939 = ~n28936 & ~n28938 ;
  assign n28940 = \b[41]  & n5595 ;
  assign n28941 = n5592 & n28940 ;
  assign n28942 = ~\a[30]  & \b[42]  ;
  assign n28943 = n5203 & n28942 ;
  assign n28944 = ~n28941 & ~n28943 ;
  assign n28945 = n28939 & n28944 ;
  assign n28946 = ~n28935 & n28945 ;
  assign n28947 = ~\a[32]  & ~n28946 ;
  assign n28948 = \a[32]  & n28945 ;
  assign n28949 = ~n28935 & n28948 ;
  assign n28950 = ~n28947 & ~n28949 ;
  assign n28951 = ~n28933 & n28950 ;
  assign n28952 = ~n28639 & ~n28950 ;
  assign n28953 = ~n28932 & n28952 ;
  assign n28954 = ~n28951 & ~n28953 ;
  assign n28955 = n6309 & n9044 ;
  assign n28956 = ~n9041 & n28955 ;
  assign n28957 = n6309 & n27054 ;
  assign n28958 = ~n9040 & n28957 ;
  assign n28959 = \b[38]  & n6778 ;
  assign n28960 = n6775 & n28959 ;
  assign n28961 = ~\a[33]  & \b[39]  ;
  assign n28962 = n6301 & n28961 ;
  assign n28963 = ~n28960 & ~n28962 ;
  assign n28964 = \b[40]  & n6307 ;
  assign n28965 = \a[33]  & \b[39]  ;
  assign n28966 = n6298 & n28965 ;
  assign n28967 = \a[35]  & ~n28966 ;
  assign n28968 = ~n28964 & n28967 ;
  assign n28969 = n28963 & n28968 ;
  assign n28970 = ~n28958 & n28969 ;
  assign n28971 = ~n28956 & n28970 ;
  assign n28972 = ~n28964 & ~n28966 ;
  assign n28973 = n28963 & n28972 ;
  assign n28974 = ~n28958 & n28973 ;
  assign n28975 = ~n28956 & n28974 ;
  assign n28976 = ~\a[35]  & ~n28975 ;
  assign n28977 = ~n28971 & ~n28976 ;
  assign n28978 = n28605 & ~n28615 ;
  assign n28979 = n28610 & ~n28978 ;
  assign n28980 = ~n28463 & ~n28491 ;
  assign n28981 = ~n28464 & ~n28980 ;
  assign n28982 = ~n28326 & ~n28457 ;
  assign n28983 = ~n28458 & ~n28982 ;
  assign n28984 = ~n28328 & ~n28399 ;
  assign n28985 = ~n28398 & ~n28984 ;
  assign n28986 = n1512 & n18516 ;
  assign n28987 = ~n1509 & n28986 ;
  assign n28988 = ~n1512 & n18516 ;
  assign n28989 = ~n1228 & n28988 ;
  assign n28990 = ~n1508 & n28989 ;
  assign n28991 = \b[16]  & n18514 ;
  assign n28992 = \a[56]  & \b[15]  ;
  assign n28993 = n19181 & n28992 ;
  assign n28994 = ~\a[57]  & \b[15]  ;
  assign n28995 = n18508 & n28994 ;
  assign n28996 = ~n28993 & ~n28995 ;
  assign n28997 = ~n28991 & n28996 ;
  assign n28998 = \b[14]  & n19183 ;
  assign n28999 = n19180 & n28998 ;
  assign n29000 = \a[59]  & ~n28999 ;
  assign n29001 = n28997 & n29000 ;
  assign n29002 = ~n28990 & n29001 ;
  assign n29003 = ~n28987 & n29002 ;
  assign n29004 = n28997 & ~n28999 ;
  assign n29005 = ~n28990 & n29004 ;
  assign n29006 = ~n28987 & n29005 ;
  assign n29007 = ~\a[59]  & ~n29006 ;
  assign n29008 = ~n29003 & ~n29007 ;
  assign n29009 = \b[13]  & n20519 ;
  assign n29010 = \a[60]  & \b[12]  ;
  assign n29011 = n20510 & n29010 ;
  assign n29012 = ~n29009 & ~n29011 ;
  assign n29013 = \b[11]  & n21315 ;
  assign n29014 = n21312 & n29013 ;
  assign n29015 = ~\a[60]  & \b[12]  ;
  assign n29016 = n20513 & n29015 ;
  assign n29017 = ~n29014 & ~n29016 ;
  assign n29018 = n29012 & n29017 ;
  assign n29019 = n28380 & n28386 ;
  assign n29020 = ~n28382 & ~n29019 ;
  assign n29021 = \b[10]  & n21958 ;
  assign n29022 = \b[9]  & n21957 ;
  assign n29023 = ~n29021 & ~n29022 ;
  assign n29024 = ~n29020 & ~n29023 ;
  assign n29025 = ~n28382 & n29023 ;
  assign n29026 = ~n29019 & n29025 ;
  assign n29027 = ~\a[62]  & ~n29026 ;
  assign n29028 = ~n29024 & n29027 ;
  assign n29029 = ~n29018 & n29028 ;
  assign n29030 = ~n948 & n20521 ;
  assign n29031 = ~n908 & n20521 ;
  assign n29032 = ~n912 & n29031 ;
  assign n29033 = ~n29030 & ~n29032 ;
  assign n29034 = ~n951 & n29028 ;
  assign n29035 = ~n29033 & n29034 ;
  assign n29036 = ~n29029 & ~n29035 ;
  assign n29037 = ~n951 & ~n29033 ;
  assign n29038 = \a[62]  & ~n29026 ;
  assign n29039 = ~n29024 & n29038 ;
  assign n29040 = n29018 & n29039 ;
  assign n29041 = ~n29037 & n29040 ;
  assign n29042 = n29036 & ~n29041 ;
  assign n29043 = ~\a[62]  & ~n29018 ;
  assign n29044 = ~\a[62]  & ~n951 ;
  assign n29045 = ~n29033 & n29044 ;
  assign n29046 = ~n29043 & ~n29045 ;
  assign n29047 = ~n29024 & ~n29026 ;
  assign n29048 = \a[62]  & n29018 ;
  assign n29049 = ~n29037 & n29048 ;
  assign n29050 = ~n29047 & ~n29049 ;
  assign n29051 = n29046 & n29050 ;
  assign n29052 = n29042 & ~n29051 ;
  assign n29053 = ~n28372 & ~n28391 ;
  assign n29054 = ~n28370 & n29053 ;
  assign n29055 = ~n28393 & ~n29054 ;
  assign n29056 = n29052 & n29055 ;
  assign n29057 = ~n29052 & ~n29055 ;
  assign n29058 = ~n29056 & ~n29057 ;
  assign n29059 = n29008 & n29058 ;
  assign n29060 = ~n29008 & ~n29058 ;
  assign n29061 = ~n29059 & ~n29060 ;
  assign n29062 = ~n28985 & n29061 ;
  assign n29063 = n28985 & ~n29061 ;
  assign n29064 = ~n29062 & ~n29063 ;
  assign n29065 = ~n2076 & n16655 ;
  assign n29066 = ~n1874 & n16655 ;
  assign n29067 = ~n1878 & n29066 ;
  assign n29068 = ~n29065 & ~n29067 ;
  assign n29069 = ~n2079 & ~n29068 ;
  assign n29070 = \b[19]  & n16653 ;
  assign n29071 = \a[53]  & \b[18]  ;
  assign n29072 = n17306 & n29071 ;
  assign n29073 = ~\a[54]  & \b[18]  ;
  assign n29074 = n16647 & n29073 ;
  assign n29075 = ~n29072 & ~n29074 ;
  assign n29076 = ~n29070 & n29075 ;
  assign n29077 = \b[17]  & n17308 ;
  assign n29078 = n17305 & n29077 ;
  assign n29079 = \a[56]  & ~n29078 ;
  assign n29080 = n29076 & n29079 ;
  assign n29081 = ~n29069 & n29080 ;
  assign n29082 = n29076 & ~n29078 ;
  assign n29083 = ~\a[56]  & ~n29082 ;
  assign n29084 = ~\a[56]  & ~n2079 ;
  assign n29085 = ~n29068 & n29084 ;
  assign n29086 = ~n29083 & ~n29085 ;
  assign n29087 = ~n29081 & n29086 ;
  assign n29088 = ~n29064 & n29087 ;
  assign n29089 = n29064 & ~n29087 ;
  assign n29090 = ~n29088 & ~n29089 ;
  assign n29091 = ~n28427 & ~n28431 ;
  assign n29092 = ~n28428 & ~n29091 ;
  assign n29093 = n2768 & n14793 ;
  assign n29094 = ~n2765 & n29093 ;
  assign n29095 = n6462 & n14793 ;
  assign n29096 = ~n2764 & n29095 ;
  assign n29097 = \b[20]  & n15517 ;
  assign n29098 = n15514 & n29097 ;
  assign n29099 = \b[22]  & n14791 ;
  assign n29100 = \a[50]  & \b[21]  ;
  assign n29101 = n15515 & n29100 ;
  assign n29102 = ~\a[51]  & \b[21]  ;
  assign n29103 = n14785 & n29102 ;
  assign n29104 = ~n29101 & ~n29103 ;
  assign n29105 = ~n29099 & n29104 ;
  assign n29106 = ~n29098 & n29105 ;
  assign n29107 = ~n29096 & n29106 ;
  assign n29108 = ~n29094 & n29107 ;
  assign n29109 = ~\a[53]  & ~n29108 ;
  assign n29110 = \a[53]  & n29106 ;
  assign n29111 = ~n29096 & n29110 ;
  assign n29112 = ~n29094 & n29111 ;
  assign n29113 = ~n29109 & ~n29112 ;
  assign n29114 = n29092 & ~n29113 ;
  assign n29115 = ~n29090 & n29114 ;
  assign n29116 = ~n29092 & ~n29113 ;
  assign n29117 = n29090 & n29116 ;
  assign n29118 = ~n29115 & ~n29117 ;
  assign n29119 = ~n29092 & n29113 ;
  assign n29120 = ~n29090 & n29119 ;
  assign n29121 = n29092 & n29113 ;
  assign n29122 = n29090 & n29121 ;
  assign n29123 = ~n29120 & ~n29122 ;
  assign n29124 = n29118 & n29123 ;
  assign n29125 = ~n28983 & ~n29124 ;
  assign n29126 = n28983 & n29124 ;
  assign n29127 = ~n29125 & ~n29126 ;
  assign n29128 = ~n3564 & n13125 ;
  assign n29129 = ~n3282 & n13125 ;
  assign n29130 = ~n3560 & n29129 ;
  assign n29131 = ~n29128 & ~n29130 ;
  assign n29132 = ~n3567 & ~n29131 ;
  assign n29133 = \b[23]  & n13794 ;
  assign n29134 = n13792 & n29133 ;
  assign n29135 = ~\a[48]  & \b[24]  ;
  assign n29136 = n13117 & n29135 ;
  assign n29137 = ~n29134 & ~n29136 ;
  assign n29138 = \b[25]  & n13123 ;
  assign n29139 = \a[48]  & \b[24]  ;
  assign n29140 = n13786 & n29139 ;
  assign n29141 = \a[50]  & ~n29140 ;
  assign n29142 = ~n29138 & n29141 ;
  assign n29143 = n29137 & n29142 ;
  assign n29144 = ~n29132 & n29143 ;
  assign n29145 = ~n29138 & ~n29140 ;
  assign n29146 = n29137 & n29145 ;
  assign n29147 = ~\a[50]  & ~n29146 ;
  assign n29148 = ~\a[50]  & ~n3567 ;
  assign n29149 = ~n29131 & n29148 ;
  assign n29150 = ~n29147 & ~n29149 ;
  assign n29151 = ~n29144 & n29150 ;
  assign n29152 = ~n29127 & n29151 ;
  assign n29153 = n29127 & ~n29151 ;
  assign n29154 = ~n29152 & ~n29153 ;
  assign n29155 = ~n28981 & ~n29154 ;
  assign n29156 = n28981 & n29154 ;
  assign n29157 = ~n29155 & ~n29156 ;
  assign n29158 = n4456 & n11572 ;
  assign n29159 = ~n18723 & n29158 ;
  assign n29160 = n11572 & n16805 ;
  assign n29161 = ~n4452 & n29160 ;
  assign n29162 = \b[26]  & n12159 ;
  assign n29163 = n12156 & n29162 ;
  assign n29164 = ~\a[45]  & \b[27]  ;
  assign n29165 = n11564 & n29164 ;
  assign n29166 = ~n29163 & ~n29165 ;
  assign n29167 = \b[28]  & n11570 ;
  assign n29168 = \a[45]  & \b[27]  ;
  assign n29169 = n11561 & n29168 ;
  assign n29170 = \a[47]  & ~n29169 ;
  assign n29171 = ~n29167 & n29170 ;
  assign n29172 = n29166 & n29171 ;
  assign n29173 = ~n29161 & n29172 ;
  assign n29174 = ~n29159 & n29173 ;
  assign n29175 = ~n29167 & ~n29169 ;
  assign n29176 = n29166 & n29175 ;
  assign n29177 = ~n29161 & n29176 ;
  assign n29178 = ~n29159 & n29177 ;
  assign n29179 = ~\a[47]  & ~n29178 ;
  assign n29180 = ~n29174 & ~n29179 ;
  assign n29181 = n29157 & ~n29180 ;
  assign n29182 = ~n29157 & n29180 ;
  assign n29183 = ~n29181 & ~n29182 ;
  assign n29184 = n28496 & ~n28506 ;
  assign n29185 = n28501 & ~n29184 ;
  assign n29186 = ~n5462 & n10082 ;
  assign n29187 = ~n5460 & n29186 ;
  assign n29188 = \b[31]  & n10080 ;
  assign n29189 = \a[41]  & \b[30]  ;
  assign n29190 = n10679 & n29189 ;
  assign n29191 = ~\a[42]  & \b[30]  ;
  assign n29192 = n10074 & n29191 ;
  assign n29193 = ~n29190 & ~n29192 ;
  assign n29194 = ~n29188 & n29193 ;
  assign n29195 = \b[29]  & n10681 ;
  assign n29196 = n10678 & n29195 ;
  assign n29197 = \a[44]  & ~n29196 ;
  assign n29198 = n29194 & n29197 ;
  assign n29199 = ~n29187 & n29198 ;
  assign n29200 = n29194 & ~n29196 ;
  assign n29201 = ~n29187 & n29200 ;
  assign n29202 = ~\a[44]  & ~n29201 ;
  assign n29203 = ~n29199 & ~n29202 ;
  assign n29204 = ~n29185 & n29203 ;
  assign n29205 = ~n29183 & n29204 ;
  assign n29206 = n29185 & n29203 ;
  assign n29207 = n29183 & n29206 ;
  assign n29208 = ~n29205 & ~n29207 ;
  assign n29209 = n29185 & ~n29203 ;
  assign n29210 = ~n29183 & n29209 ;
  assign n29211 = ~n29185 & ~n29203 ;
  assign n29212 = n29183 & n29211 ;
  assign n29213 = ~n29210 & ~n29212 ;
  assign n29214 = n29208 & n29213 ;
  assign n29215 = n6565 & n8759 ;
  assign n29216 = ~n6562 & n29215 ;
  assign n29217 = ~n6565 & n8759 ;
  assign n29218 = ~n5850 & n29217 ;
  assign n29219 = ~n6561 & n29218 ;
  assign n29220 = \b[32]  & n9301 ;
  assign n29221 = n9298 & n29220 ;
  assign n29222 = ~\a[39]  & \b[33]  ;
  assign n29223 = n8751 & n29222 ;
  assign n29224 = ~n29221 & ~n29223 ;
  assign n29225 = \b[34]  & n8757 ;
  assign n29226 = \a[39]  & \b[33]  ;
  assign n29227 = n8748 & n29226 ;
  assign n29228 = \a[41]  & ~n29227 ;
  assign n29229 = ~n29225 & n29228 ;
  assign n29230 = n29224 & n29229 ;
  assign n29231 = ~n29219 & n29230 ;
  assign n29232 = ~n29216 & n29231 ;
  assign n29233 = ~n29225 & ~n29227 ;
  assign n29234 = n29224 & n29233 ;
  assign n29235 = ~n29219 & n29234 ;
  assign n29236 = ~n29216 & n29235 ;
  assign n29237 = ~\a[41]  & ~n29236 ;
  assign n29238 = ~n29232 & ~n29237 ;
  assign n29239 = n28538 & ~n28562 ;
  assign n29240 = n28533 & ~n29239 ;
  assign n29241 = ~n29238 & ~n29240 ;
  assign n29242 = n29214 & n29241 ;
  assign n29243 = ~n29238 & n29240 ;
  assign n29244 = ~n29214 & n29243 ;
  assign n29245 = ~n29242 & ~n29244 ;
  assign n29246 = n29238 & ~n29240 ;
  assign n29247 = ~n29214 & n29246 ;
  assign n29248 = n29238 & n29240 ;
  assign n29249 = n29214 & n29248 ;
  assign n29250 = ~n29247 & ~n29249 ;
  assign n29251 = n29245 & n29250 ;
  assign n29252 = n7534 & ~n7761 ;
  assign n29253 = ~n7759 & n29252 ;
  assign n29254 = \b[35]  & n7973 ;
  assign n29255 = n7970 & n29254 ;
  assign n29256 = ~\a[36]  & \b[36]  ;
  assign n29257 = n7526 & n29256 ;
  assign n29258 = ~n29255 & ~n29257 ;
  assign n29259 = \b[37]  & n7532 ;
  assign n29260 = \a[36]  & \b[36]  ;
  assign n29261 = n17801 & n29260 ;
  assign n29262 = \a[38]  & ~n29261 ;
  assign n29263 = ~n29259 & n29262 ;
  assign n29264 = n29258 & n29263 ;
  assign n29265 = ~n29253 & n29264 ;
  assign n29266 = ~n29259 & ~n29261 ;
  assign n29267 = n29258 & n29266 ;
  assign n29268 = ~n29253 & n29267 ;
  assign n29269 = ~\a[38]  & ~n29268 ;
  assign n29270 = ~n29265 & ~n29269 ;
  assign n29271 = n28567 & ~n28600 ;
  assign n29272 = n28572 & ~n29271 ;
  assign n29273 = n29270 & n29272 ;
  assign n29274 = ~n29251 & n29273 ;
  assign n29275 = n29270 & ~n29272 ;
  assign n29276 = n29251 & n29275 ;
  assign n29277 = ~n29274 & ~n29276 ;
  assign n29278 = ~n29270 & ~n29272 ;
  assign n29279 = ~n29251 & n29278 ;
  assign n29280 = ~n29270 & n29272 ;
  assign n29281 = n29251 & n29280 ;
  assign n29282 = ~n29279 & ~n29281 ;
  assign n29283 = n29277 & n29282 ;
  assign n29284 = n28979 & ~n29283 ;
  assign n29285 = ~n28979 & n29283 ;
  assign n29286 = ~n29284 & ~n29285 ;
  assign n29287 = n28977 & n29286 ;
  assign n29288 = ~n28977 & ~n29286 ;
  assign n29289 = ~n29287 & ~n29288 ;
  assign n29290 = n28954 & ~n29289 ;
  assign n29291 = ~n28954 & n29289 ;
  assign n29292 = ~n29290 & ~n29291 ;
  assign n29293 = ~n28931 & n29292 ;
  assign n29294 = n28928 & n29293 ;
  assign n29295 = ~n28928 & ~n29292 ;
  assign n29296 = n28931 & ~n29292 ;
  assign n29297 = ~n29295 & ~n29296 ;
  assign n29298 = ~n29294 & n29297 ;
  assign n29299 = n28266 & ~n28664 ;
  assign n29300 = ~n28270 & ~n29299 ;
  assign n29301 = n3402 & ~n13524 ;
  assign n29302 = ~n13522 & n29301 ;
  assign n29303 = \b[49]  & n3400 ;
  assign n29304 = \a[24]  & \b[48]  ;
  assign n29305 = n27626 & n29304 ;
  assign n29306 = ~n29303 & ~n29305 ;
  assign n29307 = \b[47]  & n3733 ;
  assign n29308 = n3730 & n29307 ;
  assign n29309 = ~\a[24]  & \b[48]  ;
  assign n29310 = n3394 & n29309 ;
  assign n29311 = ~n29308 & ~n29310 ;
  assign n29312 = n29306 & n29311 ;
  assign n29313 = ~n29302 & n29312 ;
  assign n29314 = \a[26]  & ~n29313 ;
  assign n29315 = ~\a[26]  & n29313 ;
  assign n29316 = ~n29314 & ~n29315 ;
  assign n29317 = n29300 & n29316 ;
  assign n29318 = ~\a[26]  & ~n29313 ;
  assign n29319 = \a[26]  & n29312 ;
  assign n29320 = ~n29302 & n29319 ;
  assign n29321 = ~n29318 & ~n29320 ;
  assign n29322 = ~n29300 & n29321 ;
  assign n29323 = ~n29317 & ~n29322 ;
  assign n29324 = n29298 & n29323 ;
  assign n29325 = ~n29298 & ~n29323 ;
  assign n29326 = ~n29324 & ~n29325 ;
  assign n29327 = ~n28689 & ~n28891 ;
  assign n29328 = n28243 & n29327 ;
  assign n29329 = ~n28665 & ~n28691 ;
  assign n29330 = n29327 & n29329 ;
  assign n29331 = ~n28891 & n29329 ;
  assign n29332 = n28243 & n29331 ;
  assign n29333 = ~n29330 & ~n29332 ;
  assign n29334 = ~n29328 & n29333 ;
  assign n29335 = n29326 & n29334 ;
  assign n29336 = ~n28897 & n29335 ;
  assign n29337 = n28896 & ~n29326 ;
  assign n29338 = n28698 & n29337 ;
  assign n29339 = n28698 & n28895 ;
  assign n29340 = ~n28891 & ~n29326 ;
  assign n29341 = ~n29339 & n29340 ;
  assign n29342 = ~n29338 & ~n29341 ;
  assign n29343 = ~n29336 & n29342 ;
  assign n29344 = n28868 & n29343 ;
  assign n29345 = ~n28868 & ~n29343 ;
  assign n29346 = ~n29344 & ~n29345 ;
  assign n29347 = n28752 & n28756 ;
  assign n29348 = n28723 & n28756 ;
  assign n29349 = ~n29347 & ~n29348 ;
  assign n29350 = ~n1304 & ~n17685 ;
  assign n29351 = ~n18940 & n29350 ;
  assign n29352 = ~n18936 & n29351 ;
  assign n29353 = ~n1464 & n29352 ;
  assign n29354 = n1467 & n18940 ;
  assign n29355 = ~n18937 & n29354 ;
  assign n29356 = ~n29353 & ~n29355 ;
  assign n29357 = \b[56]  & n1652 ;
  assign n29358 = n1649 & n29357 ;
  assign n29359 = ~\a[15]  & \b[57]  ;
  assign n29360 = n1459 & n29359 ;
  assign n29361 = ~n29358 & ~n29360 ;
  assign n29362 = \b[58]  & n1465 ;
  assign n29363 = \a[15]  & \b[57]  ;
  assign n29364 = n1456 & n29363 ;
  assign n29365 = \a[17]  & ~n29364 ;
  assign n29366 = ~n29362 & n29365 ;
  assign n29367 = n29361 & n29366 ;
  assign n29368 = n29356 & n29367 ;
  assign n29369 = ~n29362 & ~n29364 ;
  assign n29370 = n29361 & n29369 ;
  assign n29371 = n29356 & n29370 ;
  assign n29372 = ~\a[17]  & ~n29371 ;
  assign n29373 = ~n29368 & ~n29372 ;
  assign n29374 = n29349 & ~n29373 ;
  assign n29375 = ~n29349 & n29373 ;
  assign n29376 = ~n29374 & ~n29375 ;
  assign n29377 = n29346 & n29376 ;
  assign n29378 = ~n29346 & n29374 ;
  assign n29379 = ~n29346 & ~n29349 ;
  assign n29380 = n29373 & n29379 ;
  assign n29381 = ~n29378 & ~n29380 ;
  assign n29382 = ~n29377 & n29381 ;
  assign n29383 = ~n28835 & n29382 ;
  assign n29384 = ~n28829 & n29383 ;
  assign n29385 = ~n28829 & ~n28835 ;
  assign n29386 = ~n29382 & ~n29385 ;
  assign n29387 = ~n29384 & ~n29386 ;
  assign n29388 = \b[62]  & n796 ;
  assign n29389 = n793 & n29388 ;
  assign n29390 = ~\a[9]  & \b[63]  ;
  assign n29391 = n638 & n29390 ;
  assign n29392 = \a[9]  & \b[63]  ;
  assign n29393 = n28143 & n29392 ;
  assign n29394 = ~n29391 & ~n29393 ;
  assign n29395 = ~n29389 & n29394 ;
  assign n29396 = ~\a[11]  & ~n29395 ;
  assign n29397 = n646 & ~n22458 ;
  assign n29398 = ~\a[11]  & n29397 ;
  assign n29399 = ~n23173 & n29398 ;
  assign n29400 = ~n29396 & ~n29399 ;
  assign n29401 = ~n23173 & n29397 ;
  assign n29402 = \a[11]  & n29395 ;
  assign n29403 = ~n29401 & n29402 ;
  assign n29404 = n29400 & ~n29403 ;
  assign n29405 = ~n28208 & ~n29404 ;
  assign n29406 = n28161 & n29405 ;
  assign n29407 = n28776 & ~n29404 ;
  assign n29408 = n28161 & n29407 ;
  assign n29409 = n28776 & n29405 ;
  assign n29410 = ~n29408 & ~n29409 ;
  assign n29411 = ~n29406 & n29410 ;
  assign n29412 = n28075 & ~n28208 ;
  assign n29413 = ~n27555 & n29412 ;
  assign n29414 = n27550 & ~n28208 ;
  assign n29415 = ~n29413 & ~n29414 ;
  assign n29416 = n29404 & n29415 ;
  assign n29417 = n28773 & n29416 ;
  assign n29418 = n29411 & ~n29417 ;
  assign n29419 = n29387 & n29418 ;
  assign n29420 = ~n29387 & ~n29418 ;
  assign n29421 = ~n29419 & ~n29420 ;
  assign n29422 = n28808 & n29421 ;
  assign n29423 = ~n28808 & ~n29421 ;
  assign n29424 = ~n29422 & ~n29423 ;
  assign n29425 = ~n28799 & n29424 ;
  assign n29426 = ~n28806 & n29425 ;
  assign n29427 = ~n28799 & ~n28806 ;
  assign n29428 = ~n29424 & ~n29427 ;
  assign n29429 = ~n29426 & ~n29428 ;
  assign n29430 = ~n29422 & ~n29426 ;
  assign n29431 = ~n29387 & n29411 ;
  assign n29432 = ~n29417 & ~n29431 ;
  assign n29433 = ~n29374 & n29375 ;
  assign n29434 = ~n29346 & ~n29374 ;
  assign n29435 = ~n29433 & ~n29434 ;
  assign n29436 = n999 & n21696 ;
  assign n29437 = ~n21693 & n29436 ;
  assign n29438 = n999 & ~n21696 ;
  assign n29439 = ~n20966 & n29438 ;
  assign n29440 = ~n21692 & n29439 ;
  assign n29441 = \b[62]  & n997 ;
  assign n29442 = \a[12]  & \b[61]  ;
  assign n29443 = n28195 & n29442 ;
  assign n29444 = ~n29441 & ~n29443 ;
  assign n29445 = \b[60]  & n1182 ;
  assign n29446 = n1179 & n29445 ;
  assign n29447 = ~\a[12]  & \b[61]  ;
  assign n29448 = n7674 & n29447 ;
  assign n29449 = ~n29446 & ~n29448 ;
  assign n29450 = n29444 & n29449 ;
  assign n29451 = ~n29440 & n29450 ;
  assign n29452 = ~n29437 & n29451 ;
  assign n29453 = \a[14]  & ~n29452 ;
  assign n29454 = ~\a[14]  & n29452 ;
  assign n29455 = ~n29453 & ~n29454 ;
  assign n29456 = n29435 & n29455 ;
  assign n29457 = ~\a[14]  & ~n29452 ;
  assign n29458 = \a[14]  & n29450 ;
  assign n29459 = ~n29440 & n29458 ;
  assign n29460 = ~n29437 & n29459 ;
  assign n29461 = ~n29457 & ~n29460 ;
  assign n29462 = ~n29349 & n29461 ;
  assign n29463 = ~n29346 & n29462 ;
  assign n29464 = n29373 & n29461 ;
  assign n29465 = ~n29349 & n29464 ;
  assign n29466 = ~n29346 & n29464 ;
  assign n29467 = ~n29465 & ~n29466 ;
  assign n29468 = ~n29463 & n29467 ;
  assign n29469 = ~n28867 & ~n29343 ;
  assign n29470 = ~n28861 & ~n28867 ;
  assign n29471 = ~n29469 & ~n29470 ;
  assign n29472 = n1467 & ~n19550 ;
  assign n29473 = ~n19548 & n29472 ;
  assign n29474 = \b[59]  & n1465 ;
  assign n29475 = \a[15]  & \b[58]  ;
  assign n29476 = n1456 & n29475 ;
  assign n29477 = ~n29474 & ~n29476 ;
  assign n29478 = \b[57]  & n1652 ;
  assign n29479 = n1649 & n29478 ;
  assign n29480 = ~\a[15]  & \b[58]  ;
  assign n29481 = n1459 & n29480 ;
  assign n29482 = ~n29479 & ~n29481 ;
  assign n29483 = n29477 & n29482 ;
  assign n29484 = ~n29473 & n29483 ;
  assign n29485 = ~\a[17]  & ~n29484 ;
  assign n29486 = \a[17]  & n29483 ;
  assign n29487 = ~n29473 & n29486 ;
  assign n29488 = ~n29485 & ~n29487 ;
  assign n29489 = ~n29471 & n29488 ;
  assign n29490 = ~n29469 & ~n29488 ;
  assign n29491 = ~n29470 & n29490 ;
  assign n29492 = ~n29489 & ~n29491 ;
  assign n29493 = n28897 & n29334 ;
  assign n29494 = ~n29326 & n29334 ;
  assign n29495 = ~n29493 & ~n29494 ;
  assign n29496 = n1965 & n17647 ;
  assign n29497 = ~n17644 & n29496 ;
  assign n29498 = n1965 & ~n17647 ;
  assign n29499 = ~n16441 & n29498 ;
  assign n29500 = ~n17643 & n29499 ;
  assign n29501 = \b[56]  & n1963 ;
  assign n29502 = \a[18]  & \b[55]  ;
  assign n29503 = n28047 & n29502 ;
  assign n29504 = ~n29501 & ~n29503 ;
  assign n29505 = \b[54]  & n2218 ;
  assign n29506 = n2216 & n29505 ;
  assign n29507 = ~\a[18]  & \b[55]  ;
  assign n29508 = n1957 & n29507 ;
  assign n29509 = ~n29506 & ~n29508 ;
  assign n29510 = n29504 & n29509 ;
  assign n29511 = ~n29500 & n29510 ;
  assign n29512 = ~n29497 & n29511 ;
  assign n29513 = \a[20]  & ~n29512 ;
  assign n29514 = ~\a[20]  & n29512 ;
  assign n29515 = ~n29513 & ~n29514 ;
  assign n29516 = n29495 & n29515 ;
  assign n29517 = ~\a[20]  & ~n29512 ;
  assign n29518 = \a[20]  & n29510 ;
  assign n29519 = ~n29500 & n29518 ;
  assign n29520 = ~n29497 & n29519 ;
  assign n29521 = ~n29517 & ~n29520 ;
  assign n29522 = ~n29495 & n29521 ;
  assign n29523 = ~n29516 & ~n29522 ;
  assign n29524 = n28928 & ~n29293 ;
  assign n29525 = n3402 & n14052 ;
  assign n29526 = ~n14049 & n29525 ;
  assign n29527 = n3402 & ~n14052 ;
  assign n29528 = ~n13519 & n29527 ;
  assign n29529 = ~n14048 & n29528 ;
  assign n29530 = \b[50]  & n3400 ;
  assign n29531 = \a[24]  & \b[49]  ;
  assign n29532 = n27626 & n29531 ;
  assign n29533 = ~n29530 & ~n29532 ;
  assign n29534 = \b[48]  & n3733 ;
  assign n29535 = n3730 & n29534 ;
  assign n29536 = ~\a[24]  & \b[49]  ;
  assign n29537 = n3394 & n29536 ;
  assign n29538 = ~n29535 & ~n29537 ;
  assign n29539 = n29533 & n29538 ;
  assign n29540 = ~n29529 & n29539 ;
  assign n29541 = ~n29526 & n29540 ;
  assign n29542 = \a[26]  & ~n29541 ;
  assign n29543 = ~\a[26]  & n29541 ;
  assign n29544 = ~n29542 & ~n29543 ;
  assign n29545 = ~n29524 & n29544 ;
  assign n29546 = ~\a[26]  & ~n29541 ;
  assign n29547 = \a[26]  & n29539 ;
  assign n29548 = ~n29529 & n29547 ;
  assign n29549 = ~n29526 & n29548 ;
  assign n29550 = ~n29546 & ~n29549 ;
  assign n29551 = n28928 & n29550 ;
  assign n29552 = ~n29293 & n29551 ;
  assign n29553 = ~n29545 & ~n29552 ;
  assign n29554 = n4249 & ~n12438 ;
  assign n29555 = ~n12436 & n29554 ;
  assign n29556 = \b[47]  & n4247 ;
  assign n29557 = \a[27]  & \b[46]  ;
  assign n29558 = n4238 & n29557 ;
  assign n29559 = ~n29556 & ~n29558 ;
  assign n29560 = \b[45]  & n4647 ;
  assign n29561 = n4644 & n29560 ;
  assign n29562 = ~\a[27]  & \b[46]  ;
  assign n29563 = n4241 & n29562 ;
  assign n29564 = ~n29561 & ~n29563 ;
  assign n29565 = n29559 & n29564 ;
  assign n29566 = ~n29555 & n29565 ;
  assign n29567 = ~\a[29]  & ~n29566 ;
  assign n29568 = \a[29]  & n29565 ;
  assign n29569 = ~n29555 & n29568 ;
  assign n29570 = n28951 & ~n29569 ;
  assign n29571 = ~n28953 & ~n29569 ;
  assign n29572 = n29289 & n29571 ;
  assign n29573 = ~n29570 & ~n29572 ;
  assign n29574 = ~n29567 & ~n29573 ;
  assign n29575 = ~n28953 & n29289 ;
  assign n29576 = ~n29567 & ~n29569 ;
  assign n29577 = ~n29575 & ~n29576 ;
  assign n29578 = ~n28951 & n29577 ;
  assign n29579 = ~n29574 & ~n29578 ;
  assign n29580 = n28977 & ~n29284 ;
  assign n29581 = n5211 & ~n28007 ;
  assign n29582 = ~n28005 & n29581 ;
  assign n29583 = \b[44]  & n5209 ;
  assign n29584 = \a[30]  & \b[43]  ;
  assign n29585 = n5200 & n29584 ;
  assign n29586 = ~n29583 & ~n29585 ;
  assign n29587 = \b[42]  & n5595 ;
  assign n29588 = n5592 & n29587 ;
  assign n29589 = ~\a[30]  & \b[43]  ;
  assign n29590 = n5203 & n29589 ;
  assign n29591 = ~n29588 & ~n29590 ;
  assign n29592 = n29586 & n29591 ;
  assign n29593 = ~n29582 & n29592 ;
  assign n29594 = ~\a[32]  & ~n29593 ;
  assign n29595 = ~n29285 & n29594 ;
  assign n29596 = ~n29580 & n29595 ;
  assign n29597 = \a[32]  & n29593 ;
  assign n29598 = ~n29285 & n29597 ;
  assign n29599 = ~n29580 & n29598 ;
  assign n29600 = ~n29596 & ~n29599 ;
  assign n29601 = \a[32]  & n29592 ;
  assign n29602 = ~n29582 & n29601 ;
  assign n29603 = n29285 & ~n29602 ;
  assign n29604 = n28977 & ~n29602 ;
  assign n29605 = ~n29284 & n29604 ;
  assign n29606 = ~n29603 & ~n29605 ;
  assign n29607 = ~n29594 & ~n29606 ;
  assign n29608 = n29600 & ~n29607 ;
  assign n29609 = ~n3022 & n14793 ;
  assign n29610 = ~n3020 & n29609 ;
  assign n29611 = \b[21]  & n15517 ;
  assign n29612 = n15514 & n29611 ;
  assign n29613 = ~\a[51]  & \b[22]  ;
  assign n29614 = n14785 & n29613 ;
  assign n29615 = ~n29612 & ~n29614 ;
  assign n29616 = \b[23]  & n14791 ;
  assign n29617 = \a[51]  & \b[22]  ;
  assign n29618 = n14782 & n29617 ;
  assign n29619 = \a[53]  & ~n29618 ;
  assign n29620 = ~n29616 & n29619 ;
  assign n29621 = n29615 & n29620 ;
  assign n29622 = ~n29610 & n29621 ;
  assign n29623 = ~n29616 & ~n29618 ;
  assign n29624 = n29615 & n29623 ;
  assign n29625 = ~n29610 & n29624 ;
  assign n29626 = ~\a[53]  & ~n29625 ;
  assign n29627 = ~n29622 & ~n29626 ;
  assign n29628 = ~n1691 & n18516 ;
  assign n29629 = ~n1511 & n18516 ;
  assign n29630 = ~n1515 & n29629 ;
  assign n29631 = ~n29628 & ~n29630 ;
  assign n29632 = ~n1694 & ~n29631 ;
  assign n29633 = \b[17]  & n18514 ;
  assign n29634 = \a[56]  & \b[16]  ;
  assign n29635 = n19181 & n29634 ;
  assign n29636 = ~\a[57]  & \b[16]  ;
  assign n29637 = n18508 & n29636 ;
  assign n29638 = ~n29635 & ~n29637 ;
  assign n29639 = ~n29633 & n29638 ;
  assign n29640 = \b[15]  & n19183 ;
  assign n29641 = n19180 & n29640 ;
  assign n29642 = \a[59]  & ~n29641 ;
  assign n29643 = n29639 & n29642 ;
  assign n29644 = ~n29632 & n29643 ;
  assign n29645 = n29639 & ~n29641 ;
  assign n29646 = ~\a[59]  & ~n29645 ;
  assign n29647 = ~\a[59]  & ~n1694 ;
  assign n29648 = ~n29631 & n29647 ;
  assign n29649 = ~n29646 & ~n29648 ;
  assign n29650 = ~n29644 & n29649 ;
  assign n29651 = ~n29026 & n29042 ;
  assign n29652 = \b[11]  & n21958 ;
  assign n29653 = \b[10]  & n21957 ;
  assign n29654 = ~n29652 & ~n29653 ;
  assign n29655 = n29023 & ~n29654 ;
  assign n29656 = ~n29023 & n29654 ;
  assign n29657 = ~n29655 & ~n29656 ;
  assign n29658 = ~n29651 & n29657 ;
  assign n29659 = n1087 & n20521 ;
  assign n29660 = ~n946 & ~n1083 ;
  assign n29661 = n29659 & ~n29660 ;
  assign n29662 = n20521 & n21340 ;
  assign n29663 = ~n1083 & n29662 ;
  assign n29664 = \b[12]  & n21315 ;
  assign n29665 = n21312 & n29664 ;
  assign n29666 = ~\a[60]  & \b[13]  ;
  assign n29667 = n20513 & n29666 ;
  assign n29668 = ~n29665 & ~n29667 ;
  assign n29669 = \b[14]  & n20519 ;
  assign n29670 = \a[60]  & \b[13]  ;
  assign n29671 = n20510 & n29670 ;
  assign n29672 = \a[62]  & ~n29671 ;
  assign n29673 = ~n29669 & n29672 ;
  assign n29674 = n29668 & n29673 ;
  assign n29675 = ~n29663 & n29674 ;
  assign n29676 = ~n29661 & n29675 ;
  assign n29677 = ~n29669 & ~n29671 ;
  assign n29678 = n29668 & n29677 ;
  assign n29679 = ~n29663 & n29678 ;
  assign n29680 = ~n29661 & n29679 ;
  assign n29681 = ~\a[62]  & ~n29680 ;
  assign n29682 = ~n29676 & ~n29681 ;
  assign n29683 = ~n29026 & ~n29657 ;
  assign n29684 = n29042 & n29683 ;
  assign n29685 = ~n29682 & ~n29684 ;
  assign n29686 = ~n29658 & n29685 ;
  assign n29687 = ~n29658 & ~n29684 ;
  assign n29688 = n29682 & ~n29687 ;
  assign n29689 = ~n29686 & ~n29688 ;
  assign n29690 = n29008 & ~n29056 ;
  assign n29691 = ~n29057 & ~n29690 ;
  assign n29692 = ~n29689 & ~n29691 ;
  assign n29693 = n29650 & n29692 ;
  assign n29694 = n29689 & ~n29691 ;
  assign n29695 = ~n29650 & n29694 ;
  assign n29696 = ~n29693 & ~n29695 ;
  assign n29697 = ~n29650 & ~n29689 ;
  assign n29698 = n29691 & n29697 ;
  assign n29699 = n29689 & n29691 ;
  assign n29700 = n29650 & n29699 ;
  assign n29701 = ~n29698 & ~n29700 ;
  assign n29702 = n29696 & n29701 ;
  assign n29703 = n2293 & n16655 ;
  assign n29704 = ~n19247 & n29703 ;
  assign n29705 = n5705 & n16655 ;
  assign n29706 = ~n2289 & n29705 ;
  assign n29707 = \b[20]  & n16653 ;
  assign n29708 = \a[53]  & \b[19]  ;
  assign n29709 = n17306 & n29708 ;
  assign n29710 = ~\a[54]  & \b[19]  ;
  assign n29711 = n16647 & n29710 ;
  assign n29712 = ~n29709 & ~n29711 ;
  assign n29713 = ~n29707 & n29712 ;
  assign n29714 = \b[18]  & n17308 ;
  assign n29715 = n17305 & n29714 ;
  assign n29716 = \a[56]  & ~n29715 ;
  assign n29717 = n29713 & n29716 ;
  assign n29718 = ~n29706 & n29717 ;
  assign n29719 = ~n29704 & n29718 ;
  assign n29720 = n29713 & ~n29715 ;
  assign n29721 = ~n29706 & n29720 ;
  assign n29722 = ~n29704 & n29721 ;
  assign n29723 = ~\a[56]  & ~n29722 ;
  assign n29724 = ~n29719 & ~n29723 ;
  assign n29725 = ~n29702 & n29724 ;
  assign n29726 = n29702 & ~n29724 ;
  assign n29727 = ~n29725 & ~n29726 ;
  assign n29728 = ~n29063 & n29087 ;
  assign n29729 = ~n29062 & ~n29728 ;
  assign n29730 = n29727 & n29729 ;
  assign n29731 = ~n29727 & ~n29729 ;
  assign n29732 = ~n29730 & ~n29731 ;
  assign n29733 = n29627 & n29732 ;
  assign n29734 = ~n29627 & ~n29732 ;
  assign n29735 = ~n29733 & ~n29734 ;
  assign n29736 = n3604 & n13125 ;
  assign n29737 = ~n19292 & n29736 ;
  assign n29738 = n12021 & n13125 ;
  assign n29739 = ~n3600 & n29738 ;
  assign n29740 = \b[24]  & n13794 ;
  assign n29741 = n13792 & n29740 ;
  assign n29742 = ~\a[48]  & \b[25]  ;
  assign n29743 = n13117 & n29742 ;
  assign n29744 = ~n29741 & ~n29743 ;
  assign n29745 = \b[26]  & n13123 ;
  assign n29746 = \a[48]  & \b[25]  ;
  assign n29747 = n13786 & n29746 ;
  assign n29748 = \a[50]  & ~n29747 ;
  assign n29749 = ~n29745 & n29748 ;
  assign n29750 = n29744 & n29749 ;
  assign n29751 = ~n29739 & n29750 ;
  assign n29752 = ~n29737 & n29751 ;
  assign n29753 = ~n29745 & ~n29747 ;
  assign n29754 = n29744 & n29753 ;
  assign n29755 = ~n29739 & n29754 ;
  assign n29756 = ~n29737 & n29755 ;
  assign n29757 = ~\a[50]  & ~n29756 ;
  assign n29758 = ~n29752 & ~n29757 ;
  assign n29759 = ~n29090 & ~n29092 ;
  assign n29760 = n29090 & n29092 ;
  assign n29761 = n29113 & ~n29760 ;
  assign n29762 = ~n29759 & ~n29761 ;
  assign n29763 = ~n29758 & ~n29762 ;
  assign n29764 = ~n29735 & n29763 ;
  assign n29765 = ~n29758 & n29762 ;
  assign n29766 = n29735 & n29765 ;
  assign n29767 = ~n29764 & ~n29766 ;
  assign n29768 = n29758 & ~n29762 ;
  assign n29769 = n29735 & n29768 ;
  assign n29770 = n29758 & n29762 ;
  assign n29771 = ~n29735 & n29770 ;
  assign n29772 = ~n29769 & ~n29771 ;
  assign n29773 = n29767 & n29772 ;
  assign n29774 = ~n29126 & n29151 ;
  assign n29775 = ~n29125 & ~n29774 ;
  assign n29776 = ~n4502 & n11572 ;
  assign n29777 = ~n4500 & n29776 ;
  assign n29778 = \b[27]  & n12159 ;
  assign n29779 = n12156 & n29778 ;
  assign n29780 = ~\a[45]  & \b[28]  ;
  assign n29781 = n11564 & n29780 ;
  assign n29782 = ~n29779 & ~n29781 ;
  assign n29783 = \b[29]  & n11570 ;
  assign n29784 = \a[45]  & \b[28]  ;
  assign n29785 = n11561 & n29784 ;
  assign n29786 = \a[47]  & ~n29785 ;
  assign n29787 = ~n29783 & n29786 ;
  assign n29788 = n29782 & n29787 ;
  assign n29789 = ~n29777 & n29788 ;
  assign n29790 = ~n29783 & ~n29785 ;
  assign n29791 = n29782 & n29790 ;
  assign n29792 = ~n29777 & n29791 ;
  assign n29793 = ~\a[47]  & ~n29792 ;
  assign n29794 = ~n29789 & ~n29793 ;
  assign n29795 = ~n29775 & ~n29794 ;
  assign n29796 = n29773 & n29795 ;
  assign n29797 = n29775 & ~n29794 ;
  assign n29798 = ~n29773 & n29797 ;
  assign n29799 = ~n29796 & ~n29798 ;
  assign n29800 = ~n29775 & n29794 ;
  assign n29801 = ~n29773 & n29800 ;
  assign n29802 = n29775 & n29794 ;
  assign n29803 = n29773 & n29802 ;
  assign n29804 = ~n29801 & ~n29803 ;
  assign n29805 = n29799 & n29804 ;
  assign n29806 = ~n29156 & n29180 ;
  assign n29807 = ~n29155 & ~n29806 ;
  assign n29808 = ~n5810 & ~n9646 ;
  assign n29809 = ~n10079 & n29808 ;
  assign n29810 = n5807 & n29809 ;
  assign n29811 = n5810 & ~n9646 ;
  assign n29812 = ~n10079 & n29811 ;
  assign n29813 = ~n5807 & n29812 ;
  assign n29814 = ~n29810 & ~n29813 ;
  assign n29815 = \b[30]  & n10681 ;
  assign n29816 = n10678 & n29815 ;
  assign n29817 = \b[32]  & n10080 ;
  assign n29818 = \a[41]  & \b[31]  ;
  assign n29819 = n10679 & n29818 ;
  assign n29820 = ~\a[42]  & \b[31]  ;
  assign n29821 = n10074 & n29820 ;
  assign n29822 = ~n29819 & ~n29821 ;
  assign n29823 = ~n29817 & n29822 ;
  assign n29824 = ~n29816 & n29823 ;
  assign n29825 = n29814 & n29824 ;
  assign n29826 = ~\a[44]  & ~n29825 ;
  assign n29827 = \a[44]  & n29824 ;
  assign n29828 = n29814 & n29827 ;
  assign n29829 = ~n29826 & ~n29828 ;
  assign n29830 = ~n29807 & n29829 ;
  assign n29831 = ~n29805 & n29830 ;
  assign n29832 = n29807 & n29829 ;
  assign n29833 = n29805 & n29832 ;
  assign n29834 = ~n29831 & ~n29833 ;
  assign n29835 = ~n29807 & ~n29829 ;
  assign n29836 = n29805 & n29835 ;
  assign n29837 = n29807 & ~n29829 ;
  assign n29838 = ~n29805 & n29837 ;
  assign n29839 = ~n29836 & ~n29838 ;
  assign n29840 = n29834 & n29839 ;
  assign n29841 = ~n29183 & ~n29185 ;
  assign n29842 = n29183 & n29185 ;
  assign n29843 = n29203 & ~n29842 ;
  assign n29844 = ~n29841 & ~n29843 ;
  assign n29845 = n29840 & n29844 ;
  assign n29846 = ~n29840 & ~n29844 ;
  assign n29847 = ~n29845 & ~n29846 ;
  assign n29848 = ~n6610 & n8759 ;
  assign n29849 = ~n6608 & n29848 ;
  assign n29850 = \b[33]  & n9301 ;
  assign n29851 = n9298 & n29850 ;
  assign n29852 = ~\a[39]  & \b[34]  ;
  assign n29853 = n8751 & n29852 ;
  assign n29854 = ~n29851 & ~n29853 ;
  assign n29855 = \b[35]  & n8757 ;
  assign n29856 = \a[39]  & \b[34]  ;
  assign n29857 = n8748 & n29856 ;
  assign n29858 = \a[41]  & ~n29857 ;
  assign n29859 = ~n29855 & n29858 ;
  assign n29860 = n29854 & n29859 ;
  assign n29861 = ~n29849 & n29860 ;
  assign n29862 = ~n29855 & ~n29857 ;
  assign n29863 = n29854 & n29862 ;
  assign n29864 = ~n29849 & n29863 ;
  assign n29865 = ~\a[41]  & ~n29864 ;
  assign n29866 = ~n29861 & ~n29865 ;
  assign n29867 = ~n29847 & n29866 ;
  assign n29868 = n29847 & ~n29866 ;
  assign n29869 = ~n29867 & ~n29868 ;
  assign n29870 = n29214 & n29240 ;
  assign n29871 = n29245 & ~n29870 ;
  assign n29872 = ~n7098 & ~n7756 ;
  assign n29873 = ~n8175 & n29872 ;
  assign n29874 = ~n8171 & n29873 ;
  assign n29875 = ~n7531 & n29874 ;
  assign n29876 = n7534 & n8175 ;
  assign n29877 = ~n8172 & n29876 ;
  assign n29878 = ~n29875 & ~n29877 ;
  assign n29879 = \b[36]  & n7973 ;
  assign n29880 = n7970 & n29879 ;
  assign n29881 = ~\a[36]  & \b[37]  ;
  assign n29882 = n7526 & n29881 ;
  assign n29883 = ~n29880 & ~n29882 ;
  assign n29884 = \b[38]  & n7532 ;
  assign n29885 = \a[36]  & \b[37]  ;
  assign n29886 = n17801 & n29885 ;
  assign n29887 = \a[38]  & ~n29886 ;
  assign n29888 = ~n29884 & n29887 ;
  assign n29889 = n29883 & n29888 ;
  assign n29890 = n29878 & n29889 ;
  assign n29891 = ~n29884 & ~n29886 ;
  assign n29892 = n29883 & n29891 ;
  assign n29893 = n29878 & n29892 ;
  assign n29894 = ~\a[38]  & ~n29893 ;
  assign n29895 = ~n29890 & ~n29894 ;
  assign n29896 = n29871 & n29895 ;
  assign n29897 = ~n29869 & n29896 ;
  assign n29898 = ~n29871 & n29895 ;
  assign n29899 = n29869 & n29898 ;
  assign n29900 = ~n29897 & ~n29899 ;
  assign n29901 = ~n29871 & ~n29895 ;
  assign n29902 = ~n29869 & n29901 ;
  assign n29903 = n29871 & ~n29895 ;
  assign n29904 = n29869 & n29903 ;
  assign n29905 = ~n29902 & ~n29904 ;
  assign n29906 = n29900 & n29905 ;
  assign n29907 = n6309 & ~n9482 ;
  assign n29908 = ~n9480 & n29907 ;
  assign n29909 = \b[39]  & n6778 ;
  assign n29910 = n6775 & n29909 ;
  assign n29911 = ~\a[33]  & \b[40]  ;
  assign n29912 = n6301 & n29911 ;
  assign n29913 = ~n29910 & ~n29912 ;
  assign n29914 = \b[41]  & n6307 ;
  assign n29915 = \a[33]  & \b[40]  ;
  assign n29916 = n6298 & n29915 ;
  assign n29917 = \a[35]  & ~n29916 ;
  assign n29918 = ~n29914 & n29917 ;
  assign n29919 = n29913 & n29918 ;
  assign n29920 = ~n29908 & n29919 ;
  assign n29921 = ~n29914 & ~n29916 ;
  assign n29922 = n29913 & n29921 ;
  assign n29923 = ~n29908 & n29922 ;
  assign n29924 = ~\a[35]  & ~n29923 ;
  assign n29925 = ~n29920 & ~n29924 ;
  assign n29926 = ~n29251 & ~n29272 ;
  assign n29927 = n29251 & n29272 ;
  assign n29928 = n29270 & ~n29927 ;
  assign n29929 = ~n29926 & ~n29928 ;
  assign n29930 = n29925 & n29929 ;
  assign n29931 = ~n29906 & n29930 ;
  assign n29932 = n29925 & ~n29929 ;
  assign n29933 = n29906 & n29932 ;
  assign n29934 = ~n29931 & ~n29933 ;
  assign n29935 = ~n29925 & ~n29929 ;
  assign n29936 = ~n29906 & n29935 ;
  assign n29937 = ~n29925 & n29929 ;
  assign n29938 = n29906 & n29937 ;
  assign n29939 = ~n29936 & ~n29938 ;
  assign n29940 = n29934 & n29939 ;
  assign n29941 = n29608 & ~n29940 ;
  assign n29942 = ~n29608 & n29940 ;
  assign n29943 = ~n29941 & ~n29942 ;
  assign n29944 = n29579 & n29943 ;
  assign n29945 = ~n29579 & ~n29943 ;
  assign n29946 = ~n29944 & ~n29945 ;
  assign n29947 = n29553 & n29946 ;
  assign n29948 = ~n29553 & ~n29946 ;
  assign n29949 = ~n29947 & ~n29948 ;
  assign n29950 = ~n29298 & ~n29317 ;
  assign n29951 = ~n29317 & n29322 ;
  assign n29952 = ~n29950 & ~n29951 ;
  assign n29953 = n2622 & ~n15246 ;
  assign n29954 = ~n15244 & n29953 ;
  assign n29955 = \b[51]  & n2912 ;
  assign n29956 = n2909 & n29955 ;
  assign n29957 = \b[53]  & n2620 ;
  assign n29958 = \a[20]  & \b[52]  ;
  assign n29959 = n2910 & n29958 ;
  assign n29960 = ~\a[21]  & \b[52]  ;
  assign n29961 = n2614 & n29960 ;
  assign n29962 = ~n29959 & ~n29961 ;
  assign n29963 = ~n29957 & n29962 ;
  assign n29964 = ~n29956 & n29963 ;
  assign n29965 = ~n29954 & n29964 ;
  assign n29966 = \a[23]  & ~n29965 ;
  assign n29967 = ~\a[23]  & n29965 ;
  assign n29968 = ~n29966 & ~n29967 ;
  assign n29969 = n29952 & n29968 ;
  assign n29970 = ~\a[23]  & ~n29965 ;
  assign n29971 = \a[23]  & n29964 ;
  assign n29972 = ~n29954 & n29971 ;
  assign n29973 = ~n29970 & ~n29972 ;
  assign n29974 = ~n29952 & n29973 ;
  assign n29975 = ~n29969 & ~n29974 ;
  assign n29976 = n29949 & n29975 ;
  assign n29977 = ~n29949 & ~n29975 ;
  assign n29978 = ~n29976 & ~n29977 ;
  assign n29979 = n29523 & n29978 ;
  assign n29980 = ~n29523 & ~n29978 ;
  assign n29981 = ~n29979 & ~n29980 ;
  assign n29982 = n29492 & n29981 ;
  assign n29983 = ~n29492 & ~n29981 ;
  assign n29984 = ~n29982 & ~n29983 ;
  assign n29985 = n29468 & n29984 ;
  assign n29986 = ~n29456 & n29985 ;
  assign n29987 = ~n29456 & n29468 ;
  assign n29988 = ~n29984 & ~n29987 ;
  assign n29989 = ~n29986 & ~n29988 ;
  assign n29990 = n28829 & ~n28835 ;
  assign n29991 = ~n28835 & ~n29382 ;
  assign n29992 = \b[63]  & n646 ;
  assign n29993 = ~n21694 & n29992 ;
  assign n29994 = ~n23171 & n29993 ;
  assign n29995 = \a[8]  & \a[10]  ;
  assign n29996 = \a[9]  & ~\a[11]  ;
  assign n29997 = n29995 & n29996 ;
  assign n29998 = ~\a[8]  & ~\a[10]  ;
  assign n29999 = ~\a[9]  & \a[11]  ;
  assign n30000 = n29998 & n29999 ;
  assign n30001 = ~n29997 & ~n30000 ;
  assign n30002 = \b[63]  & ~n30001 ;
  assign n30003 = \a[11]  & ~n30002 ;
  assign n30004 = ~n29994 & n30003 ;
  assign n30005 = ~n29994 & ~n30002 ;
  assign n30006 = ~\a[11]  & ~n30005 ;
  assign n30007 = ~n30004 & ~n30006 ;
  assign n30008 = ~n29991 & ~n30007 ;
  assign n30009 = ~n29990 & n30008 ;
  assign n30010 = n29991 & n30007 ;
  assign n30011 = ~n28835 & n30007 ;
  assign n30012 = n28829 & n30011 ;
  assign n30013 = ~n30010 & ~n30012 ;
  assign n30014 = ~n30009 & n30013 ;
  assign n30015 = n29989 & n30014 ;
  assign n30016 = ~n29989 & ~n30014 ;
  assign n30017 = ~n30015 & ~n30016 ;
  assign n30018 = n29432 & n30017 ;
  assign n30019 = ~n29432 & ~n30017 ;
  assign n30020 = ~n30018 & ~n30019 ;
  assign n30021 = ~n29430 & n30020 ;
  assign n30022 = ~n29422 & ~n30020 ;
  assign n30023 = ~n29426 & n30022 ;
  assign n30024 = ~n30021 & ~n30023 ;
  assign n30025 = ~n29422 & ~n30018 ;
  assign n30026 = ~n29426 & n30025 ;
  assign n30027 = ~n29989 & ~n30009 ;
  assign n30028 = ~n30009 & ~n30013 ;
  assign n30029 = ~n30027 & ~n30028 ;
  assign n30030 = ~n29491 & ~n29981 ;
  assign n30031 = n29470 & n29488 ;
  assign n30032 = n29469 & n29488 ;
  assign n30033 = ~n30031 & ~n30032 ;
  assign n30034 = ~n30030 & n30033 ;
  assign n30035 = n1467 & n20260 ;
  assign n30036 = ~n20257 & n30035 ;
  assign n30037 = n1467 & ~n20260 ;
  assign n30038 = ~n19545 & n30037 ;
  assign n30039 = ~n20256 & n30038 ;
  assign n30040 = \b[58]  & n1652 ;
  assign n30041 = n1649 & n30040 ;
  assign n30042 = ~\a[15]  & \b[59]  ;
  assign n30043 = n1459 & n30042 ;
  assign n30044 = ~n30041 & ~n30043 ;
  assign n30045 = \b[60]  & n1465 ;
  assign n30046 = \a[15]  & \b[59]  ;
  assign n30047 = n1456 & n30046 ;
  assign n30048 = \a[17]  & ~n30047 ;
  assign n30049 = ~n30045 & n30048 ;
  assign n30050 = n30044 & n30049 ;
  assign n30051 = ~n30039 & n30050 ;
  assign n30052 = ~n30036 & n30051 ;
  assign n30053 = ~n30045 & ~n30047 ;
  assign n30054 = n30044 & n30053 ;
  assign n30055 = ~n30039 & n30054 ;
  assign n30056 = ~n30036 & n30055 ;
  assign n30057 = ~\a[17]  & ~n30056 ;
  assign n30058 = ~n30052 & ~n30057 ;
  assign n30059 = n1965 & ~n17690 ;
  assign n30060 = ~n17688 & n30059 ;
  assign n30061 = \b[57]  & n1963 ;
  assign n30062 = \a[18]  & \b[56]  ;
  assign n30063 = n28047 & n30062 ;
  assign n30064 = ~n30061 & ~n30063 ;
  assign n30065 = \b[55]  & n2218 ;
  assign n30066 = n2216 & n30065 ;
  assign n30067 = ~\a[18]  & \b[56]  ;
  assign n30068 = n1957 & n30067 ;
  assign n30069 = ~n30066 & ~n30068 ;
  assign n30070 = n30064 & n30069 ;
  assign n30071 = ~n30060 & n30070 ;
  assign n30072 = ~\a[20]  & ~n30071 ;
  assign n30073 = \a[20]  & n30070 ;
  assign n30074 = ~n30060 & n30073 ;
  assign n30075 = ~n30072 & ~n30074 ;
  assign n30076 = ~n29516 & ~n29978 ;
  assign n30077 = ~n29516 & n29522 ;
  assign n30078 = ~n30076 & ~n30077 ;
  assign n30079 = n30075 & ~n30078 ;
  assign n30080 = n29978 & ~n30075 ;
  assign n30081 = ~n29522 & n30080 ;
  assign n30082 = n29516 & ~n30075 ;
  assign n30083 = ~n30081 & ~n30082 ;
  assign n30084 = n3402 & ~n14098 ;
  assign n30085 = ~n14096 & n30084 ;
  assign n30086 = \b[51]  & n3400 ;
  assign n30087 = \a[24]  & \b[50]  ;
  assign n30088 = n27626 & n30087 ;
  assign n30089 = ~n30086 & ~n30088 ;
  assign n30090 = \b[49]  & n3733 ;
  assign n30091 = n3730 & n30090 ;
  assign n30092 = ~\a[24]  & \b[50]  ;
  assign n30093 = n3394 & n30092 ;
  assign n30094 = ~n30091 & ~n30093 ;
  assign n30095 = n30089 & n30094 ;
  assign n30096 = ~n30085 & n30095 ;
  assign n30097 = ~\a[26]  & ~n30096 ;
  assign n30098 = \a[26]  & n30095 ;
  assign n30099 = ~n30085 & n30098 ;
  assign n30100 = ~n30097 & ~n30099 ;
  assign n30101 = ~n29545 & ~n29946 ;
  assign n30102 = ~n29545 & n29552 ;
  assign n30103 = ~n30101 & ~n30102 ;
  assign n30104 = n30100 & ~n30103 ;
  assign n30105 = ~n29552 & ~n30100 ;
  assign n30106 = n29946 & n30105 ;
  assign n30107 = n29545 & ~n30100 ;
  assign n30108 = ~n30106 & ~n30107 ;
  assign n30109 = ~n30104 & n30108 ;
  assign n30110 = ~n29578 & ~n29943 ;
  assign n30111 = n29575 & n29576 ;
  assign n30112 = n28951 & n29576 ;
  assign n30113 = ~n30111 & ~n30112 ;
  assign n30114 = ~n30110 & n30113 ;
  assign n30115 = n29600 & n29940 ;
  assign n30116 = n5211 & ~n11397 ;
  assign n30117 = ~n11395 & n30116 ;
  assign n30118 = \b[45]  & n5209 ;
  assign n30119 = \a[30]  & \b[44]  ;
  assign n30120 = n5200 & n30119 ;
  assign n30121 = ~n30118 & ~n30120 ;
  assign n30122 = \b[43]  & n5595 ;
  assign n30123 = n5592 & n30122 ;
  assign n30124 = ~\a[30]  & \b[44]  ;
  assign n30125 = n5203 & n30124 ;
  assign n30126 = ~n30123 & ~n30125 ;
  assign n30127 = n30121 & n30126 ;
  assign n30128 = ~n30117 & n30127 ;
  assign n30129 = ~\a[32]  & ~n30128 ;
  assign n30130 = \a[32]  & n30127 ;
  assign n30131 = ~n30117 & n30130 ;
  assign n30132 = ~n30129 & ~n30131 ;
  assign n30133 = ~n29607 & ~n30132 ;
  assign n30134 = ~n30115 & n30133 ;
  assign n30135 = ~n29607 & ~n30115 ;
  assign n30136 = n30132 & ~n30135 ;
  assign n30137 = ~n30134 & ~n30136 ;
  assign n30138 = n4249 & n12478 ;
  assign n30139 = ~n12475 & n30138 ;
  assign n30140 = n4249 & n28668 ;
  assign n30141 = ~n12474 & n30140 ;
  assign n30142 = \b[46]  & n4647 ;
  assign n30143 = n4644 & n30142 ;
  assign n30144 = ~\a[27]  & \b[47]  ;
  assign n30145 = n4241 & n30144 ;
  assign n30146 = ~n30143 & ~n30145 ;
  assign n30147 = \b[48]  & n4247 ;
  assign n30148 = \a[27]  & \b[47]  ;
  assign n30149 = n4238 & n30148 ;
  assign n30150 = \a[29]  & ~n30149 ;
  assign n30151 = ~n30147 & n30150 ;
  assign n30152 = n30146 & n30151 ;
  assign n30153 = ~n30141 & n30152 ;
  assign n30154 = ~n30139 & n30153 ;
  assign n30155 = ~n30147 & ~n30149 ;
  assign n30156 = n30146 & n30155 ;
  assign n30157 = ~n30141 & n30156 ;
  assign n30158 = ~n30139 & n30157 ;
  assign n30159 = ~\a[29]  & ~n30158 ;
  assign n30160 = ~n30154 & ~n30159 ;
  assign n30161 = n6309 & n9930 ;
  assign n30162 = ~n9927 & n30161 ;
  assign n30163 = n6309 & ~n9930 ;
  assign n30164 = ~n9477 & n30163 ;
  assign n30165 = ~n9926 & n30164 ;
  assign n30166 = \b[40]  & n6778 ;
  assign n30167 = n6775 & n30166 ;
  assign n30168 = ~\a[33]  & \b[41]  ;
  assign n30169 = n6301 & n30168 ;
  assign n30170 = ~n30167 & ~n30169 ;
  assign n30171 = \b[42]  & n6307 ;
  assign n30172 = \a[33]  & \b[41]  ;
  assign n30173 = n6298 & n30172 ;
  assign n30174 = \a[35]  & ~n30173 ;
  assign n30175 = ~n30171 & n30174 ;
  assign n30176 = n30170 & n30175 ;
  assign n30177 = ~n30165 & n30176 ;
  assign n30178 = ~n30162 & n30177 ;
  assign n30179 = ~n30171 & ~n30173 ;
  assign n30180 = n30170 & n30179 ;
  assign n30181 = ~n30165 & n30180 ;
  assign n30182 = ~n30162 & n30181 ;
  assign n30183 = ~\a[35]  & ~n30182 ;
  assign n30184 = ~n30178 & ~n30183 ;
  assign n30185 = n29869 & ~n29871 ;
  assign n30186 = n29905 & ~n30185 ;
  assign n30187 = n3283 & n14793 ;
  assign n30188 = ~n3280 & n30187 ;
  assign n30189 = ~n3017 & ~n3283 ;
  assign n30190 = n14793 & n30189 ;
  assign n30191 = ~n3279 & n30190 ;
  assign n30192 = \b[22]  & n15517 ;
  assign n30193 = n15514 & n30192 ;
  assign n30194 = ~\a[51]  & \b[23]  ;
  assign n30195 = n14785 & n30194 ;
  assign n30196 = ~n30193 & ~n30195 ;
  assign n30197 = \b[24]  & n14791 ;
  assign n30198 = \a[51]  & \b[23]  ;
  assign n30199 = n14782 & n30198 ;
  assign n30200 = \a[53]  & ~n30199 ;
  assign n30201 = ~n30197 & n30200 ;
  assign n30202 = n30196 & n30201 ;
  assign n30203 = ~n30191 & n30202 ;
  assign n30204 = ~n30188 & n30203 ;
  assign n30205 = ~n30197 & ~n30199 ;
  assign n30206 = n30196 & n30205 ;
  assign n30207 = ~n30191 & n30206 ;
  assign n30208 = ~n30188 & n30207 ;
  assign n30209 = ~\a[53]  & ~n30208 ;
  assign n30210 = ~n30204 & ~n30209 ;
  assign n30211 = n29650 & ~n29689 ;
  assign n30212 = ~n29691 & n30211 ;
  assign n30213 = ~n29650 & n29689 ;
  assign n30214 = ~n29691 & n30213 ;
  assign n30215 = ~n30212 & ~n30214 ;
  assign n30216 = n29701 & n29724 ;
  assign n30217 = n30215 & ~n30216 ;
  assign n30218 = ~n2520 & n16655 ;
  assign n30219 = ~n2292 & n16655 ;
  assign n30220 = ~n2516 & n30219 ;
  assign n30221 = ~n30218 & ~n30220 ;
  assign n30222 = ~n2523 & ~n30221 ;
  assign n30223 = \b[19]  & n17308 ;
  assign n30224 = n17305 & n30223 ;
  assign n30225 = \b[21]  & n16653 ;
  assign n30226 = \a[54]  & \b[20]  ;
  assign n30227 = n16644 & n30226 ;
  assign n30228 = ~\a[54]  & \b[20]  ;
  assign n30229 = n16647 & n30228 ;
  assign n30230 = ~n30227 & ~n30229 ;
  assign n30231 = ~n30225 & n30230 ;
  assign n30232 = ~n30224 & n30231 ;
  assign n30233 = ~\a[56]  & n30232 ;
  assign n30234 = ~n30222 & n30233 ;
  assign n30235 = \a[56]  & ~n30232 ;
  assign n30236 = \a[56]  & ~n2523 ;
  assign n30237 = ~n30221 & n30236 ;
  assign n30238 = ~n30235 & ~n30237 ;
  assign n30239 = ~n30234 & n30238 ;
  assign n30240 = n1875 & n18516 ;
  assign n30241 = ~n1872 & n30240 ;
  assign n30242 = n5000 & n18516 ;
  assign n30243 = ~n1871 & n30242 ;
  assign n30244 = \b[16]  & n19183 ;
  assign n30245 = n19180 & n30244 ;
  assign n30246 = \b[18]  & n18514 ;
  assign n30247 = \a[56]  & \b[17]  ;
  assign n30248 = n19181 & n30247 ;
  assign n30249 = ~\a[57]  & \b[17]  ;
  assign n30250 = n18508 & n30249 ;
  assign n30251 = ~n30248 & ~n30250 ;
  assign n30252 = ~n30246 & n30251 ;
  assign n30253 = ~n30245 & n30252 ;
  assign n30254 = ~n30243 & n30253 ;
  assign n30255 = ~n30241 & n30254 ;
  assign n30256 = ~\a[59]  & ~n30255 ;
  assign n30257 = \a[59]  & n30253 ;
  assign n30258 = ~n30243 & n30257 ;
  assign n30259 = ~n30241 & n30258 ;
  assign n30260 = ~n30256 & ~n30259 ;
  assign n30261 = \b[15]  & n20519 ;
  assign n30262 = \a[60]  & \b[14]  ;
  assign n30263 = n20510 & n30262 ;
  assign n30264 = ~n30261 & ~n30263 ;
  assign n30265 = \b[13]  & n21315 ;
  assign n30266 = n21312 & n30265 ;
  assign n30267 = ~\a[60]  & \b[14]  ;
  assign n30268 = n20513 & n30267 ;
  assign n30269 = ~n30266 & ~n30268 ;
  assign n30270 = n30264 & n30269 ;
  assign n30271 = ~\a[62]  & ~n30270 ;
  assign n30272 = ~n1230 & n20521 ;
  assign n30273 = ~n1086 & n20521 ;
  assign n30274 = ~n1226 & n30273 ;
  assign n30275 = ~n30272 & ~n30274 ;
  assign n30276 = ~\a[62]  & ~n1233 ;
  assign n30277 = ~n30275 & n30276 ;
  assign n30278 = ~n30271 & ~n30277 ;
  assign n30279 = n2648 & n21957 ;
  assign n30280 = n2832 & n21958 ;
  assign n30281 = ~n30279 & ~n30280 ;
  assign n30282 = \a[11]  & ~n29022 ;
  assign n30283 = ~n29021 & n30282 ;
  assign n30284 = n30281 & ~n30283 ;
  assign n30285 = \b[12]  & n21958 ;
  assign n30286 = \b[11]  & n21957 ;
  assign n30287 = ~n30285 & ~n30286 ;
  assign n30288 = ~n30284 & ~n30287 ;
  assign n30289 = n30284 & n30287 ;
  assign n30290 = ~n30288 & ~n30289 ;
  assign n30291 = ~n1233 & ~n30275 ;
  assign n30292 = \a[62]  & n30270 ;
  assign n30293 = ~n30291 & n30292 ;
  assign n30294 = n30290 & ~n30293 ;
  assign n30295 = n30278 & n30294 ;
  assign n30296 = ~n29026 & ~n29655 ;
  assign n30297 = n29042 & n30296 ;
  assign n30298 = ~n29656 & ~n30297 ;
  assign n30299 = ~\a[62]  & ~n30287 ;
  assign n30300 = ~n30284 & n30299 ;
  assign n30301 = ~\a[62]  & n30287 ;
  assign n30302 = n30284 & n30301 ;
  assign n30303 = ~n30300 & ~n30302 ;
  assign n30304 = ~n30270 & ~n30303 ;
  assign n30305 = ~n1233 & ~n30303 ;
  assign n30306 = ~n30275 & n30305 ;
  assign n30307 = ~n30304 & ~n30306 ;
  assign n30308 = \a[62]  & ~n30287 ;
  assign n30309 = ~n30284 & n30308 ;
  assign n30310 = \a[62]  & n30287 ;
  assign n30311 = n30284 & n30310 ;
  assign n30312 = ~n30309 & ~n30311 ;
  assign n30313 = n30270 & ~n30312 ;
  assign n30314 = ~n30291 & n30313 ;
  assign n30315 = n30307 & ~n30314 ;
  assign n30316 = n30298 & n30315 ;
  assign n30317 = ~n30295 & n30316 ;
  assign n30318 = ~n30295 & n30315 ;
  assign n30319 = ~n30298 & ~n30318 ;
  assign n30320 = ~n30317 & ~n30319 ;
  assign n30321 = ~n30260 & n30320 ;
  assign n30322 = n30260 & ~n30320 ;
  assign n30323 = ~n30321 & ~n30322 ;
  assign n30324 = ~n29644 & ~n29686 ;
  assign n30325 = n29649 & n30324 ;
  assign n30326 = ~n29688 & ~n30325 ;
  assign n30327 = ~n30323 & ~n30326 ;
  assign n30328 = n30323 & n30326 ;
  assign n30329 = ~n30327 & ~n30328 ;
  assign n30330 = ~n30239 & ~n30329 ;
  assign n30331 = n30239 & n30329 ;
  assign n30332 = ~n30330 & ~n30331 ;
  assign n30333 = n30217 & n30332 ;
  assign n30334 = ~n30217 & n30330 ;
  assign n30335 = ~n30217 & n30329 ;
  assign n30336 = n30239 & n30335 ;
  assign n30337 = ~n30334 & ~n30336 ;
  assign n30338 = ~n30333 & n30337 ;
  assign n30339 = ~n30210 & n30338 ;
  assign n30340 = n30210 & ~n30338 ;
  assign n30341 = ~n30339 & ~n30340 ;
  assign n30342 = ~n4145 & n13125 ;
  assign n30343 = ~n3603 & n13125 ;
  assign n30344 = ~n4141 & n30343 ;
  assign n30345 = ~n30342 & ~n30344 ;
  assign n30346 = ~n4148 & ~n30345 ;
  assign n30347 = \b[25]  & n13794 ;
  assign n30348 = n13792 & n30347 ;
  assign n30349 = ~\a[48]  & \b[26]  ;
  assign n30350 = n13117 & n30349 ;
  assign n30351 = ~n30348 & ~n30350 ;
  assign n30352 = \b[27]  & n13123 ;
  assign n30353 = \a[48]  & \b[26]  ;
  assign n30354 = n13786 & n30353 ;
  assign n30355 = \a[50]  & ~n30354 ;
  assign n30356 = ~n30352 & n30355 ;
  assign n30357 = n30351 & n30356 ;
  assign n30358 = ~n30346 & n30357 ;
  assign n30359 = ~n30352 & ~n30354 ;
  assign n30360 = n30351 & n30359 ;
  assign n30361 = ~\a[50]  & ~n30360 ;
  assign n30362 = ~\a[50]  & ~n4148 ;
  assign n30363 = ~n30345 & n30362 ;
  assign n30364 = ~n30361 & ~n30363 ;
  assign n30365 = ~n30358 & n30364 ;
  assign n30366 = n29627 & ~n29730 ;
  assign n30367 = ~n29731 & ~n30366 ;
  assign n30368 = ~n30365 & n30367 ;
  assign n30369 = ~n30341 & n30368 ;
  assign n30370 = ~n30365 & ~n30367 ;
  assign n30371 = n30341 & n30370 ;
  assign n30372 = ~n30369 & ~n30371 ;
  assign n30373 = n30365 & ~n30367 ;
  assign n30374 = ~n30341 & n30373 ;
  assign n30375 = n30365 & n30367 ;
  assign n30376 = n30341 & n30375 ;
  assign n30377 = ~n30374 & ~n30376 ;
  assign n30378 = n30372 & n30377 ;
  assign n30379 = ~n29735 & n29762 ;
  assign n30380 = n29767 & ~n30379 ;
  assign n30381 = ~n5105 & ~n10988 ;
  assign n30382 = ~n11569 & n30381 ;
  assign n30383 = n5102 & n30382 ;
  assign n30384 = n5105 & ~n10988 ;
  assign n30385 = ~n11569 & n30384 ;
  assign n30386 = ~n5102 & n30385 ;
  assign n30387 = ~n30383 & ~n30386 ;
  assign n30388 = \b[28]  & n12159 ;
  assign n30389 = n12156 & n30388 ;
  assign n30390 = ~\a[45]  & \b[29]  ;
  assign n30391 = n11564 & n30390 ;
  assign n30392 = ~n30389 & ~n30391 ;
  assign n30393 = \b[30]  & n11570 ;
  assign n30394 = \a[45]  & \b[29]  ;
  assign n30395 = n11561 & n30394 ;
  assign n30396 = \a[47]  & ~n30395 ;
  assign n30397 = ~n30393 & n30396 ;
  assign n30398 = n30392 & n30397 ;
  assign n30399 = n30387 & n30398 ;
  assign n30400 = ~n30393 & ~n30395 ;
  assign n30401 = n30392 & n30400 ;
  assign n30402 = n30387 & n30401 ;
  assign n30403 = ~\a[47]  & ~n30402 ;
  assign n30404 = ~n30399 & ~n30403 ;
  assign n30405 = n30380 & n30404 ;
  assign n30406 = ~n30378 & n30405 ;
  assign n30407 = ~n30380 & n30404 ;
  assign n30408 = n30378 & n30407 ;
  assign n30409 = ~n30406 & ~n30408 ;
  assign n30410 = ~n30380 & ~n30404 ;
  assign n30411 = ~n30378 & n30410 ;
  assign n30412 = n30380 & ~n30404 ;
  assign n30413 = n30378 & n30412 ;
  assign n30414 = ~n30411 & ~n30413 ;
  assign n30415 = n30409 & n30414 ;
  assign n30416 = ~n5855 & n10082 ;
  assign n30417 = ~n5853 & n30416 ;
  assign n30418 = \b[31]  & n10681 ;
  assign n30419 = n10678 & n30418 ;
  assign n30420 = \b[33]  & n10080 ;
  assign n30421 = \a[41]  & \b[32]  ;
  assign n30422 = n10679 & n30421 ;
  assign n30423 = ~\a[42]  & \b[32]  ;
  assign n30424 = n10074 & n30423 ;
  assign n30425 = ~n30422 & ~n30424 ;
  assign n30426 = ~n30420 & n30425 ;
  assign n30427 = ~n30419 & n30426 ;
  assign n30428 = ~\a[44]  & n30427 ;
  assign n30429 = ~n30417 & n30428 ;
  assign n30430 = ~n30417 & n30427 ;
  assign n30431 = \a[44]  & ~n30430 ;
  assign n30432 = ~n30429 & ~n30431 ;
  assign n30433 = ~n29773 & ~n29775 ;
  assign n30434 = n29773 & n29775 ;
  assign n30435 = n29794 & ~n30434 ;
  assign n30436 = ~n30433 & ~n30435 ;
  assign n30437 = n30432 & ~n30436 ;
  assign n30438 = n30415 & n30437 ;
  assign n30439 = n30432 & n30436 ;
  assign n30440 = ~n30415 & n30439 ;
  assign n30441 = ~n30438 & ~n30440 ;
  assign n30442 = ~n30432 & ~n30436 ;
  assign n30443 = ~n30415 & n30442 ;
  assign n30444 = ~n30432 & n30436 ;
  assign n30445 = n30415 & n30444 ;
  assign n30446 = ~n30443 & ~n30445 ;
  assign n30447 = n30441 & n30446 ;
  assign n30448 = n7337 & n8759 ;
  assign n30449 = ~n7334 & n30448 ;
  assign n30450 = n8759 & n24138 ;
  assign n30451 = ~n7333 & n30450 ;
  assign n30452 = \b[34]  & n9301 ;
  assign n30453 = n9298 & n30452 ;
  assign n30454 = ~\a[39]  & \b[35]  ;
  assign n30455 = n8751 & n30454 ;
  assign n30456 = ~n30453 & ~n30455 ;
  assign n30457 = \b[36]  & n8757 ;
  assign n30458 = \a[39]  & \b[35]  ;
  assign n30459 = n8748 & n30458 ;
  assign n30460 = \a[41]  & ~n30459 ;
  assign n30461 = ~n30457 & n30460 ;
  assign n30462 = n30456 & n30461 ;
  assign n30463 = ~n30451 & n30462 ;
  assign n30464 = ~n30449 & n30463 ;
  assign n30465 = ~n30457 & ~n30459 ;
  assign n30466 = n30456 & n30465 ;
  assign n30467 = ~n30451 & n30466 ;
  assign n30468 = ~n30449 & n30467 ;
  assign n30469 = ~\a[41]  & ~n30468 ;
  assign n30470 = ~n30464 & ~n30469 ;
  assign n30471 = n29805 & n29807 ;
  assign n30472 = n29839 & ~n30471 ;
  assign n30473 = ~n30470 & ~n30472 ;
  assign n30474 = ~n30447 & n30473 ;
  assign n30475 = ~n30470 & n30472 ;
  assign n30476 = n30447 & n30475 ;
  assign n30477 = ~n30474 & ~n30476 ;
  assign n30478 = n30470 & n30472 ;
  assign n30479 = ~n30447 & n30478 ;
  assign n30480 = n30470 & ~n30472 ;
  assign n30481 = n30447 & n30480 ;
  assign n30482 = ~n30479 & ~n30481 ;
  assign n30483 = n30477 & n30482 ;
  assign n30484 = ~n29845 & n29866 ;
  assign n30485 = ~n29846 & ~n30484 ;
  assign n30486 = n7534 & ~n8602 ;
  assign n30487 = ~n8600 & n30486 ;
  assign n30488 = \b[39]  & n7532 ;
  assign n30489 = \a[36]  & \b[38]  ;
  assign n30490 = n17801 & n30489 ;
  assign n30491 = ~n30488 & ~n30490 ;
  assign n30492 = \b[37]  & n7973 ;
  assign n30493 = n7970 & n30492 ;
  assign n30494 = ~\a[36]  & \b[38]  ;
  assign n30495 = n7526 & n30494 ;
  assign n30496 = ~n30493 & ~n30495 ;
  assign n30497 = n30491 & n30496 ;
  assign n30498 = ~n30487 & n30497 ;
  assign n30499 = ~\a[38]  & ~n30498 ;
  assign n30500 = \a[38]  & n30497 ;
  assign n30501 = ~n30487 & n30500 ;
  assign n30502 = ~n30499 & ~n30501 ;
  assign n30503 = ~n30485 & ~n30502 ;
  assign n30504 = n30483 & n30503 ;
  assign n30505 = n30485 & ~n30502 ;
  assign n30506 = ~n30483 & n30505 ;
  assign n30507 = ~n30504 & ~n30506 ;
  assign n30508 = ~n30485 & n30502 ;
  assign n30509 = ~n30483 & n30508 ;
  assign n30510 = n30485 & n30502 ;
  assign n30511 = n30483 & n30510 ;
  assign n30512 = ~n30509 & ~n30511 ;
  assign n30513 = n30507 & n30512 ;
  assign n30514 = ~n30186 & n30513 ;
  assign n30515 = n30186 & ~n30513 ;
  assign n30516 = ~n30514 & ~n30515 ;
  assign n30517 = ~n30184 & n30516 ;
  assign n30518 = n30184 & ~n30516 ;
  assign n30519 = ~n30517 & ~n30518 ;
  assign n30520 = ~n29906 & ~n29929 ;
  assign n30521 = n29906 & n29929 ;
  assign n30522 = n29925 & ~n30521 ;
  assign n30523 = ~n30520 & ~n30522 ;
  assign n30524 = ~n30519 & ~n30523 ;
  assign n30525 = n30519 & n30523 ;
  assign n30526 = ~n30524 & ~n30525 ;
  assign n30527 = ~n30160 & n30526 ;
  assign n30528 = ~n30137 & n30527 ;
  assign n30529 = ~n30160 & ~n30526 ;
  assign n30530 = n30137 & n30529 ;
  assign n30531 = ~n30528 & ~n30530 ;
  assign n30532 = ~n30114 & ~n30531 ;
  assign n30533 = n30160 & n30526 ;
  assign n30534 = ~n30137 & n30533 ;
  assign n30535 = n30160 & ~n30526 ;
  assign n30536 = n30137 & n30535 ;
  assign n30537 = ~n30534 & ~n30536 ;
  assign n30538 = n30114 & ~n30537 ;
  assign n30539 = ~n30532 & ~n30538 ;
  assign n30540 = n30137 & n30526 ;
  assign n30541 = ~n30137 & ~n30526 ;
  assign n30542 = ~n30540 & ~n30541 ;
  assign n30543 = ~n30114 & n30160 ;
  assign n30544 = ~n30542 & n30543 ;
  assign n30545 = ~n30137 & n30529 ;
  assign n30546 = n30137 & n30527 ;
  assign n30547 = ~n30545 & ~n30546 ;
  assign n30548 = n30114 & ~n30547 ;
  assign n30549 = ~n30544 & ~n30548 ;
  assign n30550 = n30539 & n30549 ;
  assign n30551 = n30109 & n30550 ;
  assign n30552 = n29949 & ~n29974 ;
  assign n30553 = n2622 & ~n16398 ;
  assign n30554 = ~n15241 & n30553 ;
  assign n30555 = ~n16404 & n30554 ;
  assign n30556 = n2622 & n16398 ;
  assign n30557 = n15241 & n30556 ;
  assign n30558 = n16400 & n30556 ;
  assign n30559 = ~n15239 & n30558 ;
  assign n30560 = ~n30557 & ~n30559 ;
  assign n30561 = ~n30555 & n30560 ;
  assign n30562 = \b[52]  & n2912 ;
  assign n30563 = n2909 & n30562 ;
  assign n30564 = \b[54]  & n2620 ;
  assign n30565 = \a[20]  & \b[53]  ;
  assign n30566 = n2910 & n30565 ;
  assign n30567 = ~\a[21]  & \b[53]  ;
  assign n30568 = n2614 & n30567 ;
  assign n30569 = ~n30566 & ~n30568 ;
  assign n30570 = ~n30564 & n30569 ;
  assign n30571 = ~n30563 & n30570 ;
  assign n30572 = n30561 & n30571 ;
  assign n30573 = ~\a[23]  & ~n30572 ;
  assign n30574 = \a[23]  & n30571 ;
  assign n30575 = n30561 & n30574 ;
  assign n30576 = ~n30573 & ~n30575 ;
  assign n30577 = ~n29969 & n30576 ;
  assign n30578 = ~n30552 & n30577 ;
  assign n30579 = ~n30551 & ~n30578 ;
  assign n30580 = ~n30109 & ~n30550 ;
  assign n30581 = n29969 & ~n30576 ;
  assign n30582 = n29949 & ~n30576 ;
  assign n30583 = ~n29974 & n30582 ;
  assign n30584 = ~n30581 & ~n30583 ;
  assign n30585 = ~n30580 & n30584 ;
  assign n30586 = n30579 & n30585 ;
  assign n30587 = ~n30551 & ~n30580 ;
  assign n30588 = n30578 & ~n30587 ;
  assign n30589 = ~n29969 & ~n30552 ;
  assign n30590 = ~n30550 & ~n30576 ;
  assign n30591 = ~n30109 & n30590 ;
  assign n30592 = n30550 & ~n30576 ;
  assign n30593 = n30109 & n30592 ;
  assign n30594 = ~n30591 & ~n30593 ;
  assign n30595 = ~n30589 & ~n30594 ;
  assign n30596 = ~n30588 & ~n30595 ;
  assign n30597 = ~n30586 & n30596 ;
  assign n30598 = n30083 & n30597 ;
  assign n30599 = ~n30079 & n30598 ;
  assign n30600 = n30075 & ~n30597 ;
  assign n30601 = ~n30078 & n30600 ;
  assign n30602 = ~n30075 & ~n30597 ;
  assign n30603 = n30078 & n30602 ;
  assign n30604 = ~n30601 & ~n30603 ;
  assign n30605 = ~n30599 & n30604 ;
  assign n30606 = n30058 & ~n30605 ;
  assign n30607 = ~n30034 & n30606 ;
  assign n30608 = ~n30058 & ~n30075 ;
  assign n30609 = ~n30597 & n30608 ;
  assign n30610 = ~n30078 & n30609 ;
  assign n30611 = ~n30058 & n30075 ;
  assign n30612 = n30597 & n30611 ;
  assign n30613 = ~n30078 & n30612 ;
  assign n30614 = ~n30610 & ~n30613 ;
  assign n30615 = ~n30597 & n30611 ;
  assign n30616 = n30078 & n30615 ;
  assign n30617 = n30597 & n30608 ;
  assign n30618 = n30078 & n30617 ;
  assign n30619 = ~n30616 & ~n30618 ;
  assign n30620 = n30614 & n30619 ;
  assign n30621 = ~n30034 & ~n30620 ;
  assign n30622 = n30058 & ~n30075 ;
  assign n30623 = ~n30597 & n30622 ;
  assign n30624 = ~n30078 & n30623 ;
  assign n30625 = n30058 & n30075 ;
  assign n30626 = n30597 & n30625 ;
  assign n30627 = ~n30078 & n30626 ;
  assign n30628 = ~n30624 & ~n30627 ;
  assign n30629 = ~n30597 & n30625 ;
  assign n30630 = n30078 & n30629 ;
  assign n30631 = n30597 & n30622 ;
  assign n30632 = n30078 & n30631 ;
  assign n30633 = ~n30630 & ~n30632 ;
  assign n30634 = n30628 & n30633 ;
  assign n30635 = n30033 & ~n30634 ;
  assign n30636 = ~n30030 & n30635 ;
  assign n30637 = ~n30078 & n30615 ;
  assign n30638 = ~n30078 & n30617 ;
  assign n30639 = ~n30637 & ~n30638 ;
  assign n30640 = n30078 & n30609 ;
  assign n30641 = n30078 & n30612 ;
  assign n30642 = ~n30640 & ~n30641 ;
  assign n30643 = n30639 & n30642 ;
  assign n30644 = n30033 & ~n30643 ;
  assign n30645 = ~n30030 & n30644 ;
  assign n30646 = ~n30636 & ~n30645 ;
  assign n30647 = ~n30621 & n30646 ;
  assign n30648 = ~n30607 & n30647 ;
  assign n30649 = ~n29456 & ~n29985 ;
  assign n30650 = n999 & ~n22461 ;
  assign n30651 = ~n22459 & n30650 ;
  assign n30652 = \b[63]  & n997 ;
  assign n30653 = \a[12]  & \b[62]  ;
  assign n30654 = n28195 & n30653 ;
  assign n30655 = ~n30652 & ~n30654 ;
  assign n30656 = \b[61]  & n1182 ;
  assign n30657 = n1179 & n30656 ;
  assign n30658 = ~\a[12]  & \b[62]  ;
  assign n30659 = n7674 & n30658 ;
  assign n30660 = ~n30657 & ~n30659 ;
  assign n30661 = n30655 & n30660 ;
  assign n30662 = ~n30651 & n30661 ;
  assign n30663 = ~\a[14]  & ~n30662 ;
  assign n30664 = \a[14]  & n30661 ;
  assign n30665 = ~n30651 & n30664 ;
  assign n30666 = ~n30663 & ~n30665 ;
  assign n30667 = ~n30649 & ~n30666 ;
  assign n30668 = n30649 & n30666 ;
  assign n30669 = ~n30667 & ~n30668 ;
  assign n30670 = n30648 & n30669 ;
  assign n30671 = ~n30648 & ~n30669 ;
  assign n30672 = ~n30670 & ~n30671 ;
  assign n30673 = n30029 & n30672 ;
  assign n30674 = ~n30029 & ~n30672 ;
  assign n30675 = ~n30673 & ~n30674 ;
  assign n30676 = ~n30019 & n30675 ;
  assign n30677 = ~n30026 & n30676 ;
  assign n30678 = ~n30019 & ~n30026 ;
  assign n30679 = ~n30675 & ~n30678 ;
  assign n30680 = ~n30677 & ~n30679 ;
  assign n30681 = ~n30673 & ~n30677 ;
  assign n30682 = ~n30648 & ~n30667 ;
  assign n30683 = ~n30668 & ~n30682 ;
  assign n30684 = n30033 & ~n30058 ;
  assign n30685 = ~n30030 & n30684 ;
  assign n30686 = ~n30636 & ~n30685 ;
  assign n30687 = ~n30621 & n30686 ;
  assign n30688 = n30584 & ~n30587 ;
  assign n30689 = n1965 & n18940 ;
  assign n30690 = ~n18937 & n30689 ;
  assign n30691 = n1965 & ~n18940 ;
  assign n30692 = ~n17685 & n30691 ;
  assign n30693 = ~n18936 & n30692 ;
  assign n30694 = \b[56]  & n2218 ;
  assign n30695 = n2216 & n30694 ;
  assign n30696 = ~\a[18]  & \b[57]  ;
  assign n30697 = n1957 & n30696 ;
  assign n30698 = ~n30695 & ~n30697 ;
  assign n30699 = \b[58]  & n1963 ;
  assign n30700 = \a[18]  & \b[57]  ;
  assign n30701 = n28047 & n30700 ;
  assign n30702 = \a[20]  & ~n30701 ;
  assign n30703 = ~n30699 & n30702 ;
  assign n30704 = n30698 & n30703 ;
  assign n30705 = ~n30693 & n30704 ;
  assign n30706 = ~n30690 & n30705 ;
  assign n30707 = ~n30699 & ~n30701 ;
  assign n30708 = n30698 & n30707 ;
  assign n30709 = ~n30693 & n30708 ;
  assign n30710 = ~n30690 & n30709 ;
  assign n30711 = ~\a[20]  & ~n30710 ;
  assign n30712 = ~n30706 & ~n30711 ;
  assign n30713 = ~n30578 & ~n30712 ;
  assign n30714 = ~n30688 & n30713 ;
  assign n30715 = n30108 & ~n30550 ;
  assign n30716 = n2622 & ~n16446 ;
  assign n30717 = ~n16444 & n30716 ;
  assign n30718 = \b[53]  & n2912 ;
  assign n30719 = n2909 & n30718 ;
  assign n30720 = \b[55]  & n2620 ;
  assign n30721 = \a[20]  & \b[54]  ;
  assign n30722 = n2910 & n30721 ;
  assign n30723 = ~\a[21]  & \b[54]  ;
  assign n30724 = n2614 & n30723 ;
  assign n30725 = ~n30722 & ~n30724 ;
  assign n30726 = ~n30720 & n30725 ;
  assign n30727 = ~n30719 & n30726 ;
  assign n30728 = ~n30717 & n30727 ;
  assign n30729 = \a[23]  & ~n30728 ;
  assign n30730 = ~\a[23]  & n30728 ;
  assign n30731 = ~n30729 & ~n30730 ;
  assign n30732 = ~n30104 & n30731 ;
  assign n30733 = ~n30715 & n30732 ;
  assign n30734 = ~\a[23]  & ~n30728 ;
  assign n30735 = \a[23]  & n30727 ;
  assign n30736 = ~n30717 & n30735 ;
  assign n30737 = n30104 & ~n30736 ;
  assign n30738 = n30108 & ~n30736 ;
  assign n30739 = ~n30550 & n30738 ;
  assign n30740 = ~n30737 & ~n30739 ;
  assign n30741 = ~n30734 & ~n30740 ;
  assign n30742 = ~n30733 & ~n30741 ;
  assign n30743 = ~n30517 & ~n30523 ;
  assign n30744 = n5211 & n11906 ;
  assign n30745 = ~n11903 & n30744 ;
  assign n30746 = n5211 & ~n11906 ;
  assign n30747 = ~n11392 & n30746 ;
  assign n30748 = ~n11902 & n30747 ;
  assign n30749 = \b[46]  & n5209 ;
  assign n30750 = \a[30]  & \b[45]  ;
  assign n30751 = n5200 & n30750 ;
  assign n30752 = ~n30749 & ~n30751 ;
  assign n30753 = \b[44]  & n5595 ;
  assign n30754 = n5592 & n30753 ;
  assign n30755 = ~\a[30]  & \b[45]  ;
  assign n30756 = n5203 & n30755 ;
  assign n30757 = ~n30754 & ~n30756 ;
  assign n30758 = n30752 & n30757 ;
  assign n30759 = ~n30748 & n30758 ;
  assign n30760 = ~n30745 & n30759 ;
  assign n30761 = \a[32]  & ~n30760 ;
  assign n30762 = ~\a[32]  & n30760 ;
  assign n30763 = ~n30761 & ~n30762 ;
  assign n30764 = ~n30518 & n30763 ;
  assign n30765 = ~n30743 & n30764 ;
  assign n30766 = ~n30518 & ~n30743 ;
  assign n30767 = ~\a[32]  & ~n30760 ;
  assign n30768 = \a[32]  & n30758 ;
  assign n30769 = ~n30748 & n30768 ;
  assign n30770 = ~n30745 & n30769 ;
  assign n30771 = ~n30767 & ~n30770 ;
  assign n30772 = ~n30766 & n30771 ;
  assign n30773 = ~n30765 & ~n30772 ;
  assign n30774 = n30186 & n30507 ;
  assign n30775 = n30512 & ~n30774 ;
  assign n30776 = ~n30339 & ~n30367 ;
  assign n30777 = ~n30340 & ~n30776 ;
  assign n30778 = n30330 & ~n30331 ;
  assign n30779 = ~n30217 & ~n30331 ;
  assign n30780 = ~n30778 & ~n30779 ;
  assign n30781 = ~n30321 & ~n30326 ;
  assign n30782 = ~n30322 & ~n30781 ;
  assign n30783 = ~n30298 & n30315 ;
  assign n30784 = n30270 & ~n30291 ;
  assign n30785 = \a[62]  & n30290 ;
  assign n30786 = ~n30784 & n30785 ;
  assign n30787 = ~\a[62]  & n30290 ;
  assign n30788 = n30784 & n30787 ;
  assign n30789 = ~n30786 & ~n30788 ;
  assign n30790 = ~n30783 & n30789 ;
  assign n30791 = n1512 & n20521 ;
  assign n30792 = ~n1509 & n30791 ;
  assign n30793 = n10165 & n20521 ;
  assign n30794 = ~n1508 & n30793 ;
  assign n30795 = \b[16]  & n20519 ;
  assign n30796 = \a[60]  & \b[15]  ;
  assign n30797 = n20510 & n30796 ;
  assign n30798 = ~n30795 & ~n30797 ;
  assign n30799 = \b[14]  & n21315 ;
  assign n30800 = n21312 & n30799 ;
  assign n30801 = ~\a[60]  & \b[15]  ;
  assign n30802 = n20513 & n30801 ;
  assign n30803 = ~n30800 & ~n30802 ;
  assign n30804 = n30798 & n30803 ;
  assign n30805 = ~n30794 & n30804 ;
  assign n30806 = ~n30792 & n30805 ;
  assign n30807 = ~n30283 & ~n30287 ;
  assign n30808 = n30281 & ~n30807 ;
  assign n30809 = \b[13]  & n21958 ;
  assign n30810 = \b[12]  & n21957 ;
  assign n30811 = ~n30809 & ~n30810 ;
  assign n30812 = ~n30808 & n30811 ;
  assign n30813 = n30281 & ~n30811 ;
  assign n30814 = ~n30807 & n30813 ;
  assign n30815 = ~\a[62]  & ~n30814 ;
  assign n30816 = ~n30812 & n30815 ;
  assign n30817 = ~n30806 & n30816 ;
  assign n30818 = \a[62]  & ~n30814 ;
  assign n30819 = ~n30812 & n30818 ;
  assign n30820 = n30804 & n30819 ;
  assign n30821 = ~n30794 & n30820 ;
  assign n30822 = ~n30792 & n30821 ;
  assign n30823 = ~n30817 & ~n30822 ;
  assign n30824 = ~\a[62]  & ~n30806 ;
  assign n30825 = ~n30812 & ~n30814 ;
  assign n30826 = \a[62]  & n30804 ;
  assign n30827 = ~n30794 & n30826 ;
  assign n30828 = ~n30792 & n30827 ;
  assign n30829 = ~n30825 & ~n30828 ;
  assign n30830 = ~n30824 & n30829 ;
  assign n30831 = n30823 & ~n30830 ;
  assign n30832 = ~n30790 & ~n30831 ;
  assign n30833 = n30790 & n30831 ;
  assign n30834 = ~n30832 & ~n30833 ;
  assign n30835 = ~n2076 & n18516 ;
  assign n30836 = ~n1874 & n18516 ;
  assign n30837 = ~n1878 & n30836 ;
  assign n30838 = ~n30835 & ~n30837 ;
  assign n30839 = ~n2079 & ~n30838 ;
  assign n30840 = \b[19]  & n18514 ;
  assign n30841 = \a[56]  & \b[18]  ;
  assign n30842 = n19181 & n30841 ;
  assign n30843 = ~\a[57]  & \b[18]  ;
  assign n30844 = n18508 & n30843 ;
  assign n30845 = ~n30842 & ~n30844 ;
  assign n30846 = ~n30840 & n30845 ;
  assign n30847 = \b[17]  & n19183 ;
  assign n30848 = n19180 & n30847 ;
  assign n30849 = \a[59]  & ~n30848 ;
  assign n30850 = n30846 & n30849 ;
  assign n30851 = ~n30839 & n30850 ;
  assign n30852 = n30846 & ~n30848 ;
  assign n30853 = ~\a[59]  & ~n30852 ;
  assign n30854 = ~\a[59]  & ~n2079 ;
  assign n30855 = ~n30838 & n30854 ;
  assign n30856 = ~n30853 & ~n30855 ;
  assign n30857 = ~n30851 & n30856 ;
  assign n30858 = n30834 & ~n30857 ;
  assign n30859 = ~n30834 & n30857 ;
  assign n30860 = ~n30858 & ~n30859 ;
  assign n30861 = ~n30782 & ~n30860 ;
  assign n30862 = n30782 & n30860 ;
  assign n30863 = ~n30861 & ~n30862 ;
  assign n30864 = n2768 & n16655 ;
  assign n30865 = ~n2765 & n30864 ;
  assign n30866 = n6462 & n16655 ;
  assign n30867 = ~n2764 & n30866 ;
  assign n30868 = \b[20]  & n17308 ;
  assign n30869 = n17305 & n30868 ;
  assign n30870 = \b[22]  & n16653 ;
  assign n30871 = \a[54]  & \b[21]  ;
  assign n30872 = n16644 & n30871 ;
  assign n30873 = ~\a[54]  & \b[21]  ;
  assign n30874 = n16647 & n30873 ;
  assign n30875 = ~n30872 & ~n30874 ;
  assign n30876 = ~n30870 & n30875 ;
  assign n30877 = ~n30869 & n30876 ;
  assign n30878 = ~n30867 & n30877 ;
  assign n30879 = ~n30865 & n30878 ;
  assign n30880 = ~\a[56]  & ~n30879 ;
  assign n30881 = \a[56]  & n30877 ;
  assign n30882 = ~n30867 & n30881 ;
  assign n30883 = ~n30865 & n30882 ;
  assign n30884 = ~n30880 & ~n30883 ;
  assign n30885 = ~n30863 & n30884 ;
  assign n30886 = n30863 & ~n30884 ;
  assign n30887 = ~n30885 & ~n30886 ;
  assign n30888 = ~n30780 & ~n30887 ;
  assign n30889 = n30780 & n30887 ;
  assign n30890 = ~n30888 & ~n30889 ;
  assign n30891 = ~n3564 & n14793 ;
  assign n30892 = ~n3282 & n14793 ;
  assign n30893 = ~n3560 & n30892 ;
  assign n30894 = ~n30891 & ~n30893 ;
  assign n30895 = ~n3567 & ~n30894 ;
  assign n30896 = \b[23]  & n15517 ;
  assign n30897 = n15514 & n30896 ;
  assign n30898 = ~\a[51]  & \b[24]  ;
  assign n30899 = n14785 & n30898 ;
  assign n30900 = ~n30897 & ~n30899 ;
  assign n30901 = \b[25]  & n14791 ;
  assign n30902 = \a[51]  & \b[24]  ;
  assign n30903 = n14782 & n30902 ;
  assign n30904 = \a[53]  & ~n30903 ;
  assign n30905 = ~n30901 & n30904 ;
  assign n30906 = n30900 & n30905 ;
  assign n30907 = ~n30895 & n30906 ;
  assign n30908 = ~n30901 & ~n30903 ;
  assign n30909 = n30900 & n30908 ;
  assign n30910 = ~\a[53]  & ~n30909 ;
  assign n30911 = ~\a[53]  & ~n3567 ;
  assign n30912 = ~n30894 & n30911 ;
  assign n30913 = ~n30910 & ~n30912 ;
  assign n30914 = ~n30907 & n30913 ;
  assign n30915 = n30890 & ~n30914 ;
  assign n30916 = ~n30890 & n30914 ;
  assign n30917 = ~n30915 & ~n30916 ;
  assign n30918 = ~n30777 & ~n30917 ;
  assign n30919 = n30777 & n30917 ;
  assign n30920 = ~n30918 & ~n30919 ;
  assign n30921 = n4456 & n13125 ;
  assign n30922 = ~n18723 & n30921 ;
  assign n30923 = n13125 & n16805 ;
  assign n30924 = ~n4452 & n30923 ;
  assign n30925 = \b[26]  & n13794 ;
  assign n30926 = n13792 & n30925 ;
  assign n30927 = ~\a[48]  & \b[27]  ;
  assign n30928 = n13117 & n30927 ;
  assign n30929 = ~n30926 & ~n30928 ;
  assign n30930 = \b[28]  & n13123 ;
  assign n30931 = \a[48]  & \b[27]  ;
  assign n30932 = n13786 & n30931 ;
  assign n30933 = \a[50]  & ~n30932 ;
  assign n30934 = ~n30930 & n30933 ;
  assign n30935 = n30929 & n30934 ;
  assign n30936 = ~n30924 & n30935 ;
  assign n30937 = ~n30922 & n30936 ;
  assign n30938 = ~n30930 & ~n30932 ;
  assign n30939 = n30929 & n30938 ;
  assign n30940 = ~n30924 & n30939 ;
  assign n30941 = ~n30922 & n30940 ;
  assign n30942 = ~\a[50]  & ~n30941 ;
  assign n30943 = ~n30937 & ~n30942 ;
  assign n30944 = ~n30920 & n30943 ;
  assign n30945 = n30920 & ~n30943 ;
  assign n30946 = ~n30944 & ~n30945 ;
  assign n30947 = ~n5459 & n11572 ;
  assign n30948 = ~n5104 & n11572 ;
  assign n30949 = ~n5455 & n30948 ;
  assign n30950 = ~n30947 & ~n30949 ;
  assign n30951 = ~n5462 & ~n30950 ;
  assign n30952 = \b[29]  & n12159 ;
  assign n30953 = n12156 & n30952 ;
  assign n30954 = ~\a[45]  & \b[30]  ;
  assign n30955 = n11564 & n30954 ;
  assign n30956 = ~n30953 & ~n30955 ;
  assign n30957 = \b[31]  & n11570 ;
  assign n30958 = \a[45]  & \b[30]  ;
  assign n30959 = n11561 & n30958 ;
  assign n30960 = \a[47]  & ~n30959 ;
  assign n30961 = ~n30957 & n30960 ;
  assign n30962 = n30956 & n30961 ;
  assign n30963 = ~n30951 & n30962 ;
  assign n30964 = ~n30957 & ~n30959 ;
  assign n30965 = n30956 & n30964 ;
  assign n30966 = ~\a[47]  & ~n30965 ;
  assign n30967 = ~\a[47]  & ~n5462 ;
  assign n30968 = ~n30950 & n30967 ;
  assign n30969 = ~n30966 & ~n30968 ;
  assign n30970 = ~n30963 & n30969 ;
  assign n30971 = n30372 & n30380 ;
  assign n30972 = n30377 & ~n30971 ;
  assign n30973 = n30970 & n30972 ;
  assign n30974 = ~n30946 & n30973 ;
  assign n30975 = n30970 & ~n30972 ;
  assign n30976 = n30946 & n30975 ;
  assign n30977 = ~n30974 & ~n30976 ;
  assign n30978 = ~n30970 & ~n30972 ;
  assign n30979 = ~n30946 & n30978 ;
  assign n30980 = ~n30970 & n30972 ;
  assign n30981 = n30946 & n30980 ;
  assign n30982 = ~n30979 & ~n30981 ;
  assign n30983 = n30977 & n30982 ;
  assign n30984 = n6565 & n10082 ;
  assign n30985 = ~n6562 & n30984 ;
  assign n30986 = ~n6565 & n10082 ;
  assign n30987 = ~n5850 & n30986 ;
  assign n30988 = ~n6561 & n30987 ;
  assign n30989 = \b[32]  & n10681 ;
  assign n30990 = n10678 & n30989 ;
  assign n30991 = \b[34]  & n10080 ;
  assign n30992 = \a[41]  & \b[33]  ;
  assign n30993 = n10679 & n30992 ;
  assign n30994 = ~\a[42]  & \b[33]  ;
  assign n30995 = n10074 & n30994 ;
  assign n30996 = ~n30993 & ~n30995 ;
  assign n30997 = ~n30991 & n30996 ;
  assign n30998 = ~n30990 & n30997 ;
  assign n30999 = ~n30988 & n30998 ;
  assign n31000 = ~n30985 & n30999 ;
  assign n31001 = ~\a[44]  & ~n31000 ;
  assign n31002 = \a[44]  & n30998 ;
  assign n31003 = ~n30988 & n31002 ;
  assign n31004 = ~n30985 & n31003 ;
  assign n31005 = ~n31001 & ~n31004 ;
  assign n31006 = n30414 & ~n30436 ;
  assign n31007 = n30409 & ~n31006 ;
  assign n31008 = ~n31005 & ~n31007 ;
  assign n31009 = ~n30983 & n31008 ;
  assign n31010 = ~n31005 & n31007 ;
  assign n31011 = n30983 & n31010 ;
  assign n31012 = ~n31009 & ~n31011 ;
  assign n31013 = n31005 & ~n31007 ;
  assign n31014 = n30983 & n31013 ;
  assign n31015 = n31005 & n31007 ;
  assign n31016 = ~n30983 & n31015 ;
  assign n31017 = ~n31014 & ~n31016 ;
  assign n31018 = n31012 & n31017 ;
  assign n31019 = ~n7761 & n8759 ;
  assign n31020 = ~n7759 & n31019 ;
  assign n31021 = \b[35]  & n9301 ;
  assign n31022 = n9298 & n31021 ;
  assign n31023 = ~\a[39]  & \b[36]  ;
  assign n31024 = n8751 & n31023 ;
  assign n31025 = ~n31022 & ~n31024 ;
  assign n31026 = \b[37]  & n8757 ;
  assign n31027 = \a[39]  & \b[36]  ;
  assign n31028 = n8748 & n31027 ;
  assign n31029 = \a[41]  & ~n31028 ;
  assign n31030 = ~n31026 & n31029 ;
  assign n31031 = n31025 & n31030 ;
  assign n31032 = ~n31020 & n31031 ;
  assign n31033 = ~n31026 & ~n31028 ;
  assign n31034 = n31025 & n31033 ;
  assign n31035 = ~n31020 & n31034 ;
  assign n31036 = ~\a[41]  & ~n31035 ;
  assign n31037 = ~n31032 & ~n31036 ;
  assign n31038 = n30441 & n30472 ;
  assign n31039 = n30446 & ~n31038 ;
  assign n31040 = n31037 & n31039 ;
  assign n31041 = ~n31018 & n31040 ;
  assign n31042 = n31037 & ~n31039 ;
  assign n31043 = n31018 & n31042 ;
  assign n31044 = ~n31041 & ~n31043 ;
  assign n31045 = ~n31037 & ~n31039 ;
  assign n31046 = ~n31018 & n31045 ;
  assign n31047 = ~n31037 & n31039 ;
  assign n31048 = n31018 & n31047 ;
  assign n31049 = ~n31046 & ~n31048 ;
  assign n31050 = n31044 & n31049 ;
  assign n31051 = n7534 & n9044 ;
  assign n31052 = ~n9041 & n31051 ;
  assign n31053 = n7534 & ~n9044 ;
  assign n31054 = ~n8597 & n31053 ;
  assign n31055 = ~n9040 & n31054 ;
  assign n31056 = \b[38]  & n7973 ;
  assign n31057 = n7970 & n31056 ;
  assign n31058 = ~\a[36]  & \b[39]  ;
  assign n31059 = n7526 & n31058 ;
  assign n31060 = ~n31057 & ~n31059 ;
  assign n31061 = \b[40]  & n7532 ;
  assign n31062 = \a[36]  & \b[39]  ;
  assign n31063 = n17801 & n31062 ;
  assign n31064 = \a[38]  & ~n31063 ;
  assign n31065 = ~n31061 & n31064 ;
  assign n31066 = n31060 & n31065 ;
  assign n31067 = ~n31055 & n31066 ;
  assign n31068 = ~n31052 & n31067 ;
  assign n31069 = ~n31061 & ~n31063 ;
  assign n31070 = n31060 & n31069 ;
  assign n31071 = ~n31055 & n31070 ;
  assign n31072 = ~n31052 & n31071 ;
  assign n31073 = ~\a[38]  & ~n31072 ;
  assign n31074 = ~n31068 & ~n31073 ;
  assign n31075 = n30477 & ~n30485 ;
  assign n31076 = n30482 & ~n31075 ;
  assign n31077 = ~n31074 & ~n31076 ;
  assign n31078 = ~n31050 & n31077 ;
  assign n31079 = ~n31074 & n31076 ;
  assign n31080 = n31050 & n31079 ;
  assign n31081 = ~n31078 & ~n31080 ;
  assign n31082 = n31074 & n31076 ;
  assign n31083 = ~n31050 & n31082 ;
  assign n31084 = n31074 & ~n31076 ;
  assign n31085 = n31050 & n31084 ;
  assign n31086 = ~n31083 & ~n31085 ;
  assign n31087 = n31081 & n31086 ;
  assign n31088 = n30775 & n31087 ;
  assign n31089 = ~n30775 & ~n31087 ;
  assign n31090 = ~n31088 & ~n31089 ;
  assign n31091 = n6309 & ~n10409 ;
  assign n31092 = ~n10407 & n31091 ;
  assign n31093 = \b[41]  & n6778 ;
  assign n31094 = n6775 & n31093 ;
  assign n31095 = ~\a[33]  & \b[42]  ;
  assign n31096 = n6301 & n31095 ;
  assign n31097 = ~n31094 & ~n31096 ;
  assign n31098 = \b[43]  & n6307 ;
  assign n31099 = \a[33]  & \b[42]  ;
  assign n31100 = n6298 & n31099 ;
  assign n31101 = \a[35]  & ~n31100 ;
  assign n31102 = ~n31098 & n31101 ;
  assign n31103 = n31097 & n31102 ;
  assign n31104 = ~n31092 & n31103 ;
  assign n31105 = ~n31098 & ~n31100 ;
  assign n31106 = n31097 & n31105 ;
  assign n31107 = ~n31092 & n31106 ;
  assign n31108 = ~\a[35]  & ~n31107 ;
  assign n31109 = ~n31104 & ~n31108 ;
  assign n31110 = n31090 & ~n31109 ;
  assign n31111 = ~n31090 & n31109 ;
  assign n31112 = ~n31110 & ~n31111 ;
  assign n31113 = n30773 & n31112 ;
  assign n31114 = ~n30773 & ~n31112 ;
  assign n31115 = ~n31113 & ~n31114 ;
  assign n31116 = ~n30134 & ~n30526 ;
  assign n31117 = n4249 & ~n13524 ;
  assign n31118 = ~n13522 & n31117 ;
  assign n31119 = \b[49]  & n4247 ;
  assign n31120 = \a[27]  & \b[48]  ;
  assign n31121 = n4238 & n31120 ;
  assign n31122 = ~n31119 & ~n31121 ;
  assign n31123 = \b[47]  & n4647 ;
  assign n31124 = n4644 & n31123 ;
  assign n31125 = ~\a[27]  & \b[48]  ;
  assign n31126 = n4241 & n31125 ;
  assign n31127 = ~n31124 & ~n31126 ;
  assign n31128 = n31122 & n31127 ;
  assign n31129 = ~n31118 & n31128 ;
  assign n31130 = \a[29]  & ~n31129 ;
  assign n31131 = ~\a[29]  & n31129 ;
  assign n31132 = ~n31130 & ~n31131 ;
  assign n31133 = ~n30136 & n31132 ;
  assign n31134 = ~n31116 & n31133 ;
  assign n31135 = ~\a[29]  & ~n31129 ;
  assign n31136 = \a[29]  & n31128 ;
  assign n31137 = ~n31118 & n31136 ;
  assign n31138 = n30136 & ~n31137 ;
  assign n31139 = ~n30134 & ~n31137 ;
  assign n31140 = ~n30526 & n31139 ;
  assign n31141 = ~n31138 & ~n31140 ;
  assign n31142 = ~n31135 & ~n31141 ;
  assign n31143 = ~n31134 & ~n31142 ;
  assign n31144 = n31115 & n31143 ;
  assign n31145 = ~n31115 & ~n31143 ;
  assign n31146 = ~n31144 & ~n31145 ;
  assign n31147 = ~n3154 & ~n14093 ;
  assign n31148 = ~n15201 & n31147 ;
  assign n31149 = ~n15197 & n31148 ;
  assign n31150 = ~n3399 & n31149 ;
  assign n31151 = n3402 & n15201 ;
  assign n31152 = ~n15198 & n31151 ;
  assign n31153 = ~n31150 & ~n31152 ;
  assign n31154 = \b[50]  & n3733 ;
  assign n31155 = n3730 & n31154 ;
  assign n31156 = ~\a[24]  & \b[51]  ;
  assign n31157 = n3394 & n31156 ;
  assign n31158 = ~n31155 & ~n31157 ;
  assign n31159 = \b[52]  & n3400 ;
  assign n31160 = \a[24]  & \b[51]  ;
  assign n31161 = n27626 & n31160 ;
  assign n31162 = \a[26]  & ~n31161 ;
  assign n31163 = ~n31159 & n31162 ;
  assign n31164 = n31158 & n31163 ;
  assign n31165 = n31153 & n31164 ;
  assign n31166 = ~n31159 & ~n31161 ;
  assign n31167 = n31158 & n31166 ;
  assign n31168 = n31153 & n31167 ;
  assign n31169 = ~\a[26]  & ~n31168 ;
  assign n31170 = ~n31165 & ~n31169 ;
  assign n31171 = ~n30114 & n30540 ;
  assign n31172 = ~n30543 & ~n31171 ;
  assign n31173 = ~n30114 & n30541 ;
  assign n31174 = ~n30137 & n30535 ;
  assign n31175 = n30137 & n30533 ;
  assign n31176 = ~n31174 & ~n31175 ;
  assign n31177 = ~n31173 & n31176 ;
  assign n31178 = n31172 & n31177 ;
  assign n31179 = ~n31170 & n31178 ;
  assign n31180 = n31146 & n31179 ;
  assign n31181 = n31170 & ~n31178 ;
  assign n31182 = n31146 & n31181 ;
  assign n31183 = ~n31180 & ~n31182 ;
  assign n31184 = ~n31146 & ~n31181 ;
  assign n31185 = ~n31179 & n31184 ;
  assign n31186 = n31183 & ~n31185 ;
  assign n31187 = ~n30742 & ~n31186 ;
  assign n31188 = n30742 & n31186 ;
  assign n31189 = ~n31187 & ~n31188 ;
  assign n31190 = ~n30578 & ~n30688 ;
  assign n31191 = n30712 & ~n31190 ;
  assign n31192 = ~n31189 & ~n31191 ;
  assign n31193 = ~n30714 & n31192 ;
  assign n31194 = n31189 & n31191 ;
  assign n31195 = ~n30712 & n31190 ;
  assign n31196 = n31189 & n31195 ;
  assign n31197 = ~n31194 & ~n31196 ;
  assign n31198 = ~n31193 & n31197 ;
  assign n31199 = n30083 & ~n30597 ;
  assign n31200 = ~n30079 & ~n31199 ;
  assign n31201 = n1467 & ~n20971 ;
  assign n31202 = ~n20969 & n31201 ;
  assign n31203 = \b[61]  & n1465 ;
  assign n31204 = \a[15]  & \b[60]  ;
  assign n31205 = n1456 & n31204 ;
  assign n31206 = ~n31203 & ~n31205 ;
  assign n31207 = \b[59]  & n1652 ;
  assign n31208 = n1649 & n31207 ;
  assign n31209 = ~\a[15]  & \b[60]  ;
  assign n31210 = n1459 & n31209 ;
  assign n31211 = ~n31208 & ~n31210 ;
  assign n31212 = n31206 & n31211 ;
  assign n31213 = ~n31202 & n31212 ;
  assign n31214 = \a[17]  & ~n31213 ;
  assign n31215 = ~\a[17]  & n31213 ;
  assign n31216 = ~n31214 & ~n31215 ;
  assign n31217 = n31200 & n31216 ;
  assign n31218 = ~\a[17]  & ~n31213 ;
  assign n31219 = \a[17]  & n31212 ;
  assign n31220 = ~n31202 & n31219 ;
  assign n31221 = ~n31218 & ~n31220 ;
  assign n31222 = ~n31200 & n31221 ;
  assign n31223 = ~n31217 & ~n31222 ;
  assign n31224 = n31198 & n31223 ;
  assign n31225 = ~n31198 & ~n31223 ;
  assign n31226 = ~n31224 & ~n31225 ;
  assign n31227 = \b[62]  & n1182 ;
  assign n31228 = n1179 & n31227 ;
  assign n31229 = ~\a[12]  & \b[63]  ;
  assign n31230 = n7674 & n31229 ;
  assign n31231 = \a[12]  & \b[63]  ;
  assign n31232 = n28195 & n31231 ;
  assign n31233 = ~n31230 & ~n31232 ;
  assign n31234 = ~n31228 & n31233 ;
  assign n31235 = ~\a[14]  & ~n31234 ;
  assign n31236 = n999 & ~n22458 ;
  assign n31237 = ~\a[14]  & n31236 ;
  assign n31238 = ~n23173 & n31237 ;
  assign n31239 = ~n31235 & ~n31238 ;
  assign n31240 = ~n23173 & n31236 ;
  assign n31241 = \a[14]  & n31234 ;
  assign n31242 = ~n31240 & n31241 ;
  assign n31243 = n31239 & ~n31242 ;
  assign n31244 = n31226 & ~n31243 ;
  assign n31245 = n30687 & n31244 ;
  assign n31246 = n31226 & n31243 ;
  assign n31247 = ~n30687 & n31246 ;
  assign n31248 = ~n31245 & ~n31247 ;
  assign n31249 = ~n31226 & ~n31243 ;
  assign n31250 = ~n30687 & n31249 ;
  assign n31251 = ~n31226 & n31243 ;
  assign n31252 = n30687 & n31251 ;
  assign n31253 = ~n31250 & ~n31252 ;
  assign n31254 = n31248 & n31253 ;
  assign n31255 = n30683 & n31254 ;
  assign n31256 = ~n30683 & ~n31254 ;
  assign n31257 = ~n31255 & ~n31256 ;
  assign n31258 = ~n30681 & n31257 ;
  assign n31259 = ~n30673 & ~n31257 ;
  assign n31260 = ~n30677 & n31259 ;
  assign n31261 = ~n31258 & ~n31260 ;
  assign n31262 = ~n30673 & ~n31255 ;
  assign n31263 = ~n30677 & n31262 ;
  assign n31264 = ~n30687 & ~n31243 ;
  assign n31265 = ~n31226 & ~n31264 ;
  assign n31266 = n30687 & n31243 ;
  assign n31267 = ~n31198 & ~n31217 ;
  assign n31268 = ~n31217 & n31222 ;
  assign n31269 = ~n31267 & ~n31268 ;
  assign n31270 = \b[63]  & n999 ;
  assign n31271 = ~n21694 & n31270 ;
  assign n31272 = ~n23171 & n31271 ;
  assign n31273 = \a[11]  & \a[13]  ;
  assign n31274 = \a[12]  & ~\a[14]  ;
  assign n31275 = n31273 & n31274 ;
  assign n31276 = ~\a[11]  & ~\a[13]  ;
  assign n31277 = ~\a[12]  & \a[14]  ;
  assign n31278 = n31276 & n31277 ;
  assign n31279 = ~n31275 & ~n31278 ;
  assign n31280 = \b[63]  & ~n31279 ;
  assign n31281 = \a[14]  & ~n31280 ;
  assign n31282 = ~n31272 & n31281 ;
  assign n31283 = ~n31272 & ~n31280 ;
  assign n31284 = ~\a[14]  & ~n31283 ;
  assign n31285 = ~n31282 & ~n31284 ;
  assign n31286 = ~n31269 & n31285 ;
  assign n31287 = n1965 & ~n19550 ;
  assign n31288 = ~n19548 & n31287 ;
  assign n31289 = \b[59]  & n1963 ;
  assign n31290 = \a[18]  & \b[58]  ;
  assign n31291 = n28047 & n31290 ;
  assign n31292 = ~n31289 & ~n31291 ;
  assign n31293 = \b[57]  & n2218 ;
  assign n31294 = n2216 & n31293 ;
  assign n31295 = ~\a[18]  & \b[58]  ;
  assign n31296 = n1957 & n31295 ;
  assign n31297 = ~n31294 & ~n31296 ;
  assign n31298 = n31292 & n31297 ;
  assign n31299 = ~n31288 & n31298 ;
  assign n31300 = ~\a[20]  & ~n31299 ;
  assign n31301 = \a[20]  & n31298 ;
  assign n31302 = ~n31288 & n31301 ;
  assign n31303 = ~n30733 & ~n31302 ;
  assign n31304 = n31186 & n31303 ;
  assign n31305 = n30741 & n31303 ;
  assign n31306 = ~n31304 & ~n31305 ;
  assign n31307 = ~n31300 & ~n31306 ;
  assign n31308 = ~n30733 & n30741 ;
  assign n31309 = ~n30733 & n31186 ;
  assign n31310 = ~n31300 & ~n31302 ;
  assign n31311 = ~n31309 & ~n31310 ;
  assign n31312 = ~n31308 & n31311 ;
  assign n31313 = ~n31307 & ~n31312 ;
  assign n31314 = ~n31146 & ~n31179 ;
  assign n31315 = ~n31181 & ~n31314 ;
  assign n31316 = n2622 & n17647 ;
  assign n31317 = ~n17644 & n31316 ;
  assign n31318 = n2622 & ~n17647 ;
  assign n31319 = ~n16441 & n31318 ;
  assign n31320 = ~n17643 & n31319 ;
  assign n31321 = \b[54]  & n2912 ;
  assign n31322 = n2909 & n31321 ;
  assign n31323 = \b[56]  & n2620 ;
  assign n31324 = \a[20]  & \b[55]  ;
  assign n31325 = n2910 & n31324 ;
  assign n31326 = ~\a[21]  & \b[55]  ;
  assign n31327 = n2614 & n31326 ;
  assign n31328 = ~n31325 & ~n31327 ;
  assign n31329 = ~n31323 & n31328 ;
  assign n31330 = ~n31322 & n31329 ;
  assign n31331 = ~n31320 & n31330 ;
  assign n31332 = ~n31317 & n31331 ;
  assign n31333 = ~\a[23]  & ~n31332 ;
  assign n31334 = \a[23]  & ~n31322 ;
  assign n31335 = n31329 & n31334 ;
  assign n31336 = ~n31320 & n31335 ;
  assign n31337 = ~n31317 & n31336 ;
  assign n31338 = ~n31333 & ~n31337 ;
  assign n31339 = ~n31315 & n31338 ;
  assign n31340 = \a[23]  & ~n31332 ;
  assign n31341 = ~\a[23]  & n31332 ;
  assign n31342 = ~n31340 & ~n31341 ;
  assign n31343 = ~n31181 & n31342 ;
  assign n31344 = ~n31314 & n31343 ;
  assign n31345 = ~n31339 & ~n31344 ;
  assign n31346 = n31115 & ~n31142 ;
  assign n31347 = n3402 & ~n15246 ;
  assign n31348 = ~n15244 & n31347 ;
  assign n31349 = \b[53]  & n3400 ;
  assign n31350 = \a[24]  & \b[52]  ;
  assign n31351 = n27626 & n31350 ;
  assign n31352 = ~n31349 & ~n31351 ;
  assign n31353 = \b[51]  & n3733 ;
  assign n31354 = n3730 & n31353 ;
  assign n31355 = ~\a[24]  & \b[52]  ;
  assign n31356 = n3394 & n31355 ;
  assign n31357 = ~n31354 & ~n31356 ;
  assign n31358 = n31352 & n31357 ;
  assign n31359 = ~n31348 & n31358 ;
  assign n31360 = ~\a[26]  & ~n31359 ;
  assign n31361 = \a[26]  & n31358 ;
  assign n31362 = ~n31348 & n31361 ;
  assign n31363 = ~n31134 & ~n31362 ;
  assign n31364 = ~n31360 & n31363 ;
  assign n31365 = ~n31346 & n31364 ;
  assign n31366 = ~n31134 & ~n31346 ;
  assign n31367 = \a[26]  & ~n31359 ;
  assign n31368 = ~\a[26]  & n31359 ;
  assign n31369 = ~n31367 & ~n31368 ;
  assign n31370 = ~n31366 & n31369 ;
  assign n31371 = ~n31365 & ~n31370 ;
  assign n31372 = ~n30765 & ~n31112 ;
  assign n31373 = ~n30765 & n30772 ;
  assign n31374 = ~n31372 & ~n31373 ;
  assign n31375 = n4249 & n14052 ;
  assign n31376 = ~n14049 & n31375 ;
  assign n31377 = n4249 & ~n14052 ;
  assign n31378 = ~n13519 & n31377 ;
  assign n31379 = ~n14048 & n31378 ;
  assign n31380 = \b[50]  & n4247 ;
  assign n31381 = \a[27]  & \b[49]  ;
  assign n31382 = n4238 & n31381 ;
  assign n31383 = ~n31380 & ~n31382 ;
  assign n31384 = \b[48]  & n4647 ;
  assign n31385 = n4644 & n31384 ;
  assign n31386 = ~\a[27]  & \b[49]  ;
  assign n31387 = n4241 & n31386 ;
  assign n31388 = ~n31385 & ~n31387 ;
  assign n31389 = n31383 & n31388 ;
  assign n31390 = ~n31379 & n31389 ;
  assign n31391 = ~n31376 & n31390 ;
  assign n31392 = \a[29]  & ~n31391 ;
  assign n31393 = ~\a[29]  & n31391 ;
  assign n31394 = ~n31392 & ~n31393 ;
  assign n31395 = n31374 & n31394 ;
  assign n31396 = ~\a[29]  & ~n31391 ;
  assign n31397 = \a[29]  & n31389 ;
  assign n31398 = ~n31379 & n31397 ;
  assign n31399 = ~n31376 & n31398 ;
  assign n31400 = ~n30765 & ~n31399 ;
  assign n31401 = ~n31112 & n31400 ;
  assign n31402 = n30772 & n31400 ;
  assign n31403 = ~n31401 & ~n31402 ;
  assign n31404 = ~n31396 & ~n31403 ;
  assign n31405 = ~n31395 & ~n31404 ;
  assign n31406 = ~n31088 & n31109 ;
  assign n31407 = n5211 & ~n12438 ;
  assign n31408 = ~n12436 & n31407 ;
  assign n31409 = \b[47]  & n5209 ;
  assign n31410 = \a[30]  & \b[46]  ;
  assign n31411 = n5200 & n31410 ;
  assign n31412 = ~n31409 & ~n31411 ;
  assign n31413 = \b[45]  & n5595 ;
  assign n31414 = n5592 & n31413 ;
  assign n31415 = ~\a[30]  & \b[46]  ;
  assign n31416 = n5203 & n31415 ;
  assign n31417 = ~n31414 & ~n31416 ;
  assign n31418 = n31412 & n31417 ;
  assign n31419 = ~n31408 & n31418 ;
  assign n31420 = ~\a[32]  & ~n31419 ;
  assign n31421 = ~n31089 & n31420 ;
  assign n31422 = ~n31406 & n31421 ;
  assign n31423 = \a[32]  & n31419 ;
  assign n31424 = ~n31089 & n31423 ;
  assign n31425 = ~n31406 & n31424 ;
  assign n31426 = ~n31422 & ~n31425 ;
  assign n31427 = \a[32]  & n31418 ;
  assign n31428 = ~n31408 & n31427 ;
  assign n31429 = n31089 & ~n31428 ;
  assign n31430 = n31109 & ~n31428 ;
  assign n31431 = ~n31088 & n31430 ;
  assign n31432 = ~n31429 & ~n31431 ;
  assign n31433 = ~n31420 & ~n31432 ;
  assign n31434 = n31426 & ~n31433 ;
  assign n31435 = ~n30983 & n31007 ;
  assign n31436 = n31012 & ~n31435 ;
  assign n31437 = ~n1694 & n20521 ;
  assign n31438 = ~n1692 & n31437 ;
  assign n31439 = \b[17]  & n20519 ;
  assign n31440 = \a[60]  & \b[16]  ;
  assign n31441 = n20510 & n31440 ;
  assign n31442 = ~n31439 & ~n31441 ;
  assign n31443 = \b[15]  & n21315 ;
  assign n31444 = n21312 & n31443 ;
  assign n31445 = ~\a[60]  & \b[16]  ;
  assign n31446 = n20513 & n31445 ;
  assign n31447 = ~n31444 & ~n31446 ;
  assign n31448 = n31442 & n31447 ;
  assign n31449 = ~n31438 & n31448 ;
  assign n31450 = ~\a[62]  & ~n31449 ;
  assign n31451 = \b[14]  & n21958 ;
  assign n31452 = \b[13]  & n21957 ;
  assign n31453 = ~n31451 & ~n31452 ;
  assign n31454 = n30811 & ~n31453 ;
  assign n31455 = ~n30811 & n31453 ;
  assign n31456 = ~n31454 & ~n31455 ;
  assign n31457 = \a[62]  & n31448 ;
  assign n31458 = ~n31438 & n31457 ;
  assign n31459 = ~n31456 & ~n31458 ;
  assign n31460 = ~n31450 & n31459 ;
  assign n31461 = ~\a[62]  & n31456 ;
  assign n31462 = ~n31449 & n31461 ;
  assign n31463 = ~n30812 & ~n30822 ;
  assign n31464 = ~n30817 & n31463 ;
  assign n31465 = \a[62]  & n31456 ;
  assign n31466 = n31448 & n31465 ;
  assign n31467 = ~n31438 & n31466 ;
  assign n31468 = ~n31464 & ~n31467 ;
  assign n31469 = ~n31462 & n31468 ;
  assign n31470 = ~n31460 & n31469 ;
  assign n31471 = ~n31462 & ~n31467 ;
  assign n31472 = ~n31460 & n31471 ;
  assign n31473 = n31464 & ~n31472 ;
  assign n31474 = ~n31470 & ~n31473 ;
  assign n31475 = n2293 & n18516 ;
  assign n31476 = ~n19247 & n31475 ;
  assign n31477 = n5705 & n18516 ;
  assign n31478 = ~n2289 & n31477 ;
  assign n31479 = \b[20]  & n18514 ;
  assign n31480 = \a[56]  & \b[19]  ;
  assign n31481 = n19181 & n31480 ;
  assign n31482 = ~\a[57]  & \b[19]  ;
  assign n31483 = n18508 & n31482 ;
  assign n31484 = ~n31481 & ~n31483 ;
  assign n31485 = ~n31479 & n31484 ;
  assign n31486 = \b[18]  & n19183 ;
  assign n31487 = n19180 & n31486 ;
  assign n31488 = \a[59]  & ~n31487 ;
  assign n31489 = n31485 & n31488 ;
  assign n31490 = ~n31478 & n31489 ;
  assign n31491 = ~n31476 & n31490 ;
  assign n31492 = n31485 & ~n31487 ;
  assign n31493 = ~n31478 & n31492 ;
  assign n31494 = ~n31476 & n31493 ;
  assign n31495 = ~\a[59]  & ~n31494 ;
  assign n31496 = ~n31491 & ~n31495 ;
  assign n31497 = n31474 & ~n31496 ;
  assign n31498 = ~n31474 & n31496 ;
  assign n31499 = ~n31497 & ~n31498 ;
  assign n31500 = ~n30833 & n30857 ;
  assign n31501 = ~n30832 & ~n31500 ;
  assign n31502 = ~n31499 & ~n31501 ;
  assign n31503 = n31499 & n31501 ;
  assign n31504 = ~n31502 & ~n31503 ;
  assign n31505 = ~n3022 & n16655 ;
  assign n31506 = ~n3020 & n31505 ;
  assign n31507 = \b[23]  & n16653 ;
  assign n31508 = \a[54]  & \b[22]  ;
  assign n31509 = n16644 & n31508 ;
  assign n31510 = ~\a[54]  & \b[22]  ;
  assign n31511 = n16647 & n31510 ;
  assign n31512 = ~n31509 & ~n31511 ;
  assign n31513 = ~n31507 & n31512 ;
  assign n31514 = \b[21]  & n17308 ;
  assign n31515 = n17305 & n31514 ;
  assign n31516 = \a[56]  & ~n31515 ;
  assign n31517 = n31513 & n31516 ;
  assign n31518 = ~n31506 & n31517 ;
  assign n31519 = n31513 & ~n31515 ;
  assign n31520 = ~n31506 & n31519 ;
  assign n31521 = ~\a[56]  & ~n31520 ;
  assign n31522 = ~n31518 & ~n31521 ;
  assign n31523 = ~n31504 & n31522 ;
  assign n31524 = n31504 & ~n31522 ;
  assign n31525 = ~n31523 & ~n31524 ;
  assign n31526 = n3604 & n14793 ;
  assign n31527 = ~n19292 & n31526 ;
  assign n31528 = ~n3604 & n14793 ;
  assign n31529 = ~n3562 & n31528 ;
  assign n31530 = ~n3600 & n31529 ;
  assign n31531 = \b[24]  & n15517 ;
  assign n31532 = n15514 & n31531 ;
  assign n31533 = ~\a[51]  & \b[25]  ;
  assign n31534 = n14785 & n31533 ;
  assign n31535 = ~n31532 & ~n31534 ;
  assign n31536 = \b[26]  & n14791 ;
  assign n31537 = \a[51]  & \b[25]  ;
  assign n31538 = n14782 & n31537 ;
  assign n31539 = \a[53]  & ~n31538 ;
  assign n31540 = ~n31536 & n31539 ;
  assign n31541 = n31535 & n31540 ;
  assign n31542 = ~n31530 & n31541 ;
  assign n31543 = ~n31527 & n31542 ;
  assign n31544 = ~n31536 & ~n31538 ;
  assign n31545 = n31535 & n31544 ;
  assign n31546 = ~n31530 & n31545 ;
  assign n31547 = ~n31527 & n31546 ;
  assign n31548 = ~\a[53]  & ~n31547 ;
  assign n31549 = ~n31543 & ~n31548 ;
  assign n31550 = ~n30862 & n30884 ;
  assign n31551 = ~n30861 & ~n31550 ;
  assign n31552 = ~n31549 & ~n31551 ;
  assign n31553 = n31525 & n31552 ;
  assign n31554 = ~n31549 & n31551 ;
  assign n31555 = ~n31525 & n31554 ;
  assign n31556 = ~n31553 & ~n31555 ;
  assign n31557 = n31549 & ~n31551 ;
  assign n31558 = ~n31525 & n31557 ;
  assign n31559 = n31549 & n31551 ;
  assign n31560 = n31525 & n31559 ;
  assign n31561 = ~n31558 & ~n31560 ;
  assign n31562 = n31556 & n31561 ;
  assign n31563 = ~n30889 & n30914 ;
  assign n31564 = ~n30888 & ~n31563 ;
  assign n31565 = n31562 & n31564 ;
  assign n31566 = ~n31562 & ~n31564 ;
  assign n31567 = ~n31565 & ~n31566 ;
  assign n31568 = ~n4502 & n13125 ;
  assign n31569 = ~n4500 & n31568 ;
  assign n31570 = \b[27]  & n13794 ;
  assign n31571 = n13792 & n31570 ;
  assign n31572 = ~\a[48]  & \b[28]  ;
  assign n31573 = n13117 & n31572 ;
  assign n31574 = ~n31571 & ~n31573 ;
  assign n31575 = \b[29]  & n13123 ;
  assign n31576 = \a[48]  & \b[28]  ;
  assign n31577 = n13786 & n31576 ;
  assign n31578 = \a[50]  & ~n31577 ;
  assign n31579 = ~n31575 & n31578 ;
  assign n31580 = n31574 & n31579 ;
  assign n31581 = ~n31569 & n31580 ;
  assign n31582 = ~n31575 & ~n31577 ;
  assign n31583 = n31574 & n31582 ;
  assign n31584 = ~n31569 & n31583 ;
  assign n31585 = ~\a[50]  & ~n31584 ;
  assign n31586 = ~n31581 & ~n31585 ;
  assign n31587 = n31567 & ~n31586 ;
  assign n31588 = ~n31567 & n31586 ;
  assign n31589 = ~n31587 & ~n31588 ;
  assign n31590 = ~n5810 & ~n10988 ;
  assign n31591 = ~n11569 & n31590 ;
  assign n31592 = n5807 & n31591 ;
  assign n31593 = n5810 & ~n10988 ;
  assign n31594 = ~n11569 & n31593 ;
  assign n31595 = ~n5807 & n31594 ;
  assign n31596 = ~n31592 & ~n31595 ;
  assign n31597 = \b[30]  & n12159 ;
  assign n31598 = n12156 & n31597 ;
  assign n31599 = ~\a[45]  & \b[31]  ;
  assign n31600 = n11564 & n31599 ;
  assign n31601 = ~n31598 & ~n31600 ;
  assign n31602 = \b[32]  & n11570 ;
  assign n31603 = \a[45]  & \b[31]  ;
  assign n31604 = n11561 & n31603 ;
  assign n31605 = \a[47]  & ~n31604 ;
  assign n31606 = ~n31602 & n31605 ;
  assign n31607 = n31601 & n31606 ;
  assign n31608 = n31596 & n31607 ;
  assign n31609 = ~n31602 & ~n31604 ;
  assign n31610 = n31601 & n31609 ;
  assign n31611 = n31596 & n31610 ;
  assign n31612 = ~\a[47]  & ~n31611 ;
  assign n31613 = ~n31608 & ~n31612 ;
  assign n31614 = ~n30919 & n30943 ;
  assign n31615 = n30918 & ~n30919 ;
  assign n31616 = ~n31614 & ~n31615 ;
  assign n31617 = n31613 & n31616 ;
  assign n31618 = ~n31589 & n31617 ;
  assign n31619 = n31613 & ~n31616 ;
  assign n31620 = n31589 & n31619 ;
  assign n31621 = ~n31618 & ~n31620 ;
  assign n31622 = ~n31613 & ~n31616 ;
  assign n31623 = ~n31589 & n31622 ;
  assign n31624 = ~n31613 & n31616 ;
  assign n31625 = n31589 & n31624 ;
  assign n31626 = ~n31623 & ~n31625 ;
  assign n31627 = n31621 & n31626 ;
  assign n31628 = ~n30946 & ~n30972 ;
  assign n31629 = ~n30943 & n30970 ;
  assign n31630 = n30920 & n31629 ;
  assign n31631 = n30943 & n30970 ;
  assign n31632 = ~n30920 & n31631 ;
  assign n31633 = ~n31630 & ~n31632 ;
  assign n31634 = ~n30975 & n31633 ;
  assign n31635 = ~n31628 & n31634 ;
  assign n31636 = ~n6610 & n10082 ;
  assign n31637 = ~n6608 & n31636 ;
  assign n31638 = \b[35]  & n10080 ;
  assign n31639 = \a[41]  & \b[34]  ;
  assign n31640 = n10679 & n31639 ;
  assign n31641 = ~\a[42]  & \b[34]  ;
  assign n31642 = n10074 & n31641 ;
  assign n31643 = ~n31640 & ~n31642 ;
  assign n31644 = ~n31638 & n31643 ;
  assign n31645 = \b[33]  & n10681 ;
  assign n31646 = n10678 & n31645 ;
  assign n31647 = \a[44]  & ~n31646 ;
  assign n31648 = n31644 & n31647 ;
  assign n31649 = ~n31637 & n31648 ;
  assign n31650 = n31644 & ~n31646 ;
  assign n31651 = ~n31637 & n31650 ;
  assign n31652 = ~\a[44]  & ~n31651 ;
  assign n31653 = ~n31649 & ~n31652 ;
  assign n31654 = ~n31635 & ~n31653 ;
  assign n31655 = ~n31627 & n31654 ;
  assign n31656 = n31635 & ~n31653 ;
  assign n31657 = n31627 & n31656 ;
  assign n31658 = ~n31655 & ~n31657 ;
  assign n31659 = n31635 & n31653 ;
  assign n31660 = ~n31627 & n31659 ;
  assign n31661 = ~n31635 & n31653 ;
  assign n31662 = n31627 & n31661 ;
  assign n31663 = ~n31660 & ~n31662 ;
  assign n31664 = n31658 & n31663 ;
  assign n31665 = n31436 & ~n31664 ;
  assign n31666 = ~n31436 & n31664 ;
  assign n31667 = ~n31665 & ~n31666 ;
  assign n31668 = n8175 & n8759 ;
  assign n31669 = ~n8172 & n31668 ;
  assign n31670 = n8759 & n25622 ;
  assign n31671 = ~n8171 & n31670 ;
  assign n31672 = \b[36]  & n9301 ;
  assign n31673 = n9298 & n31672 ;
  assign n31674 = ~\a[39]  & \b[37]  ;
  assign n31675 = n8751 & n31674 ;
  assign n31676 = ~n31673 & ~n31675 ;
  assign n31677 = \b[38]  & n8757 ;
  assign n31678 = \a[39]  & \b[37]  ;
  assign n31679 = n8748 & n31678 ;
  assign n31680 = \a[41]  & ~n31679 ;
  assign n31681 = ~n31677 & n31680 ;
  assign n31682 = n31676 & n31681 ;
  assign n31683 = ~n31671 & n31682 ;
  assign n31684 = ~n31669 & n31683 ;
  assign n31685 = ~n31677 & ~n31679 ;
  assign n31686 = n31676 & n31685 ;
  assign n31687 = ~n31671 & n31686 ;
  assign n31688 = ~n31669 & n31687 ;
  assign n31689 = ~\a[41]  & ~n31688 ;
  assign n31690 = ~n31684 & ~n31689 ;
  assign n31691 = ~n31667 & n31690 ;
  assign n31692 = n31667 & ~n31690 ;
  assign n31693 = ~n31691 & ~n31692 ;
  assign n31694 = n7534 & ~n9482 ;
  assign n31695 = ~n9480 & n31694 ;
  assign n31696 = \b[39]  & n7973 ;
  assign n31697 = n7970 & n31696 ;
  assign n31698 = ~\a[36]  & \b[40]  ;
  assign n31699 = n7526 & n31698 ;
  assign n31700 = ~n31697 & ~n31699 ;
  assign n31701 = \b[41]  & n7532 ;
  assign n31702 = \a[36]  & \b[40]  ;
  assign n31703 = n17801 & n31702 ;
  assign n31704 = \a[38]  & ~n31703 ;
  assign n31705 = ~n31701 & n31704 ;
  assign n31706 = n31700 & n31705 ;
  assign n31707 = ~n31695 & n31706 ;
  assign n31708 = ~n31701 & ~n31703 ;
  assign n31709 = n31700 & n31708 ;
  assign n31710 = ~n31695 & n31709 ;
  assign n31711 = ~\a[38]  & ~n31710 ;
  assign n31712 = ~n31707 & ~n31711 ;
  assign n31713 = ~n31018 & ~n31039 ;
  assign n31714 = n31018 & n31039 ;
  assign n31715 = n31037 & ~n31714 ;
  assign n31716 = ~n31713 & ~n31715 ;
  assign n31717 = n31712 & n31716 ;
  assign n31718 = ~n31693 & n31717 ;
  assign n31719 = n31712 & ~n31716 ;
  assign n31720 = n31693 & n31719 ;
  assign n31721 = ~n31718 & ~n31720 ;
  assign n31722 = ~n31712 & ~n31716 ;
  assign n31723 = ~n31693 & n31722 ;
  assign n31724 = ~n31712 & n31716 ;
  assign n31725 = n31693 & n31724 ;
  assign n31726 = ~n31723 & ~n31725 ;
  assign n31727 = n31721 & n31726 ;
  assign n31728 = n6309 & ~n28007 ;
  assign n31729 = ~n28005 & n31728 ;
  assign n31730 = \b[42]  & n6778 ;
  assign n31731 = n6775 & n31730 ;
  assign n31732 = ~\a[33]  & \b[43]  ;
  assign n31733 = n6301 & n31732 ;
  assign n31734 = ~n31731 & ~n31733 ;
  assign n31735 = \b[44]  & n6307 ;
  assign n31736 = \a[33]  & \b[43]  ;
  assign n31737 = n6298 & n31736 ;
  assign n31738 = \a[35]  & ~n31737 ;
  assign n31739 = ~n31735 & n31738 ;
  assign n31740 = n31734 & n31739 ;
  assign n31741 = ~n31729 & n31740 ;
  assign n31742 = ~n31735 & ~n31737 ;
  assign n31743 = n31734 & n31742 ;
  assign n31744 = ~n31729 & n31743 ;
  assign n31745 = ~\a[35]  & ~n31744 ;
  assign n31746 = ~n31741 & ~n31745 ;
  assign n31747 = ~n31050 & n31076 ;
  assign n31748 = n31081 & ~n31747 ;
  assign n31749 = n31746 & n31748 ;
  assign n31750 = ~n31727 & n31749 ;
  assign n31751 = n31746 & ~n31748 ;
  assign n31752 = n31727 & n31751 ;
  assign n31753 = ~n31750 & ~n31752 ;
  assign n31754 = ~n31746 & ~n31748 ;
  assign n31755 = ~n31727 & n31754 ;
  assign n31756 = ~n31746 & n31748 ;
  assign n31757 = n31727 & n31756 ;
  assign n31758 = ~n31755 & ~n31757 ;
  assign n31759 = n31753 & n31758 ;
  assign n31760 = n31434 & ~n31759 ;
  assign n31761 = ~n31434 & n31759 ;
  assign n31762 = ~n31760 & ~n31761 ;
  assign n31763 = n31405 & n31762 ;
  assign n31764 = ~n31405 & ~n31762 ;
  assign n31765 = ~n31763 & ~n31764 ;
  assign n31766 = n31371 & ~n31765 ;
  assign n31767 = ~n31371 & n31765 ;
  assign n31768 = ~n31766 & ~n31767 ;
  assign n31769 = n31345 & ~n31768 ;
  assign n31770 = ~n31345 & n31768 ;
  assign n31771 = ~n31769 & ~n31770 ;
  assign n31772 = n31313 & n31771 ;
  assign n31773 = ~n31313 & ~n31771 ;
  assign n31774 = ~n31772 & ~n31773 ;
  assign n31775 = ~n30714 & ~n31192 ;
  assign n31776 = n1467 & n21696 ;
  assign n31777 = ~n21693 & n31776 ;
  assign n31778 = n1467 & ~n21696 ;
  assign n31779 = ~n20966 & n31778 ;
  assign n31780 = ~n21692 & n31779 ;
  assign n31781 = \b[62]  & n1465 ;
  assign n31782 = \a[15]  & \b[61]  ;
  assign n31783 = n1456 & n31782 ;
  assign n31784 = ~n31781 & ~n31783 ;
  assign n31785 = \b[60]  & n1652 ;
  assign n31786 = n1649 & n31785 ;
  assign n31787 = ~\a[15]  & \b[61]  ;
  assign n31788 = n1459 & n31787 ;
  assign n31789 = ~n31786 & ~n31788 ;
  assign n31790 = n31784 & n31789 ;
  assign n31791 = ~n31780 & n31790 ;
  assign n31792 = ~n31777 & n31791 ;
  assign n31793 = \a[17]  & ~n31792 ;
  assign n31794 = ~\a[17]  & n31792 ;
  assign n31795 = ~n31793 & ~n31794 ;
  assign n31796 = ~n31775 & n31795 ;
  assign n31797 = ~\a[17]  & ~n31792 ;
  assign n31798 = \a[17]  & n31790 ;
  assign n31799 = ~n31780 & n31798 ;
  assign n31800 = ~n31777 & n31799 ;
  assign n31801 = ~n31797 & ~n31800 ;
  assign n31802 = ~n30714 & n31801 ;
  assign n31803 = ~n31192 & n31802 ;
  assign n31804 = ~n31796 & ~n31803 ;
  assign n31805 = n31774 & n31804 ;
  assign n31806 = ~n31774 & ~n31804 ;
  assign n31807 = ~n31805 & ~n31806 ;
  assign n31808 = n31198 & ~n31285 ;
  assign n31809 = ~n31222 & n31808 ;
  assign n31810 = n31217 & ~n31285 ;
  assign n31811 = ~n31809 & ~n31810 ;
  assign n31812 = n31807 & n31811 ;
  assign n31813 = ~n31286 & n31812 ;
  assign n31814 = ~n31285 & ~n31807 ;
  assign n31815 = n31269 & n31814 ;
  assign n31816 = n31285 & ~n31807 ;
  assign n31817 = ~n31269 & n31816 ;
  assign n31818 = ~n31815 & ~n31817 ;
  assign n31819 = ~n31813 & n31818 ;
  assign n31820 = ~n31266 & n31819 ;
  assign n31821 = ~n31265 & n31820 ;
  assign n31822 = ~n31265 & ~n31266 ;
  assign n31823 = ~n31819 & ~n31822 ;
  assign n31824 = ~n31821 & ~n31823 ;
  assign n31825 = ~n31256 & n31824 ;
  assign n31826 = ~n31263 & n31825 ;
  assign n31827 = ~n31256 & ~n31263 ;
  assign n31828 = ~n31824 & ~n31827 ;
  assign n31829 = ~n31826 & ~n31828 ;
  assign n31830 = ~n31312 & ~n31771 ;
  assign n31831 = n31308 & n31310 ;
  assign n31832 = n31309 & n31310 ;
  assign n31833 = ~n31831 & ~n31832 ;
  assign n31834 = ~n31830 & n31833 ;
  assign n31835 = ~n31344 & n31768 ;
  assign n31836 = n31339 & ~n31344 ;
  assign n31837 = ~n31835 & ~n31836 ;
  assign n31838 = n2622 & ~n17690 ;
  assign n31839 = ~n17688 & n31838 ;
  assign n31840 = \b[55]  & n2912 ;
  assign n31841 = n2909 & n31840 ;
  assign n31842 = \b[57]  & n2620 ;
  assign n31843 = \a[20]  & \b[56]  ;
  assign n31844 = n2910 & n31843 ;
  assign n31845 = ~\a[21]  & \b[56]  ;
  assign n31846 = n2614 & n31845 ;
  assign n31847 = ~n31844 & ~n31846 ;
  assign n31848 = ~n31842 & n31847 ;
  assign n31849 = ~n31841 & n31848 ;
  assign n31850 = ~n31839 & n31849 ;
  assign n31851 = ~\a[23]  & ~n31850 ;
  assign n31852 = \a[23]  & n31849 ;
  assign n31853 = ~n31839 & n31852 ;
  assign n31854 = ~n31851 & ~n31853 ;
  assign n31855 = n31837 & ~n31854 ;
  assign n31856 = ~n31344 & n31854 ;
  assign n31857 = n31768 & n31856 ;
  assign n31858 = n31339 & n31856 ;
  assign n31859 = ~n31857 & ~n31858 ;
  assign n31860 = ~n31855 & n31859 ;
  assign n31861 = n1965 & n20260 ;
  assign n31862 = ~n20257 & n31861 ;
  assign n31863 = n1965 & ~n20260 ;
  assign n31864 = ~n19545 & n31863 ;
  assign n31865 = ~n20256 & n31864 ;
  assign n31866 = \b[58]  & n2218 ;
  assign n31867 = n2216 & n31866 ;
  assign n31868 = ~\a[18]  & \b[59]  ;
  assign n31869 = n1957 & n31868 ;
  assign n31870 = ~n31867 & ~n31869 ;
  assign n31871 = \b[60]  & n1963 ;
  assign n31872 = \a[18]  & \b[59]  ;
  assign n31873 = n28047 & n31872 ;
  assign n31874 = \a[20]  & ~n31873 ;
  assign n31875 = ~n31871 & n31874 ;
  assign n31876 = n31870 & n31875 ;
  assign n31877 = ~n31865 & n31876 ;
  assign n31878 = ~n31862 & n31877 ;
  assign n31879 = ~n31871 & ~n31873 ;
  assign n31880 = n31870 & n31879 ;
  assign n31881 = ~n31865 & n31880 ;
  assign n31882 = ~n31862 & n31881 ;
  assign n31883 = ~\a[20]  & ~n31882 ;
  assign n31884 = ~n31878 & ~n31883 ;
  assign n31885 = ~n31370 & ~n31765 ;
  assign n31886 = ~n31365 & ~n31885 ;
  assign n31887 = n4249 & ~n14098 ;
  assign n31888 = ~n14096 & n31887 ;
  assign n31889 = \b[51]  & n4247 ;
  assign n31890 = \a[27]  & \b[50]  ;
  assign n31891 = n4238 & n31890 ;
  assign n31892 = ~n31889 & ~n31891 ;
  assign n31893 = \b[49]  & n4647 ;
  assign n31894 = n4644 & n31893 ;
  assign n31895 = ~\a[27]  & \b[50]  ;
  assign n31896 = n4241 & n31895 ;
  assign n31897 = ~n31894 & ~n31896 ;
  assign n31898 = n31892 & n31897 ;
  assign n31899 = ~n31888 & n31898 ;
  assign n31900 = ~\a[29]  & ~n31899 ;
  assign n31901 = \a[29]  & n31898 ;
  assign n31902 = ~n31888 & n31901 ;
  assign n31903 = ~n31900 & ~n31902 ;
  assign n31904 = ~n31395 & ~n31762 ;
  assign n31905 = ~n31404 & ~n31904 ;
  assign n31906 = n31903 & ~n31905 ;
  assign n31907 = ~n31404 & ~n31903 ;
  assign n31908 = ~n31904 & n31907 ;
  assign n31909 = ~n31906 & ~n31908 ;
  assign n31910 = n3402 & ~n16398 ;
  assign n31911 = ~n15241 & n31910 ;
  assign n31912 = ~n16404 & n31911 ;
  assign n31913 = n3402 & n16398 ;
  assign n31914 = n15241 & n31913 ;
  assign n31915 = n16400 & n31913 ;
  assign n31916 = ~n15239 & n31915 ;
  assign n31917 = ~n31914 & ~n31916 ;
  assign n31918 = ~n31912 & n31917 ;
  assign n31919 = \b[52]  & n3733 ;
  assign n31920 = n3730 & n31919 ;
  assign n31921 = ~\a[24]  & \b[53]  ;
  assign n31922 = n3394 & n31921 ;
  assign n31923 = ~n31920 & ~n31922 ;
  assign n31924 = \b[54]  & n3400 ;
  assign n31925 = \a[24]  & \b[53]  ;
  assign n31926 = n27626 & n31925 ;
  assign n31927 = \a[26]  & ~n31926 ;
  assign n31928 = ~n31924 & n31927 ;
  assign n31929 = n31923 & n31928 ;
  assign n31930 = n31918 & n31929 ;
  assign n31931 = ~n31924 & ~n31926 ;
  assign n31932 = n31923 & n31931 ;
  assign n31933 = n31918 & n31932 ;
  assign n31934 = ~\a[26]  & ~n31933 ;
  assign n31935 = ~n31930 & ~n31934 ;
  assign n31936 = ~n31693 & ~n31716 ;
  assign n31937 = n31693 & n31716 ;
  assign n31938 = n31712 & ~n31937 ;
  assign n31939 = ~n31936 & ~n31938 ;
  assign n31940 = n31525 & n31551 ;
  assign n31941 = n31556 & ~n31940 ;
  assign n31942 = ~n4148 & n14793 ;
  assign n31943 = ~n4146 & n31942 ;
  assign n31944 = \b[27]  & n14791 ;
  assign n31945 = \a[51]  & \b[26]  ;
  assign n31946 = n14782 & n31945 ;
  assign n31947 = ~n31944 & ~n31946 ;
  assign n31948 = \b[25]  & n15517 ;
  assign n31949 = n15514 & n31948 ;
  assign n31950 = ~\a[51]  & \b[26]  ;
  assign n31951 = n14785 & n31950 ;
  assign n31952 = ~n31949 & ~n31951 ;
  assign n31953 = n31947 & n31952 ;
  assign n31954 = ~n31943 & n31953 ;
  assign n31955 = ~\a[53]  & ~n31954 ;
  assign n31956 = \a[53]  & n31953 ;
  assign n31957 = ~n31943 & n31956 ;
  assign n31958 = ~n31955 & ~n31957 ;
  assign n31959 = ~n31503 & n31522 ;
  assign n31960 = ~n31502 & ~n31959 ;
  assign n31961 = ~n31470 & n31496 ;
  assign n31962 = ~n31473 & ~n31961 ;
  assign n31963 = ~n2520 & n18516 ;
  assign n31964 = ~n2292 & n18516 ;
  assign n31965 = ~n2516 & n31964 ;
  assign n31966 = ~n31963 & ~n31965 ;
  assign n31967 = ~n2523 & ~n31966 ;
  assign n31968 = \b[21]  & n18514 ;
  assign n31969 = \a[56]  & \b[20]  ;
  assign n31970 = n19181 & n31969 ;
  assign n31971 = ~\a[57]  & \b[20]  ;
  assign n31972 = n18508 & n31971 ;
  assign n31973 = ~n31970 & ~n31972 ;
  assign n31974 = ~n31968 & n31973 ;
  assign n31975 = \b[19]  & n19183 ;
  assign n31976 = n19180 & n31975 ;
  assign n31977 = \a[59]  & ~n31976 ;
  assign n31978 = n31974 & n31977 ;
  assign n31979 = ~n31967 & n31978 ;
  assign n31980 = n31974 & ~n31976 ;
  assign n31981 = ~\a[59]  & ~n31980 ;
  assign n31982 = ~\a[59]  & ~n2523 ;
  assign n31983 = ~n31966 & n31982 ;
  assign n31984 = ~n31981 & ~n31983 ;
  assign n31985 = ~n31979 & n31984 ;
  assign n31986 = ~n31454 & ~n31467 ;
  assign n31987 = ~n31462 & n31986 ;
  assign n31988 = n1875 & n20521 ;
  assign n31989 = ~n1872 & n31988 ;
  assign n31990 = ~n1875 & n20521 ;
  assign n31991 = ~n1689 & n31990 ;
  assign n31992 = ~n1871 & n31991 ;
  assign n31993 = \b[18]  & n20519 ;
  assign n31994 = \a[60]  & \b[17]  ;
  assign n31995 = n20510 & n31994 ;
  assign n31996 = ~n31993 & ~n31995 ;
  assign n31997 = \b[16]  & n21315 ;
  assign n31998 = n21312 & n31997 ;
  assign n31999 = ~\a[60]  & \b[17]  ;
  assign n32000 = n20513 & n31999 ;
  assign n32001 = ~n31998 & ~n32000 ;
  assign n32002 = n31996 & n32001 ;
  assign n32003 = ~n31992 & n32002 ;
  assign n32004 = ~n31989 & n32003 ;
  assign n32005 = ~\a[14]  & \b[14]  ;
  assign n32006 = n21957 & n32005 ;
  assign n32007 = ~\a[14]  & \b[15]  ;
  assign n32008 = n21958 & n32007 ;
  assign n32009 = ~n32006 & ~n32008 ;
  assign n32010 = \b[15]  & n21958 ;
  assign n32011 = \b[14]  & n21957 ;
  assign n32012 = \a[14]  & ~n32011 ;
  assign n32013 = ~n32010 & n32012 ;
  assign n32014 = n32009 & ~n32013 ;
  assign n32015 = ~\a[62]  & ~n30811 ;
  assign n32016 = ~n32014 & n32015 ;
  assign n32017 = ~\a[62]  & n30811 ;
  assign n32018 = n32014 & n32017 ;
  assign n32019 = ~n32016 & ~n32018 ;
  assign n32020 = ~n32004 & ~n32019 ;
  assign n32021 = \a[62]  & ~n30811 ;
  assign n32022 = ~n32014 & n32021 ;
  assign n32023 = \a[62]  & n30811 ;
  assign n32024 = n32014 & n32023 ;
  assign n32025 = ~n32022 & ~n32024 ;
  assign n32026 = n32002 & ~n32025 ;
  assign n32027 = ~n31992 & n32026 ;
  assign n32028 = ~n31989 & n32027 ;
  assign n32029 = ~n32020 & ~n32028 ;
  assign n32030 = ~\a[62]  & ~n32004 ;
  assign n32031 = n30811 & n32014 ;
  assign n32032 = ~n30811 & ~n32014 ;
  assign n32033 = ~n32031 & ~n32032 ;
  assign n32034 = \a[62]  & n32002 ;
  assign n32035 = ~n31992 & n32034 ;
  assign n32036 = ~n31989 & n32035 ;
  assign n32037 = n32033 & ~n32036 ;
  assign n32038 = ~n32030 & n32037 ;
  assign n32039 = n32029 & ~n32038 ;
  assign n32040 = ~n31987 & ~n32039 ;
  assign n32041 = n31987 & n32039 ;
  assign n32042 = ~n32040 & ~n32041 ;
  assign n32043 = n31985 & n32042 ;
  assign n32044 = ~n31985 & ~n32042 ;
  assign n32045 = ~n32043 & ~n32044 ;
  assign n32046 = n31962 & n32045 ;
  assign n32047 = ~n31962 & n32043 ;
  assign n32048 = ~n31962 & n32044 ;
  assign n32049 = ~n32047 & ~n32048 ;
  assign n32050 = ~n32046 & n32049 ;
  assign n32051 = ~n3283 & ~n16016 ;
  assign n32052 = ~n16652 & n32051 ;
  assign n32053 = n3280 & n32052 ;
  assign n32054 = n3283 & ~n16016 ;
  assign n32055 = ~n16652 & n32054 ;
  assign n32056 = ~n3280 & n32055 ;
  assign n32057 = ~n32053 & ~n32056 ;
  assign n32058 = \b[22]  & n17308 ;
  assign n32059 = n17305 & n32058 ;
  assign n32060 = \b[24]  & n16653 ;
  assign n32061 = \a[54]  & \b[23]  ;
  assign n32062 = n16644 & n32061 ;
  assign n32063 = ~\a[54]  & \b[23]  ;
  assign n32064 = n16647 & n32063 ;
  assign n32065 = ~n32062 & ~n32064 ;
  assign n32066 = ~n32060 & n32065 ;
  assign n32067 = ~n32059 & n32066 ;
  assign n32068 = n32057 & n32067 ;
  assign n32069 = ~\a[56]  & ~n32068 ;
  assign n32070 = \a[56]  & n32067 ;
  assign n32071 = n32057 & n32070 ;
  assign n32072 = ~n32069 & ~n32071 ;
  assign n32073 = ~n32050 & n32072 ;
  assign n32074 = n32050 & ~n32072 ;
  assign n32075 = ~n32073 & ~n32074 ;
  assign n32076 = ~n31960 & ~n32075 ;
  assign n32077 = n31960 & n32075 ;
  assign n32078 = ~n32076 & ~n32077 ;
  assign n32079 = ~n31958 & n32078 ;
  assign n32080 = n31958 & ~n32078 ;
  assign n32081 = ~n32079 & ~n32080 ;
  assign n32082 = n31941 & ~n32081 ;
  assign n32083 = ~n31941 & n32081 ;
  assign n32084 = ~n32082 & ~n32083 ;
  assign n32085 = ~n5105 & ~n12606 ;
  assign n32086 = ~n13122 & n32085 ;
  assign n32087 = n5102 & n32086 ;
  assign n32088 = n5105 & ~n12606 ;
  assign n32089 = ~n13122 & n32088 ;
  assign n32090 = ~n5102 & n32089 ;
  assign n32091 = ~n32087 & ~n32090 ;
  assign n32092 = \b[28]  & n13794 ;
  assign n32093 = n13792 & n32092 ;
  assign n32094 = ~\a[48]  & \b[29]  ;
  assign n32095 = n13117 & n32094 ;
  assign n32096 = ~n32093 & ~n32095 ;
  assign n32097 = \b[30]  & n13123 ;
  assign n32098 = \a[48]  & \b[29]  ;
  assign n32099 = n13786 & n32098 ;
  assign n32100 = \a[50]  & ~n32099 ;
  assign n32101 = ~n32097 & n32100 ;
  assign n32102 = n32096 & n32101 ;
  assign n32103 = n32091 & n32102 ;
  assign n32104 = ~n32097 & ~n32099 ;
  assign n32105 = n32096 & n32104 ;
  assign n32106 = n32091 & n32105 ;
  assign n32107 = ~\a[50]  & ~n32106 ;
  assign n32108 = ~n32103 & ~n32107 ;
  assign n32109 = n32084 & ~n32108 ;
  assign n32110 = ~n32084 & n32108 ;
  assign n32111 = ~n32109 & ~n32110 ;
  assign n32112 = ~n31565 & n31586 ;
  assign n32113 = ~n31566 & ~n32112 ;
  assign n32114 = ~n5855 & n11572 ;
  assign n32115 = ~n5853 & n32114 ;
  assign n32116 = \b[31]  & n12159 ;
  assign n32117 = n12156 & n32116 ;
  assign n32118 = ~\a[45]  & \b[32]  ;
  assign n32119 = n11564 & n32118 ;
  assign n32120 = ~n32117 & ~n32119 ;
  assign n32121 = \b[33]  & n11570 ;
  assign n32122 = \a[45]  & \b[32]  ;
  assign n32123 = n11561 & n32122 ;
  assign n32124 = \a[47]  & ~n32123 ;
  assign n32125 = ~n32121 & n32124 ;
  assign n32126 = n32120 & n32125 ;
  assign n32127 = ~n32115 & n32126 ;
  assign n32128 = ~n32121 & ~n32123 ;
  assign n32129 = n32120 & n32128 ;
  assign n32130 = ~n32115 & n32129 ;
  assign n32131 = ~\a[47]  & ~n32130 ;
  assign n32132 = ~n32127 & ~n32131 ;
  assign n32133 = ~n32113 & ~n32132 ;
  assign n32134 = n32111 & n32133 ;
  assign n32135 = n32113 & ~n32132 ;
  assign n32136 = ~n32111 & n32135 ;
  assign n32137 = ~n32134 & ~n32136 ;
  assign n32138 = ~n32113 & n32132 ;
  assign n32139 = ~n32111 & n32138 ;
  assign n32140 = n32113 & n32132 ;
  assign n32141 = n32111 & n32140 ;
  assign n32142 = ~n32139 & ~n32141 ;
  assign n32143 = n32137 & n32142 ;
  assign n32144 = n7337 & n10082 ;
  assign n32145 = ~n7334 & n32144 ;
  assign n32146 = ~n7337 & n10082 ;
  assign n32147 = ~n6605 & n32146 ;
  assign n32148 = ~n7333 & n32147 ;
  assign n32149 = \b[34]  & n10681 ;
  assign n32150 = n10678 & n32149 ;
  assign n32151 = \b[36]  & n10080 ;
  assign n32152 = \a[41]  & \b[35]  ;
  assign n32153 = n10679 & n32152 ;
  assign n32154 = ~\a[42]  & \b[35]  ;
  assign n32155 = n10074 & n32154 ;
  assign n32156 = ~n32153 & ~n32155 ;
  assign n32157 = ~n32151 & n32156 ;
  assign n32158 = ~n32150 & n32157 ;
  assign n32159 = ~n32148 & n32158 ;
  assign n32160 = ~n32145 & n32159 ;
  assign n32161 = ~\a[44]  & ~n32160 ;
  assign n32162 = \a[44]  & n32158 ;
  assign n32163 = ~n32148 & n32162 ;
  assign n32164 = ~n32145 & n32163 ;
  assign n32165 = ~n32161 & ~n32164 ;
  assign n32166 = ~n31589 & ~n31616 ;
  assign n32167 = n31589 & n31616 ;
  assign n32168 = n31613 & ~n32167 ;
  assign n32169 = ~n32166 & ~n32168 ;
  assign n32170 = ~n32165 & ~n32169 ;
  assign n32171 = n32143 & n32170 ;
  assign n32172 = ~n32165 & n32169 ;
  assign n32173 = ~n32143 & n32172 ;
  assign n32174 = ~n32171 & ~n32173 ;
  assign n32175 = n32165 & ~n32169 ;
  assign n32176 = ~n32143 & n32175 ;
  assign n32177 = n32165 & n32169 ;
  assign n32178 = n32143 & n32177 ;
  assign n32179 = ~n32176 & ~n32178 ;
  assign n32180 = n32174 & n32179 ;
  assign n32181 = n31627 & ~n31635 ;
  assign n32182 = ~n31627 & n31635 ;
  assign n32183 = n31653 & ~n32182 ;
  assign n32184 = ~n32181 & ~n32183 ;
  assign n32185 = ~n8602 & n8759 ;
  assign n32186 = ~n8600 & n32185 ;
  assign n32187 = \b[37]  & n9301 ;
  assign n32188 = n9298 & n32187 ;
  assign n32189 = ~\a[39]  & \b[38]  ;
  assign n32190 = n8751 & n32189 ;
  assign n32191 = ~n32188 & ~n32190 ;
  assign n32192 = \b[39]  & n8757 ;
  assign n32193 = \a[39]  & \b[38]  ;
  assign n32194 = n8748 & n32193 ;
  assign n32195 = \a[41]  & ~n32194 ;
  assign n32196 = ~n32192 & n32195 ;
  assign n32197 = n32191 & n32196 ;
  assign n32198 = ~n32186 & n32197 ;
  assign n32199 = ~n32192 & ~n32194 ;
  assign n32200 = n32191 & n32199 ;
  assign n32201 = ~n32186 & n32200 ;
  assign n32202 = ~\a[41]  & ~n32201 ;
  assign n32203 = ~n32198 & ~n32202 ;
  assign n32204 = ~n32184 & ~n32203 ;
  assign n32205 = n32180 & n32204 ;
  assign n32206 = n32184 & ~n32203 ;
  assign n32207 = ~n32180 & n32206 ;
  assign n32208 = ~n32205 & ~n32207 ;
  assign n32209 = ~n32184 & n32203 ;
  assign n32210 = ~n32180 & n32209 ;
  assign n32211 = n32184 & n32203 ;
  assign n32212 = n32180 & n32211 ;
  assign n32213 = ~n32210 & ~n32212 ;
  assign n32214 = n32208 & n32213 ;
  assign n32215 = n7534 & n9930 ;
  assign n32216 = ~n9927 & n32215 ;
  assign n32217 = n7534 & ~n9930 ;
  assign n32218 = ~n9477 & n32217 ;
  assign n32219 = ~n9926 & n32218 ;
  assign n32220 = \b[40]  & n7973 ;
  assign n32221 = n7970 & n32220 ;
  assign n32222 = ~\a[36]  & \b[41]  ;
  assign n32223 = n7526 & n32222 ;
  assign n32224 = ~n32221 & ~n32223 ;
  assign n32225 = \b[42]  & n7532 ;
  assign n32226 = \a[36]  & \b[41]  ;
  assign n32227 = n17801 & n32226 ;
  assign n32228 = \a[38]  & ~n32227 ;
  assign n32229 = ~n32225 & n32228 ;
  assign n32230 = n32224 & n32229 ;
  assign n32231 = ~n32219 & n32230 ;
  assign n32232 = ~n32216 & n32231 ;
  assign n32233 = ~n32225 & ~n32227 ;
  assign n32234 = n32224 & n32233 ;
  assign n32235 = ~n32219 & n32234 ;
  assign n32236 = ~n32216 & n32235 ;
  assign n32237 = ~\a[38]  & ~n32236 ;
  assign n32238 = ~n32232 & ~n32237 ;
  assign n32239 = ~n31666 & n31690 ;
  assign n32240 = n31665 & ~n31666 ;
  assign n32241 = ~n32239 & ~n32240 ;
  assign n32242 = ~n32238 & n32241 ;
  assign n32243 = ~n32214 & n32242 ;
  assign n32244 = ~n32238 & ~n32241 ;
  assign n32245 = n32214 & n32244 ;
  assign n32246 = ~n32243 & ~n32245 ;
  assign n32247 = n32238 & ~n32241 ;
  assign n32248 = ~n32214 & n32247 ;
  assign n32249 = n32238 & n32241 ;
  assign n32250 = n32214 & n32249 ;
  assign n32251 = ~n32248 & ~n32250 ;
  assign n32252 = n32246 & n32251 ;
  assign n32253 = ~n31939 & ~n32252 ;
  assign n32254 = n31939 & n32252 ;
  assign n32255 = ~n32253 & ~n32254 ;
  assign n32256 = n6309 & ~n11397 ;
  assign n32257 = ~n11395 & n32256 ;
  assign n32258 = \b[45]  & n6307 ;
  assign n32259 = \a[33]  & \b[44]  ;
  assign n32260 = n6298 & n32259 ;
  assign n32261 = ~n32258 & ~n32260 ;
  assign n32262 = \b[43]  & n6778 ;
  assign n32263 = n6775 & n32262 ;
  assign n32264 = ~\a[33]  & \b[44]  ;
  assign n32265 = n6301 & n32264 ;
  assign n32266 = ~n32263 & ~n32265 ;
  assign n32267 = n32261 & n32266 ;
  assign n32268 = ~n32257 & n32267 ;
  assign n32269 = ~\a[35]  & ~n32268 ;
  assign n32270 = \a[35]  & n32267 ;
  assign n32271 = ~n32257 & n32270 ;
  assign n32272 = ~n32269 & ~n32271 ;
  assign n32273 = n32255 & ~n32272 ;
  assign n32274 = ~n32255 & n32272 ;
  assign n32275 = ~n32273 & ~n32274 ;
  assign n32276 = n31727 & n31748 ;
  assign n32277 = ~n31727 & ~n31748 ;
  assign n32278 = n31746 & ~n32277 ;
  assign n32279 = ~n32276 & ~n32278 ;
  assign n32280 = ~n32275 & ~n32279 ;
  assign n32281 = n32275 & n32279 ;
  assign n32282 = ~n32280 & ~n32281 ;
  assign n32283 = n5211 & n12478 ;
  assign n32284 = ~n12475 & n32283 ;
  assign n32285 = n5211 & n28668 ;
  assign n32286 = ~n12474 & n32285 ;
  assign n32287 = \b[46]  & n5595 ;
  assign n32288 = n5592 & n32287 ;
  assign n32289 = ~\a[30]  & \b[47]  ;
  assign n32290 = n5203 & n32289 ;
  assign n32291 = ~n32288 & ~n32290 ;
  assign n32292 = \b[48]  & n5209 ;
  assign n32293 = \a[30]  & \b[47]  ;
  assign n32294 = n5200 & n32293 ;
  assign n32295 = \a[32]  & ~n32294 ;
  assign n32296 = ~n32292 & n32295 ;
  assign n32297 = n32291 & n32296 ;
  assign n32298 = ~n32286 & n32297 ;
  assign n32299 = ~n32284 & n32298 ;
  assign n32300 = ~n32292 & ~n32294 ;
  assign n32301 = n32291 & n32300 ;
  assign n32302 = ~n32286 & n32301 ;
  assign n32303 = ~n32284 & n32302 ;
  assign n32304 = ~\a[32]  & ~n32303 ;
  assign n32305 = ~n32299 & ~n32304 ;
  assign n32306 = n31426 & n31759 ;
  assign n32307 = ~n31433 & ~n32306 ;
  assign n32308 = ~n32305 & n32307 ;
  assign n32309 = ~n32282 & n32308 ;
  assign n32310 = ~n32305 & ~n32307 ;
  assign n32311 = n32282 & n32310 ;
  assign n32312 = ~n32309 & ~n32311 ;
  assign n32313 = n32305 & ~n32307 ;
  assign n32314 = ~n32282 & n32313 ;
  assign n32315 = n32305 & n32307 ;
  assign n32316 = n32282 & n32315 ;
  assign n32317 = ~n32314 & ~n32316 ;
  assign n32318 = n32312 & n32317 ;
  assign n32319 = ~n31935 & ~n32318 ;
  assign n32320 = n31909 & n32319 ;
  assign n32321 = ~n31935 & n32318 ;
  assign n32322 = ~n31909 & n32321 ;
  assign n32323 = ~n32320 & ~n32322 ;
  assign n32324 = ~n31886 & ~n32323 ;
  assign n32325 = n31935 & ~n32318 ;
  assign n32326 = n31909 & n32325 ;
  assign n32327 = n31935 & n32318 ;
  assign n32328 = ~n31909 & n32327 ;
  assign n32329 = ~n32326 & ~n32328 ;
  assign n32330 = n31886 & ~n32329 ;
  assign n32331 = ~n32324 & ~n32330 ;
  assign n32332 = n31909 & n32318 ;
  assign n32333 = ~n31909 & ~n32318 ;
  assign n32334 = ~n32332 & ~n32333 ;
  assign n32335 = ~n31886 & n31935 ;
  assign n32336 = ~n32334 & n32335 ;
  assign n32337 = ~n31909 & n32319 ;
  assign n32338 = n31909 & n32321 ;
  assign n32339 = ~n32337 & ~n32338 ;
  assign n32340 = n31886 & ~n32339 ;
  assign n32341 = ~n32336 & ~n32340 ;
  assign n32342 = n32331 & n32341 ;
  assign n32343 = n31884 & n32342 ;
  assign n32344 = ~n31860 & n32343 ;
  assign n32345 = n31884 & ~n32342 ;
  assign n32346 = n31860 & n32345 ;
  assign n32347 = ~n32344 & ~n32346 ;
  assign n32348 = n31834 & ~n32347 ;
  assign n32349 = ~n31884 & n32342 ;
  assign n32350 = ~n31860 & n32349 ;
  assign n32351 = ~n31884 & ~n32342 ;
  assign n32352 = n31860 & n32351 ;
  assign n32353 = ~n32350 & ~n32352 ;
  assign n32354 = ~n31834 & ~n32353 ;
  assign n32355 = ~n32348 & ~n32354 ;
  assign n32356 = ~n31860 & n32345 ;
  assign n32357 = n31860 & n32343 ;
  assign n32358 = ~n32356 & ~n32357 ;
  assign n32359 = ~n31834 & ~n32358 ;
  assign n32360 = ~n31860 & n32351 ;
  assign n32361 = n31860 & n32349 ;
  assign n32362 = ~n32360 & ~n32361 ;
  assign n32363 = n31834 & ~n32362 ;
  assign n32364 = ~n32359 & ~n32363 ;
  assign n32365 = n32355 & n32364 ;
  assign n32366 = n1467 & ~n22461 ;
  assign n32367 = ~n22459 & n32366 ;
  assign n32368 = \b[63]  & n1465 ;
  assign n32369 = \a[15]  & \b[62]  ;
  assign n32370 = n1456 & n32369 ;
  assign n32371 = ~n32368 & ~n32370 ;
  assign n32372 = \b[61]  & n1652 ;
  assign n32373 = n1649 & n32372 ;
  assign n32374 = ~\a[15]  & \b[62]  ;
  assign n32375 = n1459 & n32374 ;
  assign n32376 = ~n32373 & ~n32375 ;
  assign n32377 = n32371 & n32376 ;
  assign n32378 = ~n32367 & n32377 ;
  assign n32379 = ~\a[17]  & ~n32378 ;
  assign n32380 = \a[17]  & n32377 ;
  assign n32381 = ~n32367 & n32380 ;
  assign n32382 = ~n32379 & ~n32381 ;
  assign n32383 = n31796 & ~n32382 ;
  assign n32384 = ~n31803 & ~n32382 ;
  assign n32385 = n31774 & n32384 ;
  assign n32386 = ~n32383 & ~n32385 ;
  assign n32387 = n31774 & ~n31803 ;
  assign n32388 = ~n31796 & n32382 ;
  assign n32389 = ~n32387 & n32388 ;
  assign n32390 = n32386 & ~n32389 ;
  assign n32391 = n32365 & n32390 ;
  assign n32392 = ~n32365 & ~n32390 ;
  assign n32393 = ~n32391 & ~n32392 ;
  assign n32394 = n31811 & ~n32393 ;
  assign n32395 = ~n31813 & n32394 ;
  assign n32396 = n31811 & ~n31813 ;
  assign n32397 = n32393 & ~n32396 ;
  assign n32398 = ~n32395 & ~n32397 ;
  assign n32399 = n31821 & n32398 ;
  assign n32400 = n31824 & n32398 ;
  assign n32401 = ~n31256 & n32400 ;
  assign n32402 = ~n31263 & n32401 ;
  assign n32403 = ~n32399 & ~n32402 ;
  assign n32404 = ~n31821 & ~n32398 ;
  assign n32405 = ~n31826 & n32404 ;
  assign n32406 = n32403 & ~n32405 ;
  assign n32407 = ~n32365 & n32386 ;
  assign n32408 = ~n32389 & ~n32407 ;
  assign n32409 = ~n31834 & n31884 ;
  assign n32410 = n31860 & n32342 ;
  assign n32411 = ~n31834 & n32410 ;
  assign n32412 = ~n32409 & ~n32411 ;
  assign n32413 = ~n31860 & ~n32342 ;
  assign n32414 = ~n31834 & n32413 ;
  assign n32415 = n32358 & ~n32414 ;
  assign n32416 = n32412 & n32415 ;
  assign n32417 = \b[62]  & n1652 ;
  assign n32418 = n1649 & n32417 ;
  assign n32419 = ~\a[15]  & \b[63]  ;
  assign n32420 = n1459 & n32419 ;
  assign n32421 = \a[15]  & \b[63]  ;
  assign n32422 = n1456 & n32421 ;
  assign n32423 = ~n32420 & ~n32422 ;
  assign n32424 = ~n32418 & n32423 ;
  assign n32425 = ~\a[17]  & ~n32424 ;
  assign n32426 = n1467 & ~n22458 ;
  assign n32427 = ~\a[17]  & n32426 ;
  assign n32428 = ~n23173 & n32427 ;
  assign n32429 = ~n32425 & ~n32428 ;
  assign n32430 = ~n23173 & n32426 ;
  assign n32431 = \a[17]  & n32424 ;
  assign n32432 = ~n32430 & n32431 ;
  assign n32433 = n32429 & ~n32432 ;
  assign n32434 = n32416 & ~n32433 ;
  assign n32435 = ~n32416 & n32433 ;
  assign n32436 = ~n32434 & ~n32435 ;
  assign n32437 = ~n31855 & ~n32342 ;
  assign n32438 = n31859 & ~n32437 ;
  assign n32439 = n1965 & ~n20971 ;
  assign n32440 = ~n20969 & n32439 ;
  assign n32441 = \b[61]  & n1963 ;
  assign n32442 = \a[18]  & \b[60]  ;
  assign n32443 = n28047 & n32442 ;
  assign n32444 = ~n32441 & ~n32443 ;
  assign n32445 = \b[59]  & n2218 ;
  assign n32446 = n2216 & n32445 ;
  assign n32447 = ~\a[18]  & \b[60]  ;
  assign n32448 = n1957 & n32447 ;
  assign n32449 = ~n32446 & ~n32448 ;
  assign n32450 = n32444 & n32449 ;
  assign n32451 = ~n32440 & n32450 ;
  assign n32452 = ~\a[20]  & ~n32451 ;
  assign n32453 = \a[20]  & n32450 ;
  assign n32454 = ~n32440 & n32453 ;
  assign n32455 = ~n32452 & ~n32454 ;
  assign n32456 = ~n32438 & n32455 ;
  assign n32457 = \a[20]  & ~n32451 ;
  assign n32458 = ~\a[20]  & n32451 ;
  assign n32459 = ~n32457 & ~n32458 ;
  assign n32460 = n31859 & n32459 ;
  assign n32461 = ~n32437 & n32460 ;
  assign n32462 = ~n32456 & ~n32461 ;
  assign n32463 = ~n31886 & n32332 ;
  assign n32464 = ~n32335 & ~n32463 ;
  assign n32465 = ~n31886 & n32333 ;
  assign n32466 = ~n31909 & n32325 ;
  assign n32467 = n31909 & n32327 ;
  assign n32468 = ~n32466 & ~n32467 ;
  assign n32469 = ~n32465 & n32468 ;
  assign n32470 = n32464 & n32469 ;
  assign n32471 = n2622 & n18940 ;
  assign n32472 = ~n18937 & n32471 ;
  assign n32473 = n2622 & ~n18940 ;
  assign n32474 = ~n17685 & n32473 ;
  assign n32475 = ~n18936 & n32474 ;
  assign n32476 = \b[58]  & n2620 ;
  assign n32477 = \a[20]  & \b[57]  ;
  assign n32478 = n2910 & n32477 ;
  assign n32479 = ~\a[21]  & \b[57]  ;
  assign n32480 = n2614 & n32479 ;
  assign n32481 = ~n32478 & ~n32480 ;
  assign n32482 = ~n32476 & n32481 ;
  assign n32483 = \b[56]  & n2912 ;
  assign n32484 = n2909 & n32483 ;
  assign n32485 = \a[23]  & ~n32484 ;
  assign n32486 = n32482 & n32485 ;
  assign n32487 = ~n32475 & n32486 ;
  assign n32488 = ~n32472 & n32487 ;
  assign n32489 = n32482 & ~n32484 ;
  assign n32490 = ~n32475 & n32489 ;
  assign n32491 = ~n32472 & n32490 ;
  assign n32492 = ~\a[23]  & ~n32491 ;
  assign n32493 = ~n32488 & ~n32492 ;
  assign n32494 = ~n32470 & n32493 ;
  assign n32495 = n32470 & ~n32493 ;
  assign n32496 = n3402 & ~n16446 ;
  assign n32497 = ~n16444 & n32496 ;
  assign n32498 = \b[55]  & n3400 ;
  assign n32499 = \a[24]  & \b[54]  ;
  assign n32500 = n27626 & n32499 ;
  assign n32501 = ~n32498 & ~n32500 ;
  assign n32502 = \b[53]  & n3733 ;
  assign n32503 = n3730 & n32502 ;
  assign n32504 = ~\a[24]  & \b[54]  ;
  assign n32505 = n3394 & n32504 ;
  assign n32506 = ~n32503 & ~n32505 ;
  assign n32507 = n32501 & n32506 ;
  assign n32508 = ~n32497 & n32507 ;
  assign n32509 = ~\a[26]  & ~n32508 ;
  assign n32510 = \a[26]  & n32507 ;
  assign n32511 = ~n32497 & n32510 ;
  assign n32512 = n31906 & ~n32511 ;
  assign n32513 = ~n31908 & ~n32511 ;
  assign n32514 = ~n32318 & n32513 ;
  assign n32515 = ~n32512 & ~n32514 ;
  assign n32516 = ~n32509 & ~n32515 ;
  assign n32517 = ~n31908 & ~n32318 ;
  assign n32518 = \a[26]  & ~n32508 ;
  assign n32519 = ~\a[26]  & n32508 ;
  assign n32520 = ~n32518 & ~n32519 ;
  assign n32521 = ~n31906 & n32520 ;
  assign n32522 = ~n32517 & n32521 ;
  assign n32523 = ~n32516 & ~n32522 ;
  assign n32524 = ~n32273 & ~n32279 ;
  assign n32525 = ~n32274 & ~n32524 ;
  assign n32526 = n5211 & ~n13524 ;
  assign n32527 = ~n13522 & n32526 ;
  assign n32528 = \b[49]  & n5209 ;
  assign n32529 = \a[30]  & \b[48]  ;
  assign n32530 = n5200 & n32529 ;
  assign n32531 = ~n32528 & ~n32530 ;
  assign n32532 = \b[47]  & n5595 ;
  assign n32533 = n5592 & n32532 ;
  assign n32534 = ~\a[30]  & \b[48]  ;
  assign n32535 = n5203 & n32534 ;
  assign n32536 = ~n32533 & ~n32535 ;
  assign n32537 = n32531 & n32536 ;
  assign n32538 = ~n32527 & n32537 ;
  assign n32539 = ~\a[32]  & ~n32538 ;
  assign n32540 = \a[32]  & n32537 ;
  assign n32541 = ~n32527 & n32540 ;
  assign n32542 = ~n32539 & ~n32541 ;
  assign n32543 = ~n32525 & n32542 ;
  assign n32544 = ~n32274 & ~n32542 ;
  assign n32545 = ~n32524 & n32544 ;
  assign n32546 = ~n32543 & ~n32545 ;
  assign n32547 = ~n31939 & n32246 ;
  assign n32548 = n32251 & ~n32547 ;
  assign n32549 = ~n32109 & ~n32113 ;
  assign n32550 = ~n32110 & ~n32549 ;
  assign n32551 = n32043 & ~n32044 ;
  assign n32552 = ~n31962 & ~n32044 ;
  assign n32553 = ~n32551 & ~n32552 ;
  assign n32554 = ~n31987 & ~n32038 ;
  assign n32555 = n32029 & ~n32554 ;
  assign n32556 = ~n2079 & n20521 ;
  assign n32557 = ~n2077 & n32556 ;
  assign n32558 = \b[19]  & n20519 ;
  assign n32559 = \a[60]  & \b[18]  ;
  assign n32560 = n20510 & n32559 ;
  assign n32561 = ~n32558 & ~n32560 ;
  assign n32562 = \b[17]  & n21315 ;
  assign n32563 = n21312 & n32562 ;
  assign n32564 = ~\a[60]  & \b[18]  ;
  assign n32565 = n20513 & n32564 ;
  assign n32566 = ~n32563 & ~n32565 ;
  assign n32567 = n32561 & n32566 ;
  assign n32568 = ~n32557 & n32567 ;
  assign n32569 = ~n30811 & ~n32013 ;
  assign n32570 = n32009 & ~n32569 ;
  assign n32571 = \b[16]  & n21958 ;
  assign n32572 = \b[15]  & n21957 ;
  assign n32573 = ~n32571 & ~n32572 ;
  assign n32574 = ~n32570 & n32573 ;
  assign n32575 = n32009 & ~n32573 ;
  assign n32576 = ~n32569 & n32575 ;
  assign n32577 = ~\a[62]  & ~n32576 ;
  assign n32578 = ~n32574 & n32577 ;
  assign n32579 = ~n32568 & n32578 ;
  assign n32580 = \a[62]  & ~n32576 ;
  assign n32581 = ~n32574 & n32580 ;
  assign n32582 = n32567 & n32581 ;
  assign n32583 = ~n32557 & n32582 ;
  assign n32584 = ~n32579 & ~n32583 ;
  assign n32585 = ~\a[62]  & ~n32568 ;
  assign n32586 = ~n32574 & ~n32576 ;
  assign n32587 = \a[62]  & n32567 ;
  assign n32588 = ~n32557 & n32587 ;
  assign n32589 = ~n32586 & ~n32588 ;
  assign n32590 = ~n32585 & n32589 ;
  assign n32591 = n32584 & ~n32590 ;
  assign n32592 = ~n32555 & n32591 ;
  assign n32593 = n32555 & ~n32591 ;
  assign n32594 = ~n32592 & ~n32593 ;
  assign n32595 = n2768 & n18516 ;
  assign n32596 = ~n2765 & n32595 ;
  assign n32597 = ~n2518 & ~n2768 ;
  assign n32598 = n18516 & n32597 ;
  assign n32599 = ~n2764 & n32598 ;
  assign n32600 = \b[22]  & n18514 ;
  assign n32601 = \a[56]  & \b[21]  ;
  assign n32602 = n19181 & n32601 ;
  assign n32603 = ~\a[57]  & \b[21]  ;
  assign n32604 = n18508 & n32603 ;
  assign n32605 = ~n32602 & ~n32604 ;
  assign n32606 = ~n32600 & n32605 ;
  assign n32607 = \b[20]  & n19183 ;
  assign n32608 = n19180 & n32607 ;
  assign n32609 = \a[59]  & ~n32608 ;
  assign n32610 = n32606 & n32609 ;
  assign n32611 = ~n32599 & n32610 ;
  assign n32612 = ~n32596 & n32611 ;
  assign n32613 = n32606 & ~n32608 ;
  assign n32614 = ~n32599 & n32613 ;
  assign n32615 = ~n32596 & n32614 ;
  assign n32616 = ~\a[59]  & ~n32615 ;
  assign n32617 = ~n32612 & ~n32616 ;
  assign n32618 = n32594 & ~n32617 ;
  assign n32619 = ~n32594 & n32617 ;
  assign n32620 = ~n32618 & ~n32619 ;
  assign n32621 = ~n32553 & ~n32620 ;
  assign n32622 = n32553 & n32620 ;
  assign n32623 = ~n32621 & ~n32622 ;
  assign n32624 = ~n3564 & n16655 ;
  assign n32625 = ~n3282 & n16655 ;
  assign n32626 = ~n3560 & n32625 ;
  assign n32627 = ~n32624 & ~n32626 ;
  assign n32628 = ~n3567 & ~n32627 ;
  assign n32629 = \b[25]  & n16653 ;
  assign n32630 = \a[54]  & \b[24]  ;
  assign n32631 = n16644 & n32630 ;
  assign n32632 = ~\a[54]  & \b[24]  ;
  assign n32633 = n16647 & n32632 ;
  assign n32634 = ~n32631 & ~n32633 ;
  assign n32635 = ~n32629 & n32634 ;
  assign n32636 = \b[23]  & n17308 ;
  assign n32637 = n17305 & n32636 ;
  assign n32638 = \a[56]  & ~n32637 ;
  assign n32639 = n32635 & n32638 ;
  assign n32640 = ~n32628 & n32639 ;
  assign n32641 = n32635 & ~n32637 ;
  assign n32642 = ~\a[56]  & ~n32641 ;
  assign n32643 = ~\a[56]  & ~n3567 ;
  assign n32644 = ~n32627 & n32643 ;
  assign n32645 = ~n32642 & ~n32644 ;
  assign n32646 = ~n32640 & n32645 ;
  assign n32647 = ~n32623 & n32646 ;
  assign n32648 = n32623 & ~n32646 ;
  assign n32649 = ~n32647 & ~n32648 ;
  assign n32650 = n4456 & n14793 ;
  assign n32651 = ~n18723 & n32650 ;
  assign n32652 = ~n4456 & n14793 ;
  assign n32653 = ~n4143 & n32652 ;
  assign n32654 = ~n4452 & n32653 ;
  assign n32655 = \b[26]  & n15517 ;
  assign n32656 = n15514 & n32655 ;
  assign n32657 = ~\a[51]  & \b[27]  ;
  assign n32658 = n14785 & n32657 ;
  assign n32659 = ~n32656 & ~n32658 ;
  assign n32660 = \b[28]  & n14791 ;
  assign n32661 = \a[51]  & \b[27]  ;
  assign n32662 = n14782 & n32661 ;
  assign n32663 = \a[53]  & ~n32662 ;
  assign n32664 = ~n32660 & n32663 ;
  assign n32665 = n32659 & n32664 ;
  assign n32666 = ~n32654 & n32665 ;
  assign n32667 = ~n32651 & n32666 ;
  assign n32668 = ~n32660 & ~n32662 ;
  assign n32669 = n32659 & n32668 ;
  assign n32670 = ~n32654 & n32669 ;
  assign n32671 = ~n32651 & n32670 ;
  assign n32672 = ~\a[53]  & ~n32671 ;
  assign n32673 = ~n32667 & ~n32672 ;
  assign n32674 = ~n31960 & ~n32074 ;
  assign n32675 = ~n32073 & ~n32674 ;
  assign n32676 = n32673 & ~n32675 ;
  assign n32677 = ~n32649 & n32676 ;
  assign n32678 = n32673 & n32675 ;
  assign n32679 = n32649 & n32678 ;
  assign n32680 = ~n32677 & ~n32679 ;
  assign n32681 = ~n32673 & ~n32675 ;
  assign n32682 = n32649 & n32681 ;
  assign n32683 = ~n32673 & n32675 ;
  assign n32684 = ~n32649 & n32683 ;
  assign n32685 = ~n32682 & ~n32684 ;
  assign n32686 = n32680 & n32685 ;
  assign n32687 = n31941 & ~n32079 ;
  assign n32688 = ~n32080 & ~n32687 ;
  assign n32689 = n32686 & n32688 ;
  assign n32690 = ~n32686 & ~n32688 ;
  assign n32691 = ~n32689 & ~n32690 ;
  assign n32692 = ~n5459 & n13125 ;
  assign n32693 = ~n5104 & n13125 ;
  assign n32694 = ~n5455 & n32693 ;
  assign n32695 = ~n32692 & ~n32694 ;
  assign n32696 = ~n5462 & ~n32695 ;
  assign n32697 = \b[29]  & n13794 ;
  assign n32698 = n13792 & n32697 ;
  assign n32699 = ~\a[48]  & \b[30]  ;
  assign n32700 = n13117 & n32699 ;
  assign n32701 = ~n32698 & ~n32700 ;
  assign n32702 = \b[31]  & n13123 ;
  assign n32703 = \a[48]  & \b[30]  ;
  assign n32704 = n13786 & n32703 ;
  assign n32705 = \a[50]  & ~n32704 ;
  assign n32706 = ~n32702 & n32705 ;
  assign n32707 = n32701 & n32706 ;
  assign n32708 = ~n32696 & n32707 ;
  assign n32709 = ~n32702 & ~n32704 ;
  assign n32710 = n32701 & n32709 ;
  assign n32711 = ~\a[50]  & ~n32710 ;
  assign n32712 = ~\a[50]  & ~n5462 ;
  assign n32713 = ~n32695 & n32712 ;
  assign n32714 = ~n32711 & ~n32713 ;
  assign n32715 = ~n32708 & n32714 ;
  assign n32716 = ~n32691 & n32715 ;
  assign n32717 = n32691 & ~n32715 ;
  assign n32718 = ~n32716 & ~n32717 ;
  assign n32719 = ~n32550 & ~n32718 ;
  assign n32720 = n32550 & n32718 ;
  assign n32721 = ~n32719 & ~n32720 ;
  assign n32722 = n6565 & n11572 ;
  assign n32723 = ~n6562 & n32722 ;
  assign n32724 = n11572 & n22947 ;
  assign n32725 = ~n6561 & n32724 ;
  assign n32726 = \b[32]  & n12159 ;
  assign n32727 = n12156 & n32726 ;
  assign n32728 = ~\a[45]  & \b[33]  ;
  assign n32729 = n11564 & n32728 ;
  assign n32730 = ~n32727 & ~n32729 ;
  assign n32731 = \b[34]  & n11570 ;
  assign n32732 = \a[45]  & \b[33]  ;
  assign n32733 = n11561 & n32732 ;
  assign n32734 = \a[47]  & ~n32733 ;
  assign n32735 = ~n32731 & n32734 ;
  assign n32736 = n32730 & n32735 ;
  assign n32737 = ~n32725 & n32736 ;
  assign n32738 = ~n32723 & n32737 ;
  assign n32739 = ~n32731 & ~n32733 ;
  assign n32740 = n32730 & n32739 ;
  assign n32741 = ~n32725 & n32740 ;
  assign n32742 = ~n32723 & n32741 ;
  assign n32743 = ~\a[47]  & ~n32742 ;
  assign n32744 = ~n32738 & ~n32743 ;
  assign n32745 = ~n32721 & n32744 ;
  assign n32746 = n32721 & ~n32744 ;
  assign n32747 = ~n32745 & ~n32746 ;
  assign n32748 = ~n7761 & n10082 ;
  assign n32749 = ~n7759 & n32748 ;
  assign n32750 = \b[37]  & n10080 ;
  assign n32751 = \a[41]  & \b[36]  ;
  assign n32752 = n10679 & n32751 ;
  assign n32753 = ~\a[42]  & \b[36]  ;
  assign n32754 = n10074 & n32753 ;
  assign n32755 = ~n32752 & ~n32754 ;
  assign n32756 = ~n32750 & n32755 ;
  assign n32757 = \b[35]  & n10681 ;
  assign n32758 = n10678 & n32757 ;
  assign n32759 = \a[44]  & ~n32758 ;
  assign n32760 = n32756 & n32759 ;
  assign n32761 = ~n32749 & n32760 ;
  assign n32762 = n32756 & ~n32758 ;
  assign n32763 = ~n32749 & n32762 ;
  assign n32764 = ~\a[44]  & ~n32763 ;
  assign n32765 = ~n32761 & ~n32764 ;
  assign n32766 = n32137 & ~n32169 ;
  assign n32767 = n32142 & ~n32766 ;
  assign n32768 = n32765 & n32767 ;
  assign n32769 = ~n32747 & n32768 ;
  assign n32770 = n32765 & ~n32767 ;
  assign n32771 = n32747 & n32770 ;
  assign n32772 = ~n32769 & ~n32771 ;
  assign n32773 = ~n32765 & ~n32767 ;
  assign n32774 = ~n32747 & n32773 ;
  assign n32775 = ~n32765 & n32767 ;
  assign n32776 = n32747 & n32775 ;
  assign n32777 = ~n32774 & ~n32776 ;
  assign n32778 = n32772 & n32777 ;
  assign n32779 = n8759 & n9044 ;
  assign n32780 = ~n9041 & n32779 ;
  assign n32781 = n8759 & ~n9044 ;
  assign n32782 = ~n8597 & n32781 ;
  assign n32783 = ~n9040 & n32782 ;
  assign n32784 = \b[38]  & n9301 ;
  assign n32785 = n9298 & n32784 ;
  assign n32786 = ~\a[39]  & \b[39]  ;
  assign n32787 = n8751 & n32786 ;
  assign n32788 = ~n32785 & ~n32787 ;
  assign n32789 = \b[40]  & n8757 ;
  assign n32790 = \a[39]  & \b[39]  ;
  assign n32791 = n8748 & n32790 ;
  assign n32792 = \a[41]  & ~n32791 ;
  assign n32793 = ~n32789 & n32792 ;
  assign n32794 = n32788 & n32793 ;
  assign n32795 = ~n32783 & n32794 ;
  assign n32796 = ~n32780 & n32795 ;
  assign n32797 = ~n32789 & ~n32791 ;
  assign n32798 = n32788 & n32797 ;
  assign n32799 = ~n32783 & n32798 ;
  assign n32800 = ~n32780 & n32799 ;
  assign n32801 = ~\a[41]  & ~n32800 ;
  assign n32802 = ~n32796 & ~n32801 ;
  assign n32803 = n32174 & ~n32184 ;
  assign n32804 = n32179 & ~n32803 ;
  assign n32805 = ~n32802 & ~n32804 ;
  assign n32806 = ~n32778 & n32805 ;
  assign n32807 = ~n32802 & n32804 ;
  assign n32808 = n32778 & n32807 ;
  assign n32809 = ~n32806 & ~n32808 ;
  assign n32810 = n32802 & n32804 ;
  assign n32811 = ~n32778 & n32810 ;
  assign n32812 = n32802 & ~n32804 ;
  assign n32813 = n32778 & n32812 ;
  assign n32814 = ~n32811 & ~n32813 ;
  assign n32815 = n32809 & n32814 ;
  assign n32816 = n32208 & ~n32241 ;
  assign n32817 = n32213 & ~n32816 ;
  assign n32818 = n7534 & ~n10409 ;
  assign n32819 = ~n10407 & n32818 ;
  assign n32820 = \b[41]  & n7973 ;
  assign n32821 = n7970 & n32820 ;
  assign n32822 = ~\a[36]  & \b[42]  ;
  assign n32823 = n7526 & n32822 ;
  assign n32824 = ~n32821 & ~n32823 ;
  assign n32825 = \b[43]  & n7532 ;
  assign n32826 = \a[36]  & \b[42]  ;
  assign n32827 = n17801 & n32826 ;
  assign n32828 = \a[38]  & ~n32827 ;
  assign n32829 = ~n32825 & n32828 ;
  assign n32830 = n32824 & n32829 ;
  assign n32831 = ~n32819 & n32830 ;
  assign n32832 = ~n32825 & ~n32827 ;
  assign n32833 = n32824 & n32832 ;
  assign n32834 = ~n32819 & n32833 ;
  assign n32835 = ~\a[38]  & ~n32834 ;
  assign n32836 = ~n32831 & ~n32835 ;
  assign n32837 = n32817 & ~n32836 ;
  assign n32838 = ~n32815 & n32837 ;
  assign n32839 = ~n32817 & ~n32836 ;
  assign n32840 = n32815 & n32839 ;
  assign n32841 = ~n32838 & ~n32840 ;
  assign n32842 = ~n32817 & n32836 ;
  assign n32843 = ~n32815 & n32842 ;
  assign n32844 = n32817 & n32836 ;
  assign n32845 = n32815 & n32844 ;
  assign n32846 = ~n32843 & ~n32845 ;
  assign n32847 = n32841 & n32846 ;
  assign n32848 = ~n32548 & ~n32847 ;
  assign n32849 = n32548 & n32847 ;
  assign n32850 = ~n32848 & ~n32849 ;
  assign n32851 = n6309 & n11906 ;
  assign n32852 = ~n11903 & n32851 ;
  assign n32853 = n6309 & ~n11906 ;
  assign n32854 = ~n11392 & n32853 ;
  assign n32855 = ~n11902 & n32854 ;
  assign n32856 = \b[44]  & n6778 ;
  assign n32857 = n6775 & n32856 ;
  assign n32858 = ~\a[33]  & \b[45]  ;
  assign n32859 = n6301 & n32858 ;
  assign n32860 = ~n32857 & ~n32859 ;
  assign n32861 = \b[46]  & n6307 ;
  assign n32862 = \a[33]  & \b[45]  ;
  assign n32863 = n6298 & n32862 ;
  assign n32864 = \a[35]  & ~n32863 ;
  assign n32865 = ~n32861 & n32864 ;
  assign n32866 = n32860 & n32865 ;
  assign n32867 = ~n32855 & n32866 ;
  assign n32868 = ~n32852 & n32867 ;
  assign n32869 = ~n32861 & ~n32863 ;
  assign n32870 = n32860 & n32869 ;
  assign n32871 = ~n32855 & n32870 ;
  assign n32872 = ~n32852 & n32871 ;
  assign n32873 = ~\a[35]  & ~n32872 ;
  assign n32874 = ~n32868 & ~n32873 ;
  assign n32875 = ~n32850 & n32874 ;
  assign n32876 = n32850 & ~n32874 ;
  assign n32877 = ~n32875 & ~n32876 ;
  assign n32878 = n32546 & n32877 ;
  assign n32879 = ~n32546 & ~n32877 ;
  assign n32880 = ~n32878 & ~n32879 ;
  assign n32881 = n4249 & n15201 ;
  assign n32882 = ~n15198 & n32881 ;
  assign n32883 = n4249 & ~n15201 ;
  assign n32884 = ~n14093 & n32883 ;
  assign n32885 = ~n15197 & n32884 ;
  assign n32886 = \b[50]  & n4647 ;
  assign n32887 = n4644 & n32886 ;
  assign n32888 = ~\a[27]  & \b[51]  ;
  assign n32889 = n4241 & n32888 ;
  assign n32890 = ~n32887 & ~n32889 ;
  assign n32891 = \b[52]  & n4247 ;
  assign n32892 = \a[27]  & \b[51]  ;
  assign n32893 = n4238 & n32892 ;
  assign n32894 = \a[29]  & ~n32893 ;
  assign n32895 = ~n32891 & n32894 ;
  assign n32896 = n32890 & n32895 ;
  assign n32897 = ~n32885 & n32896 ;
  assign n32898 = ~n32882 & n32897 ;
  assign n32899 = ~n32891 & ~n32893 ;
  assign n32900 = n32890 & n32899 ;
  assign n32901 = ~n32885 & n32900 ;
  assign n32902 = ~n32882 & n32901 ;
  assign n32903 = ~\a[29]  & ~n32902 ;
  assign n32904 = ~n32898 & ~n32903 ;
  assign n32905 = n32281 & ~n32307 ;
  assign n32906 = ~n32313 & ~n32905 ;
  assign n32907 = n32280 & ~n32307 ;
  assign n32908 = n32279 & n32305 ;
  assign n32909 = n32275 & n32908 ;
  assign n32910 = ~n32279 & n32305 ;
  assign n32911 = ~n32275 & n32910 ;
  assign n32912 = ~n32909 & ~n32911 ;
  assign n32913 = ~n32907 & n32912 ;
  assign n32914 = n32906 & n32913 ;
  assign n32915 = ~n32904 & n32914 ;
  assign n32916 = n32904 & ~n32914 ;
  assign n32917 = ~n32915 & ~n32916 ;
  assign n32918 = n32880 & n32917 ;
  assign n32919 = ~n32880 & n32915 ;
  assign n32920 = ~n32880 & n32916 ;
  assign n32921 = ~n32919 & ~n32920 ;
  assign n32922 = ~n32918 & n32921 ;
  assign n32923 = n32523 & n32922 ;
  assign n32924 = ~n32523 & ~n32922 ;
  assign n32925 = ~n32923 & ~n32924 ;
  assign n32926 = ~n32495 & n32925 ;
  assign n32927 = ~n32494 & n32926 ;
  assign n32928 = n32495 & ~n32925 ;
  assign n32929 = n32494 & ~n32925 ;
  assign n32930 = ~n32928 & ~n32929 ;
  assign n32931 = ~n32927 & n32930 ;
  assign n32932 = n32462 & n32931 ;
  assign n32933 = ~n32462 & ~n32931 ;
  assign n32934 = ~n32932 & ~n32933 ;
  assign n32935 = ~n32436 & n32934 ;
  assign n32936 = n32436 & ~n32934 ;
  assign n32937 = ~n32935 & ~n32936 ;
  assign n32938 = ~n32408 & n32937 ;
  assign n32939 = n32408 & ~n32937 ;
  assign n32940 = ~n32938 & ~n32939 ;
  assign n32941 = ~n32397 & n32940 ;
  assign n32942 = ~n32399 & n32941 ;
  assign n32943 = ~n32402 & n32942 ;
  assign n32944 = ~n32397 & ~n32399 ;
  assign n32945 = ~n32402 & n32944 ;
  assign n32946 = ~n32940 & ~n32945 ;
  assign n32947 = ~n32943 & ~n32946 ;
  assign n32948 = ~n32397 & ~n32939 ;
  assign n32949 = ~n32399 & n32948 ;
  assign n32950 = ~n32402 & n32949 ;
  assign n32951 = n1965 & n21696 ;
  assign n32952 = ~n21693 & n32951 ;
  assign n32953 = n1965 & ~n21696 ;
  assign n32954 = ~n20966 & n32953 ;
  assign n32955 = ~n21692 & n32954 ;
  assign n32956 = \b[62]  & n1963 ;
  assign n32957 = \a[18]  & \b[61]  ;
  assign n32958 = n28047 & n32957 ;
  assign n32959 = ~n32956 & ~n32958 ;
  assign n32960 = \b[60]  & n2218 ;
  assign n32961 = n2216 & n32960 ;
  assign n32962 = ~\a[18]  & \b[61]  ;
  assign n32963 = n1957 & n32962 ;
  assign n32964 = ~n32961 & ~n32963 ;
  assign n32965 = n32959 & n32964 ;
  assign n32966 = ~n32955 & n32965 ;
  assign n32967 = ~n32952 & n32966 ;
  assign n32968 = ~\a[20]  & ~n32967 ;
  assign n32969 = \a[20]  & ~n32958 ;
  assign n32970 = ~n32956 & n32969 ;
  assign n32971 = n32964 & n32970 ;
  assign n32972 = ~n32955 & n32971 ;
  assign n32973 = ~n32952 & n32972 ;
  assign n32974 = ~n32968 & ~n32973 ;
  assign n32975 = ~n32495 & n32974 ;
  assign n32976 = ~n32927 & n32975 ;
  assign n32977 = ~n32495 & ~n32925 ;
  assign n32978 = n32494 & ~n32495 ;
  assign n32979 = ~n32977 & ~n32978 ;
  assign n32980 = \a[20]  & ~n32967 ;
  assign n32981 = ~\a[20]  & n32967 ;
  assign n32982 = ~n32980 & ~n32981 ;
  assign n32983 = n32979 & n32982 ;
  assign n32984 = ~n32976 & ~n32983 ;
  assign n32985 = n3402 & n17647 ;
  assign n32986 = ~n17644 & n32985 ;
  assign n32987 = n3402 & ~n17647 ;
  assign n32988 = ~n16441 & n32987 ;
  assign n32989 = ~n17643 & n32988 ;
  assign n32990 = \b[56]  & n3400 ;
  assign n32991 = \a[24]  & \b[55]  ;
  assign n32992 = n27626 & n32991 ;
  assign n32993 = ~n32990 & ~n32992 ;
  assign n32994 = \b[54]  & n3733 ;
  assign n32995 = n3730 & n32994 ;
  assign n32996 = ~\a[24]  & \b[55]  ;
  assign n32997 = n3394 & n32996 ;
  assign n32998 = ~n32995 & ~n32997 ;
  assign n32999 = n32993 & n32998 ;
  assign n33000 = ~n32989 & n32999 ;
  assign n33001 = ~n32986 & n33000 ;
  assign n33002 = ~\a[26]  & ~n33001 ;
  assign n33003 = \a[26]  & ~n32992 ;
  assign n33004 = ~n32990 & n33003 ;
  assign n33005 = n32998 & n33004 ;
  assign n33006 = ~n32989 & n33005 ;
  assign n33007 = ~n32986 & n33006 ;
  assign n33008 = ~n33002 & ~n33007 ;
  assign n33009 = ~n32915 & n33008 ;
  assign n33010 = ~n32918 & n33009 ;
  assign n33011 = ~n32915 & n32916 ;
  assign n33012 = ~n32880 & ~n32915 ;
  assign n33013 = ~n33011 & ~n33012 ;
  assign n33014 = \a[26]  & ~n33001 ;
  assign n33015 = ~\a[26]  & n33001 ;
  assign n33016 = ~n33014 & ~n33015 ;
  assign n33017 = n33013 & n33016 ;
  assign n33018 = ~n33010 & ~n33017 ;
  assign n33019 = ~n32849 & n32874 ;
  assign n33020 = ~n32848 & ~n33019 ;
  assign n33021 = n5211 & n14052 ;
  assign n33022 = ~n14049 & n33021 ;
  assign n33023 = n5211 & ~n14052 ;
  assign n33024 = ~n13519 & n33023 ;
  assign n33025 = ~n14048 & n33024 ;
  assign n33026 = \b[50]  & n5209 ;
  assign n33027 = \a[30]  & \b[49]  ;
  assign n33028 = n5200 & n33027 ;
  assign n33029 = ~n33026 & ~n33028 ;
  assign n33030 = \b[48]  & n5595 ;
  assign n33031 = n5592 & n33030 ;
  assign n33032 = ~\a[30]  & \b[49]  ;
  assign n33033 = n5203 & n33032 ;
  assign n33034 = ~n33031 & ~n33033 ;
  assign n33035 = n33029 & n33034 ;
  assign n33036 = ~n33025 & n33035 ;
  assign n33037 = ~n33022 & n33036 ;
  assign n33038 = ~\a[32]  & ~n33037 ;
  assign n33039 = \a[32]  & ~n33028 ;
  assign n33040 = ~n33026 & n33039 ;
  assign n33041 = n33034 & n33040 ;
  assign n33042 = ~n33025 & n33041 ;
  assign n33043 = ~n33022 & n33042 ;
  assign n33044 = ~n33038 & ~n33043 ;
  assign n33045 = ~n33020 & n33044 ;
  assign n33046 = \a[32]  & ~n33037 ;
  assign n33047 = ~\a[32]  & n33037 ;
  assign n33048 = ~n33046 & ~n33047 ;
  assign n33049 = ~n32848 & n33048 ;
  assign n33050 = ~n33019 & n33049 ;
  assign n33051 = ~n33045 & ~n33050 ;
  assign n33052 = n8759 & ~n9482 ;
  assign n33053 = ~n9480 & n33052 ;
  assign n33054 = \b[39]  & n9301 ;
  assign n33055 = n9298 & n33054 ;
  assign n33056 = ~\a[39]  & \b[40]  ;
  assign n33057 = n8751 & n33056 ;
  assign n33058 = ~n33055 & ~n33057 ;
  assign n33059 = \b[41]  & n8757 ;
  assign n33060 = \a[39]  & \b[40]  ;
  assign n33061 = n8748 & n33060 ;
  assign n33062 = \a[41]  & ~n33061 ;
  assign n33063 = ~n33059 & n33062 ;
  assign n33064 = n33058 & n33063 ;
  assign n33065 = ~n33053 & n33064 ;
  assign n33066 = ~n33059 & ~n33061 ;
  assign n33067 = n33058 & n33066 ;
  assign n33068 = ~n33053 & n33067 ;
  assign n33069 = ~\a[41]  & ~n33068 ;
  assign n33070 = ~n33065 & ~n33069 ;
  assign n33071 = ~n32747 & ~n32767 ;
  assign n33072 = n32747 & n32767 ;
  assign n33073 = n32765 & ~n33072 ;
  assign n33074 = ~n33071 & ~n33073 ;
  assign n33075 = n3604 & n16655 ;
  assign n33076 = ~n19292 & n33075 ;
  assign n33077 = n12021 & n16655 ;
  assign n33078 = ~n3600 & n33077 ;
  assign n33079 = \b[26]  & n16653 ;
  assign n33080 = \a[54]  & \b[25]  ;
  assign n33081 = n16644 & n33080 ;
  assign n33082 = ~\a[54]  & \b[25]  ;
  assign n33083 = n16647 & n33082 ;
  assign n33084 = ~n33081 & ~n33083 ;
  assign n33085 = ~n33079 & n33084 ;
  assign n33086 = \b[24]  & n17308 ;
  assign n33087 = n17305 & n33086 ;
  assign n33088 = \a[56]  & ~n33087 ;
  assign n33089 = n33085 & n33088 ;
  assign n33090 = ~n33078 & n33089 ;
  assign n33091 = ~n33076 & n33090 ;
  assign n33092 = n33085 & ~n33087 ;
  assign n33093 = ~n33078 & n33092 ;
  assign n33094 = ~n33076 & n33093 ;
  assign n33095 = ~\a[56]  & ~n33094 ;
  assign n33096 = ~n33091 & ~n33095 ;
  assign n33097 = ~n32574 & ~n32583 ;
  assign n33098 = ~n32579 & n33097 ;
  assign n33099 = n2293 & n20521 ;
  assign n33100 = ~n19247 & n33099 ;
  assign n33101 = ~n2293 & n20521 ;
  assign n33102 = ~n2074 & n33101 ;
  assign n33103 = ~n2289 & n33102 ;
  assign n33104 = \b[20]  & n20519 ;
  assign n33105 = \a[60]  & \b[19]  ;
  assign n33106 = n20510 & n33105 ;
  assign n33107 = ~n33104 & ~n33106 ;
  assign n33108 = \b[18]  & n21315 ;
  assign n33109 = n21312 & n33108 ;
  assign n33110 = ~\a[60]  & \b[19]  ;
  assign n33111 = n20513 & n33110 ;
  assign n33112 = ~n33109 & ~n33111 ;
  assign n33113 = n33107 & n33112 ;
  assign n33114 = ~n33103 & n33113 ;
  assign n33115 = ~n33100 & n33114 ;
  assign n33116 = \b[17]  & n21958 ;
  assign n33117 = \b[16]  & n21957 ;
  assign n33118 = ~n33116 & ~n33117 ;
  assign n33119 = n32573 & ~n33118 ;
  assign n33120 = ~n32573 & n33118 ;
  assign n33121 = ~n33119 & ~n33120 ;
  assign n33122 = ~\a[62]  & n33121 ;
  assign n33123 = ~n33115 & n33122 ;
  assign n33124 = \a[62]  & n33121 ;
  assign n33125 = n33113 & n33124 ;
  assign n33126 = ~n33103 & n33125 ;
  assign n33127 = ~n33100 & n33126 ;
  assign n33128 = ~n33123 & ~n33127 ;
  assign n33129 = ~\a[62]  & ~n33115 ;
  assign n33130 = \a[62]  & n33113 ;
  assign n33131 = ~n33103 & n33130 ;
  assign n33132 = ~n33100 & n33131 ;
  assign n33133 = ~n33121 & ~n33132 ;
  assign n33134 = ~n33129 & n33133 ;
  assign n33135 = n33128 & ~n33134 ;
  assign n33136 = n33098 & ~n33135 ;
  assign n33137 = ~n33098 & n33135 ;
  assign n33138 = ~n33136 & ~n33137 ;
  assign n33139 = ~n3022 & n18516 ;
  assign n33140 = ~n3020 & n33139 ;
  assign n33141 = \b[23]  & n18514 ;
  assign n33142 = \a[56]  & \b[22]  ;
  assign n33143 = n19181 & n33142 ;
  assign n33144 = ~\a[57]  & \b[22]  ;
  assign n33145 = n18508 & n33144 ;
  assign n33146 = ~n33143 & ~n33145 ;
  assign n33147 = ~n33141 & n33146 ;
  assign n33148 = \b[21]  & n19183 ;
  assign n33149 = n19180 & n33148 ;
  assign n33150 = \a[59]  & ~n33149 ;
  assign n33151 = n33147 & n33150 ;
  assign n33152 = ~n33140 & n33151 ;
  assign n33153 = n33147 & ~n33149 ;
  assign n33154 = ~n33140 & n33153 ;
  assign n33155 = ~\a[59]  & ~n33154 ;
  assign n33156 = ~n33152 & ~n33155 ;
  assign n33157 = n33138 & ~n33156 ;
  assign n33158 = ~n33138 & n33156 ;
  assign n33159 = ~n32592 & n32617 ;
  assign n33160 = ~n32593 & ~n33159 ;
  assign n33161 = ~n33158 & n33160 ;
  assign n33162 = ~n33157 & n33161 ;
  assign n33163 = ~n33156 & ~n33160 ;
  assign n33164 = n33138 & n33163 ;
  assign n33165 = ~n33138 & ~n33160 ;
  assign n33166 = n33156 & n33165 ;
  assign n33167 = ~n33164 & ~n33166 ;
  assign n33168 = ~n33162 & n33167 ;
  assign n33169 = ~n33096 & ~n33168 ;
  assign n33170 = n33096 & n33168 ;
  assign n33171 = ~n33169 & ~n33170 ;
  assign n33172 = ~n32622 & n32646 ;
  assign n33173 = ~n32621 & ~n33172 ;
  assign n33174 = ~n33171 & n33173 ;
  assign n33175 = n33171 & ~n33173 ;
  assign n33176 = ~n33174 & ~n33175 ;
  assign n33177 = ~n4502 & n14793 ;
  assign n33178 = ~n4500 & n33177 ;
  assign n33179 = \b[27]  & n15517 ;
  assign n33180 = n15514 & n33179 ;
  assign n33181 = ~\a[51]  & \b[28]  ;
  assign n33182 = n14785 & n33181 ;
  assign n33183 = ~n33180 & ~n33182 ;
  assign n33184 = \b[29]  & n14791 ;
  assign n33185 = \a[51]  & \b[28]  ;
  assign n33186 = n14782 & n33185 ;
  assign n33187 = \a[53]  & ~n33186 ;
  assign n33188 = ~n33184 & n33187 ;
  assign n33189 = n33183 & n33188 ;
  assign n33190 = ~n33178 & n33189 ;
  assign n33191 = ~n33184 & ~n33186 ;
  assign n33192 = n33183 & n33191 ;
  assign n33193 = ~n33178 & n33192 ;
  assign n33194 = ~\a[53]  & ~n33193 ;
  assign n33195 = ~n33190 & ~n33194 ;
  assign n33196 = n33176 & ~n33195 ;
  assign n33197 = ~n33176 & n33195 ;
  assign n33198 = ~n33196 & ~n33197 ;
  assign n33199 = ~n5810 & ~n12606 ;
  assign n33200 = ~n13122 & n33199 ;
  assign n33201 = n5807 & n33200 ;
  assign n33202 = n5810 & ~n12606 ;
  assign n33203 = ~n13122 & n33202 ;
  assign n33204 = ~n5807 & n33203 ;
  assign n33205 = ~n33201 & ~n33204 ;
  assign n33206 = \b[30]  & n13794 ;
  assign n33207 = n13792 & n33206 ;
  assign n33208 = ~\a[48]  & \b[31]  ;
  assign n33209 = n13117 & n33208 ;
  assign n33210 = ~n33207 & ~n33209 ;
  assign n33211 = \b[32]  & n13123 ;
  assign n33212 = \a[48]  & \b[31]  ;
  assign n33213 = n13786 & n33212 ;
  assign n33214 = \a[50]  & ~n33213 ;
  assign n33215 = ~n33211 & n33214 ;
  assign n33216 = n33210 & n33215 ;
  assign n33217 = n33205 & n33216 ;
  assign n33218 = ~n33211 & ~n33213 ;
  assign n33219 = n33210 & n33218 ;
  assign n33220 = n33205 & n33219 ;
  assign n33221 = ~\a[50]  & ~n33220 ;
  assign n33222 = ~n33217 & ~n33221 ;
  assign n33223 = n32649 & n32675 ;
  assign n33224 = n32685 & ~n33223 ;
  assign n33225 = n33222 & ~n33224 ;
  assign n33226 = ~n33198 & n33225 ;
  assign n33227 = n33222 & n33224 ;
  assign n33228 = n33198 & n33227 ;
  assign n33229 = ~n33226 & ~n33228 ;
  assign n33230 = ~n33222 & n33224 ;
  assign n33231 = ~n33198 & n33230 ;
  assign n33232 = ~n33222 & ~n33224 ;
  assign n33233 = n33198 & n33232 ;
  assign n33234 = ~n33231 & ~n33233 ;
  assign n33235 = n33229 & n33234 ;
  assign n33236 = ~n32689 & n32715 ;
  assign n33237 = ~n32690 & ~n33236 ;
  assign n33238 = ~n6607 & n11572 ;
  assign n33239 = ~n6564 & n11572 ;
  assign n33240 = ~n6603 & n33239 ;
  assign n33241 = ~n33238 & ~n33240 ;
  assign n33242 = ~n6610 & ~n33241 ;
  assign n33243 = \b[33]  & n12159 ;
  assign n33244 = n12156 & n33243 ;
  assign n33245 = ~\a[45]  & \b[34]  ;
  assign n33246 = n11564 & n33245 ;
  assign n33247 = ~n33244 & ~n33246 ;
  assign n33248 = \b[35]  & n11570 ;
  assign n33249 = \a[45]  & \b[34]  ;
  assign n33250 = n11561 & n33249 ;
  assign n33251 = \a[47]  & ~n33250 ;
  assign n33252 = ~n33248 & n33251 ;
  assign n33253 = n33247 & n33252 ;
  assign n33254 = ~n33242 & n33253 ;
  assign n33255 = ~n33248 & ~n33250 ;
  assign n33256 = n33247 & n33255 ;
  assign n33257 = ~\a[47]  & ~n33256 ;
  assign n33258 = ~\a[47]  & ~n6610 ;
  assign n33259 = ~n33241 & n33258 ;
  assign n33260 = ~n33257 & ~n33259 ;
  assign n33261 = ~n33254 & n33260 ;
  assign n33262 = ~n33237 & ~n33261 ;
  assign n33263 = ~n33235 & n33262 ;
  assign n33264 = n33237 & ~n33261 ;
  assign n33265 = n33235 & n33264 ;
  assign n33266 = ~n33263 & ~n33265 ;
  assign n33267 = n33237 & n33261 ;
  assign n33268 = ~n33235 & n33267 ;
  assign n33269 = ~n33237 & n33261 ;
  assign n33270 = n33235 & n33269 ;
  assign n33271 = ~n33268 & ~n33270 ;
  assign n33272 = n33266 & n33271 ;
  assign n33273 = n8175 & n10082 ;
  assign n33274 = ~n8172 & n33273 ;
  assign n33275 = ~n8175 & n10082 ;
  assign n33276 = ~n7756 & n33275 ;
  assign n33277 = ~n8171 & n33276 ;
  assign n33278 = \b[36]  & n10681 ;
  assign n33279 = n10678 & n33278 ;
  assign n33280 = \b[38]  & n10080 ;
  assign n33281 = \a[41]  & \b[37]  ;
  assign n33282 = n10679 & n33281 ;
  assign n33283 = ~\a[42]  & \b[37]  ;
  assign n33284 = n10074 & n33283 ;
  assign n33285 = ~n33282 & ~n33284 ;
  assign n33286 = ~n33280 & n33285 ;
  assign n33287 = ~n33279 & n33286 ;
  assign n33288 = ~n33277 & n33287 ;
  assign n33289 = ~n33274 & n33288 ;
  assign n33290 = ~\a[44]  & ~n33289 ;
  assign n33291 = \a[44]  & n33287 ;
  assign n33292 = ~n33277 & n33291 ;
  assign n33293 = ~n33274 & n33292 ;
  assign n33294 = ~n33290 & ~n33293 ;
  assign n33295 = ~n32720 & n32744 ;
  assign n33296 = n32719 & ~n32720 ;
  assign n33297 = ~n33295 & ~n33296 ;
  assign n33298 = ~n33294 & n33297 ;
  assign n33299 = ~n33272 & n33298 ;
  assign n33300 = ~n33294 & ~n33297 ;
  assign n33301 = n33272 & n33300 ;
  assign n33302 = ~n33299 & ~n33301 ;
  assign n33303 = n33294 & ~n33297 ;
  assign n33304 = ~n33272 & n33303 ;
  assign n33305 = n33294 & n33297 ;
  assign n33306 = n33272 & n33305 ;
  assign n33307 = ~n33304 & ~n33306 ;
  assign n33308 = n33302 & n33307 ;
  assign n33309 = n33074 & n33308 ;
  assign n33310 = ~n33074 & ~n33308 ;
  assign n33311 = ~n33309 & ~n33310 ;
  assign n33312 = n33070 & n33311 ;
  assign n33313 = ~n33070 & ~n33311 ;
  assign n33314 = ~n33312 & ~n33313 ;
  assign n33315 = n7534 & ~n28007 ;
  assign n33316 = ~n28005 & n33315 ;
  assign n33317 = \b[42]  & n7973 ;
  assign n33318 = n7970 & n33317 ;
  assign n33319 = ~\a[36]  & \b[43]  ;
  assign n33320 = n7526 & n33319 ;
  assign n33321 = ~n33318 & ~n33320 ;
  assign n33322 = \b[44]  & n7532 ;
  assign n33323 = \a[36]  & \b[43]  ;
  assign n33324 = n17801 & n33323 ;
  assign n33325 = \a[38]  & ~n33324 ;
  assign n33326 = ~n33322 & n33325 ;
  assign n33327 = n33321 & n33326 ;
  assign n33328 = ~n33316 & n33327 ;
  assign n33329 = ~n33322 & ~n33324 ;
  assign n33330 = n33321 & n33329 ;
  assign n33331 = ~n33316 & n33330 ;
  assign n33332 = ~\a[38]  & ~n33331 ;
  assign n33333 = ~n33328 & ~n33332 ;
  assign n33334 = ~n32778 & n32804 ;
  assign n33335 = n32809 & ~n33334 ;
  assign n33336 = ~n33333 & n33335 ;
  assign n33337 = ~n33314 & n33336 ;
  assign n33338 = ~n33333 & ~n33335 ;
  assign n33339 = n33314 & n33338 ;
  assign n33340 = ~n33337 & ~n33339 ;
  assign n33341 = n33333 & ~n33335 ;
  assign n33342 = ~n33314 & n33341 ;
  assign n33343 = n33333 & n33335 ;
  assign n33344 = n33314 & n33343 ;
  assign n33345 = ~n33342 & ~n33344 ;
  assign n33346 = n33340 & n33345 ;
  assign n33347 = ~n32815 & ~n32817 ;
  assign n33348 = n32815 & n32817 ;
  assign n33349 = n32836 & ~n33348 ;
  assign n33350 = ~n33347 & ~n33349 ;
  assign n33351 = n6309 & ~n12438 ;
  assign n33352 = ~n12436 & n33351 ;
  assign n33353 = \b[45]  & n6778 ;
  assign n33354 = n6775 & n33353 ;
  assign n33355 = ~\a[33]  & \b[46]  ;
  assign n33356 = n6301 & n33355 ;
  assign n33357 = ~n33354 & ~n33356 ;
  assign n33358 = \b[47]  & n6307 ;
  assign n33359 = \a[33]  & \b[46]  ;
  assign n33360 = n6298 & n33359 ;
  assign n33361 = \a[35]  & ~n33360 ;
  assign n33362 = ~n33358 & n33361 ;
  assign n33363 = n33357 & n33362 ;
  assign n33364 = ~n33352 & n33363 ;
  assign n33365 = ~n33358 & ~n33360 ;
  assign n33366 = n33357 & n33365 ;
  assign n33367 = ~n33352 & n33366 ;
  assign n33368 = ~\a[35]  & ~n33367 ;
  assign n33369 = ~n33364 & ~n33368 ;
  assign n33370 = ~n33350 & ~n33369 ;
  assign n33371 = n33346 & n33370 ;
  assign n33372 = n33350 & ~n33369 ;
  assign n33373 = ~n33346 & n33372 ;
  assign n33374 = ~n33371 & ~n33373 ;
  assign n33375 = ~n33350 & n33369 ;
  assign n33376 = ~n33346 & n33375 ;
  assign n33377 = n33350 & n33369 ;
  assign n33378 = n33346 & n33377 ;
  assign n33379 = ~n33376 & ~n33378 ;
  assign n33380 = n33374 & n33379 ;
  assign n33381 = n33051 & n33380 ;
  assign n33382 = ~n33051 & ~n33380 ;
  assign n33383 = ~n33381 & ~n33382 ;
  assign n33384 = ~n32545 & ~n32877 ;
  assign n33385 = n32274 & n32542 ;
  assign n33386 = n32524 & n32542 ;
  assign n33387 = ~n33385 & ~n33386 ;
  assign n33388 = n4249 & ~n15246 ;
  assign n33389 = ~n15244 & n33388 ;
  assign n33390 = \b[53]  & n4247 ;
  assign n33391 = \a[27]  & \b[52]  ;
  assign n33392 = n4238 & n33391 ;
  assign n33393 = ~n33390 & ~n33392 ;
  assign n33394 = \b[51]  & n4647 ;
  assign n33395 = n4644 & n33394 ;
  assign n33396 = ~\a[27]  & \b[52]  ;
  assign n33397 = n4241 & n33396 ;
  assign n33398 = ~n33395 & ~n33397 ;
  assign n33399 = n33393 & n33398 ;
  assign n33400 = ~n33389 & n33399 ;
  assign n33401 = ~\a[29]  & ~n33400 ;
  assign n33402 = n33387 & n33401 ;
  assign n33403 = ~n33384 & n33402 ;
  assign n33404 = \a[29]  & n33400 ;
  assign n33405 = n33387 & n33404 ;
  assign n33406 = ~n33384 & n33405 ;
  assign n33407 = ~n33403 & ~n33406 ;
  assign n33408 = \a[29]  & n33399 ;
  assign n33409 = ~n33389 & n33408 ;
  assign n33410 = ~n33387 & ~n33409 ;
  assign n33411 = ~n32545 & ~n33409 ;
  assign n33412 = ~n32877 & n33411 ;
  assign n33413 = ~n33410 & ~n33412 ;
  assign n33414 = ~n33401 & ~n33413 ;
  assign n33415 = n33407 & ~n33414 ;
  assign n33416 = n33383 & n33415 ;
  assign n33417 = ~n33383 & ~n33415 ;
  assign n33418 = ~n33416 & ~n33417 ;
  assign n33419 = n33018 & n33418 ;
  assign n33420 = ~n33018 & ~n33418 ;
  assign n33421 = ~n33419 & ~n33420 ;
  assign n33422 = ~n32522 & ~n32922 ;
  assign n33423 = n32516 & ~n32522 ;
  assign n33424 = ~n33422 & ~n33423 ;
  assign n33425 = n2622 & ~n19550 ;
  assign n33426 = ~n19548 & n33425 ;
  assign n33427 = \b[57]  & n2912 ;
  assign n33428 = n2909 & n33427 ;
  assign n33429 = \b[59]  & n2620 ;
  assign n33430 = \a[20]  & \b[58]  ;
  assign n33431 = n2910 & n33430 ;
  assign n33432 = ~\a[21]  & \b[58]  ;
  assign n33433 = n2614 & n33432 ;
  assign n33434 = ~n33431 & ~n33433 ;
  assign n33435 = ~n33429 & n33434 ;
  assign n33436 = ~n33428 & n33435 ;
  assign n33437 = ~n33426 & n33436 ;
  assign n33438 = \a[23]  & ~n33437 ;
  assign n33439 = ~\a[23]  & n33437 ;
  assign n33440 = ~n33438 & ~n33439 ;
  assign n33441 = n33424 & n33440 ;
  assign n33442 = ~\a[23]  & ~n33437 ;
  assign n33443 = \a[23]  & n33436 ;
  assign n33444 = ~n33426 & n33443 ;
  assign n33445 = ~n32522 & ~n33444 ;
  assign n33446 = ~n32922 & n33445 ;
  assign n33447 = n32516 & n33445 ;
  assign n33448 = ~n33446 & ~n33447 ;
  assign n33449 = ~n33442 & ~n33448 ;
  assign n33450 = ~n33441 & ~n33449 ;
  assign n33451 = n33421 & n33450 ;
  assign n33452 = ~n33421 & ~n33450 ;
  assign n33453 = ~n33451 & ~n33452 ;
  assign n33454 = ~n32984 & ~n33453 ;
  assign n33455 = n32984 & n33453 ;
  assign n33456 = ~n33454 & ~n33455 ;
  assign n33457 = ~n32461 & ~n32931 ;
  assign n33458 = n32456 & ~n32461 ;
  assign n33459 = ~n33457 & ~n33458 ;
  assign n33460 = \b[63]  & n1467 ;
  assign n33461 = ~n21694 & n33460 ;
  assign n33462 = ~n23171 & n33461 ;
  assign n33463 = \a[14]  & \a[16]  ;
  assign n33464 = \a[15]  & ~\a[17]  ;
  assign n33465 = n33463 & n33464 ;
  assign n33466 = ~\a[14]  & ~\a[16]  ;
  assign n33467 = ~\a[15]  & \a[17]  ;
  assign n33468 = n33466 & n33467 ;
  assign n33469 = ~n33465 & ~n33468 ;
  assign n33470 = \b[63]  & ~n33469 ;
  assign n33471 = \a[17]  & ~n33470 ;
  assign n33472 = ~n33462 & n33471 ;
  assign n33473 = ~n33462 & ~n33470 ;
  assign n33474 = ~\a[17]  & ~n33473 ;
  assign n33475 = ~n33472 & ~n33474 ;
  assign n33476 = n33459 & ~n33475 ;
  assign n33477 = ~n32461 & n33475 ;
  assign n33478 = ~n32931 & n33477 ;
  assign n33479 = n32456 & n33477 ;
  assign n33480 = ~n33478 & ~n33479 ;
  assign n33481 = ~n33476 & n33480 ;
  assign n33482 = n33456 & n33481 ;
  assign n33483 = ~n33456 & ~n33481 ;
  assign n33484 = ~n33482 & ~n33483 ;
  assign n33485 = ~n32434 & ~n32934 ;
  assign n33486 = ~n32435 & ~n33485 ;
  assign n33487 = n33484 & n33486 ;
  assign n33488 = ~n33484 & ~n33486 ;
  assign n33489 = ~n33487 & ~n33488 ;
  assign n33490 = ~n32938 & n33489 ;
  assign n33491 = ~n32950 & n33490 ;
  assign n33492 = ~n32938 & ~n32950 ;
  assign n33493 = ~n33489 & ~n33492 ;
  assign n33494 = ~n33491 & ~n33493 ;
  assign n33495 = ~n33487 & ~n33491 ;
  assign n33496 = ~n33476 & ~n33480 ;
  assign n33497 = ~n33456 & ~n33476 ;
  assign n33498 = ~n33496 & ~n33497 ;
  assign n33499 = ~n32983 & ~n33453 ;
  assign n33500 = n32976 & ~n32983 ;
  assign n33501 = ~n33499 & ~n33500 ;
  assign n33502 = n1965 & ~n22461 ;
  assign n33503 = ~n22459 & n33502 ;
  assign n33504 = \b[63]  & n1963 ;
  assign n33505 = \a[18]  & \b[62]  ;
  assign n33506 = n28047 & n33505 ;
  assign n33507 = ~n33504 & ~n33506 ;
  assign n33508 = \b[61]  & n2218 ;
  assign n33509 = n2216 & n33508 ;
  assign n33510 = ~\a[18]  & \b[62]  ;
  assign n33511 = n1957 & n33510 ;
  assign n33512 = ~n33509 & ~n33511 ;
  assign n33513 = n33507 & n33512 ;
  assign n33514 = ~n33503 & n33513 ;
  assign n33515 = ~\a[20]  & ~n33514 ;
  assign n33516 = \a[20]  & n33513 ;
  assign n33517 = ~n33503 & n33516 ;
  assign n33518 = ~n33515 & ~n33517 ;
  assign n33519 = n33501 & ~n33518 ;
  assign n33520 = ~n33501 & n33518 ;
  assign n33521 = ~n33519 & ~n33520 ;
  assign n33522 = n3402 & ~n17690 ;
  assign n33523 = ~n17688 & n33522 ;
  assign n33524 = \b[57]  & n3400 ;
  assign n33525 = \a[24]  & \b[56]  ;
  assign n33526 = n27626 & n33525 ;
  assign n33527 = ~n33524 & ~n33526 ;
  assign n33528 = \b[55]  & n3733 ;
  assign n33529 = n3730 & n33528 ;
  assign n33530 = ~\a[24]  & \b[56]  ;
  assign n33531 = n3394 & n33530 ;
  assign n33532 = ~n33529 & ~n33531 ;
  assign n33533 = n33527 & n33532 ;
  assign n33534 = ~n33523 & n33533 ;
  assign n33535 = ~\a[26]  & ~n33534 ;
  assign n33536 = \a[26]  & n33533 ;
  assign n33537 = ~n33523 & n33536 ;
  assign n33538 = ~n33535 & ~n33537 ;
  assign n33539 = ~n33017 & ~n33418 ;
  assign n33540 = n33010 & ~n33017 ;
  assign n33541 = ~n33539 & ~n33540 ;
  assign n33542 = ~n33538 & n33541 ;
  assign n33543 = n33538 & ~n33541 ;
  assign n33544 = ~n33542 & ~n33543 ;
  assign n33545 = ~n33314 & ~n33335 ;
  assign n33546 = n33340 & ~n33545 ;
  assign n33547 = n33198 & ~n33224 ;
  assign n33548 = n33222 & ~n33547 ;
  assign n33549 = ~n33198 & n33224 ;
  assign n33550 = ~n5852 & n13125 ;
  assign n33551 = ~n5809 & n13125 ;
  assign n33552 = ~n5848 & n33551 ;
  assign n33553 = ~n33550 & ~n33552 ;
  assign n33554 = ~n5855 & ~n33553 ;
  assign n33555 = \b[31]  & n13794 ;
  assign n33556 = n13792 & n33555 ;
  assign n33557 = ~\a[48]  & \b[32]  ;
  assign n33558 = n13117 & n33557 ;
  assign n33559 = ~n33556 & ~n33558 ;
  assign n33560 = \b[33]  & n13123 ;
  assign n33561 = \a[48]  & \b[32]  ;
  assign n33562 = n13786 & n33561 ;
  assign n33563 = \a[50]  & ~n33562 ;
  assign n33564 = ~n33560 & n33563 ;
  assign n33565 = n33559 & n33564 ;
  assign n33566 = ~n33554 & n33565 ;
  assign n33567 = ~n33560 & ~n33562 ;
  assign n33568 = n33559 & n33567 ;
  assign n33569 = ~\a[50]  & ~n33568 ;
  assign n33570 = ~\a[50]  & ~n5855 ;
  assign n33571 = ~n33553 & n33570 ;
  assign n33572 = ~n33569 & ~n33571 ;
  assign n33573 = ~n33566 & n33572 ;
  assign n33574 = ~n33549 & ~n33573 ;
  assign n33575 = ~n33548 & n33574 ;
  assign n33576 = n33549 & n33573 ;
  assign n33577 = n33222 & n33573 ;
  assign n33578 = ~n33547 & n33577 ;
  assign n33579 = ~n33576 & ~n33578 ;
  assign n33580 = ~n33575 & n33579 ;
  assign n33581 = n7337 & n11572 ;
  assign n33582 = ~n7334 & n33581 ;
  assign n33583 = n11572 & n24138 ;
  assign n33584 = ~n7333 & n33583 ;
  assign n33585 = \b[34]  & n12159 ;
  assign n33586 = n12156 & n33585 ;
  assign n33587 = ~\a[45]  & \b[35]  ;
  assign n33588 = n11564 & n33587 ;
  assign n33589 = ~n33586 & ~n33588 ;
  assign n33590 = \b[36]  & n11570 ;
  assign n33591 = \a[45]  & \b[35]  ;
  assign n33592 = n11561 & n33591 ;
  assign n33593 = \a[47]  & ~n33592 ;
  assign n33594 = ~n33590 & n33593 ;
  assign n33595 = n33589 & n33594 ;
  assign n33596 = ~n33584 & n33595 ;
  assign n33597 = ~n33582 & n33596 ;
  assign n33598 = ~n33590 & ~n33592 ;
  assign n33599 = n33589 & n33598 ;
  assign n33600 = ~n33584 & n33599 ;
  assign n33601 = ~n33582 & n33600 ;
  assign n33602 = ~\a[47]  & ~n33601 ;
  assign n33603 = ~n33597 & ~n33602 ;
  assign n33604 = ~n33137 & ~n33152 ;
  assign n33605 = ~n33155 & n33604 ;
  assign n33606 = ~n33136 & ~n33605 ;
  assign n33607 = ~n3283 & ~n17912 ;
  assign n33608 = ~n18513 & n33607 ;
  assign n33609 = n3280 & n33608 ;
  assign n33610 = n3283 & ~n17912 ;
  assign n33611 = ~n18513 & n33610 ;
  assign n33612 = ~n3280 & n33611 ;
  assign n33613 = ~n33609 & ~n33612 ;
  assign n33614 = \b[22]  & n19183 ;
  assign n33615 = n19180 & n33614 ;
  assign n33616 = \b[24]  & n18514 ;
  assign n33617 = \a[56]  & \b[23]  ;
  assign n33618 = n19181 & n33617 ;
  assign n33619 = ~\a[57]  & \b[23]  ;
  assign n33620 = n18508 & n33619 ;
  assign n33621 = ~n33618 & ~n33620 ;
  assign n33622 = ~n33616 & n33621 ;
  assign n33623 = ~n33615 & n33622 ;
  assign n33624 = n33613 & n33623 ;
  assign n33625 = ~\a[59]  & ~n33624 ;
  assign n33626 = \a[59]  & n33623 ;
  assign n33627 = n33613 & n33626 ;
  assign n33628 = ~n33625 & ~n33627 ;
  assign n33629 = ~n33120 & ~n33127 ;
  assign n33630 = ~n33123 & n33629 ;
  assign n33631 = ~n2523 & n20521 ;
  assign n33632 = ~n2521 & n33631 ;
  assign n33633 = \b[21]  & n20519 ;
  assign n33634 = \a[60]  & \b[20]  ;
  assign n33635 = n20510 & n33634 ;
  assign n33636 = ~n33633 & ~n33635 ;
  assign n33637 = \b[19]  & n21315 ;
  assign n33638 = n21312 & n33637 ;
  assign n33639 = ~\a[60]  & \b[20]  ;
  assign n33640 = n20513 & n33639 ;
  assign n33641 = ~n33638 & ~n33640 ;
  assign n33642 = n33636 & n33641 ;
  assign n33643 = ~n33632 & n33642 ;
  assign n33644 = ~\a[17]  & \b[17]  ;
  assign n33645 = n21957 & n33644 ;
  assign n33646 = ~\a[17]  & \b[18]  ;
  assign n33647 = n21958 & n33646 ;
  assign n33648 = ~n33645 & ~n33647 ;
  assign n33649 = \b[18]  & n21958 ;
  assign n33650 = \b[17]  & n21957 ;
  assign n33651 = \a[17]  & ~n33650 ;
  assign n33652 = ~n33649 & n33651 ;
  assign n33653 = n33648 & ~n33652 ;
  assign n33654 = ~\a[62]  & ~n33118 ;
  assign n33655 = ~n33653 & n33654 ;
  assign n33656 = ~\a[62]  & n33118 ;
  assign n33657 = n33653 & n33656 ;
  assign n33658 = ~n33655 & ~n33657 ;
  assign n33659 = ~n33643 & ~n33658 ;
  assign n33660 = \a[62]  & ~n33118 ;
  assign n33661 = ~n33653 & n33660 ;
  assign n33662 = \a[62]  & n33118 ;
  assign n33663 = n33653 & n33662 ;
  assign n33664 = ~n33661 & ~n33663 ;
  assign n33665 = n33642 & ~n33664 ;
  assign n33666 = ~n33632 & n33665 ;
  assign n33667 = ~n33659 & ~n33666 ;
  assign n33668 = ~\a[62]  & ~n33643 ;
  assign n33669 = ~n33118 & ~n33653 ;
  assign n33670 = n33118 & n33653 ;
  assign n33671 = ~n33669 & ~n33670 ;
  assign n33672 = \a[62]  & n33642 ;
  assign n33673 = ~n33632 & n33672 ;
  assign n33674 = n33671 & ~n33673 ;
  assign n33675 = ~n33668 & n33674 ;
  assign n33676 = n33667 & ~n33675 ;
  assign n33677 = ~n33630 & ~n33676 ;
  assign n33678 = n33630 & ~n33666 ;
  assign n33679 = ~n33659 & n33678 ;
  assign n33680 = ~n33675 & n33679 ;
  assign n33681 = ~n33677 & ~n33680 ;
  assign n33682 = n33628 & n33681 ;
  assign n33683 = ~n33628 & ~n33681 ;
  assign n33684 = ~n33682 & ~n33683 ;
  assign n33685 = n33606 & n33684 ;
  assign n33686 = ~n33606 & ~n33684 ;
  assign n33687 = ~n33685 & ~n33686 ;
  assign n33688 = ~n4145 & n16655 ;
  assign n33689 = ~n3603 & n16655 ;
  assign n33690 = ~n4141 & n33689 ;
  assign n33691 = ~n33688 & ~n33690 ;
  assign n33692 = ~n4148 & ~n33691 ;
  assign n33693 = \b[25]  & n17308 ;
  assign n33694 = n17305 & n33693 ;
  assign n33695 = \b[27]  & n16653 ;
  assign n33696 = \a[54]  & \b[26]  ;
  assign n33697 = n16644 & n33696 ;
  assign n33698 = ~\a[54]  & \b[26]  ;
  assign n33699 = n16647 & n33698 ;
  assign n33700 = ~n33697 & ~n33699 ;
  assign n33701 = ~n33695 & n33700 ;
  assign n33702 = ~n33694 & n33701 ;
  assign n33703 = ~\a[56]  & n33702 ;
  assign n33704 = ~n33692 & n33703 ;
  assign n33705 = \a[56]  & ~n33702 ;
  assign n33706 = \a[56]  & ~n4148 ;
  assign n33707 = ~n33691 & n33706 ;
  assign n33708 = ~n33705 & ~n33707 ;
  assign n33709 = ~n33704 & n33708 ;
  assign n33710 = n33157 & ~n33160 ;
  assign n33711 = n33158 & ~n33160 ;
  assign n33712 = ~n33710 & ~n33711 ;
  assign n33713 = n33096 & ~n33162 ;
  assign n33714 = n33712 & ~n33713 ;
  assign n33715 = ~n33709 & ~n33714 ;
  assign n33716 = n33709 & n33712 ;
  assign n33717 = ~n33713 & n33716 ;
  assign n33718 = ~n33715 & ~n33717 ;
  assign n33719 = ~n33687 & ~n33718 ;
  assign n33720 = n33687 & ~n33717 ;
  assign n33721 = ~n33715 & n33720 ;
  assign n33722 = ~n5105 & ~n14276 ;
  assign n33723 = ~n14790 & n33722 ;
  assign n33724 = n5102 & n33723 ;
  assign n33725 = n5105 & ~n14276 ;
  assign n33726 = ~n14790 & n33725 ;
  assign n33727 = ~n5102 & n33726 ;
  assign n33728 = ~n33724 & ~n33727 ;
  assign n33729 = \b[28]  & n15517 ;
  assign n33730 = n15514 & n33729 ;
  assign n33731 = ~\a[51]  & \b[29]  ;
  assign n33732 = n14785 & n33731 ;
  assign n33733 = ~n33730 & ~n33732 ;
  assign n33734 = \b[30]  & n14791 ;
  assign n33735 = \a[51]  & \b[29]  ;
  assign n33736 = n14782 & n33735 ;
  assign n33737 = \a[53]  & ~n33736 ;
  assign n33738 = ~n33734 & n33737 ;
  assign n33739 = n33733 & n33738 ;
  assign n33740 = n33728 & n33739 ;
  assign n33741 = ~n33734 & ~n33736 ;
  assign n33742 = n33733 & n33741 ;
  assign n33743 = n33728 & n33742 ;
  assign n33744 = ~\a[53]  & ~n33743 ;
  assign n33745 = ~n33740 & ~n33744 ;
  assign n33746 = ~n33721 & ~n33745 ;
  assign n33747 = ~n33719 & n33746 ;
  assign n33748 = ~n33719 & ~n33721 ;
  assign n33749 = n33745 & ~n33748 ;
  assign n33750 = ~n33747 & ~n33749 ;
  assign n33751 = ~n33174 & n33195 ;
  assign n33752 = ~n33175 & ~n33751 ;
  assign n33753 = ~n33750 & ~n33752 ;
  assign n33754 = ~n33747 & n33752 ;
  assign n33755 = ~n33749 & n33754 ;
  assign n33756 = ~n33753 & ~n33755 ;
  assign n33757 = ~n33603 & n33756 ;
  assign n33758 = ~n33580 & n33757 ;
  assign n33759 = ~n33603 & ~n33756 ;
  assign n33760 = n33580 & n33759 ;
  assign n33761 = ~n33758 & ~n33760 ;
  assign n33762 = n33603 & ~n33756 ;
  assign n33763 = ~n33580 & n33762 ;
  assign n33764 = n33603 & n33756 ;
  assign n33765 = n33580 & n33764 ;
  assign n33766 = ~n33763 & ~n33765 ;
  assign n33767 = n33761 & n33766 ;
  assign n33768 = n33235 & ~n33237 ;
  assign n33769 = ~n33235 & n33237 ;
  assign n33770 = n33261 & ~n33769 ;
  assign n33771 = ~n33768 & ~n33770 ;
  assign n33772 = ~n8602 & n10082 ;
  assign n33773 = ~n8600 & n33772 ;
  assign n33774 = \b[37]  & n10681 ;
  assign n33775 = n10678 & n33774 ;
  assign n33776 = \b[39]  & n10080 ;
  assign n33777 = \a[41]  & \b[38]  ;
  assign n33778 = n10679 & n33777 ;
  assign n33779 = ~\a[42]  & \b[38]  ;
  assign n33780 = n10074 & n33779 ;
  assign n33781 = ~n33778 & ~n33780 ;
  assign n33782 = ~n33776 & n33781 ;
  assign n33783 = ~n33775 & n33782 ;
  assign n33784 = ~n33773 & n33783 ;
  assign n33785 = ~\a[44]  & ~n33784 ;
  assign n33786 = \a[44]  & n33783 ;
  assign n33787 = ~n33773 & n33786 ;
  assign n33788 = ~n33785 & ~n33787 ;
  assign n33789 = ~n33771 & ~n33788 ;
  assign n33790 = n33767 & n33789 ;
  assign n33791 = n33771 & ~n33788 ;
  assign n33792 = ~n33767 & n33791 ;
  assign n33793 = ~n33790 & ~n33792 ;
  assign n33794 = ~n33771 & n33788 ;
  assign n33795 = ~n33767 & n33794 ;
  assign n33796 = n33771 & n33788 ;
  assign n33797 = n33767 & n33796 ;
  assign n33798 = ~n33795 & ~n33797 ;
  assign n33799 = n33793 & n33798 ;
  assign n33800 = n8759 & n9930 ;
  assign n33801 = ~n9927 & n33800 ;
  assign n33802 = n8759 & n11358 ;
  assign n33803 = ~n9926 & n33802 ;
  assign n33804 = \b[40]  & n9301 ;
  assign n33805 = n9298 & n33804 ;
  assign n33806 = ~\a[39]  & \b[41]  ;
  assign n33807 = n8751 & n33806 ;
  assign n33808 = ~n33805 & ~n33807 ;
  assign n33809 = \b[42]  & n8757 ;
  assign n33810 = \a[39]  & \b[41]  ;
  assign n33811 = n8748 & n33810 ;
  assign n33812 = \a[41]  & ~n33811 ;
  assign n33813 = ~n33809 & n33812 ;
  assign n33814 = n33808 & n33813 ;
  assign n33815 = ~n33803 & n33814 ;
  assign n33816 = ~n33801 & n33815 ;
  assign n33817 = ~n33809 & ~n33811 ;
  assign n33818 = n33808 & n33817 ;
  assign n33819 = ~n33803 & n33818 ;
  assign n33820 = ~n33801 & n33819 ;
  assign n33821 = ~\a[41]  & ~n33820 ;
  assign n33822 = ~n33816 & ~n33821 ;
  assign n33823 = n33272 & n33297 ;
  assign n33824 = n33302 & ~n33823 ;
  assign n33825 = ~n33822 & ~n33824 ;
  assign n33826 = ~n33799 & n33825 ;
  assign n33827 = ~n33822 & n33824 ;
  assign n33828 = n33799 & n33827 ;
  assign n33829 = ~n33826 & ~n33828 ;
  assign n33830 = n33822 & n33824 ;
  assign n33831 = ~n33799 & n33830 ;
  assign n33832 = n33822 & ~n33824 ;
  assign n33833 = n33799 & n33832 ;
  assign n33834 = ~n33831 & ~n33833 ;
  assign n33835 = n33829 & n33834 ;
  assign n33836 = n33070 & ~n33309 ;
  assign n33837 = ~n33310 & ~n33836 ;
  assign n33838 = n7534 & ~n11397 ;
  assign n33839 = ~n11395 & n33838 ;
  assign n33840 = \b[45]  & n7532 ;
  assign n33841 = \a[36]  & \b[44]  ;
  assign n33842 = n17801 & n33841 ;
  assign n33843 = ~n33840 & ~n33842 ;
  assign n33844 = \b[43]  & n7973 ;
  assign n33845 = n7970 & n33844 ;
  assign n33846 = ~\a[36]  & \b[44]  ;
  assign n33847 = n7526 & n33846 ;
  assign n33848 = ~n33845 & ~n33847 ;
  assign n33849 = n33843 & n33848 ;
  assign n33850 = ~n33839 & n33849 ;
  assign n33851 = ~\a[38]  & ~n33850 ;
  assign n33852 = \a[38]  & n33849 ;
  assign n33853 = ~n33839 & n33852 ;
  assign n33854 = ~n33851 & ~n33853 ;
  assign n33855 = n33837 & ~n33854 ;
  assign n33856 = ~n33835 & n33855 ;
  assign n33857 = ~n33837 & ~n33854 ;
  assign n33858 = n33835 & n33857 ;
  assign n33859 = ~n33856 & ~n33858 ;
  assign n33860 = ~n33837 & n33854 ;
  assign n33861 = ~n33835 & n33860 ;
  assign n33862 = n33837 & n33854 ;
  assign n33863 = n33835 & n33862 ;
  assign n33864 = ~n33861 & ~n33863 ;
  assign n33865 = n33859 & n33864 ;
  assign n33866 = n33546 & ~n33865 ;
  assign n33867 = ~n33546 & n33865 ;
  assign n33868 = ~n33866 & ~n33867 ;
  assign n33869 = n6309 & n12478 ;
  assign n33870 = ~n12475 & n33869 ;
  assign n33871 = n6309 & n28668 ;
  assign n33872 = ~n12474 & n33871 ;
  assign n33873 = \b[46]  & n6778 ;
  assign n33874 = n6775 & n33873 ;
  assign n33875 = ~\a[33]  & \b[47]  ;
  assign n33876 = n6301 & n33875 ;
  assign n33877 = ~n33874 & ~n33876 ;
  assign n33878 = \b[48]  & n6307 ;
  assign n33879 = \a[33]  & \b[47]  ;
  assign n33880 = n6298 & n33879 ;
  assign n33881 = \a[35]  & ~n33880 ;
  assign n33882 = ~n33878 & n33881 ;
  assign n33883 = n33877 & n33882 ;
  assign n33884 = ~n33872 & n33883 ;
  assign n33885 = ~n33870 & n33884 ;
  assign n33886 = ~n33878 & ~n33880 ;
  assign n33887 = n33877 & n33886 ;
  assign n33888 = ~n33872 & n33887 ;
  assign n33889 = ~n33870 & n33888 ;
  assign n33890 = ~\a[35]  & ~n33889 ;
  assign n33891 = ~n33885 & ~n33890 ;
  assign n33892 = n33868 & ~n33891 ;
  assign n33893 = ~n33868 & n33891 ;
  assign n33894 = ~n33892 & ~n33893 ;
  assign n33895 = ~n33346 & ~n33350 ;
  assign n33896 = n33346 & n33350 ;
  assign n33897 = n33369 & ~n33896 ;
  assign n33898 = ~n33895 & ~n33897 ;
  assign n33899 = ~n33894 & ~n33898 ;
  assign n33900 = n33894 & n33898 ;
  assign n33901 = ~n33899 & ~n33900 ;
  assign n33902 = n5211 & ~n14098 ;
  assign n33903 = ~n14096 & n33902 ;
  assign n33904 = \b[51]  & n5209 ;
  assign n33905 = \a[30]  & \b[50]  ;
  assign n33906 = n5200 & n33905 ;
  assign n33907 = ~n33904 & ~n33906 ;
  assign n33908 = \b[49]  & n5595 ;
  assign n33909 = n5592 & n33908 ;
  assign n33910 = ~\a[30]  & \b[50]  ;
  assign n33911 = n5203 & n33910 ;
  assign n33912 = ~n33909 & ~n33911 ;
  assign n33913 = n33907 & n33912 ;
  assign n33914 = ~n33903 & n33913 ;
  assign n33915 = ~\a[32]  & ~n33914 ;
  assign n33916 = \a[32]  & n33913 ;
  assign n33917 = ~n33903 & n33916 ;
  assign n33918 = ~n33915 & ~n33917 ;
  assign n33919 = ~n33045 & n33380 ;
  assign n33920 = ~n32848 & n33038 ;
  assign n33921 = ~n33019 & n33920 ;
  assign n33922 = \a[32]  & n33037 ;
  assign n33923 = ~n32848 & n33922 ;
  assign n33924 = ~n33019 & n33923 ;
  assign n33925 = ~n33921 & ~n33924 ;
  assign n33926 = ~n33919 & n33925 ;
  assign n33927 = ~n33918 & ~n33926 ;
  assign n33928 = n33918 & ~n33921 ;
  assign n33929 = ~n33924 & n33928 ;
  assign n33930 = ~n33919 & n33929 ;
  assign n33931 = ~n33927 & ~n33930 ;
  assign n33932 = n33901 & n33931 ;
  assign n33933 = ~n33901 & ~n33931 ;
  assign n33934 = ~n33932 & ~n33933 ;
  assign n33935 = n33383 & ~n33414 ;
  assign n33936 = n33407 & ~n33935 ;
  assign n33937 = n4249 & ~n16398 ;
  assign n33938 = ~n15241 & n33937 ;
  assign n33939 = ~n16404 & n33938 ;
  assign n33940 = n4249 & n16398 ;
  assign n33941 = n15241 & n33940 ;
  assign n33942 = n16400 & n33940 ;
  assign n33943 = ~n15239 & n33942 ;
  assign n33944 = ~n33941 & ~n33943 ;
  assign n33945 = ~n33939 & n33944 ;
  assign n33946 = \b[52]  & n4647 ;
  assign n33947 = n4644 & n33946 ;
  assign n33948 = ~\a[27]  & \b[53]  ;
  assign n33949 = n4241 & n33948 ;
  assign n33950 = ~n33947 & ~n33949 ;
  assign n33951 = \b[54]  & n4247 ;
  assign n33952 = \a[27]  & \b[53]  ;
  assign n33953 = n4238 & n33952 ;
  assign n33954 = \a[29]  & ~n33953 ;
  assign n33955 = ~n33951 & n33954 ;
  assign n33956 = n33950 & n33955 ;
  assign n33957 = n33945 & n33956 ;
  assign n33958 = ~n33951 & ~n33953 ;
  assign n33959 = n33950 & n33958 ;
  assign n33960 = n33945 & n33959 ;
  assign n33961 = ~\a[29]  & ~n33960 ;
  assign n33962 = ~n33957 & ~n33961 ;
  assign n33963 = ~n33936 & ~n33962 ;
  assign n33964 = n33407 & n33962 ;
  assign n33965 = ~n33935 & n33964 ;
  assign n33966 = ~n33963 & ~n33965 ;
  assign n33967 = ~n33934 & ~n33966 ;
  assign n33968 = n33934 & n33966 ;
  assign n33969 = ~n33967 & ~n33968 ;
  assign n33970 = n33544 & n33969 ;
  assign n33971 = ~n33544 & ~n33969 ;
  assign n33972 = ~n33970 & ~n33971 ;
  assign n33973 = n33421 & ~n33449 ;
  assign n33974 = ~n33441 & ~n33973 ;
  assign n33975 = n2622 & n20260 ;
  assign n33976 = ~n20257 & n33975 ;
  assign n33977 = n2622 & ~n20260 ;
  assign n33978 = ~n19545 & n33977 ;
  assign n33979 = ~n20256 & n33978 ;
  assign n33980 = \b[58]  & n2912 ;
  assign n33981 = n2909 & n33980 ;
  assign n33982 = \b[60]  & n2620 ;
  assign n33983 = \a[20]  & \b[59]  ;
  assign n33984 = n2910 & n33983 ;
  assign n33985 = ~\a[21]  & \b[59]  ;
  assign n33986 = n2614 & n33985 ;
  assign n33987 = ~n33984 & ~n33986 ;
  assign n33988 = ~n33982 & n33987 ;
  assign n33989 = ~n33981 & n33988 ;
  assign n33990 = ~n33979 & n33989 ;
  assign n33991 = ~n33976 & n33990 ;
  assign n33992 = ~\a[23]  & ~n33991 ;
  assign n33993 = \a[23]  & n33989 ;
  assign n33994 = ~n33979 & n33993 ;
  assign n33995 = ~n33976 & n33994 ;
  assign n33996 = ~n33992 & ~n33995 ;
  assign n33997 = ~n33974 & ~n33996 ;
  assign n33998 = ~n33441 & n33996 ;
  assign n33999 = ~n33973 & n33998 ;
  assign n34000 = ~n33997 & ~n33999 ;
  assign n34001 = ~n33972 & ~n34000 ;
  assign n34002 = n33972 & n34000 ;
  assign n34003 = ~n34001 & ~n34002 ;
  assign n34004 = n33521 & n34003 ;
  assign n34005 = ~n33521 & ~n34003 ;
  assign n34006 = ~n34004 & ~n34005 ;
  assign n34007 = n33498 & n34006 ;
  assign n34008 = ~n33498 & ~n34006 ;
  assign n34009 = ~n34007 & ~n34008 ;
  assign n34010 = ~n33495 & n34009 ;
  assign n34011 = ~n33487 & ~n34009 ;
  assign n34012 = ~n33491 & n34011 ;
  assign n34013 = ~n34010 & ~n34012 ;
  assign n34014 = ~n33487 & ~n34007 ;
  assign n34015 = ~n33491 & n34014 ;
  assign n34016 = ~n33519 & ~n34003 ;
  assign n34017 = ~n33520 & ~n34016 ;
  assign n34018 = ~n33972 & ~n33997 ;
  assign n34019 = \b[62]  & n2218 ;
  assign n34020 = n2216 & n34019 ;
  assign n34021 = ~\a[18]  & \b[63]  ;
  assign n34022 = n1957 & n34021 ;
  assign n34023 = \a[18]  & \b[63]  ;
  assign n34024 = n28047 & n34023 ;
  assign n34025 = ~n34022 & ~n34024 ;
  assign n34026 = ~n34020 & n34025 ;
  assign n34027 = ~\a[20]  & ~n34026 ;
  assign n34028 = n1965 & ~n22458 ;
  assign n34029 = ~\a[20]  & n34028 ;
  assign n34030 = ~n23173 & n34029 ;
  assign n34031 = ~n34027 & ~n34030 ;
  assign n34032 = ~n23173 & n34028 ;
  assign n34033 = \a[20]  & n34026 ;
  assign n34034 = ~n34032 & n34033 ;
  assign n34035 = n34031 & ~n34034 ;
  assign n34036 = ~n33999 & ~n34035 ;
  assign n34037 = ~n34018 & n34036 ;
  assign n34038 = ~n33999 & ~n34018 ;
  assign n34039 = n34035 & ~n34038 ;
  assign n34040 = ~n34037 & ~n34039 ;
  assign n34041 = ~n33542 & ~n33969 ;
  assign n34042 = ~n33543 & ~n34041 ;
  assign n34043 = n2622 & ~n20971 ;
  assign n34044 = ~n20969 & n34043 ;
  assign n34045 = \b[59]  & n2912 ;
  assign n34046 = n2909 & n34045 ;
  assign n34047 = \b[61]  & n2620 ;
  assign n34048 = \a[20]  & \b[60]  ;
  assign n34049 = n2910 & n34048 ;
  assign n34050 = ~\a[21]  & \b[60]  ;
  assign n34051 = n2614 & n34050 ;
  assign n34052 = ~n34049 & ~n34051 ;
  assign n34053 = ~n34047 & n34052 ;
  assign n34054 = ~n34046 & n34053 ;
  assign n34055 = ~n34044 & n34054 ;
  assign n34056 = ~\a[23]  & ~n34055 ;
  assign n34057 = \a[23]  & n34054 ;
  assign n34058 = ~n34044 & n34057 ;
  assign n34059 = ~n34056 & ~n34058 ;
  assign n34060 = ~n34042 & n34059 ;
  assign n34061 = ~n33543 & ~n34059 ;
  assign n34062 = ~n34041 & n34061 ;
  assign n34063 = ~n34060 & ~n34062 ;
  assign n34064 = n3402 & n18940 ;
  assign n34065 = ~n18937 & n34064 ;
  assign n34066 = n3402 & ~n18940 ;
  assign n34067 = ~n17685 & n34066 ;
  assign n34068 = ~n18936 & n34067 ;
  assign n34069 = \b[56]  & n3733 ;
  assign n34070 = n3730 & n34069 ;
  assign n34071 = ~\a[24]  & \b[57]  ;
  assign n34072 = n3394 & n34071 ;
  assign n34073 = ~n34070 & ~n34072 ;
  assign n34074 = \b[58]  & n3400 ;
  assign n34075 = \a[24]  & \b[57]  ;
  assign n34076 = n27626 & n34075 ;
  assign n34077 = \a[26]  & ~n34076 ;
  assign n34078 = ~n34074 & n34077 ;
  assign n34079 = n34073 & n34078 ;
  assign n34080 = ~n34068 & n34079 ;
  assign n34081 = ~n34065 & n34080 ;
  assign n34082 = ~n34074 & ~n34076 ;
  assign n34083 = n34073 & n34082 ;
  assign n34084 = ~n34068 & n34083 ;
  assign n34085 = ~n34065 & n34084 ;
  assign n34086 = ~\a[26]  & ~n34085 ;
  assign n34087 = ~n34081 & ~n34086 ;
  assign n34088 = ~n33934 & ~n33963 ;
  assign n34089 = ~n33965 & ~n34088 ;
  assign n34090 = n34087 & ~n34089 ;
  assign n34091 = ~n33965 & ~n34087 ;
  assign n34092 = ~n34088 & n34091 ;
  assign n34093 = n33901 & ~n33930 ;
  assign n34094 = n4249 & ~n16446 ;
  assign n34095 = ~n16444 & n34094 ;
  assign n34096 = \b[55]  & n4247 ;
  assign n34097 = \a[27]  & \b[54]  ;
  assign n34098 = n4238 & n34097 ;
  assign n34099 = ~n34096 & ~n34098 ;
  assign n34100 = \b[53]  & n4647 ;
  assign n34101 = n4644 & n34100 ;
  assign n34102 = ~\a[27]  & \b[54]  ;
  assign n34103 = n4241 & n34102 ;
  assign n34104 = ~n34101 & ~n34103 ;
  assign n34105 = n34099 & n34104 ;
  assign n34106 = ~n34095 & n34105 ;
  assign n34107 = ~\a[29]  & ~n34106 ;
  assign n34108 = \a[29]  & n34105 ;
  assign n34109 = ~n34095 & n34108 ;
  assign n34110 = ~n34107 & ~n34109 ;
  assign n34111 = ~n33927 & n34110 ;
  assign n34112 = ~n34093 & n34111 ;
  assign n34113 = ~n33927 & ~n34093 ;
  assign n34114 = \a[29]  & ~n34106 ;
  assign n34115 = ~\a[29]  & n34106 ;
  assign n34116 = ~n34114 & ~n34115 ;
  assign n34117 = ~n34113 & n34116 ;
  assign n34118 = ~n34112 & ~n34117 ;
  assign n34119 = ~n33892 & ~n33898 ;
  assign n34120 = ~n33893 & ~n34119 ;
  assign n34121 = n5211 & n15201 ;
  assign n34122 = ~n15198 & n34121 ;
  assign n34123 = n5211 & ~n15201 ;
  assign n34124 = ~n14093 & n34123 ;
  assign n34125 = ~n15197 & n34124 ;
  assign n34126 = \b[52]  & n5209 ;
  assign n34127 = \a[30]  & \b[51]  ;
  assign n34128 = n5200 & n34127 ;
  assign n34129 = ~n34126 & ~n34128 ;
  assign n34130 = \b[50]  & n5595 ;
  assign n34131 = n5592 & n34130 ;
  assign n34132 = ~\a[30]  & \b[51]  ;
  assign n34133 = n5203 & n34132 ;
  assign n34134 = ~n34131 & ~n34133 ;
  assign n34135 = n34129 & n34134 ;
  assign n34136 = ~n34125 & n34135 ;
  assign n34137 = ~n34122 & n34136 ;
  assign n34138 = ~\a[32]  & ~n34137 ;
  assign n34139 = \a[32]  & ~n34128 ;
  assign n34140 = ~n34126 & n34139 ;
  assign n34141 = n34134 & n34140 ;
  assign n34142 = ~n34125 & n34141 ;
  assign n34143 = ~n34122 & n34142 ;
  assign n34144 = ~n34138 & ~n34143 ;
  assign n34145 = ~n34120 & n34144 ;
  assign n34146 = \a[32]  & ~n34137 ;
  assign n34147 = ~\a[32]  & n34137 ;
  assign n34148 = ~n34146 & ~n34147 ;
  assign n34149 = ~n33893 & n34148 ;
  assign n34150 = ~n34119 & n34149 ;
  assign n34151 = ~n34145 & ~n34150 ;
  assign n34152 = n33546 & n33859 ;
  assign n34153 = n33864 & ~n34152 ;
  assign n34154 = n4456 & n16655 ;
  assign n34155 = ~n18723 & n34154 ;
  assign n34156 = n16655 & n16805 ;
  assign n34157 = ~n4452 & n34156 ;
  assign n34158 = \b[26]  & n17308 ;
  assign n34159 = n17305 & n34158 ;
  assign n34160 = \b[28]  & n16653 ;
  assign n34161 = \a[54]  & \b[27]  ;
  assign n34162 = n16644 & n34161 ;
  assign n34163 = ~\a[54]  & \b[27]  ;
  assign n34164 = n16647 & n34163 ;
  assign n34165 = ~n34162 & ~n34164 ;
  assign n34166 = ~n34160 & n34165 ;
  assign n34167 = ~n34159 & n34166 ;
  assign n34168 = ~n34157 & n34167 ;
  assign n34169 = ~n34155 & n34168 ;
  assign n34170 = ~\a[56]  & ~n34169 ;
  assign n34171 = \a[56]  & n34167 ;
  assign n34172 = ~n34157 & n34171 ;
  assign n34173 = ~n34155 & n34172 ;
  assign n34174 = ~n34170 & ~n34173 ;
  assign n34175 = ~n33606 & ~n33683 ;
  assign n34176 = ~n33682 & ~n34175 ;
  assign n34177 = n2768 & n20521 ;
  assign n34178 = ~n2765 & n34177 ;
  assign n34179 = n20521 & n32597 ;
  assign n34180 = ~n2764 & n34179 ;
  assign n34181 = \b[22]  & n20519 ;
  assign n34182 = \a[60]  & \b[21]  ;
  assign n34183 = n20510 & n34182 ;
  assign n34184 = ~n34181 & ~n34183 ;
  assign n34185 = \b[20]  & n21315 ;
  assign n34186 = n21312 & n34185 ;
  assign n34187 = ~\a[60]  & \b[21]  ;
  assign n34188 = n20513 & n34187 ;
  assign n34189 = ~n34186 & ~n34188 ;
  assign n34190 = n34184 & n34189 ;
  assign n34191 = ~n34180 & n34190 ;
  assign n34192 = ~n34178 & n34191 ;
  assign n34193 = ~\a[62]  & ~n34192 ;
  assign n34194 = n33118 & n33648 ;
  assign n34195 = n33648 & n33652 ;
  assign n34196 = ~n34194 & ~n34195 ;
  assign n34197 = \b[19]  & n21958 ;
  assign n34198 = \b[18]  & n21957 ;
  assign n34199 = ~n34197 & ~n34198 ;
  assign n34200 = ~n34196 & ~n34199 ;
  assign n34201 = n34196 & n34199 ;
  assign n34202 = ~n34200 & ~n34201 ;
  assign n34203 = \a[62]  & n34190 ;
  assign n34204 = ~n34180 & n34203 ;
  assign n34205 = ~n34178 & n34204 ;
  assign n34206 = ~n34202 & ~n34205 ;
  assign n34207 = ~n34193 & n34206 ;
  assign n34208 = ~\a[62]  & n34202 ;
  assign n34209 = ~n34192 & n34208 ;
  assign n34210 = \a[62]  & ~n34199 ;
  assign n34211 = n34196 & n34210 ;
  assign n34212 = \a[62]  & n34199 ;
  assign n34213 = ~n34196 & n34212 ;
  assign n34214 = ~n34211 & ~n34213 ;
  assign n34215 = n34190 & ~n34214 ;
  assign n34216 = ~n34180 & n34215 ;
  assign n34217 = ~n34178 & n34216 ;
  assign n34218 = ~n34209 & ~n34217 ;
  assign n34219 = ~n34207 & n34218 ;
  assign n34220 = ~n33630 & ~n33675 ;
  assign n34221 = n33667 & ~n34220 ;
  assign n34222 = n34219 & ~n34221 ;
  assign n34223 = ~n34219 & n34221 ;
  assign n34224 = ~n34222 & ~n34223 ;
  assign n34225 = \b[23]  & n19183 ;
  assign n34226 = n19180 & n34225 ;
  assign n34227 = \b[25]  & n18514 ;
  assign n34228 = \a[56]  & \b[24]  ;
  assign n34229 = n19181 & n34228 ;
  assign n34230 = ~\a[57]  & \b[24]  ;
  assign n34231 = n18508 & n34230 ;
  assign n34232 = ~n34229 & ~n34231 ;
  assign n34233 = ~n34227 & n34232 ;
  assign n34234 = ~n34226 & n34233 ;
  assign n34235 = ~\a[59]  & ~n34234 ;
  assign n34236 = ~n3564 & n18516 ;
  assign n34237 = ~n3282 & n18516 ;
  assign n34238 = ~n3560 & n34237 ;
  assign n34239 = ~n34236 & ~n34238 ;
  assign n34240 = ~\a[59]  & ~n3567 ;
  assign n34241 = ~n34239 & n34240 ;
  assign n34242 = ~n34235 & ~n34241 ;
  assign n34243 = ~n3567 & ~n34239 ;
  assign n34244 = \a[59]  & ~n34226 ;
  assign n34245 = n34233 & n34244 ;
  assign n34246 = ~n34243 & n34245 ;
  assign n34247 = n34242 & ~n34246 ;
  assign n34248 = ~n34224 & n34247 ;
  assign n34249 = n34224 & ~n34247 ;
  assign n34250 = ~n34248 & ~n34249 ;
  assign n34251 = n34176 & n34250 ;
  assign n34252 = ~n34176 & ~n34250 ;
  assign n34253 = ~n34251 & ~n34252 ;
  assign n34254 = n34174 & ~n34253 ;
  assign n34255 = ~n34174 & n34253 ;
  assign n34256 = ~n34254 & ~n34255 ;
  assign n34257 = n33687 & n33709 ;
  assign n34258 = ~n33687 & ~n33709 ;
  assign n34259 = ~n34257 & n34258 ;
  assign n34260 = ~n33714 & ~n34257 ;
  assign n34261 = ~n34259 & ~n34260 ;
  assign n34262 = n34256 & n34261 ;
  assign n34263 = ~n34256 & ~n34261 ;
  assign n34264 = ~n34262 & ~n34263 ;
  assign n34265 = ~n5462 & n14793 ;
  assign n34266 = ~n5460 & n34265 ;
  assign n34267 = \b[29]  & n15517 ;
  assign n34268 = n15514 & n34267 ;
  assign n34269 = ~\a[51]  & \b[30]  ;
  assign n34270 = n14785 & n34269 ;
  assign n34271 = ~n34268 & ~n34270 ;
  assign n34272 = \b[31]  & n14791 ;
  assign n34273 = \a[51]  & \b[30]  ;
  assign n34274 = n14782 & n34273 ;
  assign n34275 = \a[53]  & ~n34274 ;
  assign n34276 = ~n34272 & n34275 ;
  assign n34277 = n34271 & n34276 ;
  assign n34278 = ~n34266 & n34277 ;
  assign n34279 = ~n34272 & ~n34274 ;
  assign n34280 = n34271 & n34279 ;
  assign n34281 = ~n34266 & n34280 ;
  assign n34282 = ~\a[53]  & ~n34281 ;
  assign n34283 = ~n34278 & ~n34282 ;
  assign n34284 = ~n34264 & n34283 ;
  assign n34285 = n34264 & ~n34283 ;
  assign n34286 = ~n34284 & ~n34285 ;
  assign n34287 = ~n33747 & ~n33752 ;
  assign n34288 = ~n33749 & ~n34287 ;
  assign n34289 = n6565 & n13125 ;
  assign n34290 = ~n6562 & n34289 ;
  assign n34291 = n13125 & n22947 ;
  assign n34292 = ~n6561 & n34291 ;
  assign n34293 = \b[32]  & n13794 ;
  assign n34294 = n13792 & n34293 ;
  assign n34295 = ~\a[48]  & \b[33]  ;
  assign n34296 = n13117 & n34295 ;
  assign n34297 = ~n34294 & ~n34296 ;
  assign n34298 = \b[34]  & n13123 ;
  assign n34299 = \a[48]  & \b[33]  ;
  assign n34300 = n13786 & n34299 ;
  assign n34301 = \a[50]  & ~n34300 ;
  assign n34302 = ~n34298 & n34301 ;
  assign n34303 = n34297 & n34302 ;
  assign n34304 = ~n34292 & n34303 ;
  assign n34305 = ~n34290 & n34304 ;
  assign n34306 = ~n34298 & ~n34300 ;
  assign n34307 = n34297 & n34306 ;
  assign n34308 = ~n34292 & n34307 ;
  assign n34309 = ~n34290 & n34308 ;
  assign n34310 = ~\a[50]  & ~n34309 ;
  assign n34311 = ~n34305 & ~n34310 ;
  assign n34312 = n34288 & ~n34311 ;
  assign n34313 = ~n34286 & n34312 ;
  assign n34314 = ~n34288 & ~n34311 ;
  assign n34315 = n34286 & n34314 ;
  assign n34316 = ~n34313 & ~n34315 ;
  assign n34317 = ~n34288 & n34311 ;
  assign n34318 = ~n34286 & n34317 ;
  assign n34319 = n34288 & n34311 ;
  assign n34320 = n34286 & n34319 ;
  assign n34321 = ~n34318 & ~n34320 ;
  assign n34322 = n34316 & n34321 ;
  assign n34323 = ~n33575 & ~n33756 ;
  assign n34324 = n33579 & ~n34323 ;
  assign n34325 = ~n34322 & ~n34324 ;
  assign n34326 = n34322 & n34324 ;
  assign n34327 = ~n34325 & ~n34326 ;
  assign n34328 = ~n7758 & n11572 ;
  assign n34329 = ~n7336 & n11572 ;
  assign n34330 = ~n7754 & n34329 ;
  assign n34331 = ~n34328 & ~n34330 ;
  assign n34332 = ~n7761 & ~n34331 ;
  assign n34333 = \b[35]  & n12159 ;
  assign n34334 = n12156 & n34333 ;
  assign n34335 = ~\a[45]  & \b[36]  ;
  assign n34336 = n11564 & n34335 ;
  assign n34337 = ~n34334 & ~n34336 ;
  assign n34338 = \b[37]  & n11570 ;
  assign n34339 = \a[45]  & \b[36]  ;
  assign n34340 = n11561 & n34339 ;
  assign n34341 = \a[47]  & ~n34340 ;
  assign n34342 = ~n34338 & n34341 ;
  assign n34343 = n34337 & n34342 ;
  assign n34344 = ~n34332 & n34343 ;
  assign n34345 = ~n34338 & ~n34340 ;
  assign n34346 = n34337 & n34345 ;
  assign n34347 = ~\a[47]  & ~n34346 ;
  assign n34348 = ~\a[47]  & ~n7761 ;
  assign n34349 = ~n34331 & n34348 ;
  assign n34350 = ~n34347 & ~n34349 ;
  assign n34351 = ~n34344 & n34350 ;
  assign n34352 = ~n34327 & n34351 ;
  assign n34353 = n34327 & ~n34351 ;
  assign n34354 = ~n34352 & ~n34353 ;
  assign n34355 = n9044 & n10082 ;
  assign n34356 = ~n9041 & n34355 ;
  assign n34357 = ~n9044 & n10082 ;
  assign n34358 = ~n8597 & n34357 ;
  assign n34359 = ~n9040 & n34358 ;
  assign n34360 = \b[38]  & n10681 ;
  assign n34361 = n10678 & n34360 ;
  assign n34362 = \b[40]  & n10080 ;
  assign n34363 = \a[41]  & \b[39]  ;
  assign n34364 = n10679 & n34363 ;
  assign n34365 = ~\a[42]  & \b[39]  ;
  assign n34366 = n10074 & n34365 ;
  assign n34367 = ~n34364 & ~n34366 ;
  assign n34368 = ~n34362 & n34367 ;
  assign n34369 = ~n34361 & n34368 ;
  assign n34370 = ~n34359 & n34369 ;
  assign n34371 = ~n34356 & n34370 ;
  assign n34372 = ~\a[44]  & ~n34371 ;
  assign n34373 = \a[44]  & n34369 ;
  assign n34374 = ~n34359 & n34373 ;
  assign n34375 = ~n34356 & n34374 ;
  assign n34376 = ~n34372 & ~n34375 ;
  assign n34377 = n33761 & ~n33771 ;
  assign n34378 = n33766 & ~n34377 ;
  assign n34379 = ~n34376 & n34378 ;
  assign n34380 = ~n34354 & n34379 ;
  assign n34381 = ~n34376 & ~n34378 ;
  assign n34382 = n34354 & n34381 ;
  assign n34383 = ~n34380 & ~n34382 ;
  assign n34384 = n34376 & ~n34378 ;
  assign n34385 = ~n34354 & n34384 ;
  assign n34386 = n34376 & n34378 ;
  assign n34387 = n34354 & n34386 ;
  assign n34388 = ~n34385 & ~n34387 ;
  assign n34389 = n34383 & n34388 ;
  assign n34390 = n33793 & n33824 ;
  assign n34391 = n33798 & ~n34390 ;
  assign n34392 = n8759 & ~n10409 ;
  assign n34393 = ~n10407 & n34392 ;
  assign n34394 = \b[41]  & n9301 ;
  assign n34395 = n9298 & n34394 ;
  assign n34396 = ~\a[39]  & \b[42]  ;
  assign n34397 = n8751 & n34396 ;
  assign n34398 = ~n34395 & ~n34397 ;
  assign n34399 = \b[43]  & n8757 ;
  assign n34400 = \a[39]  & \b[42]  ;
  assign n34401 = n8748 & n34400 ;
  assign n34402 = \a[41]  & ~n34401 ;
  assign n34403 = ~n34399 & n34402 ;
  assign n34404 = n34398 & n34403 ;
  assign n34405 = ~n34393 & n34404 ;
  assign n34406 = ~n34399 & ~n34401 ;
  assign n34407 = n34398 & n34406 ;
  assign n34408 = ~n34393 & n34407 ;
  assign n34409 = ~\a[41]  & ~n34408 ;
  assign n34410 = ~n34405 & ~n34409 ;
  assign n34411 = n34391 & ~n34410 ;
  assign n34412 = ~n34389 & n34411 ;
  assign n34413 = ~n34391 & ~n34410 ;
  assign n34414 = n34389 & n34413 ;
  assign n34415 = ~n34412 & ~n34414 ;
  assign n34416 = ~n34391 & n34410 ;
  assign n34417 = ~n34389 & n34416 ;
  assign n34418 = n34391 & n34410 ;
  assign n34419 = n34389 & n34418 ;
  assign n34420 = ~n34417 & ~n34419 ;
  assign n34421 = n34415 & n34420 ;
  assign n34422 = n33829 & ~n33837 ;
  assign n34423 = n33834 & ~n34422 ;
  assign n34424 = n7534 & n11906 ;
  assign n34425 = ~n11903 & n34424 ;
  assign n34426 = n7534 & ~n11906 ;
  assign n34427 = ~n11392 & n34426 ;
  assign n34428 = ~n11902 & n34427 ;
  assign n34429 = \b[44]  & n7973 ;
  assign n34430 = n7970 & n34429 ;
  assign n34431 = ~\a[36]  & \b[45]  ;
  assign n34432 = n7526 & n34431 ;
  assign n34433 = ~n34430 & ~n34432 ;
  assign n34434 = \b[46]  & n7532 ;
  assign n34435 = \a[36]  & \b[45]  ;
  assign n34436 = n17801 & n34435 ;
  assign n34437 = \a[38]  & ~n34436 ;
  assign n34438 = ~n34434 & n34437 ;
  assign n34439 = n34433 & n34438 ;
  assign n34440 = ~n34428 & n34439 ;
  assign n34441 = ~n34425 & n34440 ;
  assign n34442 = ~n34434 & ~n34436 ;
  assign n34443 = n34433 & n34442 ;
  assign n34444 = ~n34428 & n34443 ;
  assign n34445 = ~n34425 & n34444 ;
  assign n34446 = ~\a[38]  & ~n34445 ;
  assign n34447 = ~n34441 & ~n34446 ;
  assign n34448 = ~n34423 & n34447 ;
  assign n34449 = ~n34421 & n34448 ;
  assign n34450 = n34423 & n34447 ;
  assign n34451 = n34421 & n34450 ;
  assign n34452 = ~n34449 & ~n34451 ;
  assign n34453 = n34423 & ~n34447 ;
  assign n34454 = ~n34421 & n34453 ;
  assign n34455 = ~n34423 & ~n34447 ;
  assign n34456 = n34421 & n34455 ;
  assign n34457 = ~n34454 & ~n34456 ;
  assign n34458 = n34452 & n34457 ;
  assign n34459 = ~n34153 & ~n34458 ;
  assign n34460 = n34153 & n34458 ;
  assign n34461 = ~n34459 & ~n34460 ;
  assign n34462 = n6309 & ~n13524 ;
  assign n34463 = ~n13522 & n34462 ;
  assign n34464 = \b[47]  & n6778 ;
  assign n34465 = n6775 & n34464 ;
  assign n34466 = ~\a[33]  & \b[48]  ;
  assign n34467 = n6301 & n34466 ;
  assign n34468 = ~n34465 & ~n34467 ;
  assign n34469 = \b[49]  & n6307 ;
  assign n34470 = \a[33]  & \b[48]  ;
  assign n34471 = n6298 & n34470 ;
  assign n34472 = \a[35]  & ~n34471 ;
  assign n34473 = ~n34469 & n34472 ;
  assign n34474 = n34468 & n34473 ;
  assign n34475 = ~n34463 & n34474 ;
  assign n34476 = ~n34469 & ~n34471 ;
  assign n34477 = n34468 & n34476 ;
  assign n34478 = ~n34463 & n34477 ;
  assign n34479 = ~\a[35]  & ~n34478 ;
  assign n34480 = ~n34475 & ~n34479 ;
  assign n34481 = n34461 & ~n34480 ;
  assign n34482 = ~n34461 & n34480 ;
  assign n34483 = ~n34481 & ~n34482 ;
  assign n34484 = n34151 & n34483 ;
  assign n34485 = ~n34151 & ~n34483 ;
  assign n34486 = ~n34484 & ~n34485 ;
  assign n34487 = n34118 & n34486 ;
  assign n34488 = ~n34118 & ~n34486 ;
  assign n34489 = ~n34487 & ~n34488 ;
  assign n34490 = ~n34092 & n34489 ;
  assign n34491 = ~n34090 & n34490 ;
  assign n34492 = n34090 & ~n34489 ;
  assign n34493 = ~n34087 & n34089 ;
  assign n34494 = ~n34489 & n34493 ;
  assign n34495 = ~n34492 & ~n34494 ;
  assign n34496 = ~n34491 & n34495 ;
  assign n34497 = n34063 & n34496 ;
  assign n34498 = ~n34063 & ~n34496 ;
  assign n34499 = ~n34497 & ~n34498 ;
  assign n34500 = n34040 & n34499 ;
  assign n34501 = ~n34040 & ~n34499 ;
  assign n34502 = ~n34500 & ~n34501 ;
  assign n34503 = n34017 & n34502 ;
  assign n34504 = ~n34017 & ~n34502 ;
  assign n34505 = ~n34503 & ~n34504 ;
  assign n34506 = ~n34008 & n34505 ;
  assign n34507 = ~n34015 & n34506 ;
  assign n34508 = ~n34008 & ~n34015 ;
  assign n34509 = ~n34505 & ~n34508 ;
  assign n34510 = ~n34507 & ~n34509 ;
  assign n34511 = ~n34503 & ~n34507 ;
  assign n34512 = ~n34037 & ~n34499 ;
  assign n34513 = ~n34039 & ~n34512 ;
  assign n34514 = ~n34062 & ~n34496 ;
  assign n34515 = \b[63]  & n1965 ;
  assign n34516 = ~n21694 & n34515 ;
  assign n34517 = ~n23171 & n34516 ;
  assign n34518 = \a[17]  & \a[19]  ;
  assign n34519 = \a[18]  & ~\a[20]  ;
  assign n34520 = n34518 & n34519 ;
  assign n34521 = ~\a[17]  & ~\a[19]  ;
  assign n34522 = ~\a[18]  & \a[20]  ;
  assign n34523 = n34521 & n34522 ;
  assign n34524 = ~n34520 & ~n34523 ;
  assign n34525 = \b[63]  & ~n34524 ;
  assign n34526 = \a[20]  & ~n34525 ;
  assign n34527 = ~n34517 & n34526 ;
  assign n34528 = ~n34517 & ~n34525 ;
  assign n34529 = ~\a[20]  & ~n34528 ;
  assign n34530 = ~n34527 & ~n34529 ;
  assign n34531 = ~n34060 & ~n34530 ;
  assign n34532 = ~n34514 & n34531 ;
  assign n34533 = n34060 & n34530 ;
  assign n34534 = ~n34062 & n34530 ;
  assign n34535 = ~n34496 & n34534 ;
  assign n34536 = ~n34533 & ~n34535 ;
  assign n34537 = ~n34532 & n34536 ;
  assign n34538 = ~n34092 & ~n34489 ;
  assign n34539 = n34090 & ~n34092 ;
  assign n34540 = ~n34538 & ~n34539 ;
  assign n34541 = n2622 & n21696 ;
  assign n34542 = ~n21693 & n34541 ;
  assign n34543 = n2622 & ~n21696 ;
  assign n34544 = ~n20966 & n34543 ;
  assign n34545 = ~n21692 & n34544 ;
  assign n34546 = \b[60]  & n2912 ;
  assign n34547 = n2909 & n34546 ;
  assign n34548 = \b[62]  & n2620 ;
  assign n34549 = \a[20]  & \b[61]  ;
  assign n34550 = n2910 & n34549 ;
  assign n34551 = ~\a[21]  & \b[61]  ;
  assign n34552 = n2614 & n34551 ;
  assign n34553 = ~n34550 & ~n34552 ;
  assign n34554 = ~n34548 & n34553 ;
  assign n34555 = ~n34547 & n34554 ;
  assign n34556 = ~n34545 & n34555 ;
  assign n34557 = ~n34542 & n34556 ;
  assign n34558 = \a[23]  & ~n34557 ;
  assign n34559 = ~\a[23]  & n34557 ;
  assign n34560 = ~n34558 & ~n34559 ;
  assign n34561 = n34540 & n34560 ;
  assign n34562 = ~\a[23]  & ~n34557 ;
  assign n34563 = \a[23]  & n34555 ;
  assign n34564 = ~n34545 & n34563 ;
  assign n34565 = ~n34542 & n34564 ;
  assign n34566 = ~n34562 & ~n34565 ;
  assign n34567 = ~n34540 & n34566 ;
  assign n34568 = ~n34561 & ~n34567 ;
  assign n34569 = ~n34117 & ~n34486 ;
  assign n34570 = ~n33927 & n34114 ;
  assign n34571 = ~n34093 & n34570 ;
  assign n34572 = ~n33927 & n34115 ;
  assign n34573 = ~n34093 & n34572 ;
  assign n34574 = ~n34571 & ~n34573 ;
  assign n34575 = ~n34569 & n34574 ;
  assign n34576 = n3402 & ~n19550 ;
  assign n34577 = ~n19548 & n34576 ;
  assign n34578 = \b[59]  & n3400 ;
  assign n34579 = \a[24]  & \b[58]  ;
  assign n34580 = n27626 & n34579 ;
  assign n34581 = ~n34578 & ~n34580 ;
  assign n34582 = \b[57]  & n3733 ;
  assign n34583 = n3730 & n34582 ;
  assign n34584 = ~\a[24]  & \b[58]  ;
  assign n34585 = n3394 & n34584 ;
  assign n34586 = ~n34583 & ~n34585 ;
  assign n34587 = n34581 & n34586 ;
  assign n34588 = ~n34577 & n34587 ;
  assign n34589 = ~\a[26]  & ~n34588 ;
  assign n34590 = \a[26]  & n34587 ;
  assign n34591 = ~n34577 & n34590 ;
  assign n34592 = ~n34589 & ~n34591 ;
  assign n34593 = ~n34575 & n34592 ;
  assign n34594 = ~n34569 & ~n34592 ;
  assign n34595 = n34574 & n34594 ;
  assign n34596 = ~n34593 & ~n34595 ;
  assign n34597 = n5211 & ~n15246 ;
  assign n34598 = ~n15244 & n34597 ;
  assign n34599 = \b[53]  & n5209 ;
  assign n34600 = \a[30]  & \b[52]  ;
  assign n34601 = n5200 & n34600 ;
  assign n34602 = ~n34599 & ~n34601 ;
  assign n34603 = \b[51]  & n5595 ;
  assign n34604 = n5592 & n34603 ;
  assign n34605 = ~\a[30]  & \b[52]  ;
  assign n34606 = n5203 & n34605 ;
  assign n34607 = ~n34604 & ~n34606 ;
  assign n34608 = n34602 & n34607 ;
  assign n34609 = ~n34598 & n34608 ;
  assign n34610 = ~\a[32]  & ~n34609 ;
  assign n34611 = \a[32]  & n34608 ;
  assign n34612 = ~n34598 & n34611 ;
  assign n34613 = n34459 & ~n34612 ;
  assign n34614 = n34480 & ~n34612 ;
  assign n34615 = ~n34460 & n34614 ;
  assign n34616 = ~n34613 & ~n34615 ;
  assign n34617 = ~n34610 & ~n34616 ;
  assign n34618 = ~n34460 & n34480 ;
  assign n34619 = ~n34610 & ~n34612 ;
  assign n34620 = ~n34618 & ~n34619 ;
  assign n34621 = ~n34459 & n34620 ;
  assign n34622 = ~n34617 & ~n34621 ;
  assign n34623 = n8759 & ~n28007 ;
  assign n34624 = ~n28005 & n34623 ;
  assign n34625 = \b[42]  & n9301 ;
  assign n34626 = n9298 & n34625 ;
  assign n34627 = ~\a[39]  & \b[43]  ;
  assign n34628 = n8751 & n34627 ;
  assign n34629 = ~n34626 & ~n34628 ;
  assign n34630 = \b[44]  & n8757 ;
  assign n34631 = \a[39]  & \b[43]  ;
  assign n34632 = n8748 & n34631 ;
  assign n34633 = \a[41]  & ~n34632 ;
  assign n34634 = ~n34630 & n34633 ;
  assign n34635 = n34629 & n34634 ;
  assign n34636 = ~n34624 & n34635 ;
  assign n34637 = ~n34630 & ~n34632 ;
  assign n34638 = n34629 & n34637 ;
  assign n34639 = ~n34624 & n34638 ;
  assign n34640 = ~\a[41]  & ~n34639 ;
  assign n34641 = ~n34636 & ~n34640 ;
  assign n34642 = n34354 & n34378 ;
  assign n34643 = n34383 & ~n34642 ;
  assign n34644 = ~n5810 & ~n14276 ;
  assign n34645 = ~n14790 & n34644 ;
  assign n34646 = n5807 & n34645 ;
  assign n34647 = n5810 & ~n14276 ;
  assign n34648 = ~n14790 & n34647 ;
  assign n34649 = ~n5807 & n34648 ;
  assign n34650 = ~n34646 & ~n34649 ;
  assign n34651 = \b[30]  & n15517 ;
  assign n34652 = n15514 & n34651 ;
  assign n34653 = ~\a[51]  & \b[31]  ;
  assign n34654 = n14785 & n34653 ;
  assign n34655 = ~n34652 & ~n34654 ;
  assign n34656 = \b[32]  & n14791 ;
  assign n34657 = \a[51]  & \b[31]  ;
  assign n34658 = n14782 & n34657 ;
  assign n34659 = \a[53]  & ~n34658 ;
  assign n34660 = ~n34656 & n34659 ;
  assign n34661 = n34655 & n34660 ;
  assign n34662 = n34650 & n34661 ;
  assign n34663 = ~n34656 & ~n34658 ;
  assign n34664 = n34655 & n34663 ;
  assign n34665 = n34650 & n34664 ;
  assign n34666 = ~\a[53]  & ~n34665 ;
  assign n34667 = ~n34662 & ~n34666 ;
  assign n34668 = n34174 & ~n34251 ;
  assign n34669 = ~n34251 & n34252 ;
  assign n34670 = ~n34668 & ~n34669 ;
  assign n34671 = n3604 & n18516 ;
  assign n34672 = ~n19292 & n34671 ;
  assign n34673 = n12021 & n18516 ;
  assign n34674 = ~n3600 & n34673 ;
  assign n34675 = \b[26]  & n18514 ;
  assign n34676 = \a[56]  & \b[25]  ;
  assign n34677 = n19181 & n34676 ;
  assign n34678 = ~\a[57]  & \b[25]  ;
  assign n34679 = n18508 & n34678 ;
  assign n34680 = ~n34677 & ~n34679 ;
  assign n34681 = ~n34675 & n34680 ;
  assign n34682 = \b[24]  & n19183 ;
  assign n34683 = n19180 & n34682 ;
  assign n34684 = \a[59]  & ~n34683 ;
  assign n34685 = n34681 & n34684 ;
  assign n34686 = ~n34674 & n34685 ;
  assign n34687 = ~n34672 & n34686 ;
  assign n34688 = n34681 & ~n34683 ;
  assign n34689 = ~n34674 & n34688 ;
  assign n34690 = ~n34672 & n34689 ;
  assign n34691 = ~\a[59]  & ~n34690 ;
  assign n34692 = ~n34687 & ~n34691 ;
  assign n34693 = ~n3022 & n20521 ;
  assign n34694 = ~n3020 & n34693 ;
  assign n34695 = \b[23]  & n20519 ;
  assign n34696 = \a[60]  & \b[22]  ;
  assign n34697 = n20510 & n34696 ;
  assign n34698 = ~n34695 & ~n34697 ;
  assign n34699 = \b[21]  & n21315 ;
  assign n34700 = n21312 & n34699 ;
  assign n34701 = ~\a[60]  & \b[22]  ;
  assign n34702 = n20513 & n34701 ;
  assign n34703 = ~n34700 & ~n34702 ;
  assign n34704 = n34698 & n34703 ;
  assign n34705 = ~n34694 & n34704 ;
  assign n34706 = ~\a[62]  & ~n34705 ;
  assign n34707 = \b[20]  & n21958 ;
  assign n34708 = \b[19]  & n21957 ;
  assign n34709 = ~n34707 & ~n34708 ;
  assign n34710 = ~n34199 & n34709 ;
  assign n34711 = n34199 & ~n34709 ;
  assign n34712 = ~n34710 & ~n34711 ;
  assign n34713 = \a[62]  & n34704 ;
  assign n34714 = ~n34694 & n34713 ;
  assign n34715 = ~n34712 & ~n34714 ;
  assign n34716 = ~n34706 & n34715 ;
  assign n34717 = ~\a[62]  & n34712 ;
  assign n34718 = ~n34705 & n34717 ;
  assign n34719 = ~n34201 & ~n34217 ;
  assign n34720 = ~n34209 & n34719 ;
  assign n34721 = \a[62]  & n34712 ;
  assign n34722 = n34704 & n34721 ;
  assign n34723 = ~n34694 & n34722 ;
  assign n34724 = ~n34720 & ~n34723 ;
  assign n34725 = ~n34718 & n34724 ;
  assign n34726 = ~n34716 & n34725 ;
  assign n34727 = ~n34718 & ~n34723 ;
  assign n34728 = ~n34716 & n34727 ;
  assign n34729 = n34720 & ~n34728 ;
  assign n34730 = ~n34726 & ~n34729 ;
  assign n34731 = n34692 & n34730 ;
  assign n34732 = ~n34692 & ~n34730 ;
  assign n34733 = ~n34731 & ~n34732 ;
  assign n34734 = ~n34223 & ~n34242 ;
  assign n34735 = n34234 & ~n34243 ;
  assign n34736 = \a[59]  & n34735 ;
  assign n34737 = ~n34223 & n34736 ;
  assign n34738 = ~n34734 & ~n34737 ;
  assign n34739 = ~n34222 & n34738 ;
  assign n34740 = ~n34733 & ~n34739 ;
  assign n34741 = n34733 & n34739 ;
  assign n34742 = ~n34740 & ~n34741 ;
  assign n34743 = ~n4499 & n16655 ;
  assign n34744 = ~n4455 & n16655 ;
  assign n34745 = ~n4495 & n34744 ;
  assign n34746 = ~n34743 & ~n34745 ;
  assign n34747 = ~n4502 & ~n34746 ;
  assign n34748 = \b[29]  & n16653 ;
  assign n34749 = \a[54]  & \b[28]  ;
  assign n34750 = n16644 & n34749 ;
  assign n34751 = ~\a[54]  & \b[28]  ;
  assign n34752 = n16647 & n34751 ;
  assign n34753 = ~n34750 & ~n34752 ;
  assign n34754 = ~n34748 & n34753 ;
  assign n34755 = \b[27]  & n17308 ;
  assign n34756 = n17305 & n34755 ;
  assign n34757 = \a[56]  & ~n34756 ;
  assign n34758 = n34754 & n34757 ;
  assign n34759 = ~n34747 & n34758 ;
  assign n34760 = n34754 & ~n34756 ;
  assign n34761 = ~\a[56]  & ~n34760 ;
  assign n34762 = ~\a[56]  & ~n4502 ;
  assign n34763 = ~n34746 & n34762 ;
  assign n34764 = ~n34761 & ~n34763 ;
  assign n34765 = ~n34759 & n34764 ;
  assign n34766 = ~n34742 & n34765 ;
  assign n34767 = n34742 & ~n34765 ;
  assign n34768 = ~n34766 & ~n34767 ;
  assign n34769 = n34670 & n34768 ;
  assign n34770 = ~n34670 & ~n34768 ;
  assign n34771 = ~n34769 & ~n34770 ;
  assign n34772 = n34667 & n34771 ;
  assign n34773 = ~n34667 & ~n34771 ;
  assign n34774 = ~n34772 & ~n34773 ;
  assign n34775 = ~n6610 & n13125 ;
  assign n34776 = ~n6608 & n34775 ;
  assign n34777 = \b[33]  & n13794 ;
  assign n34778 = n13792 & n34777 ;
  assign n34779 = ~\a[48]  & \b[34]  ;
  assign n34780 = n13117 & n34779 ;
  assign n34781 = ~n34778 & ~n34780 ;
  assign n34782 = \b[35]  & n13123 ;
  assign n34783 = \a[48]  & \b[34]  ;
  assign n34784 = n13786 & n34783 ;
  assign n34785 = \a[50]  & ~n34784 ;
  assign n34786 = ~n34782 & n34785 ;
  assign n34787 = n34781 & n34786 ;
  assign n34788 = ~n34776 & n34787 ;
  assign n34789 = ~n34782 & ~n34784 ;
  assign n34790 = n34781 & n34789 ;
  assign n34791 = ~n34776 & n34790 ;
  assign n34792 = ~\a[50]  & ~n34791 ;
  assign n34793 = ~n34788 & ~n34792 ;
  assign n34794 = ~n34262 & n34283 ;
  assign n34795 = ~n34263 & ~n34794 ;
  assign n34796 = n34793 & ~n34795 ;
  assign n34797 = ~n34774 & n34796 ;
  assign n34798 = n34793 & n34795 ;
  assign n34799 = n34774 & n34798 ;
  assign n34800 = ~n34797 & ~n34799 ;
  assign n34801 = ~n34793 & n34795 ;
  assign n34802 = ~n34774 & n34801 ;
  assign n34803 = ~n34793 & ~n34795 ;
  assign n34804 = n34774 & n34803 ;
  assign n34805 = ~n34802 & ~n34804 ;
  assign n34806 = n34800 & n34805 ;
  assign n34807 = n8175 & n11572 ;
  assign n34808 = ~n8172 & n34807 ;
  assign n34809 = n11572 & n25622 ;
  assign n34810 = ~n8171 & n34809 ;
  assign n34811 = \b[36]  & n12159 ;
  assign n34812 = n12156 & n34811 ;
  assign n34813 = ~\a[45]  & \b[37]  ;
  assign n34814 = n11564 & n34813 ;
  assign n34815 = ~n34812 & ~n34814 ;
  assign n34816 = \b[38]  & n11570 ;
  assign n34817 = \a[45]  & \b[37]  ;
  assign n34818 = n11561 & n34817 ;
  assign n34819 = \a[47]  & ~n34818 ;
  assign n34820 = ~n34816 & n34819 ;
  assign n34821 = n34815 & n34820 ;
  assign n34822 = ~n34810 & n34821 ;
  assign n34823 = ~n34808 & n34822 ;
  assign n34824 = ~n34816 & ~n34818 ;
  assign n34825 = n34815 & n34824 ;
  assign n34826 = ~n34810 & n34825 ;
  assign n34827 = ~n34808 & n34826 ;
  assign n34828 = ~\a[47]  & ~n34827 ;
  assign n34829 = ~n34823 & ~n34828 ;
  assign n34830 = ~n34286 & ~n34288 ;
  assign n34831 = n34286 & n34288 ;
  assign n34832 = n34311 & ~n34831 ;
  assign n34833 = ~n34830 & ~n34832 ;
  assign n34834 = ~n34829 & ~n34833 ;
  assign n34835 = ~n34806 & n34834 ;
  assign n34836 = ~n34829 & n34833 ;
  assign n34837 = n34806 & n34836 ;
  assign n34838 = ~n34835 & ~n34837 ;
  assign n34839 = n34829 & ~n34833 ;
  assign n34840 = n34806 & n34839 ;
  assign n34841 = n34829 & n34833 ;
  assign n34842 = ~n34806 & n34841 ;
  assign n34843 = ~n34840 & ~n34842 ;
  assign n34844 = n34838 & n34843 ;
  assign n34845 = ~n9479 & n10082 ;
  assign n34846 = ~n9043 & n10082 ;
  assign n34847 = ~n9475 & n34846 ;
  assign n34848 = ~n34845 & ~n34847 ;
  assign n34849 = ~n9482 & ~n34848 ;
  assign n34850 = \b[41]  & n10080 ;
  assign n34851 = \a[41]  & \b[40]  ;
  assign n34852 = n10679 & n34851 ;
  assign n34853 = ~\a[42]  & \b[40]  ;
  assign n34854 = n10074 & n34853 ;
  assign n34855 = ~n34852 & ~n34854 ;
  assign n34856 = ~n34850 & n34855 ;
  assign n34857 = \b[39]  & n10681 ;
  assign n34858 = n10678 & n34857 ;
  assign n34859 = \a[44]  & ~n34858 ;
  assign n34860 = n34856 & n34859 ;
  assign n34861 = ~n34849 & n34860 ;
  assign n34862 = n34856 & ~n34858 ;
  assign n34863 = ~\a[44]  & ~n34862 ;
  assign n34864 = ~\a[44]  & ~n9482 ;
  assign n34865 = ~n34848 & n34864 ;
  assign n34866 = ~n34863 & ~n34865 ;
  assign n34867 = ~n34861 & n34866 ;
  assign n34868 = ~n34326 & n34351 ;
  assign n34869 = ~n34325 & ~n34868 ;
  assign n34870 = n34867 & n34869 ;
  assign n34871 = ~n34844 & n34870 ;
  assign n34872 = n34867 & ~n34869 ;
  assign n34873 = n34844 & n34872 ;
  assign n34874 = ~n34871 & ~n34873 ;
  assign n34875 = ~n34867 & ~n34869 ;
  assign n34876 = ~n34844 & n34875 ;
  assign n34877 = ~n34867 & n34869 ;
  assign n34878 = n34844 & n34877 ;
  assign n34879 = ~n34876 & ~n34878 ;
  assign n34880 = n34874 & n34879 ;
  assign n34881 = ~n34643 & ~n34880 ;
  assign n34882 = n34643 & n34880 ;
  assign n34883 = ~n34881 & ~n34882 ;
  assign n34884 = ~n34641 & n34883 ;
  assign n34885 = n34641 & ~n34883 ;
  assign n34886 = ~n34884 & ~n34885 ;
  assign n34887 = ~n34389 & ~n34391 ;
  assign n34888 = n34389 & n34391 ;
  assign n34889 = n34410 & ~n34888 ;
  assign n34890 = ~n34887 & ~n34889 ;
  assign n34891 = n7534 & ~n12438 ;
  assign n34892 = ~n12436 & n34891 ;
  assign n34893 = \b[45]  & n7973 ;
  assign n34894 = n7970 & n34893 ;
  assign n34895 = ~\a[36]  & \b[46]  ;
  assign n34896 = n7526 & n34895 ;
  assign n34897 = ~n34894 & ~n34896 ;
  assign n34898 = \b[47]  & n7532 ;
  assign n34899 = \a[36]  & \b[46]  ;
  assign n34900 = n17801 & n34899 ;
  assign n34901 = \a[38]  & ~n34900 ;
  assign n34902 = ~n34898 & n34901 ;
  assign n34903 = n34897 & n34902 ;
  assign n34904 = ~n34892 & n34903 ;
  assign n34905 = ~n34898 & ~n34900 ;
  assign n34906 = n34897 & n34905 ;
  assign n34907 = ~n34892 & n34906 ;
  assign n34908 = ~\a[38]  & ~n34907 ;
  assign n34909 = ~n34904 & ~n34908 ;
  assign n34910 = ~n34890 & ~n34909 ;
  assign n34911 = n34886 & n34910 ;
  assign n34912 = n34890 & ~n34909 ;
  assign n34913 = ~n34886 & n34912 ;
  assign n34914 = ~n34911 & ~n34913 ;
  assign n34915 = ~n34890 & n34909 ;
  assign n34916 = ~n34886 & n34915 ;
  assign n34917 = n34890 & n34909 ;
  assign n34918 = n34886 & n34917 ;
  assign n34919 = ~n34916 & ~n34918 ;
  assign n34920 = n34914 & n34919 ;
  assign n34921 = ~n34421 & ~n34423 ;
  assign n34922 = n34421 & n34423 ;
  assign n34923 = n34447 & ~n34922 ;
  assign n34924 = ~n34921 & ~n34923 ;
  assign n34925 = n6309 & n14052 ;
  assign n34926 = ~n14049 & n34925 ;
  assign n34927 = n6309 & ~n14052 ;
  assign n34928 = ~n13519 & n34927 ;
  assign n34929 = ~n14048 & n34928 ;
  assign n34930 = \b[48]  & n6778 ;
  assign n34931 = n6775 & n34930 ;
  assign n34932 = ~\a[33]  & \b[49]  ;
  assign n34933 = n6301 & n34932 ;
  assign n34934 = ~n34931 & ~n34933 ;
  assign n34935 = \b[50]  & n6307 ;
  assign n34936 = \a[33]  & \b[49]  ;
  assign n34937 = n6298 & n34936 ;
  assign n34938 = \a[35]  & ~n34937 ;
  assign n34939 = ~n34935 & n34938 ;
  assign n34940 = n34934 & n34939 ;
  assign n34941 = ~n34929 & n34940 ;
  assign n34942 = ~n34926 & n34941 ;
  assign n34943 = ~n34935 & ~n34937 ;
  assign n34944 = n34934 & n34943 ;
  assign n34945 = ~n34929 & n34944 ;
  assign n34946 = ~n34926 & n34945 ;
  assign n34947 = ~\a[35]  & ~n34946 ;
  assign n34948 = ~n34942 & ~n34947 ;
  assign n34949 = ~n34924 & ~n34948 ;
  assign n34950 = n34920 & n34949 ;
  assign n34951 = n34924 & ~n34948 ;
  assign n34952 = ~n34920 & n34951 ;
  assign n34953 = ~n34950 & ~n34952 ;
  assign n34954 = ~n34924 & n34948 ;
  assign n34955 = ~n34920 & n34954 ;
  assign n34956 = n34924 & n34948 ;
  assign n34957 = n34920 & n34956 ;
  assign n34958 = ~n34955 & ~n34957 ;
  assign n34959 = n34953 & n34958 ;
  assign n34960 = n34622 & n34959 ;
  assign n34961 = ~n34622 & ~n34959 ;
  assign n34962 = ~n34960 & ~n34961 ;
  assign n34963 = ~n34145 & n34483 ;
  assign n34964 = ~n33893 & n34138 ;
  assign n34965 = ~n34119 & n34964 ;
  assign n34966 = \a[32]  & n34137 ;
  assign n34967 = ~n33893 & n34966 ;
  assign n34968 = ~n34119 & n34967 ;
  assign n34969 = ~n34965 & ~n34968 ;
  assign n34970 = ~n34963 & n34969 ;
  assign n34971 = n4249 & n17647 ;
  assign n34972 = ~n17644 & n34971 ;
  assign n34973 = n4249 & ~n17647 ;
  assign n34974 = ~n16441 & n34973 ;
  assign n34975 = ~n17643 & n34974 ;
  assign n34976 = \b[56]  & n4247 ;
  assign n34977 = \a[27]  & \b[55]  ;
  assign n34978 = n4238 & n34977 ;
  assign n34979 = ~n34976 & ~n34978 ;
  assign n34980 = \b[54]  & n4647 ;
  assign n34981 = n4644 & n34980 ;
  assign n34982 = ~\a[27]  & \b[55]  ;
  assign n34983 = n4241 & n34982 ;
  assign n34984 = ~n34981 & ~n34983 ;
  assign n34985 = n34979 & n34984 ;
  assign n34986 = ~n34975 & n34985 ;
  assign n34987 = ~n34972 & n34986 ;
  assign n34988 = \a[29]  & ~n34987 ;
  assign n34989 = ~\a[29]  & n34987 ;
  assign n34990 = ~n34988 & ~n34989 ;
  assign n34991 = ~n34970 & n34990 ;
  assign n34992 = ~\a[29]  & ~n34987 ;
  assign n34993 = \a[29]  & n34985 ;
  assign n34994 = ~n34975 & n34993 ;
  assign n34995 = ~n34972 & n34994 ;
  assign n34996 = ~n34965 & ~n34995 ;
  assign n34997 = ~n34968 & n34996 ;
  assign n34998 = ~n34963 & n34997 ;
  assign n34999 = ~n34992 & n34998 ;
  assign n35000 = ~n34991 & ~n34999 ;
  assign n35001 = n34962 & n35000 ;
  assign n35002 = ~n34962 & ~n35000 ;
  assign n35003 = ~n35001 & ~n35002 ;
  assign n35004 = n34596 & n35003 ;
  assign n35005 = ~n34596 & ~n35003 ;
  assign n35006 = ~n35004 & ~n35005 ;
  assign n35007 = n34568 & ~n35006 ;
  assign n35008 = ~n34568 & n35006 ;
  assign n35009 = ~n35007 & ~n35008 ;
  assign n35010 = n34537 & ~n35009 ;
  assign n35011 = ~n34537 & n35009 ;
  assign n35012 = ~n35010 & ~n35011 ;
  assign n35013 = n34513 & n35012 ;
  assign n35014 = ~n34513 & ~n35012 ;
  assign n35015 = ~n35013 & ~n35014 ;
  assign n35016 = ~n34511 & n35015 ;
  assign n35017 = ~n34503 & ~n35015 ;
  assign n35018 = ~n34507 & n35017 ;
  assign n35019 = ~n35016 & ~n35018 ;
  assign n35020 = ~n34503 & ~n35013 ;
  assign n35021 = ~n34507 & n35020 ;
  assign n35022 = ~n34532 & ~n35010 ;
  assign n35023 = ~n34595 & ~n35003 ;
  assign n35024 = ~n34593 & ~n35023 ;
  assign n35025 = n34962 & ~n34999 ;
  assign n35026 = ~n34991 & ~n35025 ;
  assign n35027 = n4249 & ~n17690 ;
  assign n35028 = ~n17688 & n35027 ;
  assign n35029 = \b[57]  & n4247 ;
  assign n35030 = \a[27]  & \b[56]  ;
  assign n35031 = n4238 & n35030 ;
  assign n35032 = ~n35029 & ~n35031 ;
  assign n35033 = \b[55]  & n4647 ;
  assign n35034 = n4644 & n35033 ;
  assign n35035 = ~\a[27]  & \b[56]  ;
  assign n35036 = n4241 & n35035 ;
  assign n35037 = ~n35034 & ~n35036 ;
  assign n35038 = n35032 & n35037 ;
  assign n35039 = ~n35028 & n35038 ;
  assign n35040 = ~\a[29]  & ~n35039 ;
  assign n35041 = \a[29]  & n35038 ;
  assign n35042 = ~n35028 & n35041 ;
  assign n35043 = ~n35040 & ~n35042 ;
  assign n35044 = ~n35026 & ~n35043 ;
  assign n35045 = ~n34991 & n35043 ;
  assign n35046 = ~n35025 & n35045 ;
  assign n35047 = ~n35044 & ~n35046 ;
  assign n35048 = n3402 & n20260 ;
  assign n35049 = ~n20257 & n35048 ;
  assign n35050 = n3402 & ~n20260 ;
  assign n35051 = ~n19545 & n35050 ;
  assign n35052 = ~n20256 & n35051 ;
  assign n35053 = \b[58]  & n3733 ;
  assign n35054 = n3730 & n35053 ;
  assign n35055 = ~\a[24]  & \b[59]  ;
  assign n35056 = n3394 & n35055 ;
  assign n35057 = ~n35054 & ~n35056 ;
  assign n35058 = \b[60]  & n3400 ;
  assign n35059 = \a[24]  & \b[59]  ;
  assign n35060 = n27626 & n35059 ;
  assign n35061 = \a[26]  & ~n35060 ;
  assign n35062 = ~n35058 & n35061 ;
  assign n35063 = n35057 & n35062 ;
  assign n35064 = ~n35052 & n35063 ;
  assign n35065 = ~n35049 & n35064 ;
  assign n35066 = ~n35058 & ~n35060 ;
  assign n35067 = n35057 & n35066 ;
  assign n35068 = ~n35052 & n35067 ;
  assign n35069 = ~n35049 & n35068 ;
  assign n35070 = ~\a[26]  & ~n35069 ;
  assign n35071 = ~n35065 & ~n35070 ;
  assign n35072 = n34920 & n34924 ;
  assign n35073 = n34953 & ~n35072 ;
  assign n35074 = n34774 & ~n34795 ;
  assign n35075 = ~n34774 & n34795 ;
  assign n35076 = n34793 & ~n35075 ;
  assign n35077 = ~n35074 & ~n35076 ;
  assign n35078 = n34667 & ~n34769 ;
  assign n35079 = ~n5852 & n14793 ;
  assign n35080 = ~n5809 & n14793 ;
  assign n35081 = ~n5848 & n35080 ;
  assign n35082 = ~n35079 & ~n35081 ;
  assign n35083 = ~n5855 & ~n35082 ;
  assign n35084 = \b[31]  & n15517 ;
  assign n35085 = n15514 & n35084 ;
  assign n35086 = ~\a[51]  & \b[32]  ;
  assign n35087 = n14785 & n35086 ;
  assign n35088 = ~n35085 & ~n35087 ;
  assign n35089 = \b[33]  & n14791 ;
  assign n35090 = \a[51]  & \b[32]  ;
  assign n35091 = n14782 & n35090 ;
  assign n35092 = \a[53]  & ~n35091 ;
  assign n35093 = ~n35089 & n35092 ;
  assign n35094 = n35088 & n35093 ;
  assign n35095 = ~n35083 & n35094 ;
  assign n35096 = ~n35089 & ~n35091 ;
  assign n35097 = n35088 & n35096 ;
  assign n35098 = ~\a[53]  & ~n35097 ;
  assign n35099 = ~\a[53]  & ~n5855 ;
  assign n35100 = ~n35082 & n35099 ;
  assign n35101 = ~n35098 & ~n35100 ;
  assign n35102 = ~n35095 & n35101 ;
  assign n35103 = ~n34770 & ~n35102 ;
  assign n35104 = ~n35078 & n35103 ;
  assign n35105 = n34770 & n35102 ;
  assign n35106 = n34667 & n35102 ;
  assign n35107 = ~n34769 & n35106 ;
  assign n35108 = ~n35105 & ~n35107 ;
  assign n35109 = ~n35104 & n35108 ;
  assign n35110 = n7337 & n13125 ;
  assign n35111 = ~n7334 & n35110 ;
  assign n35112 = ~n7337 & n13125 ;
  assign n35113 = ~n6605 & n35112 ;
  assign n35114 = ~n7333 & n35113 ;
  assign n35115 = \b[34]  & n13794 ;
  assign n35116 = n13792 & n35115 ;
  assign n35117 = ~\a[48]  & \b[35]  ;
  assign n35118 = n13117 & n35117 ;
  assign n35119 = ~n35116 & ~n35118 ;
  assign n35120 = \b[36]  & n13123 ;
  assign n35121 = \a[48]  & \b[35]  ;
  assign n35122 = n13786 & n35121 ;
  assign n35123 = \a[50]  & ~n35122 ;
  assign n35124 = ~n35120 & n35123 ;
  assign n35125 = n35119 & n35124 ;
  assign n35126 = ~n35114 & n35125 ;
  assign n35127 = ~n35111 & n35126 ;
  assign n35128 = ~n35120 & ~n35122 ;
  assign n35129 = n35119 & n35128 ;
  assign n35130 = ~n35114 & n35129 ;
  assign n35131 = ~n35111 & n35130 ;
  assign n35132 = ~\a[50]  & ~n35131 ;
  assign n35133 = ~n35127 & ~n35132 ;
  assign n35134 = ~n34740 & n34765 ;
  assign n35135 = ~n34741 & ~n35134 ;
  assign n35136 = ~n4145 & n18516 ;
  assign n35137 = ~n3603 & n18516 ;
  assign n35138 = ~n4141 & n35137 ;
  assign n35139 = ~n35136 & ~n35138 ;
  assign n35140 = ~n4148 & ~n35139 ;
  assign n35141 = \b[27]  & n18514 ;
  assign n35142 = \a[56]  & \b[26]  ;
  assign n35143 = n19181 & n35142 ;
  assign n35144 = ~\a[57]  & \b[26]  ;
  assign n35145 = n18508 & n35144 ;
  assign n35146 = ~n35143 & ~n35145 ;
  assign n35147 = ~n35141 & n35146 ;
  assign n35148 = \b[25]  & n19183 ;
  assign n35149 = n19180 & n35148 ;
  assign n35150 = \a[59]  & ~n35149 ;
  assign n35151 = n35147 & n35150 ;
  assign n35152 = ~n35140 & n35151 ;
  assign n35153 = n35147 & ~n35149 ;
  assign n35154 = ~\a[59]  & ~n35153 ;
  assign n35155 = ~\a[59]  & ~n4148 ;
  assign n35156 = ~n35139 & n35155 ;
  assign n35157 = ~n35154 & ~n35156 ;
  assign n35158 = ~n35152 & n35157 ;
  assign n35159 = n34692 & ~n34726 ;
  assign n35160 = ~n34729 & ~n35159 ;
  assign n35161 = ~n34710 & ~n34723 ;
  assign n35162 = ~n34718 & n35161 ;
  assign n35163 = ~n3283 & ~n19861 ;
  assign n35164 = ~n20518 & n35163 ;
  assign n35165 = n3280 & n35164 ;
  assign n35166 = n3283 & ~n19861 ;
  assign n35167 = ~n20518 & n35166 ;
  assign n35168 = ~n3280 & n35167 ;
  assign n35169 = ~n35165 & ~n35168 ;
  assign n35170 = \b[24]  & n20519 ;
  assign n35171 = \a[60]  & \b[23]  ;
  assign n35172 = n20510 & n35171 ;
  assign n35173 = ~n35170 & ~n35172 ;
  assign n35174 = \b[22]  & n21315 ;
  assign n35175 = n21312 & n35174 ;
  assign n35176 = ~\a[60]  & \b[23]  ;
  assign n35177 = n20513 & n35176 ;
  assign n35178 = ~n35175 & ~n35177 ;
  assign n35179 = n35173 & n35178 ;
  assign n35180 = n35169 & n35179 ;
  assign n35181 = ~\a[20]  & \b[20]  ;
  assign n35182 = n21957 & n35181 ;
  assign n35183 = ~\a[20]  & \b[21]  ;
  assign n35184 = n21958 & n35183 ;
  assign n35185 = ~n35182 & ~n35184 ;
  assign n35186 = \b[21]  & n21958 ;
  assign n35187 = \b[20]  & n21957 ;
  assign n35188 = \a[20]  & ~n35187 ;
  assign n35189 = ~n35186 & n35188 ;
  assign n35190 = n35185 & ~n35189 ;
  assign n35191 = ~\a[62]  & ~n34709 ;
  assign n35192 = ~n35190 & n35191 ;
  assign n35193 = ~\a[62]  & n34709 ;
  assign n35194 = n35190 & n35193 ;
  assign n35195 = ~n35192 & ~n35194 ;
  assign n35196 = ~n35180 & ~n35195 ;
  assign n35197 = \a[62]  & ~n34709 ;
  assign n35198 = ~n35190 & n35197 ;
  assign n35199 = \a[62]  & n34709 ;
  assign n35200 = n35190 & n35199 ;
  assign n35201 = ~n35198 & ~n35200 ;
  assign n35202 = n35179 & ~n35201 ;
  assign n35203 = n35169 & n35202 ;
  assign n35204 = ~n35196 & ~n35203 ;
  assign n35205 = ~\a[62]  & ~n35180 ;
  assign n35206 = ~n34709 & ~n35190 ;
  assign n35207 = n34709 & n35190 ;
  assign n35208 = ~n35206 & ~n35207 ;
  assign n35209 = \a[62]  & n35179 ;
  assign n35210 = n35169 & n35209 ;
  assign n35211 = n35208 & ~n35210 ;
  assign n35212 = ~n35205 & n35211 ;
  assign n35213 = n35204 & ~n35212 ;
  assign n35214 = ~n35162 & ~n35213 ;
  assign n35215 = n35162 & n35213 ;
  assign n35216 = ~n35214 & ~n35215 ;
  assign n35217 = ~n35160 & n35216 ;
  assign n35218 = n35158 & n35217 ;
  assign n35219 = ~n35160 & ~n35216 ;
  assign n35220 = ~n35158 & n35219 ;
  assign n35221 = ~n35218 & ~n35220 ;
  assign n35222 = ~n35158 & ~n35216 ;
  assign n35223 = n35158 & n35216 ;
  assign n35224 = n35160 & ~n35223 ;
  assign n35225 = ~n35222 & n35224 ;
  assign n35226 = n35221 & ~n35225 ;
  assign n35227 = ~n5105 & ~n16016 ;
  assign n35228 = ~n16652 & n35227 ;
  assign n35229 = n5102 & n35228 ;
  assign n35230 = n5105 & ~n16016 ;
  assign n35231 = ~n16652 & n35230 ;
  assign n35232 = ~n5102 & n35231 ;
  assign n35233 = ~n35229 & ~n35232 ;
  assign n35234 = \b[28]  & n17308 ;
  assign n35235 = n17305 & n35234 ;
  assign n35236 = \b[30]  & n16653 ;
  assign n35237 = \a[54]  & \b[29]  ;
  assign n35238 = n16644 & n35237 ;
  assign n35239 = ~\a[54]  & \b[29]  ;
  assign n35240 = n16647 & n35239 ;
  assign n35241 = ~n35238 & ~n35240 ;
  assign n35242 = ~n35236 & n35241 ;
  assign n35243 = ~n35235 & n35242 ;
  assign n35244 = n35233 & n35243 ;
  assign n35245 = ~\a[56]  & ~n35244 ;
  assign n35246 = \a[56]  & n35243 ;
  assign n35247 = n35233 & n35246 ;
  assign n35248 = ~n35245 & ~n35247 ;
  assign n35249 = n35226 & ~n35248 ;
  assign n35250 = ~n35226 & n35248 ;
  assign n35251 = ~n35249 & ~n35250 ;
  assign n35252 = ~n35135 & ~n35251 ;
  assign n35253 = n35135 & n35251 ;
  assign n35254 = ~n35252 & ~n35253 ;
  assign n35255 = ~n35133 & n35254 ;
  assign n35256 = ~n35109 & n35255 ;
  assign n35257 = ~n35133 & ~n35254 ;
  assign n35258 = n35109 & n35257 ;
  assign n35259 = ~n35256 & ~n35258 ;
  assign n35260 = n35133 & ~n35254 ;
  assign n35261 = ~n35109 & n35260 ;
  assign n35262 = n35133 & n35254 ;
  assign n35263 = n35109 & n35262 ;
  assign n35264 = ~n35261 & ~n35263 ;
  assign n35265 = n35259 & n35264 ;
  assign n35266 = ~n35077 & ~n35265 ;
  assign n35267 = n35077 & n35265 ;
  assign n35268 = ~n35266 & ~n35267 ;
  assign n35269 = ~n8599 & n11572 ;
  assign n35270 = ~n8174 & n11572 ;
  assign n35271 = ~n8595 & n35270 ;
  assign n35272 = ~n35269 & ~n35271 ;
  assign n35273 = ~n8602 & ~n35272 ;
  assign n35274 = \b[37]  & n12159 ;
  assign n35275 = n12156 & n35274 ;
  assign n35276 = ~\a[45]  & \b[38]  ;
  assign n35277 = n11564 & n35276 ;
  assign n35278 = ~n35275 & ~n35277 ;
  assign n35279 = \b[39]  & n11570 ;
  assign n35280 = \a[45]  & \b[38]  ;
  assign n35281 = n11561 & n35280 ;
  assign n35282 = \a[47]  & ~n35281 ;
  assign n35283 = ~n35279 & n35282 ;
  assign n35284 = n35278 & n35283 ;
  assign n35285 = ~n35273 & n35284 ;
  assign n35286 = ~n35279 & ~n35281 ;
  assign n35287 = n35278 & n35286 ;
  assign n35288 = ~\a[47]  & ~n35287 ;
  assign n35289 = ~\a[47]  & ~n8602 ;
  assign n35290 = ~n35272 & n35289 ;
  assign n35291 = ~n35288 & ~n35290 ;
  assign n35292 = ~n35285 & n35291 ;
  assign n35293 = n35268 & ~n35292 ;
  assign n35294 = ~n35268 & n35292 ;
  assign n35295 = ~n35293 & ~n35294 ;
  assign n35296 = ~n34806 & n34833 ;
  assign n35297 = n34838 & ~n35296 ;
  assign n35298 = ~n9646 & ~n9930 ;
  assign n35299 = ~n10079 & n35298 ;
  assign n35300 = n9927 & n35299 ;
  assign n35301 = ~n9646 & n9930 ;
  assign n35302 = ~n10079 & n35301 ;
  assign n35303 = ~n9927 & n35302 ;
  assign n35304 = ~n35300 & ~n35303 ;
  assign n35305 = \b[40]  & n10681 ;
  assign n35306 = n10678 & n35305 ;
  assign n35307 = \b[42]  & n10080 ;
  assign n35308 = \a[41]  & \b[41]  ;
  assign n35309 = n10679 & n35308 ;
  assign n35310 = ~\a[42]  & \b[41]  ;
  assign n35311 = n10074 & n35310 ;
  assign n35312 = ~n35309 & ~n35311 ;
  assign n35313 = ~n35307 & n35312 ;
  assign n35314 = ~n35306 & n35313 ;
  assign n35315 = n35304 & n35314 ;
  assign n35316 = ~\a[44]  & ~n35315 ;
  assign n35317 = \a[44]  & n35314 ;
  assign n35318 = n35304 & n35317 ;
  assign n35319 = ~n35316 & ~n35318 ;
  assign n35320 = ~n35297 & ~n35319 ;
  assign n35321 = ~n35295 & n35320 ;
  assign n35322 = n35297 & ~n35319 ;
  assign n35323 = n35295 & n35322 ;
  assign n35324 = ~n35321 & ~n35323 ;
  assign n35325 = n35297 & n35319 ;
  assign n35326 = ~n35295 & n35325 ;
  assign n35327 = ~n35297 & n35319 ;
  assign n35328 = n35295 & n35327 ;
  assign n35329 = ~n35326 & ~n35328 ;
  assign n35330 = n35324 & n35329 ;
  assign n35331 = ~n34844 & ~n34869 ;
  assign n35332 = n34844 & n34869 ;
  assign n35333 = n34867 & ~n35332 ;
  assign n35334 = ~n35331 & ~n35333 ;
  assign n35335 = n8759 & ~n11397 ;
  assign n35336 = ~n11395 & n35335 ;
  assign n35337 = \b[43]  & n9301 ;
  assign n35338 = n9298 & n35337 ;
  assign n35339 = ~\a[39]  & \b[44]  ;
  assign n35340 = n8751 & n35339 ;
  assign n35341 = ~n35338 & ~n35340 ;
  assign n35342 = \b[45]  & n8757 ;
  assign n35343 = \a[39]  & \b[44]  ;
  assign n35344 = n8748 & n35343 ;
  assign n35345 = \a[41]  & ~n35344 ;
  assign n35346 = ~n35342 & n35345 ;
  assign n35347 = n35341 & n35346 ;
  assign n35348 = ~n35336 & n35347 ;
  assign n35349 = ~n35342 & ~n35344 ;
  assign n35350 = n35341 & n35349 ;
  assign n35351 = ~n35336 & n35350 ;
  assign n35352 = ~\a[41]  & ~n35351 ;
  assign n35353 = ~n35348 & ~n35352 ;
  assign n35354 = n35334 & ~n35353 ;
  assign n35355 = ~n35330 & n35354 ;
  assign n35356 = ~n35334 & ~n35353 ;
  assign n35357 = n35330 & n35356 ;
  assign n35358 = ~n35355 & ~n35357 ;
  assign n35359 = ~n35334 & n35353 ;
  assign n35360 = ~n35330 & n35359 ;
  assign n35361 = n35334 & n35353 ;
  assign n35362 = n35330 & n35361 ;
  assign n35363 = ~n35360 & ~n35362 ;
  assign n35364 = n35358 & n35363 ;
  assign n35365 = n34641 & ~n34881 ;
  assign n35366 = ~n34881 & n34882 ;
  assign n35367 = ~n35365 & ~n35366 ;
  assign n35368 = n7534 & n12478 ;
  assign n35369 = ~n12475 & n35368 ;
  assign n35370 = n7534 & n28668 ;
  assign n35371 = ~n12474 & n35370 ;
  assign n35372 = \b[46]  & n7973 ;
  assign n35373 = n7970 & n35372 ;
  assign n35374 = ~\a[36]  & \b[47]  ;
  assign n35375 = n7526 & n35374 ;
  assign n35376 = ~n35373 & ~n35375 ;
  assign n35377 = \b[48]  & n7532 ;
  assign n35378 = \a[36]  & \b[47]  ;
  assign n35379 = n17801 & n35378 ;
  assign n35380 = \a[38]  & ~n35379 ;
  assign n35381 = ~n35377 & n35380 ;
  assign n35382 = n35376 & n35381 ;
  assign n35383 = ~n35371 & n35382 ;
  assign n35384 = ~n35369 & n35383 ;
  assign n35385 = ~n35377 & ~n35379 ;
  assign n35386 = n35376 & n35385 ;
  assign n35387 = ~n35371 & n35386 ;
  assign n35388 = ~n35369 & n35387 ;
  assign n35389 = ~\a[38]  & ~n35388 ;
  assign n35390 = ~n35384 & ~n35389 ;
  assign n35391 = n35367 & ~n35390 ;
  assign n35392 = ~n35364 & n35391 ;
  assign n35393 = ~n35367 & ~n35390 ;
  assign n35394 = n35364 & n35393 ;
  assign n35395 = ~n35392 & ~n35394 ;
  assign n35396 = ~n35367 & n35390 ;
  assign n35397 = ~n35364 & n35396 ;
  assign n35398 = n35367 & n35390 ;
  assign n35399 = n35364 & n35398 ;
  assign n35400 = ~n35397 & ~n35399 ;
  assign n35401 = n35395 & n35400 ;
  assign n35402 = ~n34886 & ~n34890 ;
  assign n35403 = n34886 & n34890 ;
  assign n35404 = n34909 & ~n35403 ;
  assign n35405 = ~n35402 & ~n35404 ;
  assign n35406 = ~n35401 & ~n35405 ;
  assign n35407 = n35401 & n35405 ;
  assign n35408 = ~n35406 & ~n35407 ;
  assign n35409 = n6309 & ~n14098 ;
  assign n35410 = ~n14096 & n35409 ;
  assign n35411 = \b[51]  & n6307 ;
  assign n35412 = \a[33]  & \b[50]  ;
  assign n35413 = n6298 & n35412 ;
  assign n35414 = ~n35411 & ~n35413 ;
  assign n35415 = \b[49]  & n6778 ;
  assign n35416 = n6775 & n35415 ;
  assign n35417 = ~\a[33]  & \b[50]  ;
  assign n35418 = n6301 & n35417 ;
  assign n35419 = ~n35416 & ~n35418 ;
  assign n35420 = n35414 & n35419 ;
  assign n35421 = ~n35410 & n35420 ;
  assign n35422 = ~\a[35]  & ~n35421 ;
  assign n35423 = \a[35]  & n35420 ;
  assign n35424 = ~n35410 & n35423 ;
  assign n35425 = ~n35422 & ~n35424 ;
  assign n35426 = ~n35408 & n35425 ;
  assign n35427 = n35408 & ~n35425 ;
  assign n35428 = ~n35426 & ~n35427 ;
  assign n35429 = n35073 & ~n35428 ;
  assign n35430 = ~n35073 & n35428 ;
  assign n35431 = ~n35429 & ~n35430 ;
  assign n35432 = ~n34621 & ~n34959 ;
  assign n35433 = n34618 & n34619 ;
  assign n35434 = n34459 & n34619 ;
  assign n35435 = ~n35433 & ~n35434 ;
  assign n35436 = n5211 & ~n16398 ;
  assign n35437 = ~n15241 & n35436 ;
  assign n35438 = ~n16404 & n35437 ;
  assign n35439 = n5211 & n16398 ;
  assign n35440 = n15241 & n35439 ;
  assign n35441 = n16400 & n35439 ;
  assign n35442 = ~n15239 & n35441 ;
  assign n35443 = ~n35440 & ~n35442 ;
  assign n35444 = ~n35438 & n35443 ;
  assign n35445 = \b[52]  & n5595 ;
  assign n35446 = n5592 & n35445 ;
  assign n35447 = ~\a[30]  & \b[53]  ;
  assign n35448 = n5203 & n35447 ;
  assign n35449 = ~n35446 & ~n35448 ;
  assign n35450 = \b[54]  & n5209 ;
  assign n35451 = \a[30]  & \b[53]  ;
  assign n35452 = n5200 & n35451 ;
  assign n35453 = \a[32]  & ~n35452 ;
  assign n35454 = ~n35450 & n35453 ;
  assign n35455 = n35449 & n35454 ;
  assign n35456 = n35444 & n35455 ;
  assign n35457 = ~n35450 & ~n35452 ;
  assign n35458 = n35449 & n35457 ;
  assign n35459 = n35444 & n35458 ;
  assign n35460 = ~\a[32]  & ~n35459 ;
  assign n35461 = ~n35456 & ~n35460 ;
  assign n35462 = n35435 & ~n35461 ;
  assign n35463 = ~n35432 & n35462 ;
  assign n35464 = ~n35432 & n35435 ;
  assign n35465 = n35461 & ~n35464 ;
  assign n35466 = ~n35463 & ~n35465 ;
  assign n35467 = ~n35431 & ~n35466 ;
  assign n35468 = n35431 & n35466 ;
  assign n35469 = ~n35467 & ~n35468 ;
  assign n35470 = ~n35071 & n35469 ;
  assign n35471 = ~n35047 & n35470 ;
  assign n35472 = ~n35071 & ~n35469 ;
  assign n35473 = n35047 & n35472 ;
  assign n35474 = ~n35471 & ~n35473 ;
  assign n35475 = ~n35024 & ~n35474 ;
  assign n35476 = n35071 & n35469 ;
  assign n35477 = ~n35047 & n35476 ;
  assign n35478 = n35071 & ~n35469 ;
  assign n35479 = n35047 & n35478 ;
  assign n35480 = ~n35477 & ~n35479 ;
  assign n35481 = n35024 & ~n35480 ;
  assign n35482 = ~n35475 & ~n35481 ;
  assign n35483 = n35047 & n35469 ;
  assign n35484 = ~n35047 & ~n35469 ;
  assign n35485 = ~n35483 & ~n35484 ;
  assign n35486 = ~n35024 & n35071 ;
  assign n35487 = ~n35485 & n35486 ;
  assign n35488 = ~n35047 & n35472 ;
  assign n35489 = n35047 & n35470 ;
  assign n35490 = ~n35488 & ~n35489 ;
  assign n35491 = n35024 & ~n35490 ;
  assign n35492 = ~n35487 & ~n35491 ;
  assign n35493 = n35482 & n35492 ;
  assign n35494 = ~n34561 & ~n35006 ;
  assign n35495 = ~n34561 & n34567 ;
  assign n35496 = ~n35494 & ~n35495 ;
  assign n35497 = n2622 & ~n22461 ;
  assign n35498 = ~n22459 & n35497 ;
  assign n35499 = \b[61]  & n2912 ;
  assign n35500 = n2909 & n35499 ;
  assign n35501 = \b[63]  & n2620 ;
  assign n35502 = \a[20]  & \b[62]  ;
  assign n35503 = n2910 & n35502 ;
  assign n35504 = ~\a[21]  & \b[62]  ;
  assign n35505 = n2614 & n35504 ;
  assign n35506 = ~n35503 & ~n35505 ;
  assign n35507 = ~n35501 & n35506 ;
  assign n35508 = ~n35500 & n35507 ;
  assign n35509 = ~n35498 & n35508 ;
  assign n35510 = ~\a[23]  & ~n35509 ;
  assign n35511 = \a[23]  & n35508 ;
  assign n35512 = ~n35498 & n35511 ;
  assign n35513 = ~n35510 & ~n35512 ;
  assign n35514 = n35496 & ~n35513 ;
  assign n35515 = ~n35496 & n35513 ;
  assign n35516 = ~n35514 & ~n35515 ;
  assign n35517 = n35493 & n35516 ;
  assign n35518 = ~n35493 & ~n35516 ;
  assign n35519 = ~n35517 & ~n35518 ;
  assign n35520 = n35022 & ~n35519 ;
  assign n35521 = ~n35022 & n35519 ;
  assign n35522 = ~n35520 & ~n35521 ;
  assign n35523 = ~n35014 & n35522 ;
  assign n35524 = ~n35021 & n35523 ;
  assign n35525 = ~n35014 & ~n35021 ;
  assign n35526 = ~n35522 & ~n35525 ;
  assign n35527 = ~n35524 & ~n35526 ;
  assign n35528 = ~n35493 & ~n35514 ;
  assign n35529 = ~n35515 & ~n35528 ;
  assign n35530 = ~n35024 & n35483 ;
  assign n35531 = ~n35486 & ~n35530 ;
  assign n35532 = ~n35024 & n35484 ;
  assign n35533 = ~n35047 & n35478 ;
  assign n35534 = n35047 & n35476 ;
  assign n35535 = ~n35533 & ~n35534 ;
  assign n35536 = ~n35532 & n35535 ;
  assign n35537 = n35531 & n35536 ;
  assign n35538 = \b[62]  & n2912 ;
  assign n35539 = n2909 & n35538 ;
  assign n35540 = \a[20]  & \b[63]  ;
  assign n35541 = n2910 & n35540 ;
  assign n35542 = ~\a[21]  & \b[63]  ;
  assign n35543 = n2614 & n35542 ;
  assign n35544 = ~n35541 & ~n35543 ;
  assign n35545 = ~n35539 & n35544 ;
  assign n35546 = ~\a[23]  & ~n35545 ;
  assign n35547 = n2622 & ~n22458 ;
  assign n35548 = ~\a[23]  & n35547 ;
  assign n35549 = ~n23173 & n35548 ;
  assign n35550 = ~n35546 & ~n35549 ;
  assign n35551 = ~n23173 & n35547 ;
  assign n35552 = \a[23]  & n35545 ;
  assign n35553 = ~n35551 & n35552 ;
  assign n35554 = n35550 & ~n35553 ;
  assign n35555 = n35537 & ~n35554 ;
  assign n35556 = ~n35537 & n35554 ;
  assign n35557 = ~n35555 & ~n35556 ;
  assign n35558 = ~n35044 & ~n35469 ;
  assign n35559 = ~n35046 & ~n35558 ;
  assign n35560 = n3402 & ~n20971 ;
  assign n35561 = ~n20969 & n35560 ;
  assign n35562 = \b[61]  & n3400 ;
  assign n35563 = \a[24]  & \b[60]  ;
  assign n35564 = n27626 & n35563 ;
  assign n35565 = ~n35562 & ~n35564 ;
  assign n35566 = \b[59]  & n3733 ;
  assign n35567 = n3730 & n35566 ;
  assign n35568 = ~\a[24]  & \b[60]  ;
  assign n35569 = n3394 & n35568 ;
  assign n35570 = ~n35567 & ~n35569 ;
  assign n35571 = n35565 & n35570 ;
  assign n35572 = ~n35561 & n35571 ;
  assign n35573 = ~\a[26]  & ~n35572 ;
  assign n35574 = \a[26]  & n35571 ;
  assign n35575 = ~n35561 & n35574 ;
  assign n35576 = ~n35573 & ~n35575 ;
  assign n35577 = ~n35559 & n35576 ;
  assign n35578 = ~n35046 & ~n35576 ;
  assign n35579 = ~n35558 & n35578 ;
  assign n35580 = ~n35577 & ~n35579 ;
  assign n35581 = ~n35073 & ~n35461 ;
  assign n35582 = ~n35428 & n35581 ;
  assign n35583 = n35073 & ~n35461 ;
  assign n35584 = n35428 & n35583 ;
  assign n35585 = ~n35582 & ~n35584 ;
  assign n35586 = ~n35463 & ~n35464 ;
  assign n35587 = n35585 & n35586 ;
  assign n35588 = ~n35073 & n35461 ;
  assign n35589 = ~n35428 & n35588 ;
  assign n35590 = n35073 & n35461 ;
  assign n35591 = n35428 & n35590 ;
  assign n35592 = ~n35589 & ~n35591 ;
  assign n35593 = ~n35463 & n35464 ;
  assign n35594 = n35592 & n35593 ;
  assign n35595 = ~n35587 & ~n35594 ;
  assign n35596 = n4249 & n18940 ;
  assign n35597 = ~n18937 & n35596 ;
  assign n35598 = n4249 & ~n18940 ;
  assign n35599 = ~n17685 & n35598 ;
  assign n35600 = ~n18936 & n35599 ;
  assign n35601 = \b[56]  & n4647 ;
  assign n35602 = n4644 & n35601 ;
  assign n35603 = ~\a[27]  & \b[57]  ;
  assign n35604 = n4241 & n35603 ;
  assign n35605 = ~n35602 & ~n35604 ;
  assign n35606 = \b[58]  & n4247 ;
  assign n35607 = \a[27]  & \b[57]  ;
  assign n35608 = n4238 & n35607 ;
  assign n35609 = \a[29]  & ~n35608 ;
  assign n35610 = ~n35606 & n35609 ;
  assign n35611 = n35605 & n35610 ;
  assign n35612 = ~n35600 & n35611 ;
  assign n35613 = ~n35597 & n35612 ;
  assign n35614 = ~n35606 & ~n35608 ;
  assign n35615 = n35605 & n35614 ;
  assign n35616 = ~n35600 & n35615 ;
  assign n35617 = ~n35597 & n35616 ;
  assign n35618 = ~\a[29]  & ~n35617 ;
  assign n35619 = ~n35613 & ~n35618 ;
  assign n35620 = ~n35595 & n35619 ;
  assign n35621 = n35595 & ~n35619 ;
  assign n35622 = n35073 & ~n35427 ;
  assign n35623 = n5211 & ~n16446 ;
  assign n35624 = ~n16444 & n35623 ;
  assign n35625 = \b[55]  & n5209 ;
  assign n35626 = \a[30]  & \b[54]  ;
  assign n35627 = n5200 & n35626 ;
  assign n35628 = ~n35625 & ~n35627 ;
  assign n35629 = \b[53]  & n5595 ;
  assign n35630 = n5592 & n35629 ;
  assign n35631 = ~\a[30]  & \b[54]  ;
  assign n35632 = n5203 & n35631 ;
  assign n35633 = ~n35630 & ~n35632 ;
  assign n35634 = n35628 & n35633 ;
  assign n35635 = ~n35624 & n35634 ;
  assign n35636 = \a[32]  & ~n35635 ;
  assign n35637 = ~\a[32]  & n35635 ;
  assign n35638 = ~n35636 & ~n35637 ;
  assign n35639 = ~n35426 & n35638 ;
  assign n35640 = ~n35622 & n35639 ;
  assign n35641 = ~n35426 & ~n35622 ;
  assign n35642 = ~\a[32]  & ~n35635 ;
  assign n35643 = \a[32]  & n35634 ;
  assign n35644 = ~n35624 & n35643 ;
  assign n35645 = ~n35642 & ~n35644 ;
  assign n35646 = ~n35641 & n35645 ;
  assign n35647 = ~n35640 & ~n35646 ;
  assign n35648 = n35395 & ~n35405 ;
  assign n35649 = n35400 & ~n35648 ;
  assign n35650 = n9044 & n11572 ;
  assign n35651 = ~n9041 & n35650 ;
  assign n35652 = n11572 & n27054 ;
  assign n35653 = ~n9040 & n35652 ;
  assign n35654 = \b[38]  & n12159 ;
  assign n35655 = n12156 & n35654 ;
  assign n35656 = ~\a[45]  & \b[39]  ;
  assign n35657 = n11564 & n35656 ;
  assign n35658 = ~n35655 & ~n35657 ;
  assign n35659 = \b[40]  & n11570 ;
  assign n35660 = \a[45]  & \b[39]  ;
  assign n35661 = n11561 & n35660 ;
  assign n35662 = \a[47]  & ~n35661 ;
  assign n35663 = ~n35659 & n35662 ;
  assign n35664 = n35658 & n35663 ;
  assign n35665 = ~n35653 & n35664 ;
  assign n35666 = ~n35651 & n35665 ;
  assign n35667 = ~n35659 & ~n35661 ;
  assign n35668 = n35658 & n35667 ;
  assign n35669 = ~n35653 & n35668 ;
  assign n35670 = ~n35651 & n35669 ;
  assign n35671 = ~\a[47]  & ~n35670 ;
  assign n35672 = ~n35666 & ~n35671 ;
  assign n35673 = ~n35077 & n35259 ;
  assign n35674 = n35264 & ~n35673 ;
  assign n35675 = ~n35135 & ~n35249 ;
  assign n35676 = ~n35250 & ~n35675 ;
  assign n35677 = n35158 & ~n35160 ;
  assign n35678 = ~n35217 & ~n35677 ;
  assign n35679 = ~n35223 & n35678 ;
  assign n35680 = n4456 & n18516 ;
  assign n35681 = ~n18723 & n35680 ;
  assign n35682 = n16805 & n18516 ;
  assign n35683 = ~n4452 & n35682 ;
  assign n35684 = \b[28]  & n18514 ;
  assign n35685 = \a[56]  & \b[27]  ;
  assign n35686 = n19181 & n35685 ;
  assign n35687 = ~\a[57]  & \b[27]  ;
  assign n35688 = n18508 & n35687 ;
  assign n35689 = ~n35686 & ~n35688 ;
  assign n35690 = ~n35684 & n35689 ;
  assign n35691 = \b[26]  & n19183 ;
  assign n35692 = n19180 & n35691 ;
  assign n35693 = \a[59]  & ~n35692 ;
  assign n35694 = n35690 & n35693 ;
  assign n35695 = ~n35683 & n35694 ;
  assign n35696 = ~n35681 & n35695 ;
  assign n35697 = n35690 & ~n35692 ;
  assign n35698 = ~n35683 & n35697 ;
  assign n35699 = ~n35681 & n35698 ;
  assign n35700 = ~\a[59]  & ~n35699 ;
  assign n35701 = ~n35696 & ~n35700 ;
  assign n35702 = ~n35162 & ~n35212 ;
  assign n35703 = n35204 & ~n35702 ;
  assign n35704 = \b[25]  & n20519 ;
  assign n35705 = \a[60]  & \b[24]  ;
  assign n35706 = n20510 & n35705 ;
  assign n35707 = ~n35704 & ~n35706 ;
  assign n35708 = \b[23]  & n21315 ;
  assign n35709 = n21312 & n35708 ;
  assign n35710 = ~\a[60]  & \b[24]  ;
  assign n35711 = n20513 & n35710 ;
  assign n35712 = ~n35709 & ~n35711 ;
  assign n35713 = n35707 & n35712 ;
  assign n35714 = ~n34709 & ~n35189 ;
  assign n35715 = n35185 & ~n35714 ;
  assign n35716 = \b[22]  & n21958 ;
  assign n35717 = \b[21]  & n21957 ;
  assign n35718 = ~n35716 & ~n35717 ;
  assign n35719 = ~n35715 & n35718 ;
  assign n35720 = n35185 & ~n35718 ;
  assign n35721 = ~n35714 & n35720 ;
  assign n35722 = ~\a[62]  & ~n35721 ;
  assign n35723 = ~n35719 & n35722 ;
  assign n35724 = ~n35713 & n35723 ;
  assign n35725 = ~n3564 & n20521 ;
  assign n35726 = ~n3282 & n20521 ;
  assign n35727 = ~n3560 & n35726 ;
  assign n35728 = ~n35725 & ~n35727 ;
  assign n35729 = ~n3567 & n35723 ;
  assign n35730 = ~n35728 & n35729 ;
  assign n35731 = ~n35724 & ~n35730 ;
  assign n35732 = ~n3567 & ~n35728 ;
  assign n35733 = \a[62]  & ~n35721 ;
  assign n35734 = ~n35719 & n35733 ;
  assign n35735 = n35713 & n35734 ;
  assign n35736 = ~n35732 & n35735 ;
  assign n35737 = n35731 & ~n35736 ;
  assign n35738 = ~\a[62]  & ~n35713 ;
  assign n35739 = ~\a[62]  & ~n3567 ;
  assign n35740 = ~n35728 & n35739 ;
  assign n35741 = ~n35738 & ~n35740 ;
  assign n35742 = ~n35719 & ~n35721 ;
  assign n35743 = \a[62]  & n35713 ;
  assign n35744 = ~n35732 & n35743 ;
  assign n35745 = ~n35742 & ~n35744 ;
  assign n35746 = n35741 & n35745 ;
  assign n35747 = n35737 & ~n35746 ;
  assign n35748 = ~n35703 & n35747 ;
  assign n35749 = n35703 & ~n35747 ;
  assign n35750 = ~n35748 & ~n35749 ;
  assign n35751 = n35701 & n35750 ;
  assign n35752 = ~n35701 & ~n35750 ;
  assign n35753 = ~n35751 & ~n35752 ;
  assign n35754 = n35679 & ~n35753 ;
  assign n35755 = ~n35679 & n35753 ;
  assign n35756 = ~n35754 & ~n35755 ;
  assign n35757 = ~n5459 & n16655 ;
  assign n35758 = ~n5104 & n16655 ;
  assign n35759 = ~n5455 & n35758 ;
  assign n35760 = ~n35757 & ~n35759 ;
  assign n35761 = ~n5462 & ~n35760 ;
  assign n35762 = \b[31]  & n16653 ;
  assign n35763 = \a[54]  & \b[30]  ;
  assign n35764 = n16644 & n35763 ;
  assign n35765 = ~\a[54]  & \b[30]  ;
  assign n35766 = n16647 & n35765 ;
  assign n35767 = ~n35764 & ~n35766 ;
  assign n35768 = ~n35762 & n35767 ;
  assign n35769 = \b[29]  & n17308 ;
  assign n35770 = n17305 & n35769 ;
  assign n35771 = \a[56]  & ~n35770 ;
  assign n35772 = n35768 & n35771 ;
  assign n35773 = ~n35761 & n35772 ;
  assign n35774 = n35768 & ~n35770 ;
  assign n35775 = ~\a[56]  & ~n35774 ;
  assign n35776 = ~\a[56]  & ~n5462 ;
  assign n35777 = ~n35760 & n35776 ;
  assign n35778 = ~n35775 & ~n35777 ;
  assign n35779 = ~n35773 & n35778 ;
  assign n35780 = n35756 & ~n35779 ;
  assign n35781 = ~n35756 & n35779 ;
  assign n35782 = ~n35780 & ~n35781 ;
  assign n35783 = ~n35676 & ~n35782 ;
  assign n35784 = n35676 & n35782 ;
  assign n35785 = ~n35783 & ~n35784 ;
  assign n35786 = n6565 & n14793 ;
  assign n35787 = ~n6562 & n35786 ;
  assign n35788 = n14793 & n22947 ;
  assign n35789 = ~n6561 & n35788 ;
  assign n35790 = \b[32]  & n15517 ;
  assign n35791 = n15514 & n35790 ;
  assign n35792 = ~\a[51]  & \b[33]  ;
  assign n35793 = n14785 & n35792 ;
  assign n35794 = ~n35791 & ~n35793 ;
  assign n35795 = \b[34]  & n14791 ;
  assign n35796 = \a[51]  & \b[33]  ;
  assign n35797 = n14782 & n35796 ;
  assign n35798 = \a[53]  & ~n35797 ;
  assign n35799 = ~n35795 & n35798 ;
  assign n35800 = n35794 & n35799 ;
  assign n35801 = ~n35789 & n35800 ;
  assign n35802 = ~n35787 & n35801 ;
  assign n35803 = ~n35795 & ~n35797 ;
  assign n35804 = n35794 & n35803 ;
  assign n35805 = ~n35789 & n35804 ;
  assign n35806 = ~n35787 & n35805 ;
  assign n35807 = ~\a[53]  & ~n35806 ;
  assign n35808 = ~n35802 & ~n35807 ;
  assign n35809 = ~n35785 & n35808 ;
  assign n35810 = n35785 & ~n35808 ;
  assign n35811 = ~n35809 & ~n35810 ;
  assign n35812 = ~n35104 & ~n35254 ;
  assign n35813 = n35108 & ~n35812 ;
  assign n35814 = ~n7761 & n13125 ;
  assign n35815 = ~n7759 & n35814 ;
  assign n35816 = \b[35]  & n13794 ;
  assign n35817 = n13792 & n35816 ;
  assign n35818 = ~\a[48]  & \b[36]  ;
  assign n35819 = n13117 & n35818 ;
  assign n35820 = ~n35817 & ~n35819 ;
  assign n35821 = \b[37]  & n13123 ;
  assign n35822 = \a[48]  & \b[36]  ;
  assign n35823 = n13786 & n35822 ;
  assign n35824 = \a[50]  & ~n35823 ;
  assign n35825 = ~n35821 & n35824 ;
  assign n35826 = n35820 & n35825 ;
  assign n35827 = ~n35815 & n35826 ;
  assign n35828 = ~n35821 & ~n35823 ;
  assign n35829 = n35820 & n35828 ;
  assign n35830 = ~n35815 & n35829 ;
  assign n35831 = ~\a[50]  & ~n35830 ;
  assign n35832 = ~n35827 & ~n35831 ;
  assign n35833 = ~n35813 & n35832 ;
  assign n35834 = ~n35811 & n35833 ;
  assign n35835 = n35813 & n35832 ;
  assign n35836 = n35811 & n35835 ;
  assign n35837 = ~n35834 & ~n35836 ;
  assign n35838 = ~n35813 & ~n35832 ;
  assign n35839 = n35811 & n35838 ;
  assign n35840 = n35813 & ~n35832 ;
  assign n35841 = ~n35811 & n35840 ;
  assign n35842 = ~n35839 & ~n35841 ;
  assign n35843 = n35837 & n35842 ;
  assign n35844 = n35674 & n35843 ;
  assign n35845 = ~n35674 & ~n35843 ;
  assign n35846 = ~n35844 & ~n35845 ;
  assign n35847 = ~n35672 & n35846 ;
  assign n35848 = n35672 & ~n35846 ;
  assign n35849 = ~n35847 & ~n35848 ;
  assign n35850 = ~n35293 & n35297 ;
  assign n35851 = ~n35294 & ~n35850 ;
  assign n35852 = n10082 & ~n10409 ;
  assign n35853 = ~n10407 & n35852 ;
  assign n35854 = \b[43]  & n10080 ;
  assign n35855 = \a[41]  & \b[42]  ;
  assign n35856 = n10679 & n35855 ;
  assign n35857 = ~\a[42]  & \b[42]  ;
  assign n35858 = n10074 & n35857 ;
  assign n35859 = ~n35856 & ~n35858 ;
  assign n35860 = ~n35854 & n35859 ;
  assign n35861 = \b[41]  & n10681 ;
  assign n35862 = n10678 & n35861 ;
  assign n35863 = \a[44]  & ~n35862 ;
  assign n35864 = n35860 & n35863 ;
  assign n35865 = ~n35853 & n35864 ;
  assign n35866 = n35860 & ~n35862 ;
  assign n35867 = ~n35853 & n35866 ;
  assign n35868 = ~\a[44]  & ~n35867 ;
  assign n35869 = ~n35865 & ~n35868 ;
  assign n35870 = n35851 & ~n35869 ;
  assign n35871 = ~n35849 & n35870 ;
  assign n35872 = ~n35851 & ~n35869 ;
  assign n35873 = n35849 & n35872 ;
  assign n35874 = ~n35871 & ~n35873 ;
  assign n35875 = ~n35851 & n35869 ;
  assign n35876 = ~n35849 & n35875 ;
  assign n35877 = n35851 & n35869 ;
  assign n35878 = n35849 & n35877 ;
  assign n35879 = ~n35876 & ~n35878 ;
  assign n35880 = n35874 & n35879 ;
  assign n35881 = n35324 & ~n35334 ;
  assign n35882 = n35329 & ~n35881 ;
  assign n35883 = n8759 & n11906 ;
  assign n35884 = ~n11903 & n35883 ;
  assign n35885 = n8759 & n13483 ;
  assign n35886 = ~n11902 & n35885 ;
  assign n35887 = \b[44]  & n9301 ;
  assign n35888 = n9298 & n35887 ;
  assign n35889 = ~\a[39]  & \b[45]  ;
  assign n35890 = n8751 & n35889 ;
  assign n35891 = ~n35888 & ~n35890 ;
  assign n35892 = \b[46]  & n8757 ;
  assign n35893 = \a[39]  & \b[45]  ;
  assign n35894 = n8748 & n35893 ;
  assign n35895 = \a[41]  & ~n35894 ;
  assign n35896 = ~n35892 & n35895 ;
  assign n35897 = n35891 & n35896 ;
  assign n35898 = ~n35886 & n35897 ;
  assign n35899 = ~n35884 & n35898 ;
  assign n35900 = ~n35892 & ~n35894 ;
  assign n35901 = n35891 & n35900 ;
  assign n35902 = ~n35886 & n35901 ;
  assign n35903 = ~n35884 & n35902 ;
  assign n35904 = ~\a[41]  & ~n35903 ;
  assign n35905 = ~n35899 & ~n35904 ;
  assign n35906 = ~n35882 & n35905 ;
  assign n35907 = ~n35880 & n35906 ;
  assign n35908 = n35882 & n35905 ;
  assign n35909 = n35880 & n35908 ;
  assign n35910 = ~n35907 & ~n35909 ;
  assign n35911 = n35882 & ~n35905 ;
  assign n35912 = ~n35880 & n35911 ;
  assign n35913 = ~n35882 & ~n35905 ;
  assign n35914 = n35880 & n35913 ;
  assign n35915 = ~n35912 & ~n35914 ;
  assign n35916 = n35910 & n35915 ;
  assign n35917 = n35358 & ~n35367 ;
  assign n35918 = n35363 & ~n35917 ;
  assign n35919 = n7534 & ~n13524 ;
  assign n35920 = ~n13522 & n35919 ;
  assign n35921 = \b[47]  & n7973 ;
  assign n35922 = n7970 & n35921 ;
  assign n35923 = ~\a[36]  & \b[48]  ;
  assign n35924 = n7526 & n35923 ;
  assign n35925 = ~n35922 & ~n35924 ;
  assign n35926 = \b[49]  & n7532 ;
  assign n35927 = \a[36]  & \b[48]  ;
  assign n35928 = n17801 & n35927 ;
  assign n35929 = \a[38]  & ~n35928 ;
  assign n35930 = ~n35926 & n35929 ;
  assign n35931 = n35925 & n35930 ;
  assign n35932 = ~n35920 & n35931 ;
  assign n35933 = ~n35926 & ~n35928 ;
  assign n35934 = n35925 & n35933 ;
  assign n35935 = ~n35920 & n35934 ;
  assign n35936 = ~\a[38]  & ~n35935 ;
  assign n35937 = ~n35932 & ~n35936 ;
  assign n35938 = n35918 & ~n35937 ;
  assign n35939 = ~n35916 & n35938 ;
  assign n35940 = ~n35918 & ~n35937 ;
  assign n35941 = n35916 & n35940 ;
  assign n35942 = ~n35939 & ~n35941 ;
  assign n35943 = ~n35918 & n35937 ;
  assign n35944 = ~n35916 & n35943 ;
  assign n35945 = n35918 & n35937 ;
  assign n35946 = n35916 & n35945 ;
  assign n35947 = ~n35944 & ~n35946 ;
  assign n35948 = n35942 & n35947 ;
  assign n35949 = ~n35649 & ~n35948 ;
  assign n35950 = n35649 & n35948 ;
  assign n35951 = ~n35949 & ~n35950 ;
  assign n35952 = n6309 & n15201 ;
  assign n35953 = ~n15198 & n35952 ;
  assign n35954 = n6309 & ~n15201 ;
  assign n35955 = ~n14093 & n35954 ;
  assign n35956 = ~n15197 & n35955 ;
  assign n35957 = \b[50]  & n6778 ;
  assign n35958 = n6775 & n35957 ;
  assign n35959 = ~\a[33]  & \b[51]  ;
  assign n35960 = n6301 & n35959 ;
  assign n35961 = ~n35958 & ~n35960 ;
  assign n35962 = \b[52]  & n6307 ;
  assign n35963 = \a[33]  & \b[51]  ;
  assign n35964 = n6298 & n35963 ;
  assign n35965 = \a[35]  & ~n35964 ;
  assign n35966 = ~n35962 & n35965 ;
  assign n35967 = n35961 & n35966 ;
  assign n35968 = ~n35956 & n35967 ;
  assign n35969 = ~n35953 & n35968 ;
  assign n35970 = ~n35962 & ~n35964 ;
  assign n35971 = n35961 & n35970 ;
  assign n35972 = ~n35956 & n35971 ;
  assign n35973 = ~n35953 & n35972 ;
  assign n35974 = ~\a[35]  & ~n35973 ;
  assign n35975 = ~n35969 & ~n35974 ;
  assign n35976 = ~n35951 & n35975 ;
  assign n35977 = n35951 & ~n35975 ;
  assign n35978 = ~n35976 & ~n35977 ;
  assign n35979 = n35647 & n35978 ;
  assign n35980 = ~n35647 & ~n35978 ;
  assign n35981 = ~n35979 & ~n35980 ;
  assign n35982 = ~n35621 & n35981 ;
  assign n35983 = ~n35620 & n35982 ;
  assign n35984 = n35621 & ~n35981 ;
  assign n35985 = n35620 & ~n35981 ;
  assign n35986 = ~n35984 & ~n35985 ;
  assign n35987 = ~n35983 & n35986 ;
  assign n35988 = n35580 & n35987 ;
  assign n35989 = ~n35580 & ~n35987 ;
  assign n35990 = ~n35988 & ~n35989 ;
  assign n35991 = ~n35557 & n35990 ;
  assign n35992 = n35557 & ~n35990 ;
  assign n35993 = ~n35991 & ~n35992 ;
  assign n35994 = ~n35529 & n35993 ;
  assign n35995 = n35529 & ~n35993 ;
  assign n35996 = ~n35994 & ~n35995 ;
  assign n35997 = n35521 & n35996 ;
  assign n35998 = ~n35521 & ~n35996 ;
  assign n35999 = ~n35997 & ~n35998 ;
  assign n36000 = ~n35524 & n35999 ;
  assign n36001 = ~n35996 & ~n35997 ;
  assign n36002 = n35524 & n36001 ;
  assign n36003 = ~n36000 & ~n36002 ;
  assign n36004 = n35524 & n35996 ;
  assign n36005 = ~n35995 & ~n35997 ;
  assign n36006 = ~n36004 & n36005 ;
  assign n36007 = ~n35579 & ~n35987 ;
  assign n36008 = n35046 & n35576 ;
  assign n36009 = n35558 & n35576 ;
  assign n36010 = ~n36008 & ~n36009 ;
  assign n36011 = \b[63]  & n2622 ;
  assign n36012 = ~n21694 & n36011 ;
  assign n36013 = ~n23171 & n36012 ;
  assign n36014 = \a[20]  & \a[22]  ;
  assign n36015 = \a[21]  & ~\a[23]  ;
  assign n36016 = n36014 & n36015 ;
  assign n36017 = ~\a[20]  & ~\a[22]  ;
  assign n36018 = ~\a[21]  & \a[23]  ;
  assign n36019 = n36017 & n36018 ;
  assign n36020 = ~n36016 & ~n36019 ;
  assign n36021 = \b[63]  & ~n36020 ;
  assign n36022 = \a[23]  & ~n36021 ;
  assign n36023 = ~n36013 & n36022 ;
  assign n36024 = ~n36013 & ~n36021 ;
  assign n36025 = ~\a[23]  & ~n36024 ;
  assign n36026 = ~n36023 & ~n36025 ;
  assign n36027 = n36010 & ~n36026 ;
  assign n36028 = ~n36007 & n36027 ;
  assign n36029 = ~n36010 & n36026 ;
  assign n36030 = ~n35579 & n36026 ;
  assign n36031 = ~n35987 & n36030 ;
  assign n36032 = ~n36029 & ~n36031 ;
  assign n36033 = ~n36028 & n36032 ;
  assign n36034 = n3402 & n21696 ;
  assign n36035 = ~n21693 & n36034 ;
  assign n36036 = n3402 & ~n21696 ;
  assign n36037 = ~n20966 & n36036 ;
  assign n36038 = ~n21692 & n36037 ;
  assign n36039 = \b[62]  & n3400 ;
  assign n36040 = \a[24]  & \b[61]  ;
  assign n36041 = n27626 & n36040 ;
  assign n36042 = ~n36039 & ~n36041 ;
  assign n36043 = \b[60]  & n3733 ;
  assign n36044 = n3730 & n36043 ;
  assign n36045 = ~\a[24]  & \b[61]  ;
  assign n36046 = n3394 & n36045 ;
  assign n36047 = ~n36044 & ~n36046 ;
  assign n36048 = n36042 & n36047 ;
  assign n36049 = ~n36038 & n36048 ;
  assign n36050 = ~n36035 & n36049 ;
  assign n36051 = ~\a[26]  & ~n36050 ;
  assign n36052 = \a[26]  & ~n36041 ;
  assign n36053 = ~n36039 & n36052 ;
  assign n36054 = n36047 & n36053 ;
  assign n36055 = ~n36038 & n36054 ;
  assign n36056 = ~n36035 & n36055 ;
  assign n36057 = ~n36051 & ~n36056 ;
  assign n36058 = ~n35621 & n36057 ;
  assign n36059 = ~n35983 & n36058 ;
  assign n36060 = ~n35621 & ~n35981 ;
  assign n36061 = n35620 & ~n35621 ;
  assign n36062 = ~n36060 & ~n36061 ;
  assign n36063 = \a[26]  & ~n36050 ;
  assign n36064 = ~\a[26]  & n36050 ;
  assign n36065 = ~n36063 & ~n36064 ;
  assign n36066 = n36062 & n36065 ;
  assign n36067 = ~n36059 & ~n36066 ;
  assign n36068 = ~n35640 & ~n35978 ;
  assign n36069 = ~n35640 & n35646 ;
  assign n36070 = ~n36068 & ~n36069 ;
  assign n36071 = n4249 & ~n19550 ;
  assign n36072 = ~n19548 & n36071 ;
  assign n36073 = \b[59]  & n4247 ;
  assign n36074 = \a[27]  & \b[58]  ;
  assign n36075 = n4238 & n36074 ;
  assign n36076 = ~n36073 & ~n36075 ;
  assign n36077 = \b[57]  & n4647 ;
  assign n36078 = n4644 & n36077 ;
  assign n36079 = ~\a[27]  & \b[58]  ;
  assign n36080 = n4241 & n36079 ;
  assign n36081 = ~n36078 & ~n36080 ;
  assign n36082 = n36076 & n36081 ;
  assign n36083 = ~n36072 & n36082 ;
  assign n36084 = \a[29]  & ~n36083 ;
  assign n36085 = ~\a[29]  & n36083 ;
  assign n36086 = ~n36084 & ~n36085 ;
  assign n36087 = n36070 & n36086 ;
  assign n36088 = ~\a[29]  & ~n36083 ;
  assign n36089 = \a[29]  & n36082 ;
  assign n36090 = ~n36072 & n36089 ;
  assign n36091 = ~n35640 & ~n36090 ;
  assign n36092 = ~n35978 & n36091 ;
  assign n36093 = n35646 & n36091 ;
  assign n36094 = ~n36092 & ~n36093 ;
  assign n36095 = ~n36088 & ~n36094 ;
  assign n36096 = ~n36087 & ~n36095 ;
  assign n36097 = ~n35950 & n35975 ;
  assign n36098 = ~n35949 & ~n36097 ;
  assign n36099 = n5211 & n17647 ;
  assign n36100 = ~n17644 & n36099 ;
  assign n36101 = n5211 & ~n17647 ;
  assign n36102 = ~n16441 & n36101 ;
  assign n36103 = ~n17643 & n36102 ;
  assign n36104 = \b[56]  & n5209 ;
  assign n36105 = \a[30]  & \b[55]  ;
  assign n36106 = n5200 & n36105 ;
  assign n36107 = ~n36104 & ~n36106 ;
  assign n36108 = \b[54]  & n5595 ;
  assign n36109 = n5592 & n36108 ;
  assign n36110 = ~\a[30]  & \b[55]  ;
  assign n36111 = n5203 & n36110 ;
  assign n36112 = ~n36109 & ~n36111 ;
  assign n36113 = n36107 & n36112 ;
  assign n36114 = ~n36103 & n36113 ;
  assign n36115 = ~n36100 & n36114 ;
  assign n36116 = ~\a[32]  & ~n36115 ;
  assign n36117 = \a[32]  & ~n36106 ;
  assign n36118 = ~n36104 & n36117 ;
  assign n36119 = n36112 & n36118 ;
  assign n36120 = ~n36103 & n36119 ;
  assign n36121 = ~n36100 & n36120 ;
  assign n36122 = ~n36116 & ~n36121 ;
  assign n36123 = ~n36098 & n36122 ;
  assign n36124 = \a[32]  & ~n36115 ;
  assign n36125 = ~\a[32]  & n36115 ;
  assign n36126 = ~n36124 & ~n36125 ;
  assign n36127 = ~n35949 & n36126 ;
  assign n36128 = ~n36097 & n36127 ;
  assign n36129 = ~n36123 & ~n36128 ;
  assign n36130 = ~n9479 & n11572 ;
  assign n36131 = ~n9043 & n11572 ;
  assign n36132 = ~n9475 & n36131 ;
  assign n36133 = ~n36130 & ~n36132 ;
  assign n36134 = ~n9482 & ~n36133 ;
  assign n36135 = \b[39]  & n12159 ;
  assign n36136 = n12156 & n36135 ;
  assign n36137 = ~\a[45]  & \b[40]  ;
  assign n36138 = n11564 & n36137 ;
  assign n36139 = ~n36136 & ~n36138 ;
  assign n36140 = \b[41]  & n11570 ;
  assign n36141 = \a[45]  & \b[40]  ;
  assign n36142 = n11561 & n36141 ;
  assign n36143 = \a[47]  & ~n36142 ;
  assign n36144 = ~n36140 & n36143 ;
  assign n36145 = n36139 & n36144 ;
  assign n36146 = ~n36134 & n36145 ;
  assign n36147 = ~n36140 & ~n36142 ;
  assign n36148 = n36139 & n36147 ;
  assign n36149 = ~\a[47]  & ~n36148 ;
  assign n36150 = ~\a[47]  & ~n9482 ;
  assign n36151 = ~n36133 & n36150 ;
  assign n36152 = ~n36149 & ~n36151 ;
  assign n36153 = ~n36146 & n36152 ;
  assign n36154 = ~n35811 & ~n35813 ;
  assign n36155 = n35811 & n35813 ;
  assign n36156 = n35832 & ~n36155 ;
  assign n36157 = ~n36154 & ~n36156 ;
  assign n36158 = ~n6610 & n14793 ;
  assign n36159 = ~n6608 & n36158 ;
  assign n36160 = \b[33]  & n15517 ;
  assign n36161 = n15514 & n36160 ;
  assign n36162 = ~\a[51]  & \b[34]  ;
  assign n36163 = n14785 & n36162 ;
  assign n36164 = ~n36161 & ~n36163 ;
  assign n36165 = \b[35]  & n14791 ;
  assign n36166 = \a[51]  & \b[34]  ;
  assign n36167 = n14782 & n36166 ;
  assign n36168 = \a[53]  & ~n36167 ;
  assign n36169 = ~n36165 & n36168 ;
  assign n36170 = n36164 & n36169 ;
  assign n36171 = ~n36159 & n36170 ;
  assign n36172 = ~n36165 & ~n36167 ;
  assign n36173 = n36164 & n36172 ;
  assign n36174 = ~n36159 & n36173 ;
  assign n36175 = ~\a[53]  & ~n36174 ;
  assign n36176 = ~n36171 & ~n36175 ;
  assign n36177 = n35701 & ~n35748 ;
  assign n36178 = ~n35749 & ~n36177 ;
  assign n36179 = ~n4499 & n18516 ;
  assign n36180 = ~n4455 & n18516 ;
  assign n36181 = ~n4495 & n36180 ;
  assign n36182 = ~n36179 & ~n36181 ;
  assign n36183 = ~n4502 & ~n36182 ;
  assign n36184 = \b[29]  & n18514 ;
  assign n36185 = \a[56]  & \b[28]  ;
  assign n36186 = n19181 & n36185 ;
  assign n36187 = ~\a[57]  & \b[28]  ;
  assign n36188 = n18508 & n36187 ;
  assign n36189 = ~n36186 & ~n36188 ;
  assign n36190 = ~n36184 & n36189 ;
  assign n36191 = \b[27]  & n19183 ;
  assign n36192 = n19180 & n36191 ;
  assign n36193 = \a[59]  & ~n36192 ;
  assign n36194 = n36190 & n36193 ;
  assign n36195 = ~n36183 & n36194 ;
  assign n36196 = n36190 & ~n36192 ;
  assign n36197 = ~\a[59]  & ~n36196 ;
  assign n36198 = ~\a[59]  & ~n4502 ;
  assign n36199 = ~n36182 & n36198 ;
  assign n36200 = ~n36197 & ~n36199 ;
  assign n36201 = ~n36195 & n36200 ;
  assign n36202 = ~n35719 & n35737 ;
  assign n36203 = n3604 & n20521 ;
  assign n36204 = ~n19292 & n36203 ;
  assign n36205 = n12021 & n20521 ;
  assign n36206 = ~n3600 & n36205 ;
  assign n36207 = \b[26]  & n20519 ;
  assign n36208 = \a[60]  & \b[25]  ;
  assign n36209 = n20510 & n36208 ;
  assign n36210 = ~n36207 & ~n36209 ;
  assign n36211 = \b[24]  & n21315 ;
  assign n36212 = n21312 & n36211 ;
  assign n36213 = ~\a[60]  & \b[25]  ;
  assign n36214 = n20513 & n36213 ;
  assign n36215 = ~n36212 & ~n36214 ;
  assign n36216 = n36210 & n36215 ;
  assign n36217 = ~n36206 & n36216 ;
  assign n36218 = ~n36204 & n36217 ;
  assign n36219 = \b[23]  & n21958 ;
  assign n36220 = \b[22]  & n21957 ;
  assign n36221 = ~n36219 & ~n36220 ;
  assign n36222 = ~n35718 & n36221 ;
  assign n36223 = n35718 & ~n36221 ;
  assign n36224 = ~n36222 & ~n36223 ;
  assign n36225 = ~\a[62]  & n36224 ;
  assign n36226 = ~n36218 & n36225 ;
  assign n36227 = \a[62]  & n36224 ;
  assign n36228 = n36216 & n36227 ;
  assign n36229 = ~n36206 & n36228 ;
  assign n36230 = ~n36204 & n36229 ;
  assign n36231 = ~n36226 & ~n36230 ;
  assign n36232 = ~\a[62]  & ~n36218 ;
  assign n36233 = \a[62]  & n36216 ;
  assign n36234 = ~n36206 & n36233 ;
  assign n36235 = ~n36204 & n36234 ;
  assign n36236 = ~n36224 & ~n36235 ;
  assign n36237 = ~n36232 & n36236 ;
  assign n36238 = n36231 & ~n36237 ;
  assign n36239 = ~n36202 & n36238 ;
  assign n36240 = n36202 & ~n36238 ;
  assign n36241 = ~n36239 & ~n36240 ;
  assign n36242 = ~n36201 & n36241 ;
  assign n36243 = ~n36178 & n36242 ;
  assign n36244 = n36201 & ~n36241 ;
  assign n36245 = ~n36178 & n36244 ;
  assign n36246 = ~n36243 & ~n36245 ;
  assign n36247 = n36178 & ~n36244 ;
  assign n36248 = ~n36242 & n36247 ;
  assign n36249 = n36246 & ~n36248 ;
  assign n36250 = ~n5810 & ~n16016 ;
  assign n36251 = ~n16652 & n36250 ;
  assign n36252 = n5807 & n36251 ;
  assign n36253 = n5810 & ~n16016 ;
  assign n36254 = ~n16652 & n36253 ;
  assign n36255 = ~n5807 & n36254 ;
  assign n36256 = ~n36252 & ~n36255 ;
  assign n36257 = \b[32]  & n16653 ;
  assign n36258 = \a[54]  & \b[31]  ;
  assign n36259 = n16644 & n36258 ;
  assign n36260 = ~\a[54]  & \b[31]  ;
  assign n36261 = n16647 & n36260 ;
  assign n36262 = ~n36259 & ~n36261 ;
  assign n36263 = ~n36257 & n36262 ;
  assign n36264 = \b[30]  & n17308 ;
  assign n36265 = n17305 & n36264 ;
  assign n36266 = \a[56]  & ~n36265 ;
  assign n36267 = n36263 & n36266 ;
  assign n36268 = n36256 & n36267 ;
  assign n36269 = n36263 & ~n36265 ;
  assign n36270 = n36256 & n36269 ;
  assign n36271 = ~\a[56]  & ~n36270 ;
  assign n36272 = ~n36268 & ~n36271 ;
  assign n36273 = ~n36249 & ~n36272 ;
  assign n36274 = n36249 & n36272 ;
  assign n36275 = ~n36273 & ~n36274 ;
  assign n36276 = ~n35754 & n35779 ;
  assign n36277 = ~n35755 & ~n36276 ;
  assign n36278 = ~n36275 & n36277 ;
  assign n36279 = n36275 & ~n36277 ;
  assign n36280 = ~n36278 & ~n36279 ;
  assign n36281 = n36176 & n36280 ;
  assign n36282 = ~n36176 & ~n36280 ;
  assign n36283 = ~n36281 & ~n36282 ;
  assign n36284 = ~n35784 & n35808 ;
  assign n36285 = ~n35783 & ~n36284 ;
  assign n36286 = n8175 & n13125 ;
  assign n36287 = ~n8172 & n36286 ;
  assign n36288 = ~n8175 & n13125 ;
  assign n36289 = ~n7756 & n36288 ;
  assign n36290 = ~n8171 & n36289 ;
  assign n36291 = \b[36]  & n13794 ;
  assign n36292 = n13792 & n36291 ;
  assign n36293 = ~\a[48]  & \b[37]  ;
  assign n36294 = n13117 & n36293 ;
  assign n36295 = ~n36292 & ~n36294 ;
  assign n36296 = \b[38]  & n13123 ;
  assign n36297 = \a[48]  & \b[37]  ;
  assign n36298 = n13786 & n36297 ;
  assign n36299 = \a[50]  & ~n36298 ;
  assign n36300 = ~n36296 & n36299 ;
  assign n36301 = n36295 & n36300 ;
  assign n36302 = ~n36290 & n36301 ;
  assign n36303 = ~n36287 & n36302 ;
  assign n36304 = ~n36296 & ~n36298 ;
  assign n36305 = n36295 & n36304 ;
  assign n36306 = ~n36290 & n36305 ;
  assign n36307 = ~n36287 & n36306 ;
  assign n36308 = ~\a[50]  & ~n36307 ;
  assign n36309 = ~n36303 & ~n36308 ;
  assign n36310 = ~n36285 & ~n36309 ;
  assign n36311 = ~n36283 & n36310 ;
  assign n36312 = n36285 & ~n36309 ;
  assign n36313 = n36283 & n36312 ;
  assign n36314 = ~n36311 & ~n36313 ;
  assign n36315 = ~n36285 & n36309 ;
  assign n36316 = n36283 & n36315 ;
  assign n36317 = n36285 & n36309 ;
  assign n36318 = ~n36283 & n36317 ;
  assign n36319 = ~n36316 & ~n36318 ;
  assign n36320 = n36314 & n36319 ;
  assign n36321 = n36157 & n36320 ;
  assign n36322 = ~n36157 & ~n36320 ;
  assign n36323 = ~n36321 & ~n36322 ;
  assign n36324 = n36153 & n36323 ;
  assign n36325 = ~n36153 & ~n36323 ;
  assign n36326 = ~n36324 & ~n36325 ;
  assign n36327 = n10082 & ~n28007 ;
  assign n36328 = ~n28005 & n36327 ;
  assign n36329 = \b[42]  & n10681 ;
  assign n36330 = n10678 & n36329 ;
  assign n36331 = \b[44]  & n10080 ;
  assign n36332 = \a[41]  & \b[43]  ;
  assign n36333 = n10679 & n36332 ;
  assign n36334 = ~\a[42]  & \b[43]  ;
  assign n36335 = n10074 & n36334 ;
  assign n36336 = ~n36333 & ~n36335 ;
  assign n36337 = ~n36331 & n36336 ;
  assign n36338 = ~n36330 & n36337 ;
  assign n36339 = ~n36328 & n36338 ;
  assign n36340 = ~\a[44]  & ~n36339 ;
  assign n36341 = \a[44]  & n36338 ;
  assign n36342 = ~n36328 & n36341 ;
  assign n36343 = ~n36340 & ~n36342 ;
  assign n36344 = n35672 & ~n35844 ;
  assign n36345 = ~n35844 & n35845 ;
  assign n36346 = ~n36344 & ~n36345 ;
  assign n36347 = ~n36343 & ~n36346 ;
  assign n36348 = ~n36326 & n36347 ;
  assign n36349 = ~n36343 & n36346 ;
  assign n36350 = n36326 & n36349 ;
  assign n36351 = ~n36348 & ~n36350 ;
  assign n36352 = n36343 & n36346 ;
  assign n36353 = ~n36326 & n36352 ;
  assign n36354 = n36343 & ~n36346 ;
  assign n36355 = n36326 & n36354 ;
  assign n36356 = ~n36353 & ~n36355 ;
  assign n36357 = n36351 & n36356 ;
  assign n36358 = ~n35849 & ~n35851 ;
  assign n36359 = n35849 & n35851 ;
  assign n36360 = n35869 & ~n36359 ;
  assign n36361 = ~n36358 & ~n36360 ;
  assign n36362 = n36357 & n36361 ;
  assign n36363 = ~n36357 & ~n36361 ;
  assign n36364 = ~n36362 & ~n36363 ;
  assign n36365 = n8759 & ~n12438 ;
  assign n36366 = ~n12436 & n36365 ;
  assign n36367 = \b[45]  & n9301 ;
  assign n36368 = n9298 & n36367 ;
  assign n36369 = ~\a[39]  & \b[46]  ;
  assign n36370 = n8751 & n36369 ;
  assign n36371 = ~n36368 & ~n36370 ;
  assign n36372 = \b[47]  & n8757 ;
  assign n36373 = \a[39]  & \b[46]  ;
  assign n36374 = n8748 & n36373 ;
  assign n36375 = \a[41]  & ~n36374 ;
  assign n36376 = ~n36372 & n36375 ;
  assign n36377 = n36371 & n36376 ;
  assign n36378 = ~n36366 & n36377 ;
  assign n36379 = ~n36372 & ~n36374 ;
  assign n36380 = n36371 & n36379 ;
  assign n36381 = ~n36366 & n36380 ;
  assign n36382 = ~\a[41]  & ~n36381 ;
  assign n36383 = ~n36378 & ~n36382 ;
  assign n36384 = n36364 & ~n36383 ;
  assign n36385 = ~n36364 & n36383 ;
  assign n36386 = ~n36384 & ~n36385 ;
  assign n36387 = ~n35880 & ~n35882 ;
  assign n36388 = n35880 & n35882 ;
  assign n36389 = n35905 & ~n36388 ;
  assign n36390 = ~n36387 & ~n36389 ;
  assign n36391 = n7534 & n14052 ;
  assign n36392 = ~n14049 & n36391 ;
  assign n36393 = n7534 & ~n14052 ;
  assign n36394 = ~n13519 & n36393 ;
  assign n36395 = ~n14048 & n36394 ;
  assign n36396 = \b[48]  & n7973 ;
  assign n36397 = n7970 & n36396 ;
  assign n36398 = ~\a[36]  & \b[49]  ;
  assign n36399 = n7526 & n36398 ;
  assign n36400 = ~n36397 & ~n36399 ;
  assign n36401 = \b[50]  & n7532 ;
  assign n36402 = \a[36]  & \b[49]  ;
  assign n36403 = n17801 & n36402 ;
  assign n36404 = \a[38]  & ~n36403 ;
  assign n36405 = ~n36401 & n36404 ;
  assign n36406 = n36400 & n36405 ;
  assign n36407 = ~n36395 & n36406 ;
  assign n36408 = ~n36392 & n36407 ;
  assign n36409 = ~n36401 & ~n36403 ;
  assign n36410 = n36400 & n36409 ;
  assign n36411 = ~n36395 & n36410 ;
  assign n36412 = ~n36392 & n36411 ;
  assign n36413 = ~\a[38]  & ~n36412 ;
  assign n36414 = ~n36408 & ~n36413 ;
  assign n36415 = ~n36390 & n36414 ;
  assign n36416 = ~n36386 & n36415 ;
  assign n36417 = n36390 & n36414 ;
  assign n36418 = n36386 & n36417 ;
  assign n36419 = ~n36416 & ~n36418 ;
  assign n36420 = ~n36390 & ~n36414 ;
  assign n36421 = n36386 & n36420 ;
  assign n36422 = n36390 & ~n36414 ;
  assign n36423 = ~n36386 & n36422 ;
  assign n36424 = ~n36421 & ~n36423 ;
  assign n36425 = n36419 & n36424 ;
  assign n36426 = n6309 & ~n15246 ;
  assign n36427 = ~n15244 & n36426 ;
  assign n36428 = \b[51]  & n6778 ;
  assign n36429 = n6775 & n36428 ;
  assign n36430 = ~\a[33]  & \b[52]  ;
  assign n36431 = n6301 & n36430 ;
  assign n36432 = ~n36429 & ~n36431 ;
  assign n36433 = \b[53]  & n6307 ;
  assign n36434 = \a[33]  & \b[52]  ;
  assign n36435 = n6298 & n36434 ;
  assign n36436 = \a[35]  & ~n36435 ;
  assign n36437 = ~n36433 & n36436 ;
  assign n36438 = n36432 & n36437 ;
  assign n36439 = ~n36427 & n36438 ;
  assign n36440 = ~n36433 & ~n36435 ;
  assign n36441 = n36432 & n36440 ;
  assign n36442 = ~n36427 & n36441 ;
  assign n36443 = ~\a[35]  & ~n36442 ;
  assign n36444 = ~n36439 & ~n36443 ;
  assign n36445 = ~n35916 & ~n35918 ;
  assign n36446 = n35916 & n35918 ;
  assign n36447 = n35937 & ~n36446 ;
  assign n36448 = ~n36445 & ~n36447 ;
  assign n36449 = n36444 & ~n36448 ;
  assign n36450 = n36425 & n36449 ;
  assign n36451 = n36444 & n36448 ;
  assign n36452 = ~n36425 & n36451 ;
  assign n36453 = ~n36450 & ~n36452 ;
  assign n36454 = ~n36444 & ~n36448 ;
  assign n36455 = ~n36425 & n36454 ;
  assign n36456 = ~n36444 & n36448 ;
  assign n36457 = n36425 & n36456 ;
  assign n36458 = ~n36455 & ~n36457 ;
  assign n36459 = n36453 & n36458 ;
  assign n36460 = n36129 & ~n36459 ;
  assign n36461 = ~n36129 & n36459 ;
  assign n36462 = ~n36460 & ~n36461 ;
  assign n36463 = n36096 & n36462 ;
  assign n36464 = ~n36096 & ~n36462 ;
  assign n36465 = ~n36463 & ~n36464 ;
  assign n36466 = n36067 & n36465 ;
  assign n36467 = ~n36067 & ~n36465 ;
  assign n36468 = ~n36466 & ~n36467 ;
  assign n36469 = n36033 & n36468 ;
  assign n36470 = ~n36033 & ~n36468 ;
  assign n36471 = ~n36469 & ~n36470 ;
  assign n36472 = ~n35555 & ~n35990 ;
  assign n36473 = ~n35556 & ~n36472 ;
  assign n36474 = n36471 & n36473 ;
  assign n36475 = ~n36471 & ~n36473 ;
  assign n36476 = ~n36474 & ~n36475 ;
  assign n36477 = n36006 & n36476 ;
  assign n36478 = ~n36006 & ~n36476 ;
  assign n36479 = ~n36477 & ~n36478 ;
  assign n36480 = ~n35995 & ~n36474 ;
  assign n36481 = ~n35997 & n36480 ;
  assign n36482 = ~n36004 & n36481 ;
  assign n36483 = ~n36028 & ~n36469 ;
  assign n36484 = ~n36066 & ~n36465 ;
  assign n36485 = n36059 & ~n36066 ;
  assign n36486 = ~n36484 & ~n36485 ;
  assign n36487 = n3402 & ~n22461 ;
  assign n36488 = ~n22459 & n36487 ;
  assign n36489 = \b[63]  & n3400 ;
  assign n36490 = \a[24]  & \b[62]  ;
  assign n36491 = n27626 & n36490 ;
  assign n36492 = ~n36489 & ~n36491 ;
  assign n36493 = \b[61]  & n3733 ;
  assign n36494 = n3730 & n36493 ;
  assign n36495 = ~\a[24]  & \b[62]  ;
  assign n36496 = n3394 & n36495 ;
  assign n36497 = ~n36494 & ~n36496 ;
  assign n36498 = n36492 & n36497 ;
  assign n36499 = ~n36488 & n36498 ;
  assign n36500 = ~\a[26]  & ~n36499 ;
  assign n36501 = \a[26]  & n36498 ;
  assign n36502 = ~n36488 & n36501 ;
  assign n36503 = ~n36500 & ~n36502 ;
  assign n36504 = n36486 & ~n36503 ;
  assign n36505 = ~n36486 & n36503 ;
  assign n36506 = ~n36504 & ~n36505 ;
  assign n36507 = ~n36087 & ~n36462 ;
  assign n36508 = ~n36087 & n36095 ;
  assign n36509 = ~n36507 & ~n36508 ;
  assign n36510 = n4249 & n20260 ;
  assign n36511 = ~n20257 & n36510 ;
  assign n36512 = n4249 & ~n20260 ;
  assign n36513 = ~n19545 & n36512 ;
  assign n36514 = ~n20256 & n36513 ;
  assign n36515 = \b[58]  & n4647 ;
  assign n36516 = n4644 & n36515 ;
  assign n36517 = ~\a[27]  & \b[59]  ;
  assign n36518 = n4241 & n36517 ;
  assign n36519 = ~n36516 & ~n36518 ;
  assign n36520 = \b[60]  & n4247 ;
  assign n36521 = \a[27]  & \b[59]  ;
  assign n36522 = n4238 & n36521 ;
  assign n36523 = \a[29]  & ~n36522 ;
  assign n36524 = ~n36520 & n36523 ;
  assign n36525 = n36519 & n36524 ;
  assign n36526 = ~n36514 & n36525 ;
  assign n36527 = ~n36511 & n36526 ;
  assign n36528 = ~n36520 & ~n36522 ;
  assign n36529 = n36519 & n36528 ;
  assign n36530 = ~n36514 & n36529 ;
  assign n36531 = ~n36511 & n36530 ;
  assign n36532 = ~\a[29]  & ~n36531 ;
  assign n36533 = ~n36527 & ~n36532 ;
  assign n36534 = n5211 & ~n17690 ;
  assign n36535 = ~n17688 & n36534 ;
  assign n36536 = \b[57]  & n5209 ;
  assign n36537 = \a[30]  & \b[56]  ;
  assign n36538 = n5200 & n36537 ;
  assign n36539 = ~n36536 & ~n36538 ;
  assign n36540 = \b[55]  & n5595 ;
  assign n36541 = n5592 & n36540 ;
  assign n36542 = ~\a[30]  & \b[56]  ;
  assign n36543 = n5203 & n36542 ;
  assign n36544 = ~n36541 & ~n36543 ;
  assign n36545 = n36539 & n36544 ;
  assign n36546 = ~n36535 & n36545 ;
  assign n36547 = ~\a[32]  & ~n36546 ;
  assign n36548 = \a[32]  & n36545 ;
  assign n36549 = ~n36535 & n36548 ;
  assign n36550 = ~n36547 & ~n36549 ;
  assign n36551 = n36123 & n36550 ;
  assign n36552 = ~n36128 & n36550 ;
  assign n36553 = n36459 & n36552 ;
  assign n36554 = ~n36551 & ~n36553 ;
  assign n36555 = ~n36128 & n36459 ;
  assign n36556 = ~n36123 & ~n36550 ;
  assign n36557 = ~n36555 & n36556 ;
  assign n36558 = n36554 & ~n36557 ;
  assign n36559 = n6309 & ~n16398 ;
  assign n36560 = ~n15241 & n36559 ;
  assign n36561 = ~n16404 & n36560 ;
  assign n36562 = n6309 & n16398 ;
  assign n36563 = n15241 & n36562 ;
  assign n36564 = n16400 & n36562 ;
  assign n36565 = ~n15239 & n36564 ;
  assign n36566 = ~n36563 & ~n36565 ;
  assign n36567 = ~n36561 & n36566 ;
  assign n36568 = \b[52]  & n6778 ;
  assign n36569 = n6775 & n36568 ;
  assign n36570 = ~\a[33]  & \b[53]  ;
  assign n36571 = n6301 & n36570 ;
  assign n36572 = ~n36569 & ~n36571 ;
  assign n36573 = \b[54]  & n6307 ;
  assign n36574 = \a[33]  & \b[53]  ;
  assign n36575 = n6298 & n36574 ;
  assign n36576 = \a[35]  & ~n36575 ;
  assign n36577 = ~n36573 & n36576 ;
  assign n36578 = n36572 & n36577 ;
  assign n36579 = n36567 & n36578 ;
  assign n36580 = ~n36573 & ~n36575 ;
  assign n36581 = n36572 & n36580 ;
  assign n36582 = n36567 & n36581 ;
  assign n36583 = ~\a[35]  & ~n36582 ;
  assign n36584 = ~n36579 & ~n36583 ;
  assign n36585 = n36386 & n36390 ;
  assign n36586 = n36424 & ~n36585 ;
  assign n36587 = ~n5105 & ~n17912 ;
  assign n36588 = ~n18513 & n36587 ;
  assign n36589 = n5102 & n36588 ;
  assign n36590 = n5105 & ~n17912 ;
  assign n36591 = ~n18513 & n36590 ;
  assign n36592 = ~n5102 & n36591 ;
  assign n36593 = ~n36589 & ~n36592 ;
  assign n36594 = \b[28]  & n19183 ;
  assign n36595 = n19180 & n36594 ;
  assign n36596 = \b[30]  & n18514 ;
  assign n36597 = \a[56]  & \b[29]  ;
  assign n36598 = n19181 & n36597 ;
  assign n36599 = ~\a[57]  & \b[29]  ;
  assign n36600 = n18508 & n36599 ;
  assign n36601 = ~n36598 & ~n36600 ;
  assign n36602 = ~n36596 & n36601 ;
  assign n36603 = ~n36595 & n36602 ;
  assign n36604 = n36593 & n36603 ;
  assign n36605 = ~\a[59]  & ~n36604 ;
  assign n36606 = \a[59]  & n36603 ;
  assign n36607 = n36593 & n36606 ;
  assign n36608 = ~n36605 & ~n36607 ;
  assign n36609 = ~n36222 & ~n36230 ;
  assign n36610 = ~n36226 & n36609 ;
  assign n36611 = ~n4148 & n20521 ;
  assign n36612 = ~n4146 & n36611 ;
  assign n36613 = \b[27]  & n20519 ;
  assign n36614 = \a[60]  & \b[26]  ;
  assign n36615 = n20510 & n36614 ;
  assign n36616 = ~n36613 & ~n36615 ;
  assign n36617 = \b[25]  & n21315 ;
  assign n36618 = n21312 & n36617 ;
  assign n36619 = ~\a[60]  & \b[26]  ;
  assign n36620 = n20513 & n36619 ;
  assign n36621 = ~n36618 & ~n36620 ;
  assign n36622 = n36616 & n36621 ;
  assign n36623 = ~n36612 & n36622 ;
  assign n36624 = ~\a[23]  & \b[23]  ;
  assign n36625 = n21957 & n36624 ;
  assign n36626 = ~\a[23]  & \b[24]  ;
  assign n36627 = n21958 & n36626 ;
  assign n36628 = ~n36625 & ~n36627 ;
  assign n36629 = \b[24]  & n21958 ;
  assign n36630 = \b[23]  & n21957 ;
  assign n36631 = \a[23]  & ~n36630 ;
  assign n36632 = ~n36629 & n36631 ;
  assign n36633 = n36628 & ~n36632 ;
  assign n36634 = ~\a[62]  & ~n36221 ;
  assign n36635 = ~n36633 & n36634 ;
  assign n36636 = ~\a[62]  & n36221 ;
  assign n36637 = n36633 & n36636 ;
  assign n36638 = ~n36635 & ~n36637 ;
  assign n36639 = ~n36623 & ~n36638 ;
  assign n36640 = \a[62]  & ~n36221 ;
  assign n36641 = ~n36633 & n36640 ;
  assign n36642 = \a[62]  & n36221 ;
  assign n36643 = n36633 & n36642 ;
  assign n36644 = ~n36641 & ~n36643 ;
  assign n36645 = n36622 & ~n36644 ;
  assign n36646 = ~n36612 & n36645 ;
  assign n36647 = ~n36639 & ~n36646 ;
  assign n36648 = ~\a[62]  & ~n36623 ;
  assign n36649 = ~n36221 & ~n36633 ;
  assign n36650 = n36221 & n36633 ;
  assign n36651 = ~n36649 & ~n36650 ;
  assign n36652 = \a[62]  & n36622 ;
  assign n36653 = ~n36612 & n36652 ;
  assign n36654 = n36651 & ~n36653 ;
  assign n36655 = ~n36648 & n36654 ;
  assign n36656 = n36647 & ~n36655 ;
  assign n36657 = ~n36610 & ~n36656 ;
  assign n36658 = n36610 & ~n36646 ;
  assign n36659 = ~n36639 & n36658 ;
  assign n36660 = ~n36655 & n36659 ;
  assign n36661 = ~n36657 & ~n36660 ;
  assign n36662 = ~n36608 & ~n36661 ;
  assign n36663 = n36608 & n36661 ;
  assign n36664 = ~n36662 & ~n36663 ;
  assign n36665 = n36201 & ~n36239 ;
  assign n36666 = ~n36240 & ~n36665 ;
  assign n36667 = ~n36664 & ~n36666 ;
  assign n36668 = n36664 & n36666 ;
  assign n36669 = ~n36667 & ~n36668 ;
  assign n36670 = ~n5852 & n16655 ;
  assign n36671 = ~n5809 & n16655 ;
  assign n36672 = ~n5848 & n36671 ;
  assign n36673 = ~n36670 & ~n36672 ;
  assign n36674 = ~n5855 & ~n36673 ;
  assign n36675 = \b[31]  & n17308 ;
  assign n36676 = n17305 & n36675 ;
  assign n36677 = \b[33]  & n16653 ;
  assign n36678 = \a[54]  & \b[32]  ;
  assign n36679 = n16644 & n36678 ;
  assign n36680 = ~\a[54]  & \b[32]  ;
  assign n36681 = n16647 & n36680 ;
  assign n36682 = ~n36679 & ~n36681 ;
  assign n36683 = ~n36677 & n36682 ;
  assign n36684 = ~n36676 & n36683 ;
  assign n36685 = ~\a[56]  & n36684 ;
  assign n36686 = ~n36674 & n36685 ;
  assign n36687 = \a[56]  & ~n36684 ;
  assign n36688 = \a[56]  & ~n5855 ;
  assign n36689 = ~n36673 & n36688 ;
  assign n36690 = ~n36687 & ~n36689 ;
  assign n36691 = ~n36686 & n36690 ;
  assign n36692 = ~n36248 & n36272 ;
  assign n36693 = n36246 & ~n36692 ;
  assign n36694 = ~n36691 & ~n36693 ;
  assign n36695 = ~n36669 & n36694 ;
  assign n36696 = n36246 & n36691 ;
  assign n36697 = ~n36692 & n36696 ;
  assign n36698 = n36669 & ~n36697 ;
  assign n36699 = ~n36694 & n36698 ;
  assign n36700 = ~n36669 & n36697 ;
  assign n36701 = ~n36699 & ~n36700 ;
  assign n36702 = ~n36695 & n36701 ;
  assign n36703 = n36176 & ~n36278 ;
  assign n36704 = ~n36279 & ~n36703 ;
  assign n36705 = n7337 & n14793 ;
  assign n36706 = ~n7334 & n36705 ;
  assign n36707 = ~n7337 & n14793 ;
  assign n36708 = ~n6605 & n36707 ;
  assign n36709 = ~n7333 & n36708 ;
  assign n36710 = \b[34]  & n15517 ;
  assign n36711 = n15514 & n36710 ;
  assign n36712 = ~\a[51]  & \b[35]  ;
  assign n36713 = n14785 & n36712 ;
  assign n36714 = ~n36711 & ~n36713 ;
  assign n36715 = \b[36]  & n14791 ;
  assign n36716 = \a[51]  & \b[35]  ;
  assign n36717 = n14782 & n36716 ;
  assign n36718 = \a[53]  & ~n36717 ;
  assign n36719 = ~n36715 & n36718 ;
  assign n36720 = n36714 & n36719 ;
  assign n36721 = ~n36709 & n36720 ;
  assign n36722 = ~n36706 & n36721 ;
  assign n36723 = ~n36715 & ~n36717 ;
  assign n36724 = n36714 & n36723 ;
  assign n36725 = ~n36709 & n36724 ;
  assign n36726 = ~n36706 & n36725 ;
  assign n36727 = ~\a[53]  & ~n36726 ;
  assign n36728 = ~n36722 & ~n36727 ;
  assign n36729 = ~n36704 & ~n36728 ;
  assign n36730 = n36702 & n36729 ;
  assign n36731 = ~n36704 & n36728 ;
  assign n36732 = ~n36702 & n36731 ;
  assign n36733 = ~n36730 & ~n36732 ;
  assign n36734 = ~n36702 & n36728 ;
  assign n36735 = ~n36695 & ~n36728 ;
  assign n36736 = n36701 & n36735 ;
  assign n36737 = n36704 & ~n36736 ;
  assign n36738 = ~n36734 & n36737 ;
  assign n36739 = n36733 & ~n36738 ;
  assign n36740 = ~n8602 & n13125 ;
  assign n36741 = ~n8600 & n36740 ;
  assign n36742 = \b[39]  & n13123 ;
  assign n36743 = \a[48]  & \b[38]  ;
  assign n36744 = n13786 & n36743 ;
  assign n36745 = ~n36742 & ~n36744 ;
  assign n36746 = \b[37]  & n13794 ;
  assign n36747 = n13792 & n36746 ;
  assign n36748 = ~\a[48]  & \b[38]  ;
  assign n36749 = n13117 & n36748 ;
  assign n36750 = ~n36747 & ~n36749 ;
  assign n36751 = n36745 & n36750 ;
  assign n36752 = ~n36741 & n36751 ;
  assign n36753 = ~\a[50]  & ~n36752 ;
  assign n36754 = \a[50]  & n36751 ;
  assign n36755 = ~n36741 & n36754 ;
  assign n36756 = ~n36753 & ~n36755 ;
  assign n36757 = n36739 & ~n36756 ;
  assign n36758 = ~n36739 & n36756 ;
  assign n36759 = ~n36757 & ~n36758 ;
  assign n36760 = n36283 & ~n36285 ;
  assign n36761 = ~n36283 & n36285 ;
  assign n36762 = n36309 & ~n36761 ;
  assign n36763 = ~n36760 & ~n36762 ;
  assign n36764 = ~n9930 & ~n10988 ;
  assign n36765 = ~n11569 & n36764 ;
  assign n36766 = n9927 & n36765 ;
  assign n36767 = n9930 & ~n10988 ;
  assign n36768 = ~n11569 & n36767 ;
  assign n36769 = ~n9927 & n36768 ;
  assign n36770 = ~n36766 & ~n36769 ;
  assign n36771 = \b[40]  & n12159 ;
  assign n36772 = n12156 & n36771 ;
  assign n36773 = ~\a[45]  & \b[41]  ;
  assign n36774 = n11564 & n36773 ;
  assign n36775 = ~n36772 & ~n36774 ;
  assign n36776 = \b[42]  & n11570 ;
  assign n36777 = \a[45]  & \b[41]  ;
  assign n36778 = n11561 & n36777 ;
  assign n36779 = \a[47]  & ~n36778 ;
  assign n36780 = ~n36776 & n36779 ;
  assign n36781 = n36775 & n36780 ;
  assign n36782 = n36770 & n36781 ;
  assign n36783 = ~n36776 & ~n36778 ;
  assign n36784 = n36775 & n36783 ;
  assign n36785 = n36770 & n36784 ;
  assign n36786 = ~\a[47]  & ~n36785 ;
  assign n36787 = ~n36782 & ~n36786 ;
  assign n36788 = ~n36763 & ~n36787 ;
  assign n36789 = n36759 & n36788 ;
  assign n36790 = n36763 & ~n36787 ;
  assign n36791 = ~n36759 & n36790 ;
  assign n36792 = ~n36789 & ~n36791 ;
  assign n36793 = ~n36763 & n36787 ;
  assign n36794 = ~n36759 & n36793 ;
  assign n36795 = n36763 & n36787 ;
  assign n36796 = n36759 & n36795 ;
  assign n36797 = ~n36794 & ~n36796 ;
  assign n36798 = n36792 & n36797 ;
  assign n36799 = n10082 & ~n11397 ;
  assign n36800 = ~n11395 & n36799 ;
  assign n36801 = \b[43]  & n10681 ;
  assign n36802 = n10678 & n36801 ;
  assign n36803 = \b[45]  & n10080 ;
  assign n36804 = \a[41]  & \b[44]  ;
  assign n36805 = n10679 & n36804 ;
  assign n36806 = ~\a[42]  & \b[44]  ;
  assign n36807 = n10074 & n36806 ;
  assign n36808 = ~n36805 & ~n36807 ;
  assign n36809 = ~n36803 & n36808 ;
  assign n36810 = ~n36802 & n36809 ;
  assign n36811 = ~\a[44]  & n36810 ;
  assign n36812 = ~n36800 & n36811 ;
  assign n36813 = ~n36800 & n36810 ;
  assign n36814 = \a[44]  & ~n36813 ;
  assign n36815 = ~n36812 & ~n36814 ;
  assign n36816 = n36153 & ~n36321 ;
  assign n36817 = ~n36322 & ~n36816 ;
  assign n36818 = n36815 & ~n36817 ;
  assign n36819 = n36798 & n36818 ;
  assign n36820 = n36815 & n36817 ;
  assign n36821 = ~n36798 & n36820 ;
  assign n36822 = ~n36819 & ~n36821 ;
  assign n36823 = ~n36815 & ~n36817 ;
  assign n36824 = ~n36798 & n36823 ;
  assign n36825 = ~n36815 & n36817 ;
  assign n36826 = n36798 & n36825 ;
  assign n36827 = ~n36824 & ~n36826 ;
  assign n36828 = n36822 & n36827 ;
  assign n36829 = ~n36326 & n36346 ;
  assign n36830 = n36351 & ~n36829 ;
  assign n36831 = n8759 & n12478 ;
  assign n36832 = ~n12475 & n36831 ;
  assign n36833 = n8759 & n28668 ;
  assign n36834 = ~n12474 & n36833 ;
  assign n36835 = \b[46]  & n9301 ;
  assign n36836 = n9298 & n36835 ;
  assign n36837 = ~\a[39]  & \b[47]  ;
  assign n36838 = n8751 & n36837 ;
  assign n36839 = ~n36836 & ~n36838 ;
  assign n36840 = \b[48]  & n8757 ;
  assign n36841 = \a[39]  & \b[47]  ;
  assign n36842 = n8748 & n36841 ;
  assign n36843 = \a[41]  & ~n36842 ;
  assign n36844 = ~n36840 & n36843 ;
  assign n36845 = n36839 & n36844 ;
  assign n36846 = ~n36834 & n36845 ;
  assign n36847 = ~n36832 & n36846 ;
  assign n36848 = ~n36840 & ~n36842 ;
  assign n36849 = n36839 & n36848 ;
  assign n36850 = ~n36834 & n36849 ;
  assign n36851 = ~n36832 & n36850 ;
  assign n36852 = ~\a[41]  & ~n36851 ;
  assign n36853 = ~n36847 & ~n36852 ;
  assign n36854 = ~n36830 & ~n36853 ;
  assign n36855 = ~n36828 & n36854 ;
  assign n36856 = n36830 & ~n36853 ;
  assign n36857 = n36828 & n36856 ;
  assign n36858 = ~n36855 & ~n36857 ;
  assign n36859 = n36830 & n36853 ;
  assign n36860 = ~n36828 & n36859 ;
  assign n36861 = ~n36830 & n36853 ;
  assign n36862 = n36828 & n36861 ;
  assign n36863 = ~n36860 & ~n36862 ;
  assign n36864 = n36858 & n36863 ;
  assign n36865 = ~n36362 & n36383 ;
  assign n36866 = ~n36363 & ~n36865 ;
  assign n36867 = n7534 & ~n14098 ;
  assign n36868 = ~n14096 & n36867 ;
  assign n36869 = \b[51]  & n7532 ;
  assign n36870 = \a[36]  & \b[50]  ;
  assign n36871 = n17801 & n36870 ;
  assign n36872 = ~n36869 & ~n36871 ;
  assign n36873 = \b[49]  & n7973 ;
  assign n36874 = n7970 & n36873 ;
  assign n36875 = ~\a[36]  & \b[50]  ;
  assign n36876 = n7526 & n36875 ;
  assign n36877 = ~n36874 & ~n36876 ;
  assign n36878 = n36872 & n36877 ;
  assign n36879 = ~n36868 & n36878 ;
  assign n36880 = ~\a[38]  & ~n36879 ;
  assign n36881 = \a[38]  & n36878 ;
  assign n36882 = ~n36868 & n36881 ;
  assign n36883 = ~n36880 & ~n36882 ;
  assign n36884 = ~n36866 & n36883 ;
  assign n36885 = ~n36864 & n36884 ;
  assign n36886 = n36866 & n36883 ;
  assign n36887 = n36864 & n36886 ;
  assign n36888 = ~n36885 & ~n36887 ;
  assign n36889 = ~n36866 & ~n36883 ;
  assign n36890 = n36864 & n36889 ;
  assign n36891 = n36866 & ~n36883 ;
  assign n36892 = ~n36864 & n36891 ;
  assign n36893 = ~n36890 & ~n36892 ;
  assign n36894 = n36888 & n36893 ;
  assign n36895 = n36586 & ~n36894 ;
  assign n36896 = ~n36586 & n36894 ;
  assign n36897 = ~n36895 & ~n36896 ;
  assign n36898 = n36584 & ~n36897 ;
  assign n36899 = ~n36584 & n36897 ;
  assign n36900 = ~n36898 & ~n36899 ;
  assign n36901 = ~n36425 & ~n36448 ;
  assign n36902 = n36425 & n36448 ;
  assign n36903 = n36444 & ~n36902 ;
  assign n36904 = ~n36901 & ~n36903 ;
  assign n36905 = n36900 & n36904 ;
  assign n36906 = ~n36900 & ~n36904 ;
  assign n36907 = ~n36905 & ~n36906 ;
  assign n36908 = n36558 & n36907 ;
  assign n36909 = ~n36558 & ~n36907 ;
  assign n36910 = ~n36908 & ~n36909 ;
  assign n36911 = ~n36533 & n36910 ;
  assign n36912 = ~n36509 & n36911 ;
  assign n36913 = n36533 & n36910 ;
  assign n36914 = n36509 & n36913 ;
  assign n36915 = ~n36912 & ~n36914 ;
  assign n36916 = ~n36509 & ~n36910 ;
  assign n36917 = n36533 & n36916 ;
  assign n36918 = ~n36533 & ~n36910 ;
  assign n36919 = n36509 & n36918 ;
  assign n36920 = ~n36917 & ~n36919 ;
  assign n36921 = n36915 & n36920 ;
  assign n36922 = n36506 & n36921 ;
  assign n36923 = ~n36506 & ~n36921 ;
  assign n36924 = ~n36922 & ~n36923 ;
  assign n36925 = ~n36483 & n36924 ;
  assign n36926 = n36483 & ~n36924 ;
  assign n36927 = ~n36925 & ~n36926 ;
  assign n36928 = ~n36475 & n36927 ;
  assign n36929 = ~n36482 & n36928 ;
  assign n36930 = ~n36475 & ~n36482 ;
  assign n36931 = ~n36927 & ~n36930 ;
  assign n36932 = ~n36929 & ~n36931 ;
  assign n36933 = ~n36925 & ~n36929 ;
  assign n36934 = ~n36504 & ~n36921 ;
  assign n36935 = ~n36505 & ~n36934 ;
  assign n36936 = ~n36899 & ~n36904 ;
  assign n36937 = n5211 & n18940 ;
  assign n36938 = ~n18937 & n36937 ;
  assign n36939 = n5211 & ~n18940 ;
  assign n36940 = ~n17685 & n36939 ;
  assign n36941 = ~n18936 & n36940 ;
  assign n36942 = \b[58]  & n5209 ;
  assign n36943 = \a[30]  & \b[57]  ;
  assign n36944 = n5200 & n36943 ;
  assign n36945 = ~n36942 & ~n36944 ;
  assign n36946 = \b[56]  & n5595 ;
  assign n36947 = n5592 & n36946 ;
  assign n36948 = ~\a[30]  & \b[57]  ;
  assign n36949 = n5203 & n36948 ;
  assign n36950 = ~n36947 & ~n36949 ;
  assign n36951 = n36945 & n36950 ;
  assign n36952 = ~n36941 & n36951 ;
  assign n36953 = ~n36938 & n36952 ;
  assign n36954 = \a[32]  & ~n36953 ;
  assign n36955 = ~\a[32]  & n36953 ;
  assign n36956 = ~n36954 & ~n36955 ;
  assign n36957 = ~n36898 & n36956 ;
  assign n36958 = ~n36936 & n36957 ;
  assign n36959 = ~n36898 & ~n36936 ;
  assign n36960 = ~\a[32]  & ~n36953 ;
  assign n36961 = \a[32]  & n36951 ;
  assign n36962 = ~n36941 & n36961 ;
  assign n36963 = ~n36938 & n36962 ;
  assign n36964 = ~n36960 & ~n36963 ;
  assign n36965 = ~n36959 & n36964 ;
  assign n36966 = ~n36958 & ~n36965 ;
  assign n36967 = n6309 & ~n16446 ;
  assign n36968 = ~n16444 & n36967 ;
  assign n36969 = \b[53]  & n6778 ;
  assign n36970 = n6775 & n36969 ;
  assign n36971 = ~\a[33]  & \b[54]  ;
  assign n36972 = n6301 & n36971 ;
  assign n36973 = ~n36970 & ~n36972 ;
  assign n36974 = \b[55]  & n6307 ;
  assign n36975 = \a[33]  & \b[54]  ;
  assign n36976 = n6298 & n36975 ;
  assign n36977 = \a[35]  & ~n36976 ;
  assign n36978 = ~n36974 & n36977 ;
  assign n36979 = n36973 & n36978 ;
  assign n36980 = ~n36968 & n36979 ;
  assign n36981 = ~n36974 & ~n36976 ;
  assign n36982 = n36973 & n36981 ;
  assign n36983 = ~n36968 & n36982 ;
  assign n36984 = ~\a[35]  & ~n36983 ;
  assign n36985 = ~n36980 & ~n36984 ;
  assign n36986 = ~n36757 & ~n36763 ;
  assign n36987 = ~n36758 & ~n36986 ;
  assign n36988 = ~n36697 & ~n36699 ;
  assign n36989 = ~n36662 & ~n36666 ;
  assign n36990 = ~n36663 & ~n36989 ;
  assign n36991 = \a[62]  & n36651 ;
  assign n36992 = ~n36623 & n36991 ;
  assign n36993 = ~\a[62]  & n36651 ;
  assign n36994 = n36623 & n36993 ;
  assign n36995 = ~n36992 & ~n36994 ;
  assign n36996 = ~n36659 & n36995 ;
  assign n36997 = n4456 & n20521 ;
  assign n36998 = ~n18723 & n36997 ;
  assign n36999 = n16805 & n20521 ;
  assign n37000 = ~n4452 & n36999 ;
  assign n37001 = \b[28]  & n20519 ;
  assign n37002 = \a[60]  & \b[27]  ;
  assign n37003 = n20510 & n37002 ;
  assign n37004 = ~n37001 & ~n37003 ;
  assign n37005 = \b[26]  & n21315 ;
  assign n37006 = n21312 & n37005 ;
  assign n37007 = ~\a[60]  & \b[27]  ;
  assign n37008 = n20513 & n37007 ;
  assign n37009 = ~n37006 & ~n37008 ;
  assign n37010 = n37004 & n37009 ;
  assign n37011 = ~n37000 & n37010 ;
  assign n37012 = ~n36998 & n37011 ;
  assign n37013 = n36628 & n36632 ;
  assign n37014 = n36221 & n36628 ;
  assign n37015 = ~n37013 & ~n37014 ;
  assign n37016 = \b[25]  & n21958 ;
  assign n37017 = \b[24]  & n21957 ;
  assign n37018 = ~n37016 & ~n37017 ;
  assign n37019 = ~\a[62]  & ~n37018 ;
  assign n37020 = n37015 & n37019 ;
  assign n37021 = ~\a[62]  & n37018 ;
  assign n37022 = ~n37015 & n37021 ;
  assign n37023 = ~n37020 & ~n37022 ;
  assign n37024 = ~n37012 & ~n37023 ;
  assign n37025 = \a[62]  & ~n37018 ;
  assign n37026 = n37015 & n37025 ;
  assign n37027 = \a[62]  & n37018 ;
  assign n37028 = ~n37015 & n37027 ;
  assign n37029 = ~n37026 & ~n37028 ;
  assign n37030 = n37010 & ~n37029 ;
  assign n37031 = ~n37000 & n37030 ;
  assign n37032 = ~n36998 & n37031 ;
  assign n37033 = ~n37024 & ~n37032 ;
  assign n37034 = ~\a[62]  & ~n37012 ;
  assign n37035 = ~n37015 & ~n37018 ;
  assign n37036 = n37015 & n37018 ;
  assign n37037 = ~n37035 & ~n37036 ;
  assign n37038 = \a[62]  & n37010 ;
  assign n37039 = ~n37000 & n37038 ;
  assign n37040 = ~n36998 & n37039 ;
  assign n37041 = ~n37037 & ~n37040 ;
  assign n37042 = ~n37034 & n37041 ;
  assign n37043 = n37033 & ~n37042 ;
  assign n37044 = n36996 & n37043 ;
  assign n37045 = ~n36996 & ~n37043 ;
  assign n37046 = ~n37044 & ~n37045 ;
  assign n37047 = ~n5459 & n18516 ;
  assign n37048 = ~n5104 & n18516 ;
  assign n37049 = ~n5455 & n37048 ;
  assign n37050 = ~n37047 & ~n37049 ;
  assign n37051 = ~n5462 & ~n37050 ;
  assign n37052 = \b[31]  & n18514 ;
  assign n37053 = \a[56]  & \b[30]  ;
  assign n37054 = n19181 & n37053 ;
  assign n37055 = ~\a[57]  & \b[30]  ;
  assign n37056 = n18508 & n37055 ;
  assign n37057 = ~n37054 & ~n37056 ;
  assign n37058 = ~n37052 & n37057 ;
  assign n37059 = \b[29]  & n19183 ;
  assign n37060 = n19180 & n37059 ;
  assign n37061 = \a[59]  & ~n37060 ;
  assign n37062 = n37058 & n37061 ;
  assign n37063 = ~n37051 & n37062 ;
  assign n37064 = n37058 & ~n37060 ;
  assign n37065 = ~\a[59]  & ~n37064 ;
  assign n37066 = ~\a[59]  & ~n5462 ;
  assign n37067 = ~n37050 & n37066 ;
  assign n37068 = ~n37065 & ~n37067 ;
  assign n37069 = ~n37063 & n37068 ;
  assign n37070 = n37046 & ~n37069 ;
  assign n37071 = ~n37046 & n37069 ;
  assign n37072 = ~n37070 & ~n37071 ;
  assign n37073 = ~n36990 & ~n37072 ;
  assign n37074 = n36990 & n37072 ;
  assign n37075 = ~n37073 & ~n37074 ;
  assign n37076 = n6565 & n16655 ;
  assign n37077 = ~n6562 & n37076 ;
  assign n37078 = ~n6565 & n16655 ;
  assign n37079 = ~n5850 & n37078 ;
  assign n37080 = ~n6561 & n37079 ;
  assign n37081 = \b[32]  & n17308 ;
  assign n37082 = n17305 & n37081 ;
  assign n37083 = \b[34]  & n16653 ;
  assign n37084 = \a[53]  & \b[33]  ;
  assign n37085 = n17306 & n37084 ;
  assign n37086 = ~\a[54]  & \b[33]  ;
  assign n37087 = n16647 & n37086 ;
  assign n37088 = ~n37085 & ~n37087 ;
  assign n37089 = ~n37083 & n37088 ;
  assign n37090 = ~n37082 & n37089 ;
  assign n37091 = ~n37080 & n37090 ;
  assign n37092 = ~n37077 & n37091 ;
  assign n37093 = ~\a[56]  & ~n37092 ;
  assign n37094 = \a[56]  & n37090 ;
  assign n37095 = ~n37080 & n37094 ;
  assign n37096 = ~n37077 & n37095 ;
  assign n37097 = ~n37093 & ~n37096 ;
  assign n37098 = ~n37075 & n37097 ;
  assign n37099 = n37075 & ~n37097 ;
  assign n37100 = ~n37098 & ~n37099 ;
  assign n37101 = n36988 & ~n37100 ;
  assign n37102 = ~n36988 & n37100 ;
  assign n37103 = ~n37101 & ~n37102 ;
  assign n37104 = ~n7758 & n14793 ;
  assign n37105 = ~n7336 & n14793 ;
  assign n37106 = ~n7754 & n37105 ;
  assign n37107 = ~n37104 & ~n37106 ;
  assign n37108 = ~n7761 & ~n37107 ;
  assign n37109 = \b[37]  & n14791 ;
  assign n37110 = \a[50]  & \b[36]  ;
  assign n37111 = n15515 & n37110 ;
  assign n37112 = ~\a[51]  & \b[36]  ;
  assign n37113 = n14785 & n37112 ;
  assign n37114 = ~n37111 & ~n37113 ;
  assign n37115 = ~n37109 & n37114 ;
  assign n37116 = \b[35]  & n15517 ;
  assign n37117 = n15514 & n37116 ;
  assign n37118 = \a[53]  & ~n37117 ;
  assign n37119 = n37115 & n37118 ;
  assign n37120 = ~n37108 & n37119 ;
  assign n37121 = n37115 & ~n37117 ;
  assign n37122 = ~\a[53]  & ~n37121 ;
  assign n37123 = ~\a[53]  & ~n7761 ;
  assign n37124 = ~n37107 & n37123 ;
  assign n37125 = ~n37122 & ~n37124 ;
  assign n37126 = ~n37120 & n37125 ;
  assign n37127 = ~n37103 & n37126 ;
  assign n37128 = n37103 & ~n37126 ;
  assign n37129 = ~n37127 & ~n37128 ;
  assign n37130 = n9044 & n13125 ;
  assign n37131 = ~n9041 & n37130 ;
  assign n37132 = ~n9044 & n13125 ;
  assign n37133 = ~n8597 & n37132 ;
  assign n37134 = ~n9040 & n37133 ;
  assign n37135 = \b[38]  & n13794 ;
  assign n37136 = n13792 & n37135 ;
  assign n37137 = \b[40]  & n13123 ;
  assign n37138 = \a[48]  & \b[39]  ;
  assign n37139 = n13786 & n37138 ;
  assign n37140 = ~\a[48]  & \b[39]  ;
  assign n37141 = n13117 & n37140 ;
  assign n37142 = ~n37139 & ~n37141 ;
  assign n37143 = ~n37137 & n37142 ;
  assign n37144 = ~n37136 & n37143 ;
  assign n37145 = ~n37134 & n37144 ;
  assign n37146 = ~n37131 & n37145 ;
  assign n37147 = ~\a[50]  & ~n37146 ;
  assign n37148 = \a[50]  & n37144 ;
  assign n37149 = ~n37134 & n37148 ;
  assign n37150 = ~n37131 & n37149 ;
  assign n37151 = ~n37147 & ~n37150 ;
  assign n37152 = ~n36704 & ~n36736 ;
  assign n37153 = ~n36734 & ~n37152 ;
  assign n37154 = ~n37151 & n37153 ;
  assign n37155 = ~n37129 & n37154 ;
  assign n37156 = ~n37151 & ~n37153 ;
  assign n37157 = n37129 & n37156 ;
  assign n37158 = ~n37155 & ~n37157 ;
  assign n37159 = n37151 & ~n37153 ;
  assign n37160 = ~n37129 & n37159 ;
  assign n37161 = n37151 & n37153 ;
  assign n37162 = n37129 & n37161 ;
  assign n37163 = ~n37160 & ~n37162 ;
  assign n37164 = n37158 & n37163 ;
  assign n37165 = n36987 & n37164 ;
  assign n37166 = ~n36987 & ~n37164 ;
  assign n37167 = ~n37165 & ~n37166 ;
  assign n37168 = ~n10406 & n11572 ;
  assign n37169 = ~n9929 & n11572 ;
  assign n37170 = ~n10402 & n37169 ;
  assign n37171 = ~n37168 & ~n37170 ;
  assign n37172 = ~n10409 & ~n37171 ;
  assign n37173 = \b[41]  & n12159 ;
  assign n37174 = n12156 & n37173 ;
  assign n37175 = ~\a[45]  & \b[42]  ;
  assign n37176 = n11564 & n37175 ;
  assign n37177 = ~n37174 & ~n37176 ;
  assign n37178 = \b[43]  & n11570 ;
  assign n37179 = \a[45]  & \b[42]  ;
  assign n37180 = n11561 & n37179 ;
  assign n37181 = \a[47]  & ~n37180 ;
  assign n37182 = ~n37178 & n37181 ;
  assign n37183 = n37177 & n37182 ;
  assign n37184 = ~n37172 & n37183 ;
  assign n37185 = ~n37178 & ~n37180 ;
  assign n37186 = n37177 & n37185 ;
  assign n37187 = ~\a[47]  & ~n37186 ;
  assign n37188 = ~\a[47]  & ~n10409 ;
  assign n37189 = ~n37171 & n37188 ;
  assign n37190 = ~n37187 & ~n37189 ;
  assign n37191 = ~n37184 & n37190 ;
  assign n37192 = n37167 & ~n37191 ;
  assign n37193 = ~n37167 & n37191 ;
  assign n37194 = ~n37192 & ~n37193 ;
  assign n37195 = n36792 & ~n36817 ;
  assign n37196 = n36797 & ~n37195 ;
  assign n37197 = n10082 & n11906 ;
  assign n37198 = ~n11903 & n37197 ;
  assign n37199 = n10082 & n13483 ;
  assign n37200 = ~n11902 & n37199 ;
  assign n37201 = \b[44]  & n10681 ;
  assign n37202 = n10678 & n37201 ;
  assign n37203 = \b[46]  & n10080 ;
  assign n37204 = \a[41]  & \b[45]  ;
  assign n37205 = n10679 & n37204 ;
  assign n37206 = ~\a[42]  & \b[45]  ;
  assign n37207 = n10074 & n37206 ;
  assign n37208 = ~n37205 & ~n37207 ;
  assign n37209 = ~n37203 & n37208 ;
  assign n37210 = ~n37202 & n37209 ;
  assign n37211 = ~n37200 & n37210 ;
  assign n37212 = ~n37198 & n37211 ;
  assign n37213 = ~\a[44]  & ~n37212 ;
  assign n37214 = \a[44]  & n37210 ;
  assign n37215 = ~n37200 & n37214 ;
  assign n37216 = ~n37198 & n37215 ;
  assign n37217 = ~n37213 & ~n37216 ;
  assign n37218 = ~n37196 & n37217 ;
  assign n37219 = ~n37194 & n37218 ;
  assign n37220 = n37196 & n37217 ;
  assign n37221 = n37194 & n37220 ;
  assign n37222 = ~n37219 & ~n37221 ;
  assign n37223 = n37196 & ~n37217 ;
  assign n37224 = ~n37194 & n37223 ;
  assign n37225 = ~n37196 & ~n37217 ;
  assign n37226 = n37194 & n37225 ;
  assign n37227 = ~n37224 & ~n37226 ;
  assign n37228 = n37222 & n37227 ;
  assign n37229 = n36822 & n36830 ;
  assign n37230 = n36827 & ~n37229 ;
  assign n37231 = n8759 & ~n13524 ;
  assign n37232 = ~n13522 & n37231 ;
  assign n37233 = \b[47]  & n9301 ;
  assign n37234 = n9298 & n37233 ;
  assign n37235 = ~\a[39]  & \b[48]  ;
  assign n37236 = n8751 & n37235 ;
  assign n37237 = ~n37234 & ~n37236 ;
  assign n37238 = \b[49]  & n8757 ;
  assign n37239 = \a[39]  & \b[48]  ;
  assign n37240 = n8748 & n37239 ;
  assign n37241 = \a[41]  & ~n37240 ;
  assign n37242 = ~n37238 & n37241 ;
  assign n37243 = n37237 & n37242 ;
  assign n37244 = ~n37232 & n37243 ;
  assign n37245 = ~n37238 & ~n37240 ;
  assign n37246 = n37237 & n37245 ;
  assign n37247 = ~n37232 & n37246 ;
  assign n37248 = ~\a[41]  & ~n37247 ;
  assign n37249 = ~n37244 & ~n37248 ;
  assign n37250 = n37230 & ~n37249 ;
  assign n37251 = ~n37228 & n37250 ;
  assign n37252 = ~n37230 & ~n37249 ;
  assign n37253 = n37228 & n37252 ;
  assign n37254 = ~n37251 & ~n37253 ;
  assign n37255 = ~n37230 & n37249 ;
  assign n37256 = ~n37228 & n37255 ;
  assign n37257 = n37230 & n37249 ;
  assign n37258 = n37228 & n37257 ;
  assign n37259 = ~n37256 & ~n37258 ;
  assign n37260 = n37254 & n37259 ;
  assign n37261 = n36858 & ~n36866 ;
  assign n37262 = n36863 & ~n37261 ;
  assign n37263 = n7534 & n15201 ;
  assign n37264 = ~n15198 & n37263 ;
  assign n37265 = n7534 & ~n15201 ;
  assign n37266 = ~n14093 & n37265 ;
  assign n37267 = ~n15197 & n37266 ;
  assign n37268 = \b[50]  & n7973 ;
  assign n37269 = n7970 & n37268 ;
  assign n37270 = ~\a[36]  & \b[51]  ;
  assign n37271 = n7526 & n37270 ;
  assign n37272 = ~n37269 & ~n37271 ;
  assign n37273 = \b[52]  & n7532 ;
  assign n37274 = \a[36]  & \b[51]  ;
  assign n37275 = n17801 & n37274 ;
  assign n37276 = \a[38]  & ~n37275 ;
  assign n37277 = ~n37273 & n37276 ;
  assign n37278 = n37272 & n37277 ;
  assign n37279 = ~n37267 & n37278 ;
  assign n37280 = ~n37264 & n37279 ;
  assign n37281 = ~n37273 & ~n37275 ;
  assign n37282 = n37272 & n37281 ;
  assign n37283 = ~n37267 & n37282 ;
  assign n37284 = ~n37264 & n37283 ;
  assign n37285 = ~\a[38]  & ~n37284 ;
  assign n37286 = ~n37280 & ~n37285 ;
  assign n37287 = ~n37262 & n37286 ;
  assign n37288 = ~n37260 & n37287 ;
  assign n37289 = n37262 & n37286 ;
  assign n37290 = n37260 & n37289 ;
  assign n37291 = ~n37288 & ~n37290 ;
  assign n37292 = n37262 & ~n37286 ;
  assign n37293 = ~n37260 & n37292 ;
  assign n37294 = ~n37262 & ~n37286 ;
  assign n37295 = n37260 & n37294 ;
  assign n37296 = ~n37293 & ~n37295 ;
  assign n37297 = n37291 & n37296 ;
  assign n37298 = n36586 & n36893 ;
  assign n37299 = n36888 & ~n37298 ;
  assign n37300 = n37297 & n37299 ;
  assign n37301 = ~n37297 & ~n37299 ;
  assign n37302 = ~n37300 & ~n37301 ;
  assign n37303 = n36985 & n37302 ;
  assign n37304 = ~n36985 & ~n37302 ;
  assign n37305 = ~n37303 & ~n37304 ;
  assign n37306 = n36966 & ~n37305 ;
  assign n37307 = ~n36966 & n37305 ;
  assign n37308 = ~n37306 & ~n37307 ;
  assign n37309 = ~n36557 & ~n36907 ;
  assign n37310 = n4249 & ~n20971 ;
  assign n37311 = ~n20969 & n37310 ;
  assign n37312 = \b[61]  & n4247 ;
  assign n37313 = \a[27]  & \b[60]  ;
  assign n37314 = n4238 & n37313 ;
  assign n37315 = ~n37312 & ~n37314 ;
  assign n37316 = \b[59]  & n4647 ;
  assign n37317 = n4644 & n37316 ;
  assign n37318 = ~\a[27]  & \b[60]  ;
  assign n37319 = n4241 & n37318 ;
  assign n37320 = ~n37317 & ~n37319 ;
  assign n37321 = n37315 & n37320 ;
  assign n37322 = ~n37311 & n37321 ;
  assign n37323 = \a[29]  & ~n37322 ;
  assign n37324 = ~\a[29]  & n37322 ;
  assign n37325 = ~n37323 & ~n37324 ;
  assign n37326 = n36554 & n37325 ;
  assign n37327 = ~n37309 & n37326 ;
  assign n37328 = ~\a[29]  & ~n37322 ;
  assign n37329 = \a[29]  & n37321 ;
  assign n37330 = ~n37311 & n37329 ;
  assign n37331 = ~n36554 & ~n37330 ;
  assign n37332 = ~n36557 & ~n37330 ;
  assign n37333 = ~n36907 & n37332 ;
  assign n37334 = ~n37331 & ~n37333 ;
  assign n37335 = ~n37328 & ~n37334 ;
  assign n37336 = ~n37327 & ~n37335 ;
  assign n37337 = n37308 & n37336 ;
  assign n37338 = ~n37308 & ~n37336 ;
  assign n37339 = ~n37337 & ~n37338 ;
  assign n37340 = \b[62]  & n3733 ;
  assign n37341 = n3730 & n37340 ;
  assign n37342 = ~\a[24]  & \b[63]  ;
  assign n37343 = n3394 & n37342 ;
  assign n37344 = \a[24]  & \b[63]  ;
  assign n37345 = n27626 & n37344 ;
  assign n37346 = ~n37343 & ~n37345 ;
  assign n37347 = ~n37341 & n37346 ;
  assign n37348 = ~\a[26]  & ~n37347 ;
  assign n37349 = n3402 & ~n22458 ;
  assign n37350 = ~\a[26]  & n37349 ;
  assign n37351 = ~n23173 & n37350 ;
  assign n37352 = ~n37348 & ~n37351 ;
  assign n37353 = ~n23173 & n37349 ;
  assign n37354 = \a[26]  & n37347 ;
  assign n37355 = ~n37353 & n37354 ;
  assign n37356 = n37352 & ~n37355 ;
  assign n37357 = n36910 & ~n37356 ;
  assign n37358 = n36509 & n37357 ;
  assign n37359 = ~n36533 & ~n37356 ;
  assign n37360 = n36910 & n37359 ;
  assign n37361 = n36509 & n37359 ;
  assign n37362 = ~n37360 & ~n37361 ;
  assign n37363 = ~n37358 & n37362 ;
  assign n37364 = ~n36910 & n37356 ;
  assign n37365 = ~n36509 & n37364 ;
  assign n37366 = n36533 & n37356 ;
  assign n37367 = ~n36910 & n37366 ;
  assign n37368 = ~n36509 & n37366 ;
  assign n37369 = ~n37367 & ~n37368 ;
  assign n37370 = ~n37365 & n37369 ;
  assign n37371 = n37363 & n37370 ;
  assign n37372 = n37339 & n37371 ;
  assign n37373 = ~n37339 & ~n37371 ;
  assign n37374 = ~n37372 & ~n37373 ;
  assign n37375 = n36935 & n37374 ;
  assign n37376 = ~n36935 & ~n37374 ;
  assign n37377 = ~n37375 & ~n37376 ;
  assign n37378 = ~n36933 & n37377 ;
  assign n37379 = ~n36925 & ~n37377 ;
  assign n37380 = ~n36929 & n37379 ;
  assign n37381 = ~n37378 & ~n37380 ;
  assign n37382 = ~n36925 & ~n37375 ;
  assign n37383 = ~n36929 & n37382 ;
  assign n37384 = ~n37339 & n37363 ;
  assign n37385 = n37370 & ~n37384 ;
  assign n37386 = ~n36958 & n37305 ;
  assign n37387 = ~n36958 & n36965 ;
  assign n37388 = ~n37386 & ~n37387 ;
  assign n37389 = n4249 & ~n21699 ;
  assign n37390 = ~n21697 & n37389 ;
  assign n37391 = \b[62]  & n4247 ;
  assign n37392 = \a[27]  & \b[61]  ;
  assign n37393 = n4238 & n37392 ;
  assign n37394 = ~n37391 & ~n37393 ;
  assign n37395 = \b[60]  & n4647 ;
  assign n37396 = n4644 & n37395 ;
  assign n37397 = ~\a[27]  & \b[61]  ;
  assign n37398 = n4241 & n37397 ;
  assign n37399 = ~n37396 & ~n37398 ;
  assign n37400 = n37394 & n37399 ;
  assign n37401 = ~n37390 & n37400 ;
  assign n37402 = ~\a[29]  & ~n37401 ;
  assign n37403 = \a[29]  & ~n37393 ;
  assign n37404 = ~n37391 & n37403 ;
  assign n37405 = n37399 & n37404 ;
  assign n37406 = ~n37390 & n37405 ;
  assign n37407 = ~n37402 & ~n37406 ;
  assign n37408 = ~n37388 & n37407 ;
  assign n37409 = \a[29]  & ~n37401 ;
  assign n37410 = ~\a[29]  & n37401 ;
  assign n37411 = ~n37409 & ~n37410 ;
  assign n37412 = n37388 & n37411 ;
  assign n37413 = ~n37408 & ~n37412 ;
  assign n37414 = n5211 & ~n19550 ;
  assign n37415 = ~n19548 & n37414 ;
  assign n37416 = \b[59]  & n5209 ;
  assign n37417 = \a[30]  & \b[58]  ;
  assign n37418 = n5200 & n37417 ;
  assign n37419 = ~n37416 & ~n37418 ;
  assign n37420 = \b[57]  & n5595 ;
  assign n37421 = n5592 & n37420 ;
  assign n37422 = ~\a[30]  & \b[58]  ;
  assign n37423 = n5203 & n37422 ;
  assign n37424 = ~n37421 & ~n37423 ;
  assign n37425 = n37419 & n37424 ;
  assign n37426 = ~n37415 & n37425 ;
  assign n37427 = ~\a[32]  & ~n37426 ;
  assign n37428 = \a[32]  & n37425 ;
  assign n37429 = ~n37415 & n37428 ;
  assign n37430 = n37301 & ~n37429 ;
  assign n37431 = n36985 & ~n37429 ;
  assign n37432 = ~n37300 & n37431 ;
  assign n37433 = ~n37430 & ~n37432 ;
  assign n37434 = ~n37427 & ~n37433 ;
  assign n37435 = n36985 & ~n37300 ;
  assign n37436 = ~n37301 & n37427 ;
  assign n37437 = ~n37435 & n37436 ;
  assign n37438 = \a[32]  & n37426 ;
  assign n37439 = ~n37301 & n37438 ;
  assign n37440 = ~n37435 & n37439 ;
  assign n37441 = ~n37437 & ~n37440 ;
  assign n37442 = ~n37434 & n37441 ;
  assign n37443 = n7534 & ~n15246 ;
  assign n37444 = ~n15244 & n37443 ;
  assign n37445 = \b[51]  & n7973 ;
  assign n37446 = n7970 & n37445 ;
  assign n37447 = ~\a[36]  & \b[52]  ;
  assign n37448 = n7526 & n37447 ;
  assign n37449 = ~n37446 & ~n37448 ;
  assign n37450 = \b[53]  & n7532 ;
  assign n37451 = \a[36]  & \b[52]  ;
  assign n37452 = n17801 & n37451 ;
  assign n37453 = \a[38]  & ~n37452 ;
  assign n37454 = ~n37450 & n37453 ;
  assign n37455 = n37449 & n37454 ;
  assign n37456 = ~n37444 & n37455 ;
  assign n37457 = ~n37450 & ~n37452 ;
  assign n37458 = n37449 & n37457 ;
  assign n37459 = ~n37444 & n37458 ;
  assign n37460 = ~\a[38]  & ~n37459 ;
  assign n37461 = ~n37456 & ~n37460 ;
  assign n37462 = ~n9482 & n13125 ;
  assign n37463 = ~n9480 & n37462 ;
  assign n37464 = \b[39]  & n13794 ;
  assign n37465 = n13792 & n37464 ;
  assign n37466 = ~\a[48]  & \b[40]  ;
  assign n37467 = n13117 & n37466 ;
  assign n37468 = ~n37465 & ~n37467 ;
  assign n37469 = \b[41]  & n13123 ;
  assign n37470 = \a[48]  & \b[40]  ;
  assign n37471 = n13786 & n37470 ;
  assign n37472 = \a[50]  & ~n37471 ;
  assign n37473 = ~n37469 & n37472 ;
  assign n37474 = n37468 & n37473 ;
  assign n37475 = ~n37463 & n37474 ;
  assign n37476 = ~n37469 & ~n37471 ;
  assign n37477 = n37468 & n37476 ;
  assign n37478 = ~n37463 & n37477 ;
  assign n37479 = ~\a[50]  & ~n37478 ;
  assign n37480 = ~n37475 & ~n37479 ;
  assign n37481 = ~n37102 & n37126 ;
  assign n37482 = ~n37101 & ~n37481 ;
  assign n37483 = ~n6610 & n16655 ;
  assign n37484 = ~n6608 & n37483 ;
  assign n37485 = \b[33]  & n17308 ;
  assign n37486 = n17305 & n37485 ;
  assign n37487 = ~\a[54]  & \b[34]  ;
  assign n37488 = n16647 & n37487 ;
  assign n37489 = ~n37486 & ~n37488 ;
  assign n37490 = \b[35]  & n16653 ;
  assign n37491 = \a[54]  & \b[34]  ;
  assign n37492 = n16644 & n37491 ;
  assign n37493 = \a[56]  & ~n37492 ;
  assign n37494 = ~n37490 & n37493 ;
  assign n37495 = n37489 & n37494 ;
  assign n37496 = ~n37484 & n37495 ;
  assign n37497 = ~n37490 & ~n37492 ;
  assign n37498 = n37489 & n37497 ;
  assign n37499 = ~n37484 & n37498 ;
  assign n37500 = ~\a[56]  & ~n37499 ;
  assign n37501 = ~n37496 & ~n37500 ;
  assign n37502 = n5810 & n18516 ;
  assign n37503 = ~n5807 & n37502 ;
  assign n37504 = ~n5457 & ~n5810 ;
  assign n37505 = n18516 & n37504 ;
  assign n37506 = ~n5806 & n37505 ;
  assign n37507 = \b[32]  & n18514 ;
  assign n37508 = \a[56]  & \b[31]  ;
  assign n37509 = n19181 & n37508 ;
  assign n37510 = ~\a[57]  & \b[31]  ;
  assign n37511 = n18508 & n37510 ;
  assign n37512 = ~n37509 & ~n37511 ;
  assign n37513 = ~n37507 & n37512 ;
  assign n37514 = \b[30]  & n19183 ;
  assign n37515 = n19180 & n37514 ;
  assign n37516 = \a[59]  & ~n37515 ;
  assign n37517 = n37513 & n37516 ;
  assign n37518 = ~n37506 & n37517 ;
  assign n37519 = ~n37503 & n37518 ;
  assign n37520 = n37513 & ~n37515 ;
  assign n37521 = ~n37506 & n37520 ;
  assign n37522 = ~n37503 & n37521 ;
  assign n37523 = ~\a[59]  & ~n37522 ;
  assign n37524 = ~n37519 & ~n37523 ;
  assign n37525 = ~n4502 & n20521 ;
  assign n37526 = ~n4500 & n37525 ;
  assign n37527 = \b[29]  & n20519 ;
  assign n37528 = \a[60]  & \b[28]  ;
  assign n37529 = n20510 & n37528 ;
  assign n37530 = ~n37527 & ~n37529 ;
  assign n37531 = \b[27]  & n21315 ;
  assign n37532 = n21312 & n37531 ;
  assign n37533 = ~\a[60]  & \b[28]  ;
  assign n37534 = n20513 & n37533 ;
  assign n37535 = ~n37532 & ~n37534 ;
  assign n37536 = n37530 & n37535 ;
  assign n37537 = ~n37526 & n37536 ;
  assign n37538 = ~\a[62]  & ~n37537 ;
  assign n37539 = \b[26]  & n21958 ;
  assign n37540 = \b[25]  & n21957 ;
  assign n37541 = ~n37539 & ~n37540 ;
  assign n37542 = ~n37018 & n37541 ;
  assign n37543 = n37018 & ~n37541 ;
  assign n37544 = ~n37542 & ~n37543 ;
  assign n37545 = \a[62]  & n37536 ;
  assign n37546 = ~n37526 & n37545 ;
  assign n37547 = ~n37544 & ~n37546 ;
  assign n37548 = ~n37538 & n37547 ;
  assign n37549 = ~\a[62]  & n37544 ;
  assign n37550 = ~n37537 & n37549 ;
  assign n37551 = ~n37032 & ~n37036 ;
  assign n37552 = ~n37024 & n37551 ;
  assign n37553 = \a[62]  & n37544 ;
  assign n37554 = n37536 & n37553 ;
  assign n37555 = ~n37526 & n37554 ;
  assign n37556 = ~n37552 & ~n37555 ;
  assign n37557 = ~n37550 & n37556 ;
  assign n37558 = ~n37548 & n37557 ;
  assign n37559 = ~n37550 & ~n37555 ;
  assign n37560 = ~n37548 & n37559 ;
  assign n37561 = n37552 & ~n37560 ;
  assign n37562 = ~n37558 & ~n37561 ;
  assign n37563 = n37524 & n37562 ;
  assign n37564 = ~n37524 & ~n37562 ;
  assign n37565 = ~n37563 & ~n37564 ;
  assign n37566 = ~n37044 & n37068 ;
  assign n37567 = ~n37063 & n37566 ;
  assign n37568 = ~n37045 & ~n37567 ;
  assign n37569 = ~n37565 & n37568 ;
  assign n37570 = n37565 & ~n37568 ;
  assign n37571 = ~n37569 & ~n37570 ;
  assign n37572 = n37501 & n37571 ;
  assign n37573 = ~n37501 & ~n37571 ;
  assign n37574 = ~n37572 & ~n37573 ;
  assign n37575 = ~n37074 & n37097 ;
  assign n37576 = ~n37073 & ~n37575 ;
  assign n37577 = n8175 & n14793 ;
  assign n37578 = ~n8172 & n37577 ;
  assign n37579 = n14793 & n25622 ;
  assign n37580 = ~n8171 & n37579 ;
  assign n37581 = \b[36]  & n15517 ;
  assign n37582 = n15514 & n37581 ;
  assign n37583 = ~\a[51]  & \b[37]  ;
  assign n37584 = n14785 & n37583 ;
  assign n37585 = ~n37582 & ~n37584 ;
  assign n37586 = \b[38]  & n14791 ;
  assign n37587 = \a[51]  & \b[37]  ;
  assign n37588 = n14782 & n37587 ;
  assign n37589 = \a[53]  & ~n37588 ;
  assign n37590 = ~n37586 & n37589 ;
  assign n37591 = n37585 & n37590 ;
  assign n37592 = ~n37580 & n37591 ;
  assign n37593 = ~n37578 & n37592 ;
  assign n37594 = ~n37586 & ~n37588 ;
  assign n37595 = n37585 & n37594 ;
  assign n37596 = ~n37580 & n37595 ;
  assign n37597 = ~n37578 & n37596 ;
  assign n37598 = ~\a[53]  & ~n37597 ;
  assign n37599 = ~n37593 & ~n37598 ;
  assign n37600 = ~n37576 & ~n37599 ;
  assign n37601 = ~n37574 & n37600 ;
  assign n37602 = n37576 & ~n37599 ;
  assign n37603 = n37574 & n37602 ;
  assign n37604 = ~n37601 & ~n37603 ;
  assign n37605 = ~n37576 & n37599 ;
  assign n37606 = n37574 & n37605 ;
  assign n37607 = n37576 & n37599 ;
  assign n37608 = ~n37574 & n37607 ;
  assign n37609 = ~n37606 & ~n37608 ;
  assign n37610 = n37604 & n37609 ;
  assign n37611 = n37482 & n37610 ;
  assign n37612 = ~n37482 & ~n37610 ;
  assign n37613 = ~n37611 & ~n37612 ;
  assign n37614 = n37480 & n37613 ;
  assign n37615 = ~n37480 & ~n37613 ;
  assign n37616 = ~n37614 & ~n37615 ;
  assign n37617 = ~n10889 & ~n10988 ;
  assign n37618 = ~n11569 & n37617 ;
  assign n37619 = n10886 & n37618 ;
  assign n37620 = n10889 & ~n10988 ;
  assign n37621 = ~n11569 & n37620 ;
  assign n37622 = ~n10886 & n37621 ;
  assign n37623 = ~n37619 & ~n37622 ;
  assign n37624 = \b[42]  & n12159 ;
  assign n37625 = n12156 & n37624 ;
  assign n37626 = ~\a[45]  & \b[43]  ;
  assign n37627 = n11564 & n37626 ;
  assign n37628 = ~n37625 & ~n37627 ;
  assign n37629 = \b[44]  & n11570 ;
  assign n37630 = \a[45]  & \b[43]  ;
  assign n37631 = n11561 & n37630 ;
  assign n37632 = \a[47]  & ~n37631 ;
  assign n37633 = ~n37629 & n37632 ;
  assign n37634 = n37628 & n37633 ;
  assign n37635 = n37623 & n37634 ;
  assign n37636 = ~n37629 & ~n37631 ;
  assign n37637 = n37628 & n37636 ;
  assign n37638 = n37623 & n37637 ;
  assign n37639 = ~\a[47]  & ~n37638 ;
  assign n37640 = ~n37635 & ~n37639 ;
  assign n37641 = n37129 & n37153 ;
  assign n37642 = n37158 & ~n37641 ;
  assign n37643 = ~n37640 & n37642 ;
  assign n37644 = ~n37616 & n37643 ;
  assign n37645 = ~n37640 & ~n37642 ;
  assign n37646 = n37616 & n37645 ;
  assign n37647 = ~n37644 & ~n37646 ;
  assign n37648 = n37640 & ~n37642 ;
  assign n37649 = ~n37616 & n37648 ;
  assign n37650 = n37640 & n37642 ;
  assign n37651 = n37616 & n37650 ;
  assign n37652 = ~n37649 & ~n37651 ;
  assign n37653 = n37647 & n37652 ;
  assign n37654 = ~n37165 & n37191 ;
  assign n37655 = ~n37166 & ~n37654 ;
  assign n37656 = n10082 & ~n12438 ;
  assign n37657 = ~n12436 & n37656 ;
  assign n37658 = \b[47]  & n10080 ;
  assign n37659 = \a[41]  & \b[46]  ;
  assign n37660 = n10679 & n37659 ;
  assign n37661 = ~\a[42]  & \b[46]  ;
  assign n37662 = n10074 & n37661 ;
  assign n37663 = ~n37660 & ~n37662 ;
  assign n37664 = ~n37658 & n37663 ;
  assign n37665 = \b[45]  & n10681 ;
  assign n37666 = n10678 & n37665 ;
  assign n37667 = \a[44]  & ~n37666 ;
  assign n37668 = n37664 & n37667 ;
  assign n37669 = ~n37657 & n37668 ;
  assign n37670 = n37664 & ~n37666 ;
  assign n37671 = ~n37657 & n37670 ;
  assign n37672 = ~\a[44]  & ~n37671 ;
  assign n37673 = ~n37669 & ~n37672 ;
  assign n37674 = ~n37655 & ~n37673 ;
  assign n37675 = n37653 & n37674 ;
  assign n37676 = n37655 & ~n37673 ;
  assign n37677 = ~n37653 & n37676 ;
  assign n37678 = ~n37675 & ~n37677 ;
  assign n37679 = ~n37655 & n37673 ;
  assign n37680 = ~n37653 & n37679 ;
  assign n37681 = n37655 & n37673 ;
  assign n37682 = n37653 & n37681 ;
  assign n37683 = ~n37680 & ~n37682 ;
  assign n37684 = n37678 & n37683 ;
  assign n37685 = ~n37194 & ~n37196 ;
  assign n37686 = ~n37191 & n37217 ;
  assign n37687 = n37167 & n37686 ;
  assign n37688 = n37191 & n37217 ;
  assign n37689 = ~n37167 & n37688 ;
  assign n37690 = ~n37687 & ~n37689 ;
  assign n37691 = ~n37218 & n37690 ;
  assign n37692 = ~n37685 & n37691 ;
  assign n37693 = n8759 & n14052 ;
  assign n37694 = ~n14049 & n37693 ;
  assign n37695 = n8759 & n15779 ;
  assign n37696 = ~n14048 & n37695 ;
  assign n37697 = \b[48]  & n9301 ;
  assign n37698 = n9298 & n37697 ;
  assign n37699 = ~\a[39]  & \b[49]  ;
  assign n37700 = n8751 & n37699 ;
  assign n37701 = ~n37698 & ~n37700 ;
  assign n37702 = \b[50]  & n8757 ;
  assign n37703 = \a[39]  & \b[49]  ;
  assign n37704 = n8748 & n37703 ;
  assign n37705 = \a[41]  & ~n37704 ;
  assign n37706 = ~n37702 & n37705 ;
  assign n37707 = n37701 & n37706 ;
  assign n37708 = ~n37696 & n37707 ;
  assign n37709 = ~n37694 & n37708 ;
  assign n37710 = ~n37702 & ~n37704 ;
  assign n37711 = n37701 & n37710 ;
  assign n37712 = ~n37696 & n37711 ;
  assign n37713 = ~n37694 & n37712 ;
  assign n37714 = ~\a[41]  & ~n37713 ;
  assign n37715 = ~n37709 & ~n37714 ;
  assign n37716 = ~n37692 & n37715 ;
  assign n37717 = ~n37684 & n37716 ;
  assign n37718 = n37692 & n37715 ;
  assign n37719 = n37684 & n37718 ;
  assign n37720 = ~n37717 & ~n37719 ;
  assign n37721 = ~n37692 & ~n37715 ;
  assign n37722 = n37684 & n37721 ;
  assign n37723 = n37692 & ~n37715 ;
  assign n37724 = ~n37684 & n37723 ;
  assign n37725 = ~n37722 & ~n37724 ;
  assign n37726 = n37720 & n37725 ;
  assign n37727 = ~n37228 & ~n37230 ;
  assign n37728 = n37228 & n37230 ;
  assign n37729 = n37249 & ~n37728 ;
  assign n37730 = ~n37727 & ~n37729 ;
  assign n37731 = n37726 & n37730 ;
  assign n37732 = ~n37726 & ~n37730 ;
  assign n37733 = ~n37731 & ~n37732 ;
  assign n37734 = n37461 & n37733 ;
  assign n37735 = ~n37461 & ~n37733 ;
  assign n37736 = ~n37734 & ~n37735 ;
  assign n37737 = ~n5952 & ~n16441 ;
  assign n37738 = ~n17647 & n37737 ;
  assign n37739 = ~n17643 & n37738 ;
  assign n37740 = ~n6306 & n37739 ;
  assign n37741 = n6309 & n17647 ;
  assign n37742 = ~n17644 & n37741 ;
  assign n37743 = ~n37740 & ~n37742 ;
  assign n37744 = \b[54]  & n6778 ;
  assign n37745 = n6775 & n37744 ;
  assign n37746 = ~\a[33]  & \b[55]  ;
  assign n37747 = n6301 & n37746 ;
  assign n37748 = ~n37745 & ~n37747 ;
  assign n37749 = \b[56]  & n6307 ;
  assign n37750 = \a[33]  & \b[55]  ;
  assign n37751 = n6298 & n37750 ;
  assign n37752 = \a[35]  & ~n37751 ;
  assign n37753 = ~n37749 & n37752 ;
  assign n37754 = n37748 & n37753 ;
  assign n37755 = n37743 & n37754 ;
  assign n37756 = ~n37749 & ~n37751 ;
  assign n37757 = n37748 & n37756 ;
  assign n37758 = n37743 & n37757 ;
  assign n37759 = ~\a[35]  & ~n37758 ;
  assign n37760 = ~n37755 & ~n37759 ;
  assign n37761 = ~n37260 & ~n37262 ;
  assign n37762 = n37260 & n37262 ;
  assign n37763 = n37286 & ~n37762 ;
  assign n37764 = ~n37761 & ~n37763 ;
  assign n37765 = n37760 & ~n37764 ;
  assign n37766 = ~n37736 & n37765 ;
  assign n37767 = n37760 & n37764 ;
  assign n37768 = n37736 & n37767 ;
  assign n37769 = ~n37766 & ~n37768 ;
  assign n37770 = ~n37760 & ~n37764 ;
  assign n37771 = n37736 & n37770 ;
  assign n37772 = ~n37760 & n37764 ;
  assign n37773 = ~n37736 & n37772 ;
  assign n37774 = ~n37771 & ~n37773 ;
  assign n37775 = n37769 & n37774 ;
  assign n37776 = n37442 & ~n37775 ;
  assign n37777 = ~n37442 & n37775 ;
  assign n37778 = ~n37776 & ~n37777 ;
  assign n37779 = ~n37413 & ~n37778 ;
  assign n37780 = n37413 & n37778 ;
  assign n37781 = ~n37779 & ~n37780 ;
  assign n37782 = n37308 & ~n37335 ;
  assign n37783 = ~n37327 & ~n37782 ;
  assign n37784 = \b[63]  & n3402 ;
  assign n37785 = ~n21694 & n37784 ;
  assign n37786 = ~n23171 & n37785 ;
  assign n37787 = \a[23]  & \a[25]  ;
  assign n37788 = \a[24]  & ~\a[26]  ;
  assign n37789 = n37787 & n37788 ;
  assign n37790 = ~\a[23]  & ~\a[25]  ;
  assign n37791 = ~\a[24]  & \a[26]  ;
  assign n37792 = n37790 & n37791 ;
  assign n37793 = ~n37789 & ~n37792 ;
  assign n37794 = \b[63]  & ~n37793 ;
  assign n37795 = \a[26]  & ~n37794 ;
  assign n37796 = ~n37786 & n37795 ;
  assign n37797 = ~n37786 & ~n37794 ;
  assign n37798 = ~\a[26]  & ~n37797 ;
  assign n37799 = ~n37796 & ~n37798 ;
  assign n37800 = ~n37783 & ~n37799 ;
  assign n37801 = ~n37327 & n37799 ;
  assign n37802 = ~n37782 & n37801 ;
  assign n37803 = ~n37800 & ~n37802 ;
  assign n37804 = n37781 & n37803 ;
  assign n37805 = ~n37781 & ~n37803 ;
  assign n37806 = ~n37804 & ~n37805 ;
  assign n37807 = n37385 & n37806 ;
  assign n37808 = ~n37385 & ~n37806 ;
  assign n37809 = ~n37807 & ~n37808 ;
  assign n37810 = ~n37376 & n37809 ;
  assign n37811 = ~n37383 & n37810 ;
  assign n37812 = ~n37376 & ~n37383 ;
  assign n37813 = ~n37809 & ~n37812 ;
  assign n37814 = ~n37811 & ~n37813 ;
  assign n37815 = ~n37800 & n37802 ;
  assign n37816 = ~n37781 & ~n37800 ;
  assign n37817 = ~n37815 & ~n37816 ;
  assign n37818 = ~n37408 & n37778 ;
  assign n37819 = n37388 & n37402 ;
  assign n37820 = \a[29]  & n37401 ;
  assign n37821 = n37388 & n37820 ;
  assign n37822 = ~n37819 & ~n37821 ;
  assign n37823 = ~n37818 & n37822 ;
  assign n37824 = n4249 & ~n22461 ;
  assign n37825 = ~n22459 & n37824 ;
  assign n37826 = \b[61]  & n4647 ;
  assign n37827 = n4644 & n37826 ;
  assign n37828 = ~\a[27]  & \b[62]  ;
  assign n37829 = n4241 & n37828 ;
  assign n37830 = ~n37827 & ~n37829 ;
  assign n37831 = \b[63]  & n4247 ;
  assign n37832 = \a[27]  & \b[62]  ;
  assign n37833 = n4238 & n37832 ;
  assign n37834 = \a[29]  & ~n37833 ;
  assign n37835 = ~n37831 & n37834 ;
  assign n37836 = n37830 & n37835 ;
  assign n37837 = ~n37825 & n37836 ;
  assign n37838 = ~n37831 & ~n37833 ;
  assign n37839 = n37830 & n37838 ;
  assign n37840 = ~n37825 & n37839 ;
  assign n37841 = ~\a[29]  & ~n37840 ;
  assign n37842 = ~n37837 & ~n37841 ;
  assign n37843 = ~n37823 & ~n37842 ;
  assign n37844 = n37823 & n37842 ;
  assign n37845 = ~n37843 & ~n37844 ;
  assign n37846 = n5211 & n20260 ;
  assign n37847 = ~n20257 & n37846 ;
  assign n37848 = n5211 & ~n20260 ;
  assign n37849 = ~n19545 & n37848 ;
  assign n37850 = ~n20256 & n37849 ;
  assign n37851 = \b[58]  & n5595 ;
  assign n37852 = n5592 & n37851 ;
  assign n37853 = ~\a[30]  & \b[59]  ;
  assign n37854 = n5203 & n37853 ;
  assign n37855 = ~n37852 & ~n37854 ;
  assign n37856 = \b[60]  & n5209 ;
  assign n37857 = \a[30]  & \b[59]  ;
  assign n37858 = n5200 & n37857 ;
  assign n37859 = \a[32]  & ~n37858 ;
  assign n37860 = ~n37856 & n37859 ;
  assign n37861 = n37855 & n37860 ;
  assign n37862 = ~n37850 & n37861 ;
  assign n37863 = ~n37847 & n37862 ;
  assign n37864 = ~n37856 & ~n37858 ;
  assign n37865 = n37855 & n37864 ;
  assign n37866 = ~n37850 & n37865 ;
  assign n37867 = ~n37847 & n37866 ;
  assign n37868 = ~\a[32]  & ~n37867 ;
  assign n37869 = ~n37863 & ~n37868 ;
  assign n37870 = n37441 & n37775 ;
  assign n37871 = ~n37434 & ~n37870 ;
  assign n37872 = ~n37542 & ~n37555 ;
  assign n37873 = ~n37550 & n37872 ;
  assign n37874 = ~\a[26]  & \b[26]  ;
  assign n37875 = n21957 & n37874 ;
  assign n37876 = ~\a[26]  & \b[27]  ;
  assign n37877 = n21958 & n37876 ;
  assign n37878 = ~n37875 & ~n37877 ;
  assign n37879 = \b[27]  & n21958 ;
  assign n37880 = \b[26]  & n21957 ;
  assign n37881 = \a[26]  & ~n37880 ;
  assign n37882 = ~n37879 & n37881 ;
  assign n37883 = n37878 & ~n37882 ;
  assign n37884 = ~n37541 & ~n37883 ;
  assign n37885 = n37541 & n37883 ;
  assign n37886 = ~n37884 & ~n37885 ;
  assign n37887 = ~n37873 & ~n37886 ;
  assign n37888 = n37873 & n37886 ;
  assign n37889 = ~n5105 & ~n19861 ;
  assign n37890 = ~n20518 & n37889 ;
  assign n37891 = n5102 & n37890 ;
  assign n37892 = n5105 & ~n19861 ;
  assign n37893 = ~n20518 & n37892 ;
  assign n37894 = ~n5102 & n37893 ;
  assign n37895 = ~n37891 & ~n37894 ;
  assign n37896 = \b[28]  & n21315 ;
  assign n37897 = n21312 & n37896 ;
  assign n37898 = ~\a[60]  & \b[29]  ;
  assign n37899 = n20513 & n37898 ;
  assign n37900 = ~n37897 & ~n37899 ;
  assign n37901 = \b[30]  & n20519 ;
  assign n37902 = \a[60]  & \b[29]  ;
  assign n37903 = n20510 & n37902 ;
  assign n37904 = \a[62]  & ~n37903 ;
  assign n37905 = ~n37901 & n37904 ;
  assign n37906 = n37900 & n37905 ;
  assign n37907 = n37895 & n37906 ;
  assign n37908 = ~n37901 & ~n37903 ;
  assign n37909 = n37900 & n37908 ;
  assign n37910 = n37895 & n37909 ;
  assign n37911 = ~\a[62]  & ~n37910 ;
  assign n37912 = ~n37907 & ~n37911 ;
  assign n37913 = ~n37888 & ~n37912 ;
  assign n37914 = ~n37887 & n37913 ;
  assign n37915 = ~n37887 & ~n37888 ;
  assign n37916 = n37912 & ~n37915 ;
  assign n37917 = ~n37914 & ~n37916 ;
  assign n37918 = ~n5855 & n18516 ;
  assign n37919 = ~n5853 & n37918 ;
  assign n37920 = \b[31]  & n19183 ;
  assign n37921 = n19180 & n37920 ;
  assign n37922 = \b[33]  & n18514 ;
  assign n37923 = \a[56]  & \b[32]  ;
  assign n37924 = n19181 & n37923 ;
  assign n37925 = ~\a[57]  & \b[32]  ;
  assign n37926 = n18508 & n37925 ;
  assign n37927 = ~n37924 & ~n37926 ;
  assign n37928 = ~n37922 & n37927 ;
  assign n37929 = ~n37921 & n37928 ;
  assign n37930 = ~\a[59]  & n37929 ;
  assign n37931 = ~n37919 & n37930 ;
  assign n37932 = ~n37919 & n37929 ;
  assign n37933 = \a[59]  & ~n37932 ;
  assign n37934 = ~n37931 & ~n37933 ;
  assign n37935 = n37524 & ~n37558 ;
  assign n37936 = ~n37561 & ~n37935 ;
  assign n37937 = ~n37934 & ~n37936 ;
  assign n37938 = n37934 & n37936 ;
  assign n37939 = ~n37937 & ~n37938 ;
  assign n37940 = ~n37917 & ~n37939 ;
  assign n37941 = n37917 & n37939 ;
  assign n37942 = ~n37940 & ~n37941 ;
  assign n37943 = n7337 & n16655 ;
  assign n37944 = ~n7334 & n37943 ;
  assign n37945 = ~n16016 & ~n16652 ;
  assign n37946 = ~n6605 & ~n7337 ;
  assign n37947 = n37945 & n37946 ;
  assign n37948 = ~n7333 & n37947 ;
  assign n37949 = \b[34]  & n17308 ;
  assign n37950 = n17305 & n37949 ;
  assign n37951 = ~\a[54]  & \b[35]  ;
  assign n37952 = n16647 & n37951 ;
  assign n37953 = ~n37950 & ~n37952 ;
  assign n37954 = \b[36]  & n16653 ;
  assign n37955 = \a[54]  & \b[35]  ;
  assign n37956 = n16644 & n37955 ;
  assign n37957 = \a[56]  & ~n37956 ;
  assign n37958 = ~n37954 & n37957 ;
  assign n37959 = n37953 & n37958 ;
  assign n37960 = ~n37948 & n37959 ;
  assign n37961 = ~n37944 & n37960 ;
  assign n37962 = ~n37954 & ~n37956 ;
  assign n37963 = n37953 & n37962 ;
  assign n37964 = ~n37948 & n37963 ;
  assign n37965 = ~n37944 & n37964 ;
  assign n37966 = ~\a[56]  & ~n37965 ;
  assign n37967 = ~n37961 & ~n37966 ;
  assign n37968 = n37942 & ~n37967 ;
  assign n37969 = ~n37942 & n37967 ;
  assign n37970 = ~n37968 & ~n37969 ;
  assign n37971 = n37501 & ~n37569 ;
  assign n37972 = ~n37570 & ~n37971 ;
  assign n37973 = ~n8599 & n14793 ;
  assign n37974 = ~n8174 & n14793 ;
  assign n37975 = ~n8595 & n37974 ;
  assign n37976 = ~n37973 & ~n37975 ;
  assign n37977 = ~n8602 & ~n37976 ;
  assign n37978 = \b[37]  & n15517 ;
  assign n37979 = n15514 & n37978 ;
  assign n37980 = ~\a[51]  & \b[38]  ;
  assign n37981 = n14785 & n37980 ;
  assign n37982 = ~n37979 & ~n37981 ;
  assign n37983 = \b[39]  & n14791 ;
  assign n37984 = \a[51]  & \b[38]  ;
  assign n37985 = n14782 & n37984 ;
  assign n37986 = \a[53]  & ~n37985 ;
  assign n37987 = ~n37983 & n37986 ;
  assign n37988 = n37982 & n37987 ;
  assign n37989 = ~n37977 & n37988 ;
  assign n37990 = ~n37983 & ~n37985 ;
  assign n37991 = n37982 & n37990 ;
  assign n37992 = ~\a[53]  & ~n37991 ;
  assign n37993 = ~\a[53]  & ~n8602 ;
  assign n37994 = ~n37976 & n37993 ;
  assign n37995 = ~n37992 & ~n37994 ;
  assign n37996 = ~n37989 & n37995 ;
  assign n37997 = n37972 & ~n37996 ;
  assign n37998 = ~n37970 & n37997 ;
  assign n37999 = ~n37972 & ~n37996 ;
  assign n38000 = n37970 & n37999 ;
  assign n38001 = ~n37998 & ~n38000 ;
  assign n38002 = ~n37972 & n37996 ;
  assign n38003 = ~n37970 & n38002 ;
  assign n38004 = n37972 & n37996 ;
  assign n38005 = n37970 & n38004 ;
  assign n38006 = ~n38003 & ~n38005 ;
  assign n38007 = n38001 & n38006 ;
  assign n38008 = n37574 & ~n37576 ;
  assign n38009 = ~n37574 & n37576 ;
  assign n38010 = n37599 & ~n38009 ;
  assign n38011 = ~n38008 & ~n38010 ;
  assign n38012 = ~n38007 & ~n38011 ;
  assign n38013 = n38007 & n38011 ;
  assign n38014 = ~n38012 & ~n38013 ;
  assign n38015 = ~n9930 & ~n12606 ;
  assign n38016 = ~n13122 & n38015 ;
  assign n38017 = n9927 & n38016 ;
  assign n38018 = n9930 & ~n12606 ;
  assign n38019 = ~n13122 & n38018 ;
  assign n38020 = ~n9927 & n38019 ;
  assign n38021 = ~n38017 & ~n38020 ;
  assign n38022 = \b[40]  & n13794 ;
  assign n38023 = n13792 & n38022 ;
  assign n38024 = ~\a[48]  & \b[41]  ;
  assign n38025 = n13117 & n38024 ;
  assign n38026 = ~n38023 & ~n38025 ;
  assign n38027 = \b[42]  & n13123 ;
  assign n38028 = \a[48]  & \b[41]  ;
  assign n38029 = n13786 & n38028 ;
  assign n38030 = \a[50]  & ~n38029 ;
  assign n38031 = ~n38027 & n38030 ;
  assign n38032 = n38026 & n38031 ;
  assign n38033 = n38021 & n38032 ;
  assign n38034 = ~n38027 & ~n38029 ;
  assign n38035 = n38026 & n38034 ;
  assign n38036 = n38021 & n38035 ;
  assign n38037 = ~\a[50]  & ~n38036 ;
  assign n38038 = ~n38033 & ~n38037 ;
  assign n38039 = n38014 & ~n38038 ;
  assign n38040 = ~n38014 & n38038 ;
  assign n38041 = ~n38039 & ~n38040 ;
  assign n38042 = ~n11397 & n11572 ;
  assign n38043 = ~n11395 & n38042 ;
  assign n38044 = \b[43]  & n12159 ;
  assign n38045 = n12156 & n38044 ;
  assign n38046 = ~\a[45]  & \b[44]  ;
  assign n38047 = n11564 & n38046 ;
  assign n38048 = ~n38045 & ~n38047 ;
  assign n38049 = \b[45]  & n11570 ;
  assign n38050 = \a[45]  & \b[44]  ;
  assign n38051 = n11561 & n38050 ;
  assign n38052 = \a[47]  & ~n38051 ;
  assign n38053 = ~n38049 & n38052 ;
  assign n38054 = n38048 & n38053 ;
  assign n38055 = ~n38043 & n38054 ;
  assign n38056 = ~n38049 & ~n38051 ;
  assign n38057 = n38048 & n38056 ;
  assign n38058 = ~n38043 & n38057 ;
  assign n38059 = ~\a[47]  & ~n38058 ;
  assign n38060 = ~n38055 & ~n38059 ;
  assign n38061 = n37480 & ~n37611 ;
  assign n38062 = ~n37612 & ~n38061 ;
  assign n38063 = ~n38060 & ~n38062 ;
  assign n38064 = n38041 & n38063 ;
  assign n38065 = ~n38060 & n38062 ;
  assign n38066 = ~n38041 & n38065 ;
  assign n38067 = ~n38064 & ~n38066 ;
  assign n38068 = n38060 & ~n38062 ;
  assign n38069 = ~n38041 & n38068 ;
  assign n38070 = n38060 & n38062 ;
  assign n38071 = n38041 & n38070 ;
  assign n38072 = ~n38069 & ~n38071 ;
  assign n38073 = n38067 & n38072 ;
  assign n38074 = ~n37616 & ~n37642 ;
  assign n38075 = n37647 & ~n38074 ;
  assign n38076 = n10082 & n12478 ;
  assign n38077 = ~n12475 & n38076 ;
  assign n38078 = n10082 & n28668 ;
  assign n38079 = ~n12474 & n38078 ;
  assign n38080 = \b[46]  & n10681 ;
  assign n38081 = n10678 & n38080 ;
  assign n38082 = \b[48]  & n10080 ;
  assign n38083 = \a[41]  & \b[47]  ;
  assign n38084 = n10679 & n38083 ;
  assign n38085 = ~\a[42]  & \b[47]  ;
  assign n38086 = n10074 & n38085 ;
  assign n38087 = ~n38084 & ~n38086 ;
  assign n38088 = ~n38082 & n38087 ;
  assign n38089 = ~n38081 & n38088 ;
  assign n38090 = ~n38079 & n38089 ;
  assign n38091 = ~n38077 & n38090 ;
  assign n38092 = ~\a[44]  & ~n38091 ;
  assign n38093 = \a[44]  & n38089 ;
  assign n38094 = ~n38079 & n38093 ;
  assign n38095 = ~n38077 & n38094 ;
  assign n38096 = ~n38092 & ~n38095 ;
  assign n38097 = ~n38075 & ~n38096 ;
  assign n38098 = ~n38073 & n38097 ;
  assign n38099 = n38075 & ~n38096 ;
  assign n38100 = n38073 & n38099 ;
  assign n38101 = ~n38098 & ~n38100 ;
  assign n38102 = n38075 & n38096 ;
  assign n38103 = ~n38073 & n38102 ;
  assign n38104 = ~n38075 & n38096 ;
  assign n38105 = n38073 & n38104 ;
  assign n38106 = ~n38103 & ~n38105 ;
  assign n38107 = n38101 & n38106 ;
  assign n38108 = ~n37653 & ~n37655 ;
  assign n38109 = n37653 & n37655 ;
  assign n38110 = n37673 & ~n38109 ;
  assign n38111 = ~n38108 & ~n38110 ;
  assign n38112 = n8759 & ~n14098 ;
  assign n38113 = ~n14096 & n38112 ;
  assign n38114 = \b[49]  & n9301 ;
  assign n38115 = n9298 & n38114 ;
  assign n38116 = ~\a[39]  & \b[50]  ;
  assign n38117 = n8751 & n38116 ;
  assign n38118 = ~n38115 & ~n38117 ;
  assign n38119 = \b[51]  & n8757 ;
  assign n38120 = \a[39]  & \b[50]  ;
  assign n38121 = n8748 & n38120 ;
  assign n38122 = \a[41]  & ~n38121 ;
  assign n38123 = ~n38119 & n38122 ;
  assign n38124 = n38118 & n38123 ;
  assign n38125 = ~n38113 & n38124 ;
  assign n38126 = ~n38119 & ~n38121 ;
  assign n38127 = n38118 & n38126 ;
  assign n38128 = ~n38113 & n38127 ;
  assign n38129 = ~\a[41]  & ~n38128 ;
  assign n38130 = ~n38125 & ~n38129 ;
  assign n38131 = ~n38111 & n38130 ;
  assign n38132 = ~n38107 & n38131 ;
  assign n38133 = n38111 & n38130 ;
  assign n38134 = n38107 & n38133 ;
  assign n38135 = ~n38132 & ~n38134 ;
  assign n38136 = ~n38111 & ~n38130 ;
  assign n38137 = n38107 & n38136 ;
  assign n38138 = n38111 & ~n38130 ;
  assign n38139 = ~n38107 & n38138 ;
  assign n38140 = ~n38137 & ~n38139 ;
  assign n38141 = n38135 & n38140 ;
  assign n38142 = ~n15241 & ~n16398 ;
  assign n38143 = n7534 & n38142 ;
  assign n38144 = ~n16404 & n38143 ;
  assign n38145 = n7534 & n16398 ;
  assign n38146 = n15241 & n38145 ;
  assign n38147 = n16400 & n38145 ;
  assign n38148 = ~n15239 & n38147 ;
  assign n38149 = ~n38146 & ~n38148 ;
  assign n38150 = ~n38144 & n38149 ;
  assign n38151 = \b[52]  & n7973 ;
  assign n38152 = n7970 & n38151 ;
  assign n38153 = ~\a[36]  & \b[53]  ;
  assign n38154 = n7526 & n38153 ;
  assign n38155 = ~n38152 & ~n38154 ;
  assign n38156 = \b[54]  & n7532 ;
  assign n38157 = \a[36]  & \b[53]  ;
  assign n38158 = n17801 & n38157 ;
  assign n38159 = \a[38]  & ~n38158 ;
  assign n38160 = ~n38156 & n38159 ;
  assign n38161 = n38155 & n38160 ;
  assign n38162 = n38150 & n38161 ;
  assign n38163 = ~n38156 & ~n38158 ;
  assign n38164 = n38155 & n38163 ;
  assign n38165 = n38150 & n38164 ;
  assign n38166 = ~\a[38]  & ~n38165 ;
  assign n38167 = ~n38162 & ~n38166 ;
  assign n38168 = n37684 & n37692 ;
  assign n38169 = n37725 & ~n38168 ;
  assign n38170 = n38167 & n38169 ;
  assign n38171 = ~n38141 & n38170 ;
  assign n38172 = n38167 & ~n38169 ;
  assign n38173 = n38141 & n38172 ;
  assign n38174 = ~n38171 & ~n38173 ;
  assign n38175 = ~n38167 & ~n38169 ;
  assign n38176 = ~n38141 & n38175 ;
  assign n38177 = ~n38167 & n38169 ;
  assign n38178 = n38141 & n38177 ;
  assign n38179 = ~n38176 & ~n38178 ;
  assign n38180 = n38174 & n38179 ;
  assign n38181 = n37461 & ~n37731 ;
  assign n38182 = ~n37732 & ~n38181 ;
  assign n38183 = n6309 & ~n17690 ;
  assign n38184 = ~n17688 & n38183 ;
  assign n38185 = \b[57]  & n6307 ;
  assign n38186 = \a[33]  & \b[56]  ;
  assign n38187 = n6298 & n38186 ;
  assign n38188 = ~n38185 & ~n38187 ;
  assign n38189 = \b[55]  & n6778 ;
  assign n38190 = n6775 & n38189 ;
  assign n38191 = ~\a[33]  & \b[56]  ;
  assign n38192 = n6301 & n38191 ;
  assign n38193 = ~n38190 & ~n38192 ;
  assign n38194 = n38188 & n38193 ;
  assign n38195 = ~n38184 & n38194 ;
  assign n38196 = ~\a[35]  & ~n38195 ;
  assign n38197 = \a[35]  & n38194 ;
  assign n38198 = ~n38184 & n38197 ;
  assign n38199 = ~n38196 & ~n38198 ;
  assign n38200 = n38182 & ~n38199 ;
  assign n38201 = ~n38180 & n38200 ;
  assign n38202 = ~n38182 & ~n38199 ;
  assign n38203 = n38180 & n38202 ;
  assign n38204 = ~n38201 & ~n38203 ;
  assign n38205 = ~n38182 & n38199 ;
  assign n38206 = ~n38180 & n38205 ;
  assign n38207 = n38182 & n38199 ;
  assign n38208 = n38180 & n38207 ;
  assign n38209 = ~n38206 & ~n38208 ;
  assign n38210 = n38204 & n38209 ;
  assign n38211 = n37736 & ~n37764 ;
  assign n38212 = ~n37736 & n37764 ;
  assign n38213 = n37760 & ~n38212 ;
  assign n38214 = ~n38211 & ~n38213 ;
  assign n38215 = ~n38210 & ~n38214 ;
  assign n38216 = n38210 & n38214 ;
  assign n38217 = ~n38215 & ~n38216 ;
  assign n38218 = n37871 & ~n38217 ;
  assign n38219 = ~n37871 & n38217 ;
  assign n38220 = ~n38218 & ~n38219 ;
  assign n38221 = ~n37869 & ~n38220 ;
  assign n38222 = n37869 & n38220 ;
  assign n38223 = ~n38221 & ~n38222 ;
  assign n38224 = n37845 & n38223 ;
  assign n38225 = ~n37845 & ~n38223 ;
  assign n38226 = ~n38224 & ~n38225 ;
  assign n38227 = ~n37817 & ~n38226 ;
  assign n38228 = n37817 & n38226 ;
  assign n38229 = ~n38227 & ~n38228 ;
  assign n38230 = n37807 & n38229 ;
  assign n38231 = n37810 & n38229 ;
  assign n38232 = ~n37383 & n38231 ;
  assign n38233 = ~n38230 & ~n38232 ;
  assign n38234 = ~n37807 & ~n38229 ;
  assign n38235 = ~n37811 & n38234 ;
  assign n38236 = n38233 & ~n38235 ;
  assign n38237 = ~n37843 & ~n38223 ;
  assign n38238 = ~n37844 & ~n38237 ;
  assign n38239 = n4249 & ~n22458 ;
  assign n38240 = ~n23173 & n38239 ;
  assign n38241 = \b[62]  & n4647 ;
  assign n38242 = n4644 & n38241 ;
  assign n38243 = \a[27]  & \b[63]  ;
  assign n38244 = n4238 & n38243 ;
  assign n38245 = ~\a[27]  & \b[63]  ;
  assign n38246 = n4241 & n38245 ;
  assign n38247 = \a[29]  & ~n38246 ;
  assign n38248 = ~n38244 & n38247 ;
  assign n38249 = ~n38242 & n38248 ;
  assign n38250 = ~n38240 & n38249 ;
  assign n38251 = ~n38244 & ~n38246 ;
  assign n38252 = ~n38242 & n38251 ;
  assign n38253 = ~n38240 & n38252 ;
  assign n38254 = ~\a[29]  & ~n38253 ;
  assign n38255 = ~n38250 & ~n38254 ;
  assign n38256 = n37869 & ~n37871 ;
  assign n38257 = ~n37434 & ~n37869 ;
  assign n38258 = ~n37870 & n38257 ;
  assign n38259 = ~n38217 & ~n38258 ;
  assign n38260 = ~n38256 & ~n38259 ;
  assign n38261 = ~n38255 & n38260 ;
  assign n38262 = n38255 & ~n38260 ;
  assign n38263 = ~n38261 & ~n38262 ;
  assign n38264 = n5211 & ~n20971 ;
  assign n38265 = ~n20969 & n38264 ;
  assign n38266 = \b[61]  & n5209 ;
  assign n38267 = \a[30]  & \b[60]  ;
  assign n38268 = n5200 & n38267 ;
  assign n38269 = ~n38266 & ~n38268 ;
  assign n38270 = \b[59]  & n5595 ;
  assign n38271 = n5592 & n38270 ;
  assign n38272 = ~\a[30]  & \b[60]  ;
  assign n38273 = n5203 & n38272 ;
  assign n38274 = ~n38271 & ~n38273 ;
  assign n38275 = n38269 & n38274 ;
  assign n38276 = ~n38265 & n38275 ;
  assign n38277 = ~\a[32]  & ~n38276 ;
  assign n38278 = \a[32]  & n38275 ;
  assign n38279 = ~n38265 & n38278 ;
  assign n38280 = ~n38209 & ~n38279 ;
  assign n38281 = n38204 & ~n38279 ;
  assign n38282 = ~n38214 & n38281 ;
  assign n38283 = ~n38280 & ~n38282 ;
  assign n38284 = ~n38277 & ~n38283 ;
  assign n38285 = n38204 & ~n38214 ;
  assign n38286 = ~n38277 & ~n38279 ;
  assign n38287 = n38209 & ~n38286 ;
  assign n38288 = ~n38285 & n38287 ;
  assign n38289 = ~n38039 & ~n38062 ;
  assign n38290 = ~n38040 & ~n38289 ;
  assign n38291 = n9044 & n14793 ;
  assign n38292 = ~n9041 & n38291 ;
  assign n38293 = n14793 & n27054 ;
  assign n38294 = ~n9040 & n38293 ;
  assign n38295 = \b[38]  & n15517 ;
  assign n38296 = n15514 & n38295 ;
  assign n38297 = ~\a[51]  & \b[39]  ;
  assign n38298 = n14785 & n38297 ;
  assign n38299 = ~n38296 & ~n38298 ;
  assign n38300 = \b[40]  & n14791 ;
  assign n38301 = \a[51]  & \b[39]  ;
  assign n38302 = n14782 & n38301 ;
  assign n38303 = \a[53]  & ~n38302 ;
  assign n38304 = ~n38300 & n38303 ;
  assign n38305 = n38299 & n38304 ;
  assign n38306 = ~n38294 & n38305 ;
  assign n38307 = ~n38292 & n38306 ;
  assign n38308 = ~n38300 & ~n38302 ;
  assign n38309 = n38299 & n38308 ;
  assign n38310 = ~n38294 & n38309 ;
  assign n38311 = ~n38292 & n38310 ;
  assign n38312 = ~\a[53]  & ~n38311 ;
  assign n38313 = ~n38307 & ~n38312 ;
  assign n38314 = ~n37968 & ~n37972 ;
  assign n38315 = ~n37969 & ~n38314 ;
  assign n38316 = n37934 & ~n37936 ;
  assign n38317 = ~n37934 & n37936 ;
  assign n38318 = ~n38316 & ~n38317 ;
  assign n38319 = n37917 & ~n38318 ;
  assign n38320 = ~n37938 & ~n38319 ;
  assign n38321 = ~n7758 & n37945 ;
  assign n38322 = ~n7336 & n37945 ;
  assign n38323 = ~n7754 & n38322 ;
  assign n38324 = ~n38321 & ~n38323 ;
  assign n38325 = ~n7761 & ~n38324 ;
  assign n38326 = \b[35]  & n17308 ;
  assign n38327 = n17305 & n38326 ;
  assign n38328 = ~\a[54]  & \b[36]  ;
  assign n38329 = n16647 & n38328 ;
  assign n38330 = ~n38327 & ~n38329 ;
  assign n38331 = \b[37]  & n16653 ;
  assign n38332 = \a[54]  & \b[36]  ;
  assign n38333 = n16644 & n38332 ;
  assign n38334 = \a[56]  & ~n38333 ;
  assign n38335 = ~n38331 & n38334 ;
  assign n38336 = n38330 & n38335 ;
  assign n38337 = ~n38325 & n38336 ;
  assign n38338 = ~n38331 & ~n38333 ;
  assign n38339 = n38330 & n38338 ;
  assign n38340 = ~\a[56]  & ~n38339 ;
  assign n38341 = ~\a[56]  & ~n7761 ;
  assign n38342 = ~n38324 & n38341 ;
  assign n38343 = ~n38340 & ~n38342 ;
  assign n38344 = ~n38337 & n38343 ;
  assign n38345 = \b[31]  & n20519 ;
  assign n38346 = \a[60]  & \b[30]  ;
  assign n38347 = n20510 & n38346 ;
  assign n38348 = ~n38345 & ~n38347 ;
  assign n38349 = \b[29]  & n21315 ;
  assign n38350 = n21312 & n38349 ;
  assign n38351 = ~\a[60]  & \b[30]  ;
  assign n38352 = n20513 & n38351 ;
  assign n38353 = ~n38350 & ~n38352 ;
  assign n38354 = n38348 & n38353 ;
  assign n38355 = ~\a[62]  & ~n38354 ;
  assign n38356 = ~n5459 & n20521 ;
  assign n38357 = ~n5104 & n20521 ;
  assign n38358 = ~n5455 & n38357 ;
  assign n38359 = ~n38356 & ~n38358 ;
  assign n38360 = ~\a[62]  & ~n5462 ;
  assign n38361 = ~n38359 & n38360 ;
  assign n38362 = ~n38355 & ~n38361 ;
  assign n38363 = ~n37541 & ~n37882 ;
  assign n38364 = \b[28]  & n21958 ;
  assign n38365 = \b[27]  & n21957 ;
  assign n38366 = ~n38364 & ~n38365 ;
  assign n38367 = n37878 & ~n38366 ;
  assign n38368 = ~n38363 & n38367 ;
  assign n38369 = n37878 & ~n38363 ;
  assign n38370 = n38366 & ~n38369 ;
  assign n38371 = ~n38368 & ~n38370 ;
  assign n38372 = ~n5462 & ~n38359 ;
  assign n38373 = \a[62]  & n38354 ;
  assign n38374 = ~n38372 & n38373 ;
  assign n38375 = ~n38371 & ~n38374 ;
  assign n38376 = n38362 & n38375 ;
  assign n38377 = ~n38362 & n38371 ;
  assign n38378 = \a[62]  & ~n38368 ;
  assign n38379 = ~n38370 & n38378 ;
  assign n38380 = n38354 & n38379 ;
  assign n38381 = ~n38372 & n38380 ;
  assign n38382 = ~n38377 & ~n38381 ;
  assign n38383 = ~n38376 & n38382 ;
  assign n38384 = ~n37887 & n37912 ;
  assign n38385 = ~n37888 & ~n38384 ;
  assign n38386 = n38383 & n38385 ;
  assign n38387 = ~n38383 & ~n38385 ;
  assign n38388 = ~n38386 & ~n38387 ;
  assign n38389 = n6565 & n18516 ;
  assign n38390 = ~n6562 & n38389 ;
  assign n38391 = n18516 & n22947 ;
  assign n38392 = ~n6561 & n38391 ;
  assign n38393 = \b[34]  & n18514 ;
  assign n38394 = \a[56]  & \b[33]  ;
  assign n38395 = n19181 & n38394 ;
  assign n38396 = ~\a[57]  & \b[33]  ;
  assign n38397 = n18508 & n38396 ;
  assign n38398 = ~n38395 & ~n38397 ;
  assign n38399 = ~n38393 & n38398 ;
  assign n38400 = \b[32]  & n19183 ;
  assign n38401 = n19180 & n38400 ;
  assign n38402 = \a[59]  & ~n38401 ;
  assign n38403 = n38399 & n38402 ;
  assign n38404 = ~n38392 & n38403 ;
  assign n38405 = ~n38390 & n38404 ;
  assign n38406 = n38399 & ~n38401 ;
  assign n38407 = ~n38392 & n38406 ;
  assign n38408 = ~n38390 & n38407 ;
  assign n38409 = ~\a[59]  & ~n38408 ;
  assign n38410 = ~n38405 & ~n38409 ;
  assign n38411 = n38388 & ~n38410 ;
  assign n38412 = ~n38388 & n38410 ;
  assign n38413 = ~n38411 & ~n38412 ;
  assign n38414 = n38344 & ~n38413 ;
  assign n38415 = ~n38320 & n38414 ;
  assign n38416 = n38344 & n38413 ;
  assign n38417 = n38320 & n38416 ;
  assign n38418 = ~n38415 & ~n38417 ;
  assign n38419 = ~n38344 & ~n38413 ;
  assign n38420 = n38320 & n38419 ;
  assign n38421 = ~n38344 & n38413 ;
  assign n38422 = ~n38320 & n38421 ;
  assign n38423 = ~n38420 & ~n38422 ;
  assign n38424 = n38418 & n38423 ;
  assign n38425 = n38315 & ~n38424 ;
  assign n38426 = ~n38315 & n38424 ;
  assign n38427 = ~n38425 & ~n38426 ;
  assign n38428 = ~n38313 & n38427 ;
  assign n38429 = n38313 & ~n38427 ;
  assign n38430 = ~n38428 & ~n38429 ;
  assign n38431 = n38001 & ~n38011 ;
  assign n38432 = n38006 & ~n38431 ;
  assign n38433 = ~n10406 & n13125 ;
  assign n38434 = ~n9929 & n13125 ;
  assign n38435 = ~n10402 & n38434 ;
  assign n38436 = ~n38433 & ~n38435 ;
  assign n38437 = ~n10409 & ~n38436 ;
  assign n38438 = \b[41]  & n13794 ;
  assign n38439 = n13792 & n38438 ;
  assign n38440 = ~\a[48]  & \b[42]  ;
  assign n38441 = n13117 & n38440 ;
  assign n38442 = ~n38439 & ~n38441 ;
  assign n38443 = \b[43]  & n13123 ;
  assign n38444 = \a[48]  & \b[42]  ;
  assign n38445 = n13786 & n38444 ;
  assign n38446 = \a[50]  & ~n38445 ;
  assign n38447 = ~n38443 & n38446 ;
  assign n38448 = n38442 & n38447 ;
  assign n38449 = ~n38437 & n38448 ;
  assign n38450 = ~n38443 & ~n38445 ;
  assign n38451 = n38442 & n38450 ;
  assign n38452 = ~\a[50]  & ~n38451 ;
  assign n38453 = ~\a[50]  & ~n10409 ;
  assign n38454 = ~n38436 & n38453 ;
  assign n38455 = ~n38452 & ~n38454 ;
  assign n38456 = ~n38449 & n38455 ;
  assign n38457 = n38432 & ~n38456 ;
  assign n38458 = ~n38430 & n38457 ;
  assign n38459 = ~n38432 & ~n38456 ;
  assign n38460 = n38430 & n38459 ;
  assign n38461 = ~n38458 & ~n38460 ;
  assign n38462 = ~n38432 & n38456 ;
  assign n38463 = ~n38430 & n38462 ;
  assign n38464 = n38432 & n38456 ;
  assign n38465 = n38430 & n38464 ;
  assign n38466 = ~n38463 & ~n38465 ;
  assign n38467 = n38461 & n38466 ;
  assign n38468 = ~n38290 & ~n38467 ;
  assign n38469 = n38290 & n38467 ;
  assign n38470 = ~n38468 & ~n38469 ;
  assign n38471 = n11572 & n11906 ;
  assign n38472 = ~n11903 & n38471 ;
  assign n38473 = n11572 & n13483 ;
  assign n38474 = ~n11902 & n38473 ;
  assign n38475 = \b[44]  & n12159 ;
  assign n38476 = n12156 & n38475 ;
  assign n38477 = ~\a[45]  & \b[45]  ;
  assign n38478 = n11564 & n38477 ;
  assign n38479 = ~n38476 & ~n38478 ;
  assign n38480 = \b[46]  & n11570 ;
  assign n38481 = \a[45]  & \b[45]  ;
  assign n38482 = n11561 & n38481 ;
  assign n38483 = \a[47]  & ~n38482 ;
  assign n38484 = ~n38480 & n38483 ;
  assign n38485 = n38479 & n38484 ;
  assign n38486 = ~n38474 & n38485 ;
  assign n38487 = ~n38472 & n38486 ;
  assign n38488 = ~n38480 & ~n38482 ;
  assign n38489 = n38479 & n38488 ;
  assign n38490 = ~n38474 & n38489 ;
  assign n38491 = ~n38472 & n38490 ;
  assign n38492 = ~\a[47]  & ~n38491 ;
  assign n38493 = ~n38487 & ~n38492 ;
  assign n38494 = ~n38470 & n38493 ;
  assign n38495 = n38470 & ~n38493 ;
  assign n38496 = ~n38494 & ~n38495 ;
  assign n38497 = n38067 & n38075 ;
  assign n38498 = n38072 & ~n38497 ;
  assign n38499 = n10082 & ~n13524 ;
  assign n38500 = ~n13522 & n38499 ;
  assign n38501 = \b[49]  & n10080 ;
  assign n38502 = \a[41]  & \b[48]  ;
  assign n38503 = n10679 & n38502 ;
  assign n38504 = ~\a[42]  & \b[48]  ;
  assign n38505 = n10074 & n38504 ;
  assign n38506 = ~n38503 & ~n38505 ;
  assign n38507 = ~n38501 & n38506 ;
  assign n38508 = \b[47]  & n10681 ;
  assign n38509 = n10678 & n38508 ;
  assign n38510 = \a[44]  & ~n38509 ;
  assign n38511 = n38507 & n38510 ;
  assign n38512 = ~n38500 & n38511 ;
  assign n38513 = n38507 & ~n38509 ;
  assign n38514 = ~n38500 & n38513 ;
  assign n38515 = ~\a[44]  & ~n38514 ;
  assign n38516 = ~n38512 & ~n38515 ;
  assign n38517 = n38498 & ~n38516 ;
  assign n38518 = ~n38496 & n38517 ;
  assign n38519 = ~n38498 & ~n38516 ;
  assign n38520 = n38496 & n38519 ;
  assign n38521 = ~n38518 & ~n38520 ;
  assign n38522 = ~n38498 & n38516 ;
  assign n38523 = ~n38496 & n38522 ;
  assign n38524 = n38498 & n38516 ;
  assign n38525 = n38496 & n38524 ;
  assign n38526 = ~n38523 & ~n38525 ;
  assign n38527 = n38521 & n38526 ;
  assign n38528 = n38101 & ~n38111 ;
  assign n38529 = n38106 & ~n38528 ;
  assign n38530 = n8759 & n15201 ;
  assign n38531 = ~n15198 & n38530 ;
  assign n38532 = n8759 & n28871 ;
  assign n38533 = ~n15197 & n38532 ;
  assign n38534 = \b[50]  & n9301 ;
  assign n38535 = n9298 & n38534 ;
  assign n38536 = ~\a[39]  & \b[51]  ;
  assign n38537 = n8751 & n38536 ;
  assign n38538 = ~n38535 & ~n38537 ;
  assign n38539 = \b[52]  & n8757 ;
  assign n38540 = \a[39]  & \b[51]  ;
  assign n38541 = n8748 & n38540 ;
  assign n38542 = \a[41]  & ~n38541 ;
  assign n38543 = ~n38539 & n38542 ;
  assign n38544 = n38538 & n38543 ;
  assign n38545 = ~n38533 & n38544 ;
  assign n38546 = ~n38531 & n38545 ;
  assign n38547 = ~n38539 & ~n38541 ;
  assign n38548 = n38538 & n38547 ;
  assign n38549 = ~n38533 & n38548 ;
  assign n38550 = ~n38531 & n38549 ;
  assign n38551 = ~\a[41]  & ~n38550 ;
  assign n38552 = ~n38546 & ~n38551 ;
  assign n38553 = ~n38529 & n38552 ;
  assign n38554 = ~n38527 & n38553 ;
  assign n38555 = n38529 & n38552 ;
  assign n38556 = n38527 & n38555 ;
  assign n38557 = ~n38554 & ~n38556 ;
  assign n38558 = n38529 & ~n38552 ;
  assign n38559 = ~n38527 & n38558 ;
  assign n38560 = ~n38529 & ~n38552 ;
  assign n38561 = n38527 & n38560 ;
  assign n38562 = ~n38559 & ~n38561 ;
  assign n38563 = n38557 & n38562 ;
  assign n38564 = n7534 & ~n16446 ;
  assign n38565 = ~n16444 & n38564 ;
  assign n38566 = \b[53]  & n7973 ;
  assign n38567 = n7970 & n38566 ;
  assign n38568 = ~\a[36]  & \b[54]  ;
  assign n38569 = n7526 & n38568 ;
  assign n38570 = ~n38567 & ~n38569 ;
  assign n38571 = \b[55]  & n7532 ;
  assign n38572 = \a[36]  & \b[54]  ;
  assign n38573 = n17801 & n38572 ;
  assign n38574 = \a[38]  & ~n38573 ;
  assign n38575 = ~n38571 & n38574 ;
  assign n38576 = n38570 & n38575 ;
  assign n38577 = ~n38565 & n38576 ;
  assign n38578 = ~n38571 & ~n38573 ;
  assign n38579 = n38570 & n38578 ;
  assign n38580 = ~n38565 & n38579 ;
  assign n38581 = ~\a[38]  & ~n38580 ;
  assign n38582 = ~n38577 & ~n38581 ;
  assign n38583 = n38140 & n38169 ;
  assign n38584 = n38135 & ~n38583 ;
  assign n38585 = n38582 & ~n38584 ;
  assign n38586 = n38563 & n38585 ;
  assign n38587 = n38582 & n38584 ;
  assign n38588 = ~n38563 & n38587 ;
  assign n38589 = ~n38586 & ~n38588 ;
  assign n38590 = ~n38582 & ~n38584 ;
  assign n38591 = ~n38563 & n38590 ;
  assign n38592 = ~n38582 & n38584 ;
  assign n38593 = n38563 & n38592 ;
  assign n38594 = ~n38591 & ~n38593 ;
  assign n38595 = n38589 & n38594 ;
  assign n38596 = n38179 & ~n38182 ;
  assign n38597 = n38174 & ~n38596 ;
  assign n38598 = ~n18937 & ~n18940 ;
  assign n38599 = n6309 & ~n19543 ;
  assign n38600 = ~n38598 & n38599 ;
  assign n38601 = \b[56]  & n6778 ;
  assign n38602 = n6775 & n38601 ;
  assign n38603 = ~\a[33]  & \b[57]  ;
  assign n38604 = n6301 & n38603 ;
  assign n38605 = ~n38602 & ~n38604 ;
  assign n38606 = \b[58]  & n6307 ;
  assign n38607 = \a[33]  & \b[57]  ;
  assign n38608 = n6298 & n38607 ;
  assign n38609 = \a[35]  & ~n38608 ;
  assign n38610 = ~n38606 & n38609 ;
  assign n38611 = n38605 & n38610 ;
  assign n38612 = ~n38600 & n38611 ;
  assign n38613 = ~n38606 & ~n38608 ;
  assign n38614 = n38605 & n38613 ;
  assign n38615 = ~n38600 & n38614 ;
  assign n38616 = ~\a[35]  & ~n38615 ;
  assign n38617 = ~n38612 & ~n38616 ;
  assign n38618 = ~n38597 & ~n38617 ;
  assign n38619 = ~n38595 & n38618 ;
  assign n38620 = n38597 & ~n38617 ;
  assign n38621 = n38595 & n38620 ;
  assign n38622 = ~n38619 & ~n38621 ;
  assign n38623 = n38597 & n38617 ;
  assign n38624 = ~n38595 & n38623 ;
  assign n38625 = ~n38597 & n38617 ;
  assign n38626 = n38595 & n38625 ;
  assign n38627 = ~n38624 & ~n38626 ;
  assign n38628 = n38622 & n38627 ;
  assign n38629 = ~n38288 & n38628 ;
  assign n38630 = ~n38284 & n38629 ;
  assign n38631 = ~n38284 & ~n38288 ;
  assign n38632 = ~n38628 & ~n38631 ;
  assign n38633 = ~n38630 & ~n38632 ;
  assign n38634 = n38263 & n38633 ;
  assign n38635 = ~n38263 & ~n38633 ;
  assign n38636 = ~n38634 & ~n38635 ;
  assign n38637 = ~n38238 & ~n38636 ;
  assign n38638 = n38238 & n38636 ;
  assign n38639 = ~n38637 & ~n38638 ;
  assign n38640 = ~n38228 & n38639 ;
  assign n38641 = ~n38230 & n38640 ;
  assign n38642 = ~n38232 & n38641 ;
  assign n38643 = ~n38228 & ~n38230 ;
  assign n38644 = ~n38232 & n38643 ;
  assign n38645 = ~n38639 & ~n38644 ;
  assign n38646 = ~n38642 & ~n38645 ;
  assign n38647 = ~n38228 & ~n38638 ;
  assign n38648 = ~n38230 & n38647 ;
  assign n38649 = ~n38232 & n38648 ;
  assign n38650 = ~n38261 & ~n38633 ;
  assign n38651 = ~n38262 & ~n38650 ;
  assign n38652 = n38595 & ~n38597 ;
  assign n38653 = ~n38595 & n38597 ;
  assign n38654 = n38617 & ~n38653 ;
  assign n38655 = ~n38652 & ~n38654 ;
  assign n38656 = n5211 & ~n21699 ;
  assign n38657 = ~n21697 & n38656 ;
  assign n38658 = \b[62]  & n5209 ;
  assign n38659 = \a[30]  & \b[61]  ;
  assign n38660 = n5200 & n38659 ;
  assign n38661 = ~n38658 & ~n38660 ;
  assign n38662 = \b[60]  & n5595 ;
  assign n38663 = n5592 & n38662 ;
  assign n38664 = ~\a[30]  & \b[61]  ;
  assign n38665 = n5203 & n38664 ;
  assign n38666 = ~n38663 & ~n38665 ;
  assign n38667 = n38661 & n38666 ;
  assign n38668 = ~n38657 & n38667 ;
  assign n38669 = ~\a[32]  & ~n38668 ;
  assign n38670 = \a[32]  & ~n38660 ;
  assign n38671 = ~n38658 & n38670 ;
  assign n38672 = n38666 & n38671 ;
  assign n38673 = ~n38657 & n38672 ;
  assign n38674 = ~n38669 & ~n38673 ;
  assign n38675 = ~n38655 & n38674 ;
  assign n38676 = ~n38652 & n38669 ;
  assign n38677 = ~n38654 & n38676 ;
  assign n38678 = \a[32]  & n38668 ;
  assign n38679 = ~n38652 & n38678 ;
  assign n38680 = ~n38654 & n38679 ;
  assign n38681 = ~n38677 & ~n38680 ;
  assign n38682 = ~n38675 & n38681 ;
  assign n38683 = n8759 & ~n15246 ;
  assign n38684 = ~n15244 & n38683 ;
  assign n38685 = \b[51]  & n9301 ;
  assign n38686 = n9298 & n38685 ;
  assign n38687 = ~\a[39]  & \b[52]  ;
  assign n38688 = n8751 & n38687 ;
  assign n38689 = ~n38686 & ~n38688 ;
  assign n38690 = \b[53]  & n8757 ;
  assign n38691 = \a[39]  & \b[52]  ;
  assign n38692 = n8748 & n38691 ;
  assign n38693 = \a[41]  & ~n38692 ;
  assign n38694 = ~n38690 & n38693 ;
  assign n38695 = n38689 & n38694 ;
  assign n38696 = ~n38684 & n38695 ;
  assign n38697 = ~n38690 & ~n38692 ;
  assign n38698 = n38689 & n38697 ;
  assign n38699 = ~n38684 & n38698 ;
  assign n38700 = ~\a[41]  & ~n38699 ;
  assign n38701 = ~n38696 & ~n38700 ;
  assign n38702 = ~n10889 & ~n12606 ;
  assign n38703 = ~n13122 & n38702 ;
  assign n38704 = n10886 & n38703 ;
  assign n38705 = n10889 & ~n12606 ;
  assign n38706 = ~n13122 & n38705 ;
  assign n38707 = ~n10886 & n38706 ;
  assign n38708 = ~n38704 & ~n38707 ;
  assign n38709 = \b[42]  & n13794 ;
  assign n38710 = n13792 & n38709 ;
  assign n38711 = ~\a[48]  & \b[43]  ;
  assign n38712 = n13117 & n38711 ;
  assign n38713 = ~n38710 & ~n38712 ;
  assign n38714 = \b[44]  & n13123 ;
  assign n38715 = \a[48]  & \b[43]  ;
  assign n38716 = n13786 & n38715 ;
  assign n38717 = \a[50]  & ~n38716 ;
  assign n38718 = ~n38714 & n38717 ;
  assign n38719 = n38713 & n38718 ;
  assign n38720 = n38708 & n38719 ;
  assign n38721 = ~n38714 & ~n38716 ;
  assign n38722 = n38713 & n38721 ;
  assign n38723 = n38708 & n38722 ;
  assign n38724 = ~\a[50]  & ~n38723 ;
  assign n38725 = ~n38720 & ~n38724 ;
  assign n38726 = n38313 & ~n38425 ;
  assign n38727 = ~n38425 & n38426 ;
  assign n38728 = ~n38726 & ~n38727 ;
  assign n38729 = ~n6610 & n18516 ;
  assign n38730 = ~n6608 & n38729 ;
  assign n38731 = \b[35]  & n18514 ;
  assign n38732 = \a[56]  & \b[34]  ;
  assign n38733 = n19181 & n38732 ;
  assign n38734 = ~\a[57]  & \b[34]  ;
  assign n38735 = n18508 & n38734 ;
  assign n38736 = ~n38733 & ~n38735 ;
  assign n38737 = ~n38731 & n38736 ;
  assign n38738 = \b[33]  & n19183 ;
  assign n38739 = n19180 & n38738 ;
  assign n38740 = \a[59]  & ~n38739 ;
  assign n38741 = n38737 & n38740 ;
  assign n38742 = ~n38730 & n38741 ;
  assign n38743 = n38737 & ~n38739 ;
  assign n38744 = ~n38730 & n38743 ;
  assign n38745 = ~\a[59]  & ~n38744 ;
  assign n38746 = ~n38742 & ~n38745 ;
  assign n38747 = ~n38370 & ~n38381 ;
  assign n38748 = ~n38377 & n38747 ;
  assign n38749 = \b[29]  & n21958 ;
  assign n38750 = \b[28]  & n21957 ;
  assign n38751 = ~n38749 & ~n38750 ;
  assign n38752 = n38366 & ~n38751 ;
  assign n38753 = ~n38366 & n38751 ;
  assign n38754 = ~n38752 & ~n38753 ;
  assign n38755 = ~n38748 & n38754 ;
  assign n38756 = n5810 & n20521 ;
  assign n38757 = ~n5807 & n38756 ;
  assign n38758 = n20521 & n37504 ;
  assign n38759 = ~n5806 & n38758 ;
  assign n38760 = \b[30]  & n21315 ;
  assign n38761 = n21312 & n38760 ;
  assign n38762 = ~\a[60]  & \b[31]  ;
  assign n38763 = n20513 & n38762 ;
  assign n38764 = ~n38761 & ~n38763 ;
  assign n38765 = \b[32]  & n20519 ;
  assign n38766 = \a[60]  & \b[31]  ;
  assign n38767 = n20510 & n38766 ;
  assign n38768 = \a[62]  & ~n38767 ;
  assign n38769 = ~n38765 & n38768 ;
  assign n38770 = n38764 & n38769 ;
  assign n38771 = ~n38759 & n38770 ;
  assign n38772 = ~n38757 & n38771 ;
  assign n38773 = ~n38765 & ~n38767 ;
  assign n38774 = n38764 & n38773 ;
  assign n38775 = ~n38759 & n38774 ;
  assign n38776 = ~n38757 & n38775 ;
  assign n38777 = ~\a[62]  & ~n38776 ;
  assign n38778 = ~n38772 & ~n38777 ;
  assign n38779 = n38748 & ~n38754 ;
  assign n38780 = ~n38778 & ~n38779 ;
  assign n38781 = ~n38755 & n38780 ;
  assign n38782 = ~n38755 & ~n38779 ;
  assign n38783 = n38778 & ~n38782 ;
  assign n38784 = ~n38781 & ~n38783 ;
  assign n38785 = ~n38386 & n38410 ;
  assign n38786 = ~n38387 & ~n38785 ;
  assign n38787 = ~n38784 & n38786 ;
  assign n38788 = ~n38746 & n38787 ;
  assign n38789 = n38784 & n38786 ;
  assign n38790 = n38746 & n38789 ;
  assign n38791 = ~n38788 & ~n38790 ;
  assign n38792 = n38746 & ~n38784 ;
  assign n38793 = ~n38786 & n38792 ;
  assign n38794 = n38784 & ~n38786 ;
  assign n38795 = ~n38746 & n38794 ;
  assign n38796 = ~n38793 & ~n38795 ;
  assign n38797 = n38791 & n38796 ;
  assign n38798 = n8175 & n16655 ;
  assign n38799 = ~n8172 & n38798 ;
  assign n38800 = n25622 & n37945 ;
  assign n38801 = ~n8171 & n38800 ;
  assign n38802 = \b[36]  & n17308 ;
  assign n38803 = n17305 & n38802 ;
  assign n38804 = ~\a[54]  & \b[37]  ;
  assign n38805 = n16647 & n38804 ;
  assign n38806 = ~n38803 & ~n38805 ;
  assign n38807 = \b[38]  & n16653 ;
  assign n38808 = \a[54]  & \b[37]  ;
  assign n38809 = n16644 & n38808 ;
  assign n38810 = \a[56]  & ~n38809 ;
  assign n38811 = ~n38807 & n38810 ;
  assign n38812 = n38806 & n38811 ;
  assign n38813 = ~n38801 & n38812 ;
  assign n38814 = ~n38799 & n38813 ;
  assign n38815 = ~n38807 & ~n38809 ;
  assign n38816 = n38806 & n38815 ;
  assign n38817 = ~n38801 & n38816 ;
  assign n38818 = ~n38799 & n38817 ;
  assign n38819 = ~\a[56]  & ~n38818 ;
  assign n38820 = ~n38814 & ~n38819 ;
  assign n38821 = n38797 & ~n38820 ;
  assign n38822 = ~n38797 & n38820 ;
  assign n38823 = ~n38821 & ~n38822 ;
  assign n38824 = ~n9479 & n14793 ;
  assign n38825 = ~n9043 & n14793 ;
  assign n38826 = ~n9475 & n38825 ;
  assign n38827 = ~n38824 & ~n38826 ;
  assign n38828 = ~n9482 & ~n38827 ;
  assign n38829 = \b[39]  & n15517 ;
  assign n38830 = n15514 & n38829 ;
  assign n38831 = ~\a[51]  & \b[40]  ;
  assign n38832 = n14785 & n38831 ;
  assign n38833 = ~n38830 & ~n38832 ;
  assign n38834 = \b[41]  & n14791 ;
  assign n38835 = \a[51]  & \b[40]  ;
  assign n38836 = n14782 & n38835 ;
  assign n38837 = \a[53]  & ~n38836 ;
  assign n38838 = ~n38834 & n38837 ;
  assign n38839 = n38833 & n38838 ;
  assign n38840 = ~n38828 & n38839 ;
  assign n38841 = ~n38834 & ~n38836 ;
  assign n38842 = n38833 & n38841 ;
  assign n38843 = ~\a[53]  & ~n38842 ;
  assign n38844 = ~\a[53]  & ~n9482 ;
  assign n38845 = ~n38827 & n38844 ;
  assign n38846 = ~n38843 & ~n38845 ;
  assign n38847 = ~n38840 & n38846 ;
  assign n38848 = n38320 & ~n38413 ;
  assign n38849 = ~n38320 & n38413 ;
  assign n38850 = n38344 & ~n38849 ;
  assign n38851 = ~n38848 & ~n38850 ;
  assign n38852 = n38847 & ~n38851 ;
  assign n38853 = n38823 & n38852 ;
  assign n38854 = n38847 & n38851 ;
  assign n38855 = ~n38823 & n38854 ;
  assign n38856 = ~n38853 & ~n38855 ;
  assign n38857 = ~n38847 & ~n38851 ;
  assign n38858 = ~n38823 & n38857 ;
  assign n38859 = ~n38847 & n38851 ;
  assign n38860 = n38823 & n38859 ;
  assign n38861 = ~n38858 & ~n38860 ;
  assign n38862 = n38856 & n38861 ;
  assign n38863 = n38728 & ~n38862 ;
  assign n38864 = ~n38728 & n38862 ;
  assign n38865 = ~n38863 & ~n38864 ;
  assign n38866 = ~n38725 & n38865 ;
  assign n38867 = n38725 & ~n38865 ;
  assign n38868 = ~n38866 & ~n38867 ;
  assign n38869 = ~n38430 & ~n38432 ;
  assign n38870 = ~n38432 & ~n38449 ;
  assign n38871 = n38313 & ~n38449 ;
  assign n38872 = ~n38427 & n38871 ;
  assign n38873 = ~n38313 & ~n38449 ;
  assign n38874 = n38427 & n38873 ;
  assign n38875 = ~n38872 & ~n38874 ;
  assign n38876 = ~n38870 & n38875 ;
  assign n38877 = n38455 & ~n38876 ;
  assign n38878 = ~n38869 & ~n38877 ;
  assign n38879 = n11572 & ~n12438 ;
  assign n38880 = ~n12436 & n38879 ;
  assign n38881 = \b[45]  & n12159 ;
  assign n38882 = n12156 & n38881 ;
  assign n38883 = ~\a[45]  & \b[46]  ;
  assign n38884 = n11564 & n38883 ;
  assign n38885 = ~n38882 & ~n38884 ;
  assign n38886 = \b[47]  & n11570 ;
  assign n38887 = \a[45]  & \b[46]  ;
  assign n38888 = n11561 & n38887 ;
  assign n38889 = \a[47]  & ~n38888 ;
  assign n38890 = ~n38886 & n38889 ;
  assign n38891 = n38885 & n38890 ;
  assign n38892 = ~n38880 & n38891 ;
  assign n38893 = ~n38886 & ~n38888 ;
  assign n38894 = n38885 & n38893 ;
  assign n38895 = ~n38880 & n38894 ;
  assign n38896 = ~\a[47]  & ~n38895 ;
  assign n38897 = ~n38892 & ~n38896 ;
  assign n38898 = ~n38878 & ~n38897 ;
  assign n38899 = n38868 & n38898 ;
  assign n38900 = n38878 & ~n38897 ;
  assign n38901 = ~n38868 & n38900 ;
  assign n38902 = ~n38899 & ~n38901 ;
  assign n38903 = ~n38878 & n38897 ;
  assign n38904 = ~n38868 & n38903 ;
  assign n38905 = n38878 & n38897 ;
  assign n38906 = n38868 & n38905 ;
  assign n38907 = ~n38904 & ~n38906 ;
  assign n38908 = n38902 & n38907 ;
  assign n38909 = ~n38469 & n38493 ;
  assign n38910 = ~n38468 & ~n38909 ;
  assign n38911 = n10082 & n14052 ;
  assign n38912 = ~n14049 & n38911 ;
  assign n38913 = n10082 & n15779 ;
  assign n38914 = ~n14048 & n38913 ;
  assign n38915 = \b[48]  & n10681 ;
  assign n38916 = n10678 & n38915 ;
  assign n38917 = \b[50]  & n10080 ;
  assign n38918 = \a[41]  & \b[49]  ;
  assign n38919 = n10679 & n38918 ;
  assign n38920 = ~\a[42]  & \b[49]  ;
  assign n38921 = n10074 & n38920 ;
  assign n38922 = ~n38919 & ~n38921 ;
  assign n38923 = ~n38917 & n38922 ;
  assign n38924 = ~n38916 & n38923 ;
  assign n38925 = ~n38914 & n38924 ;
  assign n38926 = ~n38912 & n38925 ;
  assign n38927 = ~\a[44]  & ~n38926 ;
  assign n38928 = \a[44]  & n38924 ;
  assign n38929 = ~n38914 & n38928 ;
  assign n38930 = ~n38912 & n38929 ;
  assign n38931 = ~n38927 & ~n38930 ;
  assign n38932 = ~n38910 & n38931 ;
  assign n38933 = ~n38908 & n38932 ;
  assign n38934 = n38910 & n38931 ;
  assign n38935 = n38908 & n38934 ;
  assign n38936 = ~n38933 & ~n38935 ;
  assign n38937 = ~n38910 & ~n38931 ;
  assign n38938 = n38908 & n38937 ;
  assign n38939 = n38910 & ~n38931 ;
  assign n38940 = ~n38908 & n38939 ;
  assign n38941 = ~n38938 & ~n38940 ;
  assign n38942 = n38936 & n38941 ;
  assign n38943 = ~n38496 & ~n38498 ;
  assign n38944 = n38496 & n38498 ;
  assign n38945 = n38516 & ~n38944 ;
  assign n38946 = ~n38943 & ~n38945 ;
  assign n38947 = n38942 & n38946 ;
  assign n38948 = ~n38942 & ~n38946 ;
  assign n38949 = ~n38947 & ~n38948 ;
  assign n38950 = n38701 & n38949 ;
  assign n38951 = ~n38701 & ~n38949 ;
  assign n38952 = ~n38950 & ~n38951 ;
  assign n38953 = n7534 & n17647 ;
  assign n38954 = ~n17644 & n38953 ;
  assign n38955 = n7534 & n19567 ;
  assign n38956 = ~n17643 & n38955 ;
  assign n38957 = \b[54]  & n7973 ;
  assign n38958 = n7970 & n38957 ;
  assign n38959 = ~\a[36]  & \b[55]  ;
  assign n38960 = n7526 & n38959 ;
  assign n38961 = ~n38958 & ~n38960 ;
  assign n38962 = \b[56]  & n7532 ;
  assign n38963 = \a[36]  & \b[55]  ;
  assign n38964 = n17801 & n38963 ;
  assign n38965 = \a[38]  & ~n38964 ;
  assign n38966 = ~n38962 & n38965 ;
  assign n38967 = n38961 & n38966 ;
  assign n38968 = ~n38956 & n38967 ;
  assign n38969 = ~n38954 & n38968 ;
  assign n38970 = ~n38962 & ~n38964 ;
  assign n38971 = n38961 & n38970 ;
  assign n38972 = ~n38956 & n38971 ;
  assign n38973 = ~n38954 & n38972 ;
  assign n38974 = ~\a[38]  & ~n38973 ;
  assign n38975 = ~n38969 & ~n38974 ;
  assign n38976 = ~n38527 & ~n38529 ;
  assign n38977 = n38527 & n38529 ;
  assign n38978 = n38552 & ~n38977 ;
  assign n38979 = ~n38976 & ~n38978 ;
  assign n38980 = ~n38975 & ~n38979 ;
  assign n38981 = ~n38952 & n38980 ;
  assign n38982 = ~n38975 & n38979 ;
  assign n38983 = n38952 & n38982 ;
  assign n38984 = ~n38981 & ~n38983 ;
  assign n38985 = n38975 & ~n38979 ;
  assign n38986 = n38952 & n38985 ;
  assign n38987 = n38975 & n38979 ;
  assign n38988 = ~n38952 & n38987 ;
  assign n38989 = ~n38986 & ~n38988 ;
  assign n38990 = n38984 & n38989 ;
  assign n38991 = ~n38563 & ~n38584 ;
  assign n38992 = n38563 & n38584 ;
  assign n38993 = n38582 & ~n38992 ;
  assign n38994 = ~n38991 & ~n38993 ;
  assign n38995 = n6309 & ~n19550 ;
  assign n38996 = ~n19548 & n38995 ;
  assign n38997 = \b[57]  & n6778 ;
  assign n38998 = n6775 & n38997 ;
  assign n38999 = ~\a[33]  & \b[58]  ;
  assign n39000 = n6301 & n38999 ;
  assign n39001 = ~n38998 & ~n39000 ;
  assign n39002 = \b[59]  & n6307 ;
  assign n39003 = \a[33]  & \b[58]  ;
  assign n39004 = n6298 & n39003 ;
  assign n39005 = \a[35]  & ~n39004 ;
  assign n39006 = ~n39002 & n39005 ;
  assign n39007 = n39001 & n39006 ;
  assign n39008 = ~n38996 & n39007 ;
  assign n39009 = ~n39002 & ~n39004 ;
  assign n39010 = n39001 & n39009 ;
  assign n39011 = ~n38996 & n39010 ;
  assign n39012 = ~\a[35]  & ~n39011 ;
  assign n39013 = ~n39008 & ~n39012 ;
  assign n39014 = n38994 & ~n39013 ;
  assign n39015 = ~n38990 & n39014 ;
  assign n39016 = ~n38994 & ~n39013 ;
  assign n39017 = n38990 & n39016 ;
  assign n39018 = ~n39015 & ~n39017 ;
  assign n39019 = ~n38994 & n39013 ;
  assign n39020 = ~n38990 & n39019 ;
  assign n39021 = n38994 & n39013 ;
  assign n39022 = n38990 & n39021 ;
  assign n39023 = ~n39020 & ~n39022 ;
  assign n39024 = n39018 & n39023 ;
  assign n39025 = ~n38682 & ~n39024 ;
  assign n39026 = n38682 & n39024 ;
  assign n39027 = ~n39025 & ~n39026 ;
  assign n39028 = ~n38288 & ~n38628 ;
  assign n39029 = ~n38209 & n38286 ;
  assign n39030 = n38285 & n38286 ;
  assign n39031 = ~n39029 & ~n39030 ;
  assign n39032 = ~n39028 & n39031 ;
  assign n39033 = \b[63]  & ~n21694 ;
  assign n39034 = n4249 & n39033 ;
  assign n39035 = ~n23171 & n39034 ;
  assign n39036 = \a[26]  & \a[28]  ;
  assign n39037 = \a[27]  & ~\a[29]  ;
  assign n39038 = n39036 & n39037 ;
  assign n39039 = ~\a[26]  & ~\a[28]  ;
  assign n39040 = ~\a[27]  & \a[29]  ;
  assign n39041 = n39039 & n39040 ;
  assign n39042 = ~n39038 & ~n39041 ;
  assign n39043 = \b[63]  & ~n39042 ;
  assign n39044 = \a[29]  & ~n39043 ;
  assign n39045 = ~n39035 & n39044 ;
  assign n39046 = ~n39035 & ~n39043 ;
  assign n39047 = ~\a[29]  & ~n39046 ;
  assign n39048 = ~n39045 & ~n39047 ;
  assign n39049 = n39032 & ~n39048 ;
  assign n39050 = ~n39032 & n39048 ;
  assign n39051 = ~n39049 & ~n39050 ;
  assign n39052 = n39027 & n39051 ;
  assign n39053 = ~n39027 & ~n39051 ;
  assign n39054 = ~n39052 & ~n39053 ;
  assign n39055 = n38651 & n39054 ;
  assign n39056 = ~n38651 & ~n39054 ;
  assign n39057 = ~n39055 & ~n39056 ;
  assign n39058 = ~n38637 & n39057 ;
  assign n39059 = ~n38649 & n39058 ;
  assign n39060 = ~n38637 & ~n38649 ;
  assign n39061 = ~n39057 & ~n39060 ;
  assign n39062 = ~n39059 & ~n39061 ;
  assign n39063 = ~n39055 & ~n39059 ;
  assign n39064 = ~n39049 & ~n39052 ;
  assign n39065 = ~n38952 & n38979 ;
  assign n39066 = n38984 & ~n39065 ;
  assign n39067 = ~n8599 & n37945 ;
  assign n39068 = ~n8174 & n37945 ;
  assign n39069 = ~n8595 & n39068 ;
  assign n39070 = ~n39067 & ~n39069 ;
  assign n39071 = ~n8602 & ~n39070 ;
  assign n39072 = \b[37]  & n17308 ;
  assign n39073 = n17305 & n39072 ;
  assign n39074 = ~\a[54]  & \b[38]  ;
  assign n39075 = n16647 & n39074 ;
  assign n39076 = ~n39073 & ~n39075 ;
  assign n39077 = \b[39]  & n16653 ;
  assign n39078 = \a[54]  & \b[38]  ;
  assign n39079 = n16644 & n39078 ;
  assign n39080 = \a[56]  & ~n39079 ;
  assign n39081 = ~n39077 & n39080 ;
  assign n39082 = n39076 & n39081 ;
  assign n39083 = ~n39071 & n39082 ;
  assign n39084 = ~n39077 & ~n39079 ;
  assign n39085 = n39076 & n39084 ;
  assign n39086 = ~\a[56]  & ~n39085 ;
  assign n39087 = ~\a[56]  & ~n8602 ;
  assign n39088 = ~n39070 & n39087 ;
  assign n39089 = ~n39086 & ~n39088 ;
  assign n39090 = ~n39083 & n39089 ;
  assign n39091 = n38755 & n38778 ;
  assign n39092 = n38778 & n38779 ;
  assign n39093 = ~n39091 & ~n39092 ;
  assign n39094 = n38746 & ~n38781 ;
  assign n39095 = n39093 & ~n39094 ;
  assign n39096 = n7337 & n18516 ;
  assign n39097 = ~n7334 & n39096 ;
  assign n39098 = n18516 & n37946 ;
  assign n39099 = ~n7333 & n39098 ;
  assign n39100 = \b[34]  & n19183 ;
  assign n39101 = n19180 & n39100 ;
  assign n39102 = \b[36]  & n18514 ;
  assign n39103 = \a[56]  & \b[35]  ;
  assign n39104 = n19181 & n39103 ;
  assign n39105 = ~\a[57]  & \b[35]  ;
  assign n39106 = n18508 & n39105 ;
  assign n39107 = ~n39104 & ~n39106 ;
  assign n39108 = ~n39102 & n39107 ;
  assign n39109 = ~n39101 & n39108 ;
  assign n39110 = ~n39099 & n39109 ;
  assign n39111 = ~n39097 & n39110 ;
  assign n39112 = ~\a[59]  & ~n39111 ;
  assign n39113 = \a[59]  & n39109 ;
  assign n39114 = ~n39099 & n39113 ;
  assign n39115 = ~n39097 & n39114 ;
  assign n39116 = ~n39112 & ~n39115 ;
  assign n39117 = ~n5855 & n20521 ;
  assign n39118 = ~n5853 & n39117 ;
  assign n39119 = \b[31]  & n21315 ;
  assign n39120 = n21312 & n39119 ;
  assign n39121 = ~\a[60]  & \b[32]  ;
  assign n39122 = n20513 & n39121 ;
  assign n39123 = ~n39120 & ~n39122 ;
  assign n39124 = \b[33]  & n20519 ;
  assign n39125 = \a[60]  & \b[32]  ;
  assign n39126 = n20510 & n39125 ;
  assign n39127 = \a[62]  & ~n39126 ;
  assign n39128 = ~n39124 & n39127 ;
  assign n39129 = n39123 & n39128 ;
  assign n39130 = ~n39118 & n39129 ;
  assign n39131 = ~n39124 & ~n39126 ;
  assign n39132 = n39123 & n39131 ;
  assign n39133 = ~n39118 & n39132 ;
  assign n39134 = ~\a[62]  & ~n39133 ;
  assign n39135 = ~n39130 & ~n39134 ;
  assign n39136 = ~n38370 & ~n38753 ;
  assign n39137 = ~n38381 & n39136 ;
  assign n39138 = ~n38377 & n39137 ;
  assign n39139 = ~\a[29]  & \b[29]  ;
  assign n39140 = n21957 & n39139 ;
  assign n39141 = ~\a[29]  & \b[30]  ;
  assign n39142 = n21958 & n39141 ;
  assign n39143 = ~n39140 & ~n39142 ;
  assign n39144 = \b[30]  & n21958 ;
  assign n39145 = \b[29]  & n21957 ;
  assign n39146 = \a[29]  & ~n39145 ;
  assign n39147 = ~n39144 & n39146 ;
  assign n39148 = n39143 & ~n39147 ;
  assign n39149 = ~n38751 & ~n39148 ;
  assign n39150 = n38751 & n39148 ;
  assign n39151 = ~n39149 & ~n39150 ;
  assign n39152 = ~n38752 & ~n39151 ;
  assign n39153 = ~n39138 & n39152 ;
  assign n39154 = ~n38752 & ~n39138 ;
  assign n39155 = n39151 & ~n39154 ;
  assign n39156 = ~n39153 & ~n39155 ;
  assign n39157 = n39135 & n39156 ;
  assign n39158 = ~n39135 & ~n39156 ;
  assign n39159 = ~n39157 & ~n39158 ;
  assign n39160 = ~n39116 & ~n39159 ;
  assign n39161 = n39116 & n39159 ;
  assign n39162 = ~n39160 & ~n39161 ;
  assign n39163 = n39095 & n39162 ;
  assign n39164 = ~n39095 & ~n39162 ;
  assign n39165 = ~n39163 & ~n39164 ;
  assign n39166 = n38746 & ~n38814 ;
  assign n39167 = ~n38789 & n39166 ;
  assign n39168 = ~n38746 & ~n38814 ;
  assign n39169 = ~n38787 & n39168 ;
  assign n39170 = ~n39167 & ~n39169 ;
  assign n39171 = ~n38819 & ~n39170 ;
  assign n39172 = n38796 & ~n39171 ;
  assign n39173 = n39165 & ~n39172 ;
  assign n39174 = ~n39090 & n39173 ;
  assign n39175 = ~n39165 & ~n39172 ;
  assign n39176 = n39090 & n39175 ;
  assign n39177 = ~n39174 & ~n39176 ;
  assign n39178 = n38796 & ~n39090 ;
  assign n39179 = ~n39171 & n39178 ;
  assign n39180 = ~n39165 & n39179 ;
  assign n39181 = n38796 & n39090 ;
  assign n39182 = ~n39171 & n39181 ;
  assign n39183 = n39165 & n39182 ;
  assign n39184 = ~n39180 & ~n39183 ;
  assign n39185 = ~n9930 & ~n14276 ;
  assign n39186 = ~n14790 & n39185 ;
  assign n39187 = n9927 & n39186 ;
  assign n39188 = n9930 & ~n14276 ;
  assign n39189 = ~n14790 & n39188 ;
  assign n39190 = ~n9927 & n39189 ;
  assign n39191 = ~n39187 & ~n39190 ;
  assign n39192 = \b[40]  & n15517 ;
  assign n39193 = n15514 & n39192 ;
  assign n39194 = ~\a[51]  & \b[41]  ;
  assign n39195 = n14785 & n39194 ;
  assign n39196 = ~n39193 & ~n39195 ;
  assign n39197 = \b[42]  & n14791 ;
  assign n39198 = \a[51]  & \b[41]  ;
  assign n39199 = n14782 & n39198 ;
  assign n39200 = \a[53]  & ~n39199 ;
  assign n39201 = ~n39197 & n39200 ;
  assign n39202 = n39196 & n39201 ;
  assign n39203 = n39191 & n39202 ;
  assign n39204 = ~n39197 & ~n39199 ;
  assign n39205 = n39196 & n39204 ;
  assign n39206 = n39191 & n39205 ;
  assign n39207 = ~\a[53]  & ~n39206 ;
  assign n39208 = ~n39203 & ~n39207 ;
  assign n39209 = n39184 & ~n39208 ;
  assign n39210 = n39177 & n39209 ;
  assign n39211 = n39177 & n39184 ;
  assign n39212 = n39208 & ~n39211 ;
  assign n39213 = ~n39210 & ~n39212 ;
  assign n39214 = ~n38823 & ~n38851 ;
  assign n39215 = n38823 & n38851 ;
  assign n39216 = n38847 & ~n39215 ;
  assign n39217 = ~n39214 & ~n39216 ;
  assign n39218 = ~n39213 & ~n39217 ;
  assign n39219 = ~n11397 & n13125 ;
  assign n39220 = ~n11395 & n39219 ;
  assign n39221 = \b[43]  & n13794 ;
  assign n39222 = n13792 & n39221 ;
  assign n39223 = ~\a[48]  & \b[44]  ;
  assign n39224 = n13117 & n39223 ;
  assign n39225 = ~n39222 & ~n39224 ;
  assign n39226 = \b[45]  & n13123 ;
  assign n39227 = \a[48]  & \b[44]  ;
  assign n39228 = n13786 & n39227 ;
  assign n39229 = \a[50]  & ~n39228 ;
  assign n39230 = ~n39226 & n39229 ;
  assign n39231 = n39225 & n39230 ;
  assign n39232 = ~n39220 & n39231 ;
  assign n39233 = ~n39226 & ~n39228 ;
  assign n39234 = n39225 & n39233 ;
  assign n39235 = ~n39220 & n39234 ;
  assign n39236 = ~\a[50]  & ~n39235 ;
  assign n39237 = ~n39232 & ~n39236 ;
  assign n39238 = ~n39210 & n39217 ;
  assign n39239 = ~n39212 & n39238 ;
  assign n39240 = ~n39237 & ~n39239 ;
  assign n39241 = ~n39218 & n39240 ;
  assign n39242 = ~n39217 & n39237 ;
  assign n39243 = ~n39213 & n39242 ;
  assign n39244 = n39217 & n39237 ;
  assign n39245 = n39213 & n39244 ;
  assign n39246 = ~n39243 & ~n39245 ;
  assign n39247 = ~n39241 & n39246 ;
  assign n39248 = n38725 & ~n38863 ;
  assign n39249 = ~n38863 & n38864 ;
  assign n39250 = ~n39248 & ~n39249 ;
  assign n39251 = n11572 & n12478 ;
  assign n39252 = ~n12475 & n39251 ;
  assign n39253 = n11572 & n28668 ;
  assign n39254 = ~n12474 & n39253 ;
  assign n39255 = \b[46]  & n12159 ;
  assign n39256 = n12156 & n39255 ;
  assign n39257 = ~\a[45]  & \b[47]  ;
  assign n39258 = n11564 & n39257 ;
  assign n39259 = ~n39256 & ~n39258 ;
  assign n39260 = \b[48]  & n11570 ;
  assign n39261 = \a[45]  & \b[47]  ;
  assign n39262 = n11561 & n39261 ;
  assign n39263 = \a[47]  & ~n39262 ;
  assign n39264 = ~n39260 & n39263 ;
  assign n39265 = n39259 & n39264 ;
  assign n39266 = ~n39254 & n39265 ;
  assign n39267 = ~n39252 & n39266 ;
  assign n39268 = ~n39260 & ~n39262 ;
  assign n39269 = n39259 & n39268 ;
  assign n39270 = ~n39254 & n39269 ;
  assign n39271 = ~n39252 & n39270 ;
  assign n39272 = ~\a[47]  & ~n39271 ;
  assign n39273 = ~n39267 & ~n39272 ;
  assign n39274 = n39250 & ~n39273 ;
  assign n39275 = ~n39247 & n39274 ;
  assign n39276 = ~n39250 & ~n39273 ;
  assign n39277 = n39247 & n39276 ;
  assign n39278 = ~n39275 & ~n39277 ;
  assign n39279 = ~n39250 & n39273 ;
  assign n39280 = ~n39247 & n39279 ;
  assign n39281 = n39250 & n39273 ;
  assign n39282 = n39247 & n39281 ;
  assign n39283 = ~n39280 & ~n39282 ;
  assign n39284 = n39278 & n39283 ;
  assign n39285 = ~n38868 & ~n38878 ;
  assign n39286 = n38868 & n38878 ;
  assign n39287 = n38897 & ~n39286 ;
  assign n39288 = ~n39285 & ~n39287 ;
  assign n39289 = n10082 & ~n14098 ;
  assign n39290 = ~n14096 & n39289 ;
  assign n39291 = \b[49]  & n10681 ;
  assign n39292 = n10678 & n39291 ;
  assign n39293 = \b[51]  & n10080 ;
  assign n39294 = \a[41]  & \b[50]  ;
  assign n39295 = n10679 & n39294 ;
  assign n39296 = ~\a[42]  & \b[50]  ;
  assign n39297 = n10074 & n39296 ;
  assign n39298 = ~n39295 & ~n39297 ;
  assign n39299 = ~n39293 & n39298 ;
  assign n39300 = ~n39292 & n39299 ;
  assign n39301 = ~\a[44]  & n39300 ;
  assign n39302 = ~n39290 & n39301 ;
  assign n39303 = ~n39290 & n39300 ;
  assign n39304 = \a[44]  & ~n39303 ;
  assign n39305 = ~n39302 & ~n39304 ;
  assign n39306 = ~n39288 & ~n39305 ;
  assign n39307 = ~n39284 & n39306 ;
  assign n39308 = n39288 & ~n39305 ;
  assign n39309 = n39284 & n39308 ;
  assign n39310 = ~n39307 & ~n39309 ;
  assign n39311 = ~n39288 & n39305 ;
  assign n39312 = n39284 & n39311 ;
  assign n39313 = n39288 & n39305 ;
  assign n39314 = ~n39284 & n39313 ;
  assign n39315 = ~n39312 & ~n39314 ;
  assign n39316 = n39310 & n39315 ;
  assign n39317 = n8759 & n38142 ;
  assign n39318 = ~n16404 & n39317 ;
  assign n39319 = n8759 & n16398 ;
  assign n39320 = n15241 & n39319 ;
  assign n39321 = n16400 & n39319 ;
  assign n39322 = ~n15239 & n39321 ;
  assign n39323 = ~n39320 & ~n39322 ;
  assign n39324 = ~n39318 & n39323 ;
  assign n39325 = \b[52]  & n9301 ;
  assign n39326 = n9298 & n39325 ;
  assign n39327 = ~\a[39]  & \b[53]  ;
  assign n39328 = n8751 & n39327 ;
  assign n39329 = ~n39326 & ~n39328 ;
  assign n39330 = \b[54]  & n8757 ;
  assign n39331 = \a[39]  & \b[53]  ;
  assign n39332 = n8748 & n39331 ;
  assign n39333 = \a[41]  & ~n39332 ;
  assign n39334 = ~n39330 & n39333 ;
  assign n39335 = n39329 & n39334 ;
  assign n39336 = n39324 & n39335 ;
  assign n39337 = ~n39330 & ~n39332 ;
  assign n39338 = n39329 & n39337 ;
  assign n39339 = n39324 & n39338 ;
  assign n39340 = ~\a[41]  & ~n39339 ;
  assign n39341 = ~n39336 & ~n39340 ;
  assign n39342 = n38908 & n38910 ;
  assign n39343 = n38941 & ~n39342 ;
  assign n39344 = n39341 & n39343 ;
  assign n39345 = ~n39316 & n39344 ;
  assign n39346 = n39341 & ~n39343 ;
  assign n39347 = n39316 & n39346 ;
  assign n39348 = ~n39345 & ~n39347 ;
  assign n39349 = ~n39341 & ~n39343 ;
  assign n39350 = ~n39316 & n39349 ;
  assign n39351 = ~n39341 & n39343 ;
  assign n39352 = n39316 & n39351 ;
  assign n39353 = ~n39350 & ~n39352 ;
  assign n39354 = n39348 & n39353 ;
  assign n39355 = n38701 & ~n38947 ;
  assign n39356 = ~n38948 & ~n39355 ;
  assign n39357 = n7534 & ~n17690 ;
  assign n39358 = ~n17688 & n39357 ;
  assign n39359 = \b[55]  & n7973 ;
  assign n39360 = n7970 & n39359 ;
  assign n39361 = ~\a[36]  & \b[56]  ;
  assign n39362 = n7526 & n39361 ;
  assign n39363 = ~n39360 & ~n39362 ;
  assign n39364 = \b[57]  & n7532 ;
  assign n39365 = \a[36]  & \b[56]  ;
  assign n39366 = n17801 & n39365 ;
  assign n39367 = \a[38]  & ~n39366 ;
  assign n39368 = ~n39364 & n39367 ;
  assign n39369 = n39363 & n39368 ;
  assign n39370 = ~n39358 & n39369 ;
  assign n39371 = ~n39364 & ~n39366 ;
  assign n39372 = n39363 & n39371 ;
  assign n39373 = ~n39358 & n39372 ;
  assign n39374 = ~\a[38]  & ~n39373 ;
  assign n39375 = ~n39370 & ~n39374 ;
  assign n39376 = n39356 & ~n39375 ;
  assign n39377 = ~n39354 & n39376 ;
  assign n39378 = ~n39356 & ~n39375 ;
  assign n39379 = n39354 & n39378 ;
  assign n39380 = ~n39377 & ~n39379 ;
  assign n39381 = ~n39356 & n39375 ;
  assign n39382 = ~n39354 & n39381 ;
  assign n39383 = n39356 & n39375 ;
  assign n39384 = n39354 & n39383 ;
  assign n39385 = ~n39382 & ~n39384 ;
  assign n39386 = n39380 & n39385 ;
  assign n39387 = n39066 & ~n39386 ;
  assign n39388 = ~n39066 & n39386 ;
  assign n39389 = ~n39387 & ~n39388 ;
  assign n39390 = n6309 & n20260 ;
  assign n39391 = ~n20257 & n39390 ;
  assign n39392 = n6309 & ~n20260 ;
  assign n39393 = ~n19545 & n39392 ;
  assign n39394 = ~n20256 & n39393 ;
  assign n39395 = \b[58]  & n6778 ;
  assign n39396 = n6775 & n39395 ;
  assign n39397 = ~\a[33]  & \b[59]  ;
  assign n39398 = n6301 & n39397 ;
  assign n39399 = ~n39396 & ~n39398 ;
  assign n39400 = \b[60]  & n6307 ;
  assign n39401 = \a[33]  & \b[59]  ;
  assign n39402 = n6298 & n39401 ;
  assign n39403 = \a[35]  & ~n39402 ;
  assign n39404 = ~n39400 & n39403 ;
  assign n39405 = n39399 & n39404 ;
  assign n39406 = ~n39394 & n39405 ;
  assign n39407 = ~n39391 & n39406 ;
  assign n39408 = ~n39400 & ~n39402 ;
  assign n39409 = n39399 & n39408 ;
  assign n39410 = ~n39394 & n39409 ;
  assign n39411 = ~n39391 & n39410 ;
  assign n39412 = ~\a[35]  & ~n39411 ;
  assign n39413 = ~n39407 & ~n39412 ;
  assign n39414 = n39389 & ~n39413 ;
  assign n39415 = ~n39389 & n39413 ;
  assign n39416 = ~n39414 & ~n39415 ;
  assign n39417 = ~n38990 & ~n38994 ;
  assign n39418 = n38990 & n38994 ;
  assign n39419 = n39013 & ~n39418 ;
  assign n39420 = ~n39417 & ~n39419 ;
  assign n39421 = ~n39416 & ~n39420 ;
  assign n39422 = n39416 & n39420 ;
  assign n39423 = ~n39421 & ~n39422 ;
  assign n39424 = n38681 & ~n39024 ;
  assign n39425 = n38675 & n38681 ;
  assign n39426 = ~n39424 & ~n39425 ;
  assign n39427 = ~n4909 & ~n5208 ;
  assign n39428 = ~n22461 & n39427 ;
  assign n39429 = ~n22459 & n39428 ;
  assign n39430 = \b[61]  & n5595 ;
  assign n39431 = n5592 & n39430 ;
  assign n39432 = ~\a[30]  & \b[62]  ;
  assign n39433 = n5203 & n39432 ;
  assign n39434 = ~n39431 & ~n39433 ;
  assign n39435 = \b[63]  & n5209 ;
  assign n39436 = \a[30]  & \b[62]  ;
  assign n39437 = n5200 & n39436 ;
  assign n39438 = \a[32]  & ~n39437 ;
  assign n39439 = ~n39435 & n39438 ;
  assign n39440 = n39434 & n39439 ;
  assign n39441 = ~n39429 & n39440 ;
  assign n39442 = ~n39435 & ~n39437 ;
  assign n39443 = n39434 & n39442 ;
  assign n39444 = ~n39429 & n39443 ;
  assign n39445 = ~\a[32]  & ~n39444 ;
  assign n39446 = ~n39441 & ~n39445 ;
  assign n39447 = n39426 & ~n39446 ;
  assign n39448 = ~n39426 & n39446 ;
  assign n39449 = ~n39447 & ~n39448 ;
  assign n39450 = ~n39423 & ~n39449 ;
  assign n39451 = n39423 & n39449 ;
  assign n39452 = ~n39450 & ~n39451 ;
  assign n39453 = ~n39064 & n39452 ;
  assign n39454 = n39064 & ~n39452 ;
  assign n39455 = ~n39453 & ~n39454 ;
  assign n39456 = ~n39063 & n39455 ;
  assign n39457 = ~n39055 & ~n39455 ;
  assign n39458 = ~n39059 & n39457 ;
  assign n39459 = ~n39456 & ~n39458 ;
  assign n39460 = ~n39055 & ~n39453 ;
  assign n39461 = ~n39059 & n39460 ;
  assign n39462 = ~n39423 & ~n39447 ;
  assign n39463 = ~n39448 & ~n39462 ;
  assign n39464 = ~n39414 & ~n39420 ;
  assign n39465 = ~n4909 & ~n22458 ;
  assign n39466 = ~n5208 & n39465 ;
  assign n39467 = ~n23173 & n39466 ;
  assign n39468 = \b[62]  & n5595 ;
  assign n39469 = n5592 & n39468 ;
  assign n39470 = \a[30]  & \b[63]  ;
  assign n39471 = n5200 & n39470 ;
  assign n39472 = ~\a[30]  & \b[63]  ;
  assign n39473 = n5203 & n39472 ;
  assign n39474 = \a[32]  & ~n39473 ;
  assign n39475 = ~n39471 & n39474 ;
  assign n39476 = ~n39469 & n39475 ;
  assign n39477 = ~n39467 & n39476 ;
  assign n39478 = ~n39471 & ~n39473 ;
  assign n39479 = ~n39469 & n39478 ;
  assign n39480 = ~n39467 & n39479 ;
  assign n39481 = ~\a[32]  & ~n39480 ;
  assign n39482 = ~n39477 & ~n39481 ;
  assign n39483 = ~n39415 & ~n39482 ;
  assign n39484 = ~n39464 & n39483 ;
  assign n39485 = ~n39415 & ~n39464 ;
  assign n39486 = n39482 & ~n39485 ;
  assign n39487 = ~n39484 & ~n39486 ;
  assign n39488 = n39066 & n39380 ;
  assign n39489 = n39385 & ~n39488 ;
  assign n39490 = ~n39241 & ~n39250 ;
  assign n39491 = n39246 & ~n39490 ;
  assign n39492 = ~n39090 & n39165 ;
  assign n39493 = n39184 & ~n39492 ;
  assign n39494 = ~n9044 & ~n16016 ;
  assign n39495 = ~n16652 & n39494 ;
  assign n39496 = n9041 & n39495 ;
  assign n39497 = n9044 & ~n16016 ;
  assign n39498 = ~n16652 & n39497 ;
  assign n39499 = ~n9041 & n39498 ;
  assign n39500 = ~n39496 & ~n39499 ;
  assign n39501 = \b[38]  & n17308 ;
  assign n39502 = n17305 & n39501 ;
  assign n39503 = ~\a[54]  & \b[39]  ;
  assign n39504 = n16647 & n39503 ;
  assign n39505 = ~n39502 & ~n39504 ;
  assign n39506 = \b[40]  & n16653 ;
  assign n39507 = \a[54]  & \b[39]  ;
  assign n39508 = n16644 & n39507 ;
  assign n39509 = \a[56]  & ~n39508 ;
  assign n39510 = ~n39506 & n39509 ;
  assign n39511 = n39505 & n39510 ;
  assign n39512 = n39500 & n39511 ;
  assign n39513 = ~n39506 & ~n39508 ;
  assign n39514 = n39505 & n39513 ;
  assign n39515 = n39500 & n39514 ;
  assign n39516 = ~\a[56]  & ~n39515 ;
  assign n39517 = ~n39512 & ~n39516 ;
  assign n39518 = ~n39095 & ~n39160 ;
  assign n39519 = ~n39161 & ~n39518 ;
  assign n39520 = ~n7758 & n18516 ;
  assign n39521 = ~n7336 & n18516 ;
  assign n39522 = ~n7754 & n39521 ;
  assign n39523 = ~n39520 & ~n39522 ;
  assign n39524 = ~n7761 & ~n39523 ;
  assign n39525 = \b[37]  & n18514 ;
  assign n39526 = \a[56]  & \b[36]  ;
  assign n39527 = n19181 & n39526 ;
  assign n39528 = ~\a[57]  & \b[36]  ;
  assign n39529 = n18508 & n39528 ;
  assign n39530 = ~n39527 & ~n39529 ;
  assign n39531 = ~n39525 & n39530 ;
  assign n39532 = \b[35]  & n19183 ;
  assign n39533 = n19180 & n39532 ;
  assign n39534 = \a[59]  & ~n39533 ;
  assign n39535 = n39531 & n39534 ;
  assign n39536 = ~n39524 & n39535 ;
  assign n39537 = n39531 & ~n39533 ;
  assign n39538 = ~\a[59]  & ~n39537 ;
  assign n39539 = ~\a[59]  & ~n7761 ;
  assign n39540 = ~n39523 & n39539 ;
  assign n39541 = ~n39538 & ~n39540 ;
  assign n39542 = ~n39536 & n39541 ;
  assign n39543 = n39135 & ~n39153 ;
  assign n39544 = ~n39155 & ~n39543 ;
  assign n39545 = ~n6565 & ~n19861 ;
  assign n39546 = ~n20518 & n39545 ;
  assign n39547 = n6562 & n39546 ;
  assign n39548 = n6565 & ~n19861 ;
  assign n39549 = ~n20518 & n39548 ;
  assign n39550 = ~n6562 & n39549 ;
  assign n39551 = ~n39547 & ~n39550 ;
  assign n39552 = \b[34]  & n20519 ;
  assign n39553 = \a[60]  & \b[33]  ;
  assign n39554 = n20510 & n39553 ;
  assign n39555 = ~n39552 & ~n39554 ;
  assign n39556 = \b[32]  & n21315 ;
  assign n39557 = n21312 & n39556 ;
  assign n39558 = ~\a[60]  & \b[33]  ;
  assign n39559 = n20513 & n39558 ;
  assign n39560 = ~n39557 & ~n39559 ;
  assign n39561 = n39555 & n39560 ;
  assign n39562 = n39551 & n39561 ;
  assign n39563 = ~\a[62]  & ~n39562 ;
  assign n39564 = ~n38751 & ~n39147 ;
  assign n39565 = \b[31]  & n21958 ;
  assign n39566 = \b[30]  & n21957 ;
  assign n39567 = ~n39565 & ~n39566 ;
  assign n39568 = n39143 & ~n39567 ;
  assign n39569 = ~n39564 & n39568 ;
  assign n39570 = n39143 & ~n39564 ;
  assign n39571 = n39567 & ~n39570 ;
  assign n39572 = ~n39569 & ~n39571 ;
  assign n39573 = \a[62]  & ~n39554 ;
  assign n39574 = ~n39552 & n39573 ;
  assign n39575 = n39560 & n39574 ;
  assign n39576 = n39551 & n39575 ;
  assign n39577 = ~n39572 & ~n39576 ;
  assign n39578 = ~n39563 & n39577 ;
  assign n39579 = ~\a[62]  & n39572 ;
  assign n39580 = ~n39562 & n39579 ;
  assign n39581 = \a[62]  & n39572 ;
  assign n39582 = n39562 & n39581 ;
  assign n39583 = ~n39580 & ~n39582 ;
  assign n39584 = ~n39578 & n39583 ;
  assign n39585 = n39544 & n39584 ;
  assign n39586 = ~n39544 & ~n39584 ;
  assign n39587 = ~n39585 & ~n39586 ;
  assign n39588 = n39542 & n39587 ;
  assign n39589 = ~n39542 & ~n39587 ;
  assign n39590 = ~n39588 & ~n39589 ;
  assign n39591 = n39519 & ~n39590 ;
  assign n39592 = ~n39519 & n39590 ;
  assign n39593 = ~n39591 & ~n39592 ;
  assign n39594 = ~n39517 & n39593 ;
  assign n39595 = n39517 & ~n39593 ;
  assign n39596 = ~n39594 & ~n39595 ;
  assign n39597 = ~n39493 & n39596 ;
  assign n39598 = n39493 & ~n39596 ;
  assign n39599 = ~n39597 & ~n39598 ;
  assign n39600 = ~n10406 & n14793 ;
  assign n39601 = ~n9929 & n14793 ;
  assign n39602 = ~n10402 & n39601 ;
  assign n39603 = ~n39600 & ~n39602 ;
  assign n39604 = ~n10409 & ~n39603 ;
  assign n39605 = \b[41]  & n15517 ;
  assign n39606 = n15514 & n39605 ;
  assign n39607 = ~\a[51]  & \b[42]  ;
  assign n39608 = n14785 & n39607 ;
  assign n39609 = ~n39606 & ~n39608 ;
  assign n39610 = \b[43]  & n14791 ;
  assign n39611 = \a[51]  & \b[42]  ;
  assign n39612 = n14782 & n39611 ;
  assign n39613 = \a[53]  & ~n39612 ;
  assign n39614 = ~n39610 & n39613 ;
  assign n39615 = n39609 & n39614 ;
  assign n39616 = ~n39604 & n39615 ;
  assign n39617 = ~n39610 & ~n39612 ;
  assign n39618 = n39609 & n39617 ;
  assign n39619 = ~\a[53]  & ~n39618 ;
  assign n39620 = ~\a[53]  & ~n10409 ;
  assign n39621 = ~n39603 & n39620 ;
  assign n39622 = ~n39619 & ~n39621 ;
  assign n39623 = ~n39616 & n39622 ;
  assign n39624 = n39599 & ~n39623 ;
  assign n39625 = ~n39599 & n39623 ;
  assign n39626 = ~n39624 & ~n39625 ;
  assign n39627 = ~n39210 & ~n39217 ;
  assign n39628 = ~n39212 & ~n39627 ;
  assign n39629 = n11906 & n13125 ;
  assign n39630 = ~n11903 & n39629 ;
  assign n39631 = ~n11906 & n13125 ;
  assign n39632 = ~n11392 & n39631 ;
  assign n39633 = ~n11902 & n39632 ;
  assign n39634 = \b[44]  & n13794 ;
  assign n39635 = n13792 & n39634 ;
  assign n39636 = ~\a[48]  & \b[45]  ;
  assign n39637 = n13117 & n39636 ;
  assign n39638 = ~n39635 & ~n39637 ;
  assign n39639 = \b[46]  & n13123 ;
  assign n39640 = \a[48]  & \b[45]  ;
  assign n39641 = n13786 & n39640 ;
  assign n39642 = \a[50]  & ~n39641 ;
  assign n39643 = ~n39639 & n39642 ;
  assign n39644 = n39638 & n39643 ;
  assign n39645 = ~n39633 & n39644 ;
  assign n39646 = ~n39630 & n39645 ;
  assign n39647 = ~n39639 & ~n39641 ;
  assign n39648 = n39638 & n39647 ;
  assign n39649 = ~n39633 & n39648 ;
  assign n39650 = ~n39630 & n39649 ;
  assign n39651 = ~\a[50]  & ~n39650 ;
  assign n39652 = ~n39646 & ~n39651 ;
  assign n39653 = ~n39628 & n39652 ;
  assign n39654 = ~n39626 & n39653 ;
  assign n39655 = n39628 & n39652 ;
  assign n39656 = n39626 & n39655 ;
  assign n39657 = ~n39654 & ~n39656 ;
  assign n39658 = n39628 & ~n39652 ;
  assign n39659 = ~n39626 & n39658 ;
  assign n39660 = ~n39628 & ~n39652 ;
  assign n39661 = n39626 & n39660 ;
  assign n39662 = ~n39659 & ~n39661 ;
  assign n39663 = n39657 & n39662 ;
  assign n39664 = ~n39491 & ~n39663 ;
  assign n39665 = n39491 & n39663 ;
  assign n39666 = ~n39664 & ~n39665 ;
  assign n39667 = n11572 & ~n13524 ;
  assign n39668 = ~n13522 & n39667 ;
  assign n39669 = \b[47]  & n12159 ;
  assign n39670 = n12156 & n39669 ;
  assign n39671 = ~\a[45]  & \b[48]  ;
  assign n39672 = n11564 & n39671 ;
  assign n39673 = ~n39670 & ~n39672 ;
  assign n39674 = \b[49]  & n11570 ;
  assign n39675 = \a[45]  & \b[48]  ;
  assign n39676 = n11561 & n39675 ;
  assign n39677 = \a[47]  & ~n39676 ;
  assign n39678 = ~n39674 & n39677 ;
  assign n39679 = n39673 & n39678 ;
  assign n39680 = ~n39668 & n39679 ;
  assign n39681 = ~n39674 & ~n39676 ;
  assign n39682 = n39673 & n39681 ;
  assign n39683 = ~n39668 & n39682 ;
  assign n39684 = ~\a[47]  & ~n39683 ;
  assign n39685 = ~n39680 & ~n39684 ;
  assign n39686 = n39666 & ~n39685 ;
  assign n39687 = ~n39666 & n39685 ;
  assign n39688 = ~n39686 & ~n39687 ;
  assign n39689 = n39278 & ~n39288 ;
  assign n39690 = n39283 & ~n39689 ;
  assign n39691 = n10082 & n15201 ;
  assign n39692 = ~n15198 & n39691 ;
  assign n39693 = n10082 & n28871 ;
  assign n39694 = ~n15197 & n39693 ;
  assign n39695 = \b[50]  & n10681 ;
  assign n39696 = n10678 & n39695 ;
  assign n39697 = \b[52]  & n10080 ;
  assign n39698 = \a[41]  & \b[51]  ;
  assign n39699 = n10679 & n39698 ;
  assign n39700 = ~\a[42]  & \b[51]  ;
  assign n39701 = n10074 & n39700 ;
  assign n39702 = ~n39699 & ~n39701 ;
  assign n39703 = ~n39697 & n39702 ;
  assign n39704 = ~n39696 & n39703 ;
  assign n39705 = ~n39694 & n39704 ;
  assign n39706 = ~n39692 & n39705 ;
  assign n39707 = ~\a[44]  & ~n39706 ;
  assign n39708 = \a[44]  & n39704 ;
  assign n39709 = ~n39694 & n39708 ;
  assign n39710 = ~n39692 & n39709 ;
  assign n39711 = ~n39707 & ~n39710 ;
  assign n39712 = ~n39690 & n39711 ;
  assign n39713 = ~n39688 & n39712 ;
  assign n39714 = n39690 & n39711 ;
  assign n39715 = n39688 & n39714 ;
  assign n39716 = ~n39713 & ~n39715 ;
  assign n39717 = n39690 & ~n39711 ;
  assign n39718 = ~n39688 & n39717 ;
  assign n39719 = ~n39690 & ~n39711 ;
  assign n39720 = n39688 & n39719 ;
  assign n39721 = ~n39718 & ~n39720 ;
  assign n39722 = n39716 & n39721 ;
  assign n39723 = n8759 & ~n16446 ;
  assign n39724 = ~n16444 & n39723 ;
  assign n39725 = \b[53]  & n9301 ;
  assign n39726 = n9298 & n39725 ;
  assign n39727 = ~\a[39]  & \b[54]  ;
  assign n39728 = n8751 & n39727 ;
  assign n39729 = ~n39726 & ~n39728 ;
  assign n39730 = \b[55]  & n8757 ;
  assign n39731 = \a[39]  & \b[54]  ;
  assign n39732 = n8748 & n39731 ;
  assign n39733 = \a[41]  & ~n39732 ;
  assign n39734 = ~n39730 & n39733 ;
  assign n39735 = n39729 & n39734 ;
  assign n39736 = ~n39724 & n39735 ;
  assign n39737 = ~n39730 & ~n39732 ;
  assign n39738 = n39729 & n39737 ;
  assign n39739 = ~n39724 & n39738 ;
  assign n39740 = ~\a[41]  & ~n39739 ;
  assign n39741 = ~n39736 & ~n39740 ;
  assign n39742 = n39315 & n39343 ;
  assign n39743 = n39310 & ~n39742 ;
  assign n39744 = n39741 & ~n39743 ;
  assign n39745 = n39722 & n39744 ;
  assign n39746 = n39741 & n39743 ;
  assign n39747 = ~n39722 & n39746 ;
  assign n39748 = ~n39745 & ~n39747 ;
  assign n39749 = ~n39741 & ~n39743 ;
  assign n39750 = ~n39722 & n39749 ;
  assign n39751 = ~n39741 & n39743 ;
  assign n39752 = n39722 & n39751 ;
  assign n39753 = ~n39750 & ~n39752 ;
  assign n39754 = n39748 & n39753 ;
  assign n39755 = n39353 & ~n39356 ;
  assign n39756 = n39348 & ~n39755 ;
  assign n39757 = n7534 & ~n19543 ;
  assign n39758 = ~n38598 & n39757 ;
  assign n39759 = \b[56]  & n7973 ;
  assign n39760 = n7970 & n39759 ;
  assign n39761 = ~\a[36]  & \b[57]  ;
  assign n39762 = n7526 & n39761 ;
  assign n39763 = ~n39760 & ~n39762 ;
  assign n39764 = \b[58]  & n7532 ;
  assign n39765 = \a[36]  & \b[57]  ;
  assign n39766 = n17801 & n39765 ;
  assign n39767 = \a[38]  & ~n39766 ;
  assign n39768 = ~n39764 & n39767 ;
  assign n39769 = n39763 & n39768 ;
  assign n39770 = ~n39758 & n39769 ;
  assign n39771 = ~n39764 & ~n39766 ;
  assign n39772 = n39763 & n39771 ;
  assign n39773 = ~n39758 & n39772 ;
  assign n39774 = ~\a[38]  & ~n39773 ;
  assign n39775 = ~n39770 & ~n39774 ;
  assign n39776 = ~n39756 & ~n39775 ;
  assign n39777 = ~n39754 & n39776 ;
  assign n39778 = n39756 & ~n39775 ;
  assign n39779 = n39754 & n39778 ;
  assign n39780 = ~n39777 & ~n39779 ;
  assign n39781 = n39756 & n39775 ;
  assign n39782 = ~n39754 & n39781 ;
  assign n39783 = ~n39756 & n39775 ;
  assign n39784 = n39754 & n39783 ;
  assign n39785 = ~n39782 & ~n39784 ;
  assign n39786 = n39780 & n39785 ;
  assign n39787 = ~n39489 & ~n39786 ;
  assign n39788 = n39489 & n39786 ;
  assign n39789 = ~n39787 & ~n39788 ;
  assign n39790 = n6309 & ~n20971 ;
  assign n39791 = ~n20969 & n39790 ;
  assign n39792 = \b[59]  & n6778 ;
  assign n39793 = n6775 & n39792 ;
  assign n39794 = ~\a[33]  & \b[60]  ;
  assign n39795 = n6301 & n39794 ;
  assign n39796 = ~n39793 & ~n39795 ;
  assign n39797 = \b[61]  & n6307 ;
  assign n39798 = \a[33]  & \b[60]  ;
  assign n39799 = n6298 & n39798 ;
  assign n39800 = \a[35]  & ~n39799 ;
  assign n39801 = ~n39797 & n39800 ;
  assign n39802 = n39796 & n39801 ;
  assign n39803 = ~n39791 & n39802 ;
  assign n39804 = ~n39797 & ~n39799 ;
  assign n39805 = n39796 & n39804 ;
  assign n39806 = ~n39791 & n39805 ;
  assign n39807 = ~\a[35]  & ~n39806 ;
  assign n39808 = ~n39803 & ~n39807 ;
  assign n39809 = n39789 & ~n39808 ;
  assign n39810 = ~n39789 & n39808 ;
  assign n39811 = ~n39809 & ~n39810 ;
  assign n39812 = n39487 & n39811 ;
  assign n39813 = ~n39487 & ~n39811 ;
  assign n39814 = ~n39812 & ~n39813 ;
  assign n39815 = n39463 & n39814 ;
  assign n39816 = ~n39463 & ~n39814 ;
  assign n39817 = ~n39815 & ~n39816 ;
  assign n39818 = ~n39454 & n39817 ;
  assign n39819 = ~n39461 & n39818 ;
  assign n39820 = ~n39454 & ~n39461 ;
  assign n39821 = ~n39817 & ~n39820 ;
  assign n39822 = ~n39819 & ~n39821 ;
  assign n39823 = ~n39815 & ~n39819 ;
  assign n39824 = ~n39484 & ~n39811 ;
  assign n39825 = ~n39486 & ~n39824 ;
  assign n39826 = ~n39788 & n39808 ;
  assign n39827 = ~n5208 & n39033 ;
  assign n39828 = ~n23171 & n39827 ;
  assign n39829 = ~n4909 & n39828 ;
  assign n39830 = \a[29]  & \a[31]  ;
  assign n39831 = \a[30]  & ~\a[32]  ;
  assign n39832 = n39830 & n39831 ;
  assign n39833 = ~\a[29]  & ~\a[31]  ;
  assign n39834 = ~\a[30]  & \a[32]  ;
  assign n39835 = n39833 & n39834 ;
  assign n39836 = ~n39832 & ~n39835 ;
  assign n39837 = \b[63]  & ~n39836 ;
  assign n39838 = \a[32]  & ~n39837 ;
  assign n39839 = ~n39829 & n39838 ;
  assign n39840 = ~\a[32]  & n39837 ;
  assign n39841 = ~\a[32]  & ~n4909 ;
  assign n39842 = n39828 & n39841 ;
  assign n39843 = ~n39840 & ~n39842 ;
  assign n39844 = ~n39839 & n39843 ;
  assign n39845 = ~n39787 & ~n39844 ;
  assign n39846 = ~n39826 & n39845 ;
  assign n39847 = ~n39787 & ~n39826 ;
  assign n39848 = n39844 & ~n39847 ;
  assign n39849 = ~n39846 & ~n39848 ;
  assign n39850 = ~n39722 & ~n39743 ;
  assign n39851 = n39722 & n39743 ;
  assign n39852 = n39741 & ~n39851 ;
  assign n39853 = ~n39850 & ~n39852 ;
  assign n39854 = ~n10889 & ~n14276 ;
  assign n39855 = ~n14790 & n39854 ;
  assign n39856 = n10886 & n39855 ;
  assign n39857 = n10889 & ~n14276 ;
  assign n39858 = ~n14790 & n39857 ;
  assign n39859 = ~n10886 & n39858 ;
  assign n39860 = ~n39856 & ~n39859 ;
  assign n39861 = \b[42]  & n15517 ;
  assign n39862 = n15514 & n39861 ;
  assign n39863 = ~\a[51]  & \b[43]  ;
  assign n39864 = n14785 & n39863 ;
  assign n39865 = ~n39862 & ~n39864 ;
  assign n39866 = \b[44]  & n14791 ;
  assign n39867 = \a[51]  & \b[43]  ;
  assign n39868 = n14782 & n39867 ;
  assign n39869 = \a[53]  & ~n39868 ;
  assign n39870 = ~n39866 & n39869 ;
  assign n39871 = n39865 & n39870 ;
  assign n39872 = n39860 & n39871 ;
  assign n39873 = ~n39866 & ~n39868 ;
  assign n39874 = n39865 & n39873 ;
  assign n39875 = n39860 & n39874 ;
  assign n39876 = ~\a[53]  & ~n39875 ;
  assign n39877 = ~n39872 & ~n39876 ;
  assign n39878 = n39517 & ~n39591 ;
  assign n39879 = ~n39591 & n39592 ;
  assign n39880 = ~n39878 & ~n39879 ;
  assign n39881 = ~n9479 & n37945 ;
  assign n39882 = ~n9043 & n37945 ;
  assign n39883 = ~n9475 & n39882 ;
  assign n39884 = ~n39881 & ~n39883 ;
  assign n39885 = ~n9482 & ~n39884 ;
  assign n39886 = \b[39]  & n17308 ;
  assign n39887 = n17305 & n39886 ;
  assign n39888 = ~\a[54]  & \b[40]  ;
  assign n39889 = n16647 & n39888 ;
  assign n39890 = ~n39887 & ~n39889 ;
  assign n39891 = \b[41]  & n16653 ;
  assign n39892 = \a[54]  & \b[40]  ;
  assign n39893 = n16644 & n39892 ;
  assign n39894 = \a[56]  & ~n39893 ;
  assign n39895 = ~n39891 & n39894 ;
  assign n39896 = n39890 & n39895 ;
  assign n39897 = ~n39885 & n39896 ;
  assign n39898 = ~n39891 & ~n39893 ;
  assign n39899 = n39890 & n39898 ;
  assign n39900 = ~\a[56]  & ~n39899 ;
  assign n39901 = ~\a[56]  & ~n9482 ;
  assign n39902 = ~n39884 & n39901 ;
  assign n39903 = ~n39900 & ~n39902 ;
  assign n39904 = ~n39897 & n39903 ;
  assign n39905 = ~n6610 & n20521 ;
  assign n39906 = ~n6608 & n39905 ;
  assign n39907 = \b[33]  & n21315 ;
  assign n39908 = n21312 & n39907 ;
  assign n39909 = ~\a[60]  & \b[34]  ;
  assign n39910 = n20513 & n39909 ;
  assign n39911 = ~n39908 & ~n39910 ;
  assign n39912 = \b[35]  & n20519 ;
  assign n39913 = \a[60]  & \b[34]  ;
  assign n39914 = n20510 & n39913 ;
  assign n39915 = \a[62]  & ~n39914 ;
  assign n39916 = ~n39912 & n39915 ;
  assign n39917 = n39911 & n39916 ;
  assign n39918 = ~n39906 & n39917 ;
  assign n39919 = ~n39912 & ~n39914 ;
  assign n39920 = n39911 & n39919 ;
  assign n39921 = ~n39906 & n39920 ;
  assign n39922 = ~\a[62]  & ~n39921 ;
  assign n39923 = ~n39918 & ~n39922 ;
  assign n39924 = ~\a[62]  & ~n39569 ;
  assign n39925 = ~n39562 & n39924 ;
  assign n39926 = \a[62]  & ~n39569 ;
  assign n39927 = n39562 & n39926 ;
  assign n39928 = ~n39925 & ~n39927 ;
  assign n39929 = \b[32]  & n21958 ;
  assign n39930 = \b[31]  & n21957 ;
  assign n39931 = ~n39929 & ~n39930 ;
  assign n39932 = ~n39567 & n39931 ;
  assign n39933 = n39567 & ~n39931 ;
  assign n39934 = ~n39932 & ~n39933 ;
  assign n39935 = ~n39571 & n39934 ;
  assign n39936 = n39928 & n39935 ;
  assign n39937 = ~n39571 & n39924 ;
  assign n39938 = ~n39562 & n39937 ;
  assign n39939 = ~n39571 & n39926 ;
  assign n39940 = n39562 & n39939 ;
  assign n39941 = ~n39938 & ~n39940 ;
  assign n39942 = ~n39571 & n39941 ;
  assign n39943 = ~n39934 & ~n39942 ;
  assign n39944 = ~n39936 & ~n39943 ;
  assign n39945 = ~n39923 & ~n39944 ;
  assign n39946 = n39923 & ~n39936 ;
  assign n39947 = ~n39943 & n39946 ;
  assign n39948 = ~n39945 & ~n39947 ;
  assign n39949 = n39542 & ~n39585 ;
  assign n39950 = ~n39586 & ~n39949 ;
  assign n39951 = n8175 & n18516 ;
  assign n39952 = ~n8172 & n39951 ;
  assign n39953 = n18516 & n25622 ;
  assign n39954 = ~n8171 & n39953 ;
  assign n39955 = \b[38]  & n18514 ;
  assign n39956 = \a[56]  & \b[37]  ;
  assign n39957 = n19181 & n39956 ;
  assign n39958 = ~\a[57]  & \b[37]  ;
  assign n39959 = n18508 & n39958 ;
  assign n39960 = ~n39957 & ~n39959 ;
  assign n39961 = ~n39955 & n39960 ;
  assign n39962 = \b[36]  & n19183 ;
  assign n39963 = n19180 & n39962 ;
  assign n39964 = \a[59]  & ~n39963 ;
  assign n39965 = n39961 & n39964 ;
  assign n39966 = ~n39954 & n39965 ;
  assign n39967 = ~n39952 & n39966 ;
  assign n39968 = n39961 & ~n39963 ;
  assign n39969 = ~n39954 & n39968 ;
  assign n39970 = ~n39952 & n39969 ;
  assign n39971 = ~\a[59]  & ~n39970 ;
  assign n39972 = ~n39967 & ~n39971 ;
  assign n39973 = n39950 & ~n39972 ;
  assign n39974 = ~n39948 & n39973 ;
  assign n39975 = n39950 & n39972 ;
  assign n39976 = n39948 & n39975 ;
  assign n39977 = ~n39974 & ~n39976 ;
  assign n39978 = ~n39948 & ~n39972 ;
  assign n39979 = ~n39947 & n39972 ;
  assign n39980 = ~n39945 & n39979 ;
  assign n39981 = ~n39950 & ~n39980 ;
  assign n39982 = ~n39978 & n39981 ;
  assign n39983 = n39977 & ~n39982 ;
  assign n39984 = n39904 & n39983 ;
  assign n39985 = ~n39904 & ~n39983 ;
  assign n39986 = ~n39984 & ~n39985 ;
  assign n39987 = n39880 & ~n39986 ;
  assign n39988 = ~n39880 & n39986 ;
  assign n39989 = ~n39987 & ~n39988 ;
  assign n39990 = ~n39877 & n39989 ;
  assign n39991 = n39877 & ~n39989 ;
  assign n39992 = ~n39990 & ~n39991 ;
  assign n39993 = ~n39597 & n39623 ;
  assign n39994 = ~n39598 & ~n39993 ;
  assign n39995 = ~n12438 & n13125 ;
  assign n39996 = ~n12436 & n39995 ;
  assign n39997 = \b[45]  & n13794 ;
  assign n39998 = n13792 & n39997 ;
  assign n39999 = ~\a[48]  & \b[46]  ;
  assign n40000 = n13117 & n39999 ;
  assign n40001 = ~n39998 & ~n40000 ;
  assign n40002 = \b[47]  & n13123 ;
  assign n40003 = \a[48]  & \b[46]  ;
  assign n40004 = n13786 & n40003 ;
  assign n40005 = \a[50]  & ~n40004 ;
  assign n40006 = ~n40002 & n40005 ;
  assign n40007 = n40001 & n40006 ;
  assign n40008 = ~n39996 & n40007 ;
  assign n40009 = ~n40002 & ~n40004 ;
  assign n40010 = n40001 & n40009 ;
  assign n40011 = ~n39996 & n40010 ;
  assign n40012 = ~\a[50]  & ~n40011 ;
  assign n40013 = ~n40008 & ~n40012 ;
  assign n40014 = ~n39994 & ~n40013 ;
  assign n40015 = n39992 & n40014 ;
  assign n40016 = n39994 & ~n40013 ;
  assign n40017 = ~n39992 & n40016 ;
  assign n40018 = ~n40015 & ~n40017 ;
  assign n40019 = ~n39994 & n40013 ;
  assign n40020 = ~n39992 & n40019 ;
  assign n40021 = n39994 & n40013 ;
  assign n40022 = n39992 & n40021 ;
  assign n40023 = ~n40020 & ~n40022 ;
  assign n40024 = n40018 & n40023 ;
  assign n40025 = ~n39626 & ~n39628 ;
  assign n40026 = n39626 & n39628 ;
  assign n40027 = n39652 & ~n40026 ;
  assign n40028 = ~n40025 & ~n40027 ;
  assign n40029 = ~n10988 & ~n13519 ;
  assign n40030 = ~n14052 & n40029 ;
  assign n40031 = ~n14048 & n40030 ;
  assign n40032 = ~n11569 & n40031 ;
  assign n40033 = n11572 & n14052 ;
  assign n40034 = ~n14049 & n40033 ;
  assign n40035 = ~n40032 & ~n40034 ;
  assign n40036 = \b[48]  & n12159 ;
  assign n40037 = n12156 & n40036 ;
  assign n40038 = ~\a[45]  & \b[49]  ;
  assign n40039 = n11564 & n40038 ;
  assign n40040 = ~n40037 & ~n40039 ;
  assign n40041 = \b[50]  & n11570 ;
  assign n40042 = \a[45]  & \b[49]  ;
  assign n40043 = n11561 & n40042 ;
  assign n40044 = \a[47]  & ~n40043 ;
  assign n40045 = ~n40041 & n40044 ;
  assign n40046 = n40040 & n40045 ;
  assign n40047 = n40035 & n40046 ;
  assign n40048 = ~n40041 & ~n40043 ;
  assign n40049 = n40040 & n40048 ;
  assign n40050 = n40035 & n40049 ;
  assign n40051 = ~\a[47]  & ~n40050 ;
  assign n40052 = ~n40047 & ~n40051 ;
  assign n40053 = ~n40028 & n40052 ;
  assign n40054 = ~n40024 & n40053 ;
  assign n40055 = n40028 & n40052 ;
  assign n40056 = n40024 & n40055 ;
  assign n40057 = ~n40054 & ~n40056 ;
  assign n40058 = ~n40028 & ~n40052 ;
  assign n40059 = n40024 & n40058 ;
  assign n40060 = n40028 & ~n40052 ;
  assign n40061 = ~n40024 & n40060 ;
  assign n40062 = ~n40059 & ~n40061 ;
  assign n40063 = n40057 & n40062 ;
  assign n40064 = n10082 & ~n15246 ;
  assign n40065 = ~n15244 & n40064 ;
  assign n40066 = \b[53]  & n10080 ;
  assign n40067 = \a[41]  & \b[52]  ;
  assign n40068 = n10679 & n40067 ;
  assign n40069 = ~\a[42]  & \b[52]  ;
  assign n40070 = n10074 & n40069 ;
  assign n40071 = ~n40068 & ~n40070 ;
  assign n40072 = ~n40066 & n40071 ;
  assign n40073 = \b[51]  & n10681 ;
  assign n40074 = n10678 & n40073 ;
  assign n40075 = \a[44]  & ~n40074 ;
  assign n40076 = n40072 & n40075 ;
  assign n40077 = ~n40065 & n40076 ;
  assign n40078 = n40072 & ~n40074 ;
  assign n40079 = ~n40065 & n40078 ;
  assign n40080 = ~\a[44]  & ~n40079 ;
  assign n40081 = ~n40077 & ~n40080 ;
  assign n40082 = ~n39665 & n39685 ;
  assign n40083 = ~n39664 & ~n40082 ;
  assign n40084 = n40081 & ~n40083 ;
  assign n40085 = n40063 & n40084 ;
  assign n40086 = n40081 & n40083 ;
  assign n40087 = ~n40063 & n40086 ;
  assign n40088 = ~n40085 & ~n40087 ;
  assign n40089 = ~n40081 & ~n40083 ;
  assign n40090 = ~n40063 & n40089 ;
  assign n40091 = ~n40081 & n40083 ;
  assign n40092 = n40063 & n40091 ;
  assign n40093 = ~n40090 & ~n40092 ;
  assign n40094 = n40088 & n40093 ;
  assign n40095 = n8759 & n17647 ;
  assign n40096 = ~n17644 & n40095 ;
  assign n40097 = n8759 & n19567 ;
  assign n40098 = ~n17643 & n40097 ;
  assign n40099 = \b[54]  & n9301 ;
  assign n40100 = n9298 & n40099 ;
  assign n40101 = ~\a[39]  & \b[55]  ;
  assign n40102 = n8751 & n40101 ;
  assign n40103 = ~n40100 & ~n40102 ;
  assign n40104 = \b[56]  & n8757 ;
  assign n40105 = \a[39]  & \b[55]  ;
  assign n40106 = n8748 & n40105 ;
  assign n40107 = \a[41]  & ~n40106 ;
  assign n40108 = ~n40104 & n40107 ;
  assign n40109 = n40103 & n40108 ;
  assign n40110 = ~n40098 & n40109 ;
  assign n40111 = ~n40096 & n40110 ;
  assign n40112 = ~n40104 & ~n40106 ;
  assign n40113 = n40103 & n40112 ;
  assign n40114 = ~n40098 & n40113 ;
  assign n40115 = ~n40096 & n40114 ;
  assign n40116 = ~\a[41]  & ~n40115 ;
  assign n40117 = ~n40111 & ~n40116 ;
  assign n40118 = ~n39688 & ~n39690 ;
  assign n40119 = ~n39685 & n39711 ;
  assign n40120 = n39666 & n40119 ;
  assign n40121 = n39685 & n39711 ;
  assign n40122 = ~n39666 & n40121 ;
  assign n40123 = ~n40120 & ~n40122 ;
  assign n40124 = ~n39712 & n40123 ;
  assign n40125 = ~n40118 & n40124 ;
  assign n40126 = ~n40117 & ~n40125 ;
  assign n40127 = ~n40094 & n40126 ;
  assign n40128 = ~n40117 & n40125 ;
  assign n40129 = n40094 & n40128 ;
  assign n40130 = ~n40127 & ~n40129 ;
  assign n40131 = n40117 & ~n40125 ;
  assign n40132 = n40094 & n40131 ;
  assign n40133 = n40117 & n40125 ;
  assign n40134 = ~n40094 & n40133 ;
  assign n40135 = ~n40132 & ~n40134 ;
  assign n40136 = n40130 & n40135 ;
  assign n40137 = n39853 & n40136 ;
  assign n40138 = ~n39853 & ~n40136 ;
  assign n40139 = ~n40137 & ~n40138 ;
  assign n40140 = n7534 & ~n19550 ;
  assign n40141 = ~n19548 & n40140 ;
  assign n40142 = \b[57]  & n7973 ;
  assign n40143 = n7970 & n40142 ;
  assign n40144 = ~\a[36]  & \b[58]  ;
  assign n40145 = n7526 & n40144 ;
  assign n40146 = ~n40143 & ~n40145 ;
  assign n40147 = \b[59]  & n7532 ;
  assign n40148 = \a[36]  & \b[58]  ;
  assign n40149 = n17801 & n40148 ;
  assign n40150 = \a[38]  & ~n40149 ;
  assign n40151 = ~n40147 & n40150 ;
  assign n40152 = n40146 & n40151 ;
  assign n40153 = ~n40141 & n40152 ;
  assign n40154 = ~n40147 & ~n40149 ;
  assign n40155 = n40146 & n40154 ;
  assign n40156 = ~n40141 & n40155 ;
  assign n40157 = ~\a[38]  & ~n40156 ;
  assign n40158 = ~n40153 & ~n40157 ;
  assign n40159 = n40139 & ~n40158 ;
  assign n40160 = ~n40139 & n40158 ;
  assign n40161 = ~n40159 & ~n40160 ;
  assign n40162 = n39754 & ~n39756 ;
  assign n40163 = ~n39754 & n39756 ;
  assign n40164 = n39775 & ~n40163 ;
  assign n40165 = ~n40162 & ~n40164 ;
  assign n40166 = ~n5952 & ~n20966 ;
  assign n40167 = ~n21696 & n40166 ;
  assign n40168 = ~n21692 & n40167 ;
  assign n40169 = ~n6306 & n40168 ;
  assign n40170 = n6309 & n21696 ;
  assign n40171 = ~n21693 & n40170 ;
  assign n40172 = ~n40169 & ~n40171 ;
  assign n40173 = \b[60]  & n6778 ;
  assign n40174 = n6775 & n40173 ;
  assign n40175 = ~\a[33]  & \b[61]  ;
  assign n40176 = n6301 & n40175 ;
  assign n40177 = ~n40174 & ~n40176 ;
  assign n40178 = \b[62]  & n6307 ;
  assign n40179 = \a[33]  & \b[61]  ;
  assign n40180 = n6298 & n40179 ;
  assign n40181 = \a[35]  & ~n40180 ;
  assign n40182 = ~n40178 & n40181 ;
  assign n40183 = n40177 & n40182 ;
  assign n40184 = n40172 & n40183 ;
  assign n40185 = ~n40178 & ~n40180 ;
  assign n40186 = n40177 & n40185 ;
  assign n40187 = n40172 & n40186 ;
  assign n40188 = ~\a[35]  & ~n40187 ;
  assign n40189 = ~n40184 & ~n40188 ;
  assign n40190 = ~n40165 & n40189 ;
  assign n40191 = ~n40161 & n40190 ;
  assign n40192 = n40165 & n40189 ;
  assign n40193 = n40161 & n40192 ;
  assign n40194 = ~n40191 & ~n40193 ;
  assign n40195 = ~n40165 & ~n40189 ;
  assign n40196 = n40161 & n40195 ;
  assign n40197 = n40165 & ~n40189 ;
  assign n40198 = ~n40161 & n40197 ;
  assign n40199 = ~n40196 & ~n40198 ;
  assign n40200 = n40194 & n40199 ;
  assign n40201 = n39849 & n40200 ;
  assign n40202 = ~n39849 & ~n40200 ;
  assign n40203 = ~n40201 & ~n40202 ;
  assign n40204 = n39825 & n40203 ;
  assign n40205 = ~n39825 & ~n40203 ;
  assign n40206 = ~n40204 & ~n40205 ;
  assign n40207 = ~n39823 & n40206 ;
  assign n40208 = ~n39815 & ~n40206 ;
  assign n40209 = ~n39819 & n40208 ;
  assign n40210 = ~n40207 & ~n40209 ;
  assign n40211 = ~n39815 & ~n40204 ;
  assign n40212 = ~n39819 & n40211 ;
  assign n40213 = n39904 & n39977 ;
  assign n40214 = ~n39982 & ~n40213 ;
  assign n40215 = ~n39947 & ~n39972 ;
  assign n40216 = ~n39945 & ~n40215 ;
  assign n40217 = ~n8599 & n18516 ;
  assign n40218 = ~n8174 & n18516 ;
  assign n40219 = ~n8595 & n40218 ;
  assign n40220 = ~n40217 & ~n40219 ;
  assign n40221 = ~n8602 & ~n40220 ;
  assign n40222 = \b[39]  & n18514 ;
  assign n40223 = \a[56]  & \b[38]  ;
  assign n40224 = n19181 & n40223 ;
  assign n40225 = ~\a[57]  & \b[38]  ;
  assign n40226 = n18508 & n40225 ;
  assign n40227 = ~n40224 & ~n40226 ;
  assign n40228 = ~n40222 & n40227 ;
  assign n40229 = \b[37]  & n19183 ;
  assign n40230 = n19180 & n40229 ;
  assign n40231 = \a[59]  & ~n40230 ;
  assign n40232 = n40228 & n40231 ;
  assign n40233 = ~n40221 & n40232 ;
  assign n40234 = n40228 & ~n40230 ;
  assign n40235 = ~\a[59]  & ~n40234 ;
  assign n40236 = ~\a[59]  & ~n8602 ;
  assign n40237 = ~n40220 & n40236 ;
  assign n40238 = ~n40235 & ~n40237 ;
  assign n40239 = ~n40233 & n40238 ;
  assign n40240 = ~n39571 & ~n39932 ;
  assign n40241 = n39928 & n40240 ;
  assign n40242 = ~n39933 & ~n40241 ;
  assign n40243 = ~\a[32]  & \b[32]  ;
  assign n40244 = n21957 & n40243 ;
  assign n40245 = ~\a[32]  & \b[33]  ;
  assign n40246 = n21958 & n40245 ;
  assign n40247 = ~n40244 & ~n40246 ;
  assign n40248 = \b[33]  & n21958 ;
  assign n40249 = \b[32]  & n21957 ;
  assign n40250 = \a[32]  & ~n40249 ;
  assign n40251 = ~n40248 & n40250 ;
  assign n40252 = n40247 & ~n40251 ;
  assign n40253 = ~n39931 & ~n40252 ;
  assign n40254 = n39931 & n40252 ;
  assign n40255 = ~n40253 & ~n40254 ;
  assign n40256 = ~n40242 & n40255 ;
  assign n40257 = n7337 & n20521 ;
  assign n40258 = ~n7334 & n40257 ;
  assign n40259 = n20521 & n37946 ;
  assign n40260 = ~n7333 & n40259 ;
  assign n40261 = \b[34]  & n21315 ;
  assign n40262 = n21312 & n40261 ;
  assign n40263 = ~\a[60]  & \b[35]  ;
  assign n40264 = n20513 & n40263 ;
  assign n40265 = ~n40262 & ~n40264 ;
  assign n40266 = \b[36]  & n20519 ;
  assign n40267 = \a[60]  & \b[35]  ;
  assign n40268 = n20510 & n40267 ;
  assign n40269 = \a[62]  & ~n40268 ;
  assign n40270 = ~n40266 & n40269 ;
  assign n40271 = n40265 & n40270 ;
  assign n40272 = ~n40260 & n40271 ;
  assign n40273 = ~n40258 & n40272 ;
  assign n40274 = ~n40266 & ~n40268 ;
  assign n40275 = n40265 & n40274 ;
  assign n40276 = ~n40260 & n40275 ;
  assign n40277 = ~n40258 & n40276 ;
  assign n40278 = ~\a[62]  & ~n40277 ;
  assign n40279 = ~n40273 & ~n40278 ;
  assign n40280 = ~n39933 & ~n40255 ;
  assign n40281 = ~n40241 & n40280 ;
  assign n40282 = n40279 & ~n40281 ;
  assign n40283 = ~n40256 & n40282 ;
  assign n40284 = ~n40255 & ~n40279 ;
  assign n40285 = n40242 & n40284 ;
  assign n40286 = n40255 & ~n40279 ;
  assign n40287 = ~n40242 & n40286 ;
  assign n40288 = ~n40285 & ~n40287 ;
  assign n40289 = ~n40283 & n40288 ;
  assign n40290 = ~n40239 & ~n40289 ;
  assign n40291 = n40239 & n40289 ;
  assign n40292 = ~n40290 & ~n40291 ;
  assign n40293 = ~n40216 & n40292 ;
  assign n40294 = n40216 & n40289 ;
  assign n40295 = n40239 & n40294 ;
  assign n40296 = n40216 & ~n40289 ;
  assign n40297 = ~n40239 & n40296 ;
  assign n40298 = ~n40295 & ~n40297 ;
  assign n40299 = ~n40293 & n40298 ;
  assign n40300 = ~n9930 & ~n16016 ;
  assign n40301 = ~n16652 & n40300 ;
  assign n40302 = n9927 & n40301 ;
  assign n40303 = n9930 & ~n16016 ;
  assign n40304 = ~n16652 & n40303 ;
  assign n40305 = ~n9927 & n40304 ;
  assign n40306 = ~n40302 & ~n40305 ;
  assign n40307 = \b[40]  & n17308 ;
  assign n40308 = n17305 & n40307 ;
  assign n40309 = ~\a[54]  & \b[41]  ;
  assign n40310 = n16647 & n40309 ;
  assign n40311 = ~n40308 & ~n40310 ;
  assign n40312 = \b[42]  & n16653 ;
  assign n40313 = \a[54]  & \b[41]  ;
  assign n40314 = n16644 & n40313 ;
  assign n40315 = \a[56]  & ~n40314 ;
  assign n40316 = ~n40312 & n40315 ;
  assign n40317 = n40311 & n40316 ;
  assign n40318 = n40306 & n40317 ;
  assign n40319 = ~n40312 & ~n40314 ;
  assign n40320 = n40311 & n40319 ;
  assign n40321 = n40306 & n40320 ;
  assign n40322 = ~\a[56]  & ~n40321 ;
  assign n40323 = ~n40318 & ~n40322 ;
  assign n40324 = n40299 & ~n40323 ;
  assign n40325 = ~n40299 & n40323 ;
  assign n40326 = ~n40324 & ~n40325 ;
  assign n40327 = ~n40214 & ~n40326 ;
  assign n40328 = n40214 & n40326 ;
  assign n40329 = ~n40327 & ~n40328 ;
  assign n40330 = ~n11397 & n14793 ;
  assign n40331 = ~n11395 & n40330 ;
  assign n40332 = \b[43]  & n15517 ;
  assign n40333 = n15514 & n40332 ;
  assign n40334 = ~\a[51]  & \b[44]  ;
  assign n40335 = n14785 & n40334 ;
  assign n40336 = ~n40333 & ~n40335 ;
  assign n40337 = \b[45]  & n14791 ;
  assign n40338 = \a[51]  & \b[44]  ;
  assign n40339 = n14782 & n40338 ;
  assign n40340 = \a[53]  & ~n40339 ;
  assign n40341 = ~n40337 & n40340 ;
  assign n40342 = n40336 & n40341 ;
  assign n40343 = ~n40331 & n40342 ;
  assign n40344 = ~n40337 & ~n40339 ;
  assign n40345 = n40336 & n40344 ;
  assign n40346 = ~n40331 & n40345 ;
  assign n40347 = ~\a[53]  & ~n40346 ;
  assign n40348 = ~n40343 & ~n40347 ;
  assign n40349 = n40329 & ~n40348 ;
  assign n40350 = ~n40329 & n40348 ;
  assign n40351 = ~n40349 & ~n40350 ;
  assign n40352 = n39877 & ~n39987 ;
  assign n40353 = ~n39987 & n39988 ;
  assign n40354 = ~n40352 & ~n40353 ;
  assign n40355 = ~n12478 & ~n12606 ;
  assign n40356 = ~n13122 & n40355 ;
  assign n40357 = n12475 & n40356 ;
  assign n40358 = n12478 & ~n12606 ;
  assign n40359 = ~n13122 & n40358 ;
  assign n40360 = ~n12475 & n40359 ;
  assign n40361 = ~n40357 & ~n40360 ;
  assign n40362 = \b[46]  & n13794 ;
  assign n40363 = n13792 & n40362 ;
  assign n40364 = ~\a[48]  & \b[47]  ;
  assign n40365 = n13117 & n40364 ;
  assign n40366 = ~n40363 & ~n40365 ;
  assign n40367 = \b[48]  & n13123 ;
  assign n40368 = \a[48]  & \b[47]  ;
  assign n40369 = n13786 & n40368 ;
  assign n40370 = \a[50]  & ~n40369 ;
  assign n40371 = ~n40367 & n40370 ;
  assign n40372 = n40366 & n40371 ;
  assign n40373 = n40361 & n40372 ;
  assign n40374 = ~n40367 & ~n40369 ;
  assign n40375 = n40366 & n40374 ;
  assign n40376 = n40361 & n40375 ;
  assign n40377 = ~\a[50]  & ~n40376 ;
  assign n40378 = ~n40373 & ~n40377 ;
  assign n40379 = n40354 & ~n40378 ;
  assign n40380 = ~n40351 & n40379 ;
  assign n40381 = ~n40354 & ~n40378 ;
  assign n40382 = n40351 & n40381 ;
  assign n40383 = ~n40380 & ~n40382 ;
  assign n40384 = ~n40354 & n40378 ;
  assign n40385 = ~n40351 & n40384 ;
  assign n40386 = n40354 & n40378 ;
  assign n40387 = n40351 & n40386 ;
  assign n40388 = ~n40385 & ~n40387 ;
  assign n40389 = n40383 & n40388 ;
  assign n40390 = ~n39992 & ~n39994 ;
  assign n40391 = n39992 & n39994 ;
  assign n40392 = n40013 & ~n40391 ;
  assign n40393 = ~n40390 & ~n40392 ;
  assign n40394 = n11572 & ~n14098 ;
  assign n40395 = ~n14096 & n40394 ;
  assign n40396 = \b[49]  & n12159 ;
  assign n40397 = n12156 & n40396 ;
  assign n40398 = ~\a[45]  & \b[50]  ;
  assign n40399 = n11564 & n40398 ;
  assign n40400 = ~n40397 & ~n40399 ;
  assign n40401 = \b[51]  & n11570 ;
  assign n40402 = \a[45]  & \b[50]  ;
  assign n40403 = n11561 & n40402 ;
  assign n40404 = \a[47]  & ~n40403 ;
  assign n40405 = ~n40401 & n40404 ;
  assign n40406 = n40400 & n40405 ;
  assign n40407 = ~n40395 & n40406 ;
  assign n40408 = ~n40401 & ~n40403 ;
  assign n40409 = n40400 & n40408 ;
  assign n40410 = ~n40395 & n40409 ;
  assign n40411 = ~\a[47]  & ~n40410 ;
  assign n40412 = ~n40407 & ~n40411 ;
  assign n40413 = ~n40393 & n40412 ;
  assign n40414 = ~n40389 & n40413 ;
  assign n40415 = n40393 & n40412 ;
  assign n40416 = n40389 & n40415 ;
  assign n40417 = ~n40414 & ~n40416 ;
  assign n40418 = ~n40393 & ~n40412 ;
  assign n40419 = n40389 & n40418 ;
  assign n40420 = n40393 & ~n40412 ;
  assign n40421 = ~n40389 & n40420 ;
  assign n40422 = ~n40419 & ~n40421 ;
  assign n40423 = n40417 & n40422 ;
  assign n40424 = n10082 & n38142 ;
  assign n40425 = ~n16404 & n40424 ;
  assign n40426 = n10082 & n16398 ;
  assign n40427 = n15241 & n40426 ;
  assign n40428 = n16400 & n40426 ;
  assign n40429 = ~n15239 & n40428 ;
  assign n40430 = ~n40427 & ~n40429 ;
  assign n40431 = ~n40425 & n40430 ;
  assign n40432 = \b[52]  & n10681 ;
  assign n40433 = n10678 & n40432 ;
  assign n40434 = \b[54]  & n10080 ;
  assign n40435 = \a[41]  & \b[53]  ;
  assign n40436 = n10679 & n40435 ;
  assign n40437 = ~\a[42]  & \b[53]  ;
  assign n40438 = n10074 & n40437 ;
  assign n40439 = ~n40436 & ~n40438 ;
  assign n40440 = ~n40434 & n40439 ;
  assign n40441 = ~n40433 & n40440 ;
  assign n40442 = n40431 & n40441 ;
  assign n40443 = ~\a[44]  & ~n40442 ;
  assign n40444 = \a[44]  & n40441 ;
  assign n40445 = n40431 & n40444 ;
  assign n40446 = ~n40443 & ~n40445 ;
  assign n40447 = n40024 & n40028 ;
  assign n40448 = n40062 & ~n40447 ;
  assign n40449 = n40446 & n40448 ;
  assign n40450 = ~n40423 & n40449 ;
  assign n40451 = n40446 & ~n40448 ;
  assign n40452 = n40423 & n40451 ;
  assign n40453 = ~n40450 & ~n40452 ;
  assign n40454 = ~n40446 & ~n40448 ;
  assign n40455 = ~n40423 & n40454 ;
  assign n40456 = ~n40446 & n40448 ;
  assign n40457 = n40423 & n40456 ;
  assign n40458 = ~n40455 & ~n40457 ;
  assign n40459 = n40453 & n40458 ;
  assign n40460 = ~n40063 & ~n40083 ;
  assign n40461 = n40063 & n40083 ;
  assign n40462 = n40081 & ~n40461 ;
  assign n40463 = ~n40460 & ~n40462 ;
  assign n40464 = n8759 & ~n17690 ;
  assign n40465 = ~n17688 & n40464 ;
  assign n40466 = \b[55]  & n9301 ;
  assign n40467 = n9298 & n40466 ;
  assign n40468 = ~\a[39]  & \b[56]  ;
  assign n40469 = n8751 & n40468 ;
  assign n40470 = ~n40467 & ~n40469 ;
  assign n40471 = \b[57]  & n8757 ;
  assign n40472 = \a[39]  & \b[56]  ;
  assign n40473 = n8748 & n40472 ;
  assign n40474 = \a[41]  & ~n40473 ;
  assign n40475 = ~n40471 & n40474 ;
  assign n40476 = n40470 & n40475 ;
  assign n40477 = ~n40465 & n40476 ;
  assign n40478 = ~n40471 & ~n40473 ;
  assign n40479 = n40470 & n40478 ;
  assign n40480 = ~n40465 & n40479 ;
  assign n40481 = ~\a[41]  & ~n40480 ;
  assign n40482 = ~n40477 & ~n40481 ;
  assign n40483 = n40463 & ~n40482 ;
  assign n40484 = ~n40459 & n40483 ;
  assign n40485 = ~n40463 & ~n40482 ;
  assign n40486 = n40459 & n40485 ;
  assign n40487 = ~n40484 & ~n40486 ;
  assign n40488 = ~n40463 & n40482 ;
  assign n40489 = ~n40459 & n40488 ;
  assign n40490 = n40463 & n40482 ;
  assign n40491 = n40459 & n40490 ;
  assign n40492 = ~n40489 & ~n40491 ;
  assign n40493 = n40487 & n40492 ;
  assign n40494 = ~n40094 & n40125 ;
  assign n40495 = n40130 & ~n40494 ;
  assign n40496 = n7534 & n20260 ;
  assign n40497 = ~n20257 & n40496 ;
  assign n40498 = ~n19545 & ~n20260 ;
  assign n40499 = n7534 & n40498 ;
  assign n40500 = ~n20256 & n40499 ;
  assign n40501 = \b[58]  & n7973 ;
  assign n40502 = n7970 & n40501 ;
  assign n40503 = ~\a[36]  & \b[59]  ;
  assign n40504 = n7526 & n40503 ;
  assign n40505 = ~n40502 & ~n40504 ;
  assign n40506 = \b[60]  & n7532 ;
  assign n40507 = \a[36]  & \b[59]  ;
  assign n40508 = n17801 & n40507 ;
  assign n40509 = \a[38]  & ~n40508 ;
  assign n40510 = ~n40506 & n40509 ;
  assign n40511 = n40505 & n40510 ;
  assign n40512 = ~n40500 & n40511 ;
  assign n40513 = ~n40497 & n40512 ;
  assign n40514 = ~n40506 & ~n40508 ;
  assign n40515 = n40505 & n40514 ;
  assign n40516 = ~n40500 & n40515 ;
  assign n40517 = ~n40497 & n40516 ;
  assign n40518 = ~\a[38]  & ~n40517 ;
  assign n40519 = ~n40513 & ~n40518 ;
  assign n40520 = ~n40495 & ~n40519 ;
  assign n40521 = ~n40493 & n40520 ;
  assign n40522 = n40495 & ~n40519 ;
  assign n40523 = n40493 & n40522 ;
  assign n40524 = ~n40521 & ~n40523 ;
  assign n40525 = n40495 & n40519 ;
  assign n40526 = ~n40493 & n40525 ;
  assign n40527 = ~n40495 & n40519 ;
  assign n40528 = n40493 & n40527 ;
  assign n40529 = ~n40526 & ~n40528 ;
  assign n40530 = n40524 & n40529 ;
  assign n40531 = ~n40137 & n40158 ;
  assign n40532 = ~n40138 & ~n40531 ;
  assign n40533 = ~n40530 & ~n40532 ;
  assign n40534 = n40530 & n40532 ;
  assign n40535 = ~n40533 & ~n40534 ;
  assign n40536 = n40161 & n40165 ;
  assign n40537 = n40189 & ~n40536 ;
  assign n40538 = ~n40161 & ~n40165 ;
  assign n40539 = n6309 & ~n22461 ;
  assign n40540 = ~n22459 & n40539 ;
  assign n40541 = \b[63]  & n6307 ;
  assign n40542 = \a[33]  & \b[62]  ;
  assign n40543 = n6298 & n40542 ;
  assign n40544 = ~n40541 & ~n40543 ;
  assign n40545 = \b[61]  & n6778 ;
  assign n40546 = n6775 & n40545 ;
  assign n40547 = ~\a[33]  & \b[62]  ;
  assign n40548 = n6301 & n40547 ;
  assign n40549 = ~n40546 & ~n40548 ;
  assign n40550 = n40544 & n40549 ;
  assign n40551 = ~n40540 & n40550 ;
  assign n40552 = ~\a[35]  & ~n40551 ;
  assign n40553 = \a[35]  & n40550 ;
  assign n40554 = ~n40540 & n40553 ;
  assign n40555 = ~n40552 & ~n40554 ;
  assign n40556 = ~n40538 & ~n40555 ;
  assign n40557 = ~n40537 & n40556 ;
  assign n40558 = n40538 & n40555 ;
  assign n40559 = n40189 & n40555 ;
  assign n40560 = ~n40536 & n40559 ;
  assign n40561 = ~n40558 & ~n40560 ;
  assign n40562 = ~n40557 & n40561 ;
  assign n40563 = ~n40535 & ~n40562 ;
  assign n40564 = n40535 & n40562 ;
  assign n40565 = ~n40563 & ~n40564 ;
  assign n40566 = ~n39846 & ~n40200 ;
  assign n40567 = ~n39848 & ~n40566 ;
  assign n40568 = n40565 & n40567 ;
  assign n40569 = ~n40565 & ~n40567 ;
  assign n40570 = ~n40568 & ~n40569 ;
  assign n40571 = ~n40205 & n40570 ;
  assign n40572 = ~n40212 & n40571 ;
  assign n40573 = ~n40205 & ~n40212 ;
  assign n40574 = ~n40570 & ~n40573 ;
  assign n40575 = ~n40572 & ~n40574 ;
  assign n40576 = ~n40568 & ~n40572 ;
  assign n40577 = ~n40535 & ~n40557 ;
  assign n40578 = n40561 & ~n40577 ;
  assign n40579 = n40524 & ~n40532 ;
  assign n40580 = ~n5952 & ~n22458 ;
  assign n40581 = ~n6306 & n40580 ;
  assign n40582 = ~n23173 & n40581 ;
  assign n40583 = \b[62]  & n6778 ;
  assign n40584 = n6775 & n40583 ;
  assign n40585 = \a[33]  & \b[63]  ;
  assign n40586 = n6298 & n40585 ;
  assign n40587 = ~\a[33]  & \b[63]  ;
  assign n40588 = n6301 & n40587 ;
  assign n40589 = \a[35]  & ~n40588 ;
  assign n40590 = ~n40586 & n40589 ;
  assign n40591 = ~n40584 & n40590 ;
  assign n40592 = ~n40582 & n40591 ;
  assign n40593 = ~n40586 & ~n40588 ;
  assign n40594 = ~n40584 & n40593 ;
  assign n40595 = ~n40582 & n40594 ;
  assign n40596 = ~\a[35]  & ~n40595 ;
  assign n40597 = ~n40592 & ~n40596 ;
  assign n40598 = n40529 & ~n40597 ;
  assign n40599 = ~n40579 & n40598 ;
  assign n40600 = n40529 & ~n40579 ;
  assign n40601 = n40597 & ~n40600 ;
  assign n40602 = ~n40599 & ~n40601 ;
  assign n40603 = ~n40349 & ~n40354 ;
  assign n40604 = ~n40350 & ~n40603 ;
  assign n40605 = ~n40214 & ~n40324 ;
  assign n40606 = ~n40325 & ~n40605 ;
  assign n40607 = n40216 & n40239 ;
  assign n40608 = ~n40294 & ~n40607 ;
  assign n40609 = ~n40291 & n40608 ;
  assign n40610 = ~n9044 & ~n17912 ;
  assign n40611 = ~n18513 & n40610 ;
  assign n40612 = n9041 & n40611 ;
  assign n40613 = n9044 & ~n17912 ;
  assign n40614 = ~n18513 & n40613 ;
  assign n40615 = ~n9041 & n40614 ;
  assign n40616 = ~n40612 & ~n40615 ;
  assign n40617 = \b[40]  & n18514 ;
  assign n40618 = \a[56]  & \b[39]  ;
  assign n40619 = n19181 & n40618 ;
  assign n40620 = ~\a[57]  & \b[39]  ;
  assign n40621 = n18508 & n40620 ;
  assign n40622 = ~n40619 & ~n40621 ;
  assign n40623 = ~n40617 & n40622 ;
  assign n40624 = \b[38]  & n19183 ;
  assign n40625 = n19180 & n40624 ;
  assign n40626 = \a[59]  & ~n40625 ;
  assign n40627 = n40623 & n40626 ;
  assign n40628 = n40616 & n40627 ;
  assign n40629 = n40623 & ~n40625 ;
  assign n40630 = n40616 & n40629 ;
  assign n40631 = ~\a[59]  & ~n40630 ;
  assign n40632 = ~n40628 & ~n40631 ;
  assign n40633 = ~n40256 & ~n40282 ;
  assign n40634 = \b[37]  & n20519 ;
  assign n40635 = \a[60]  & \b[36]  ;
  assign n40636 = n20510 & n40635 ;
  assign n40637 = ~n40634 & ~n40636 ;
  assign n40638 = \b[35]  & n21315 ;
  assign n40639 = n21312 & n40638 ;
  assign n40640 = ~\a[60]  & \b[36]  ;
  assign n40641 = n20513 & n40640 ;
  assign n40642 = ~n40639 & ~n40641 ;
  assign n40643 = n40637 & n40642 ;
  assign n40644 = ~\a[62]  & ~n40643 ;
  assign n40645 = ~n7758 & n20521 ;
  assign n40646 = ~n7336 & n20521 ;
  assign n40647 = ~n7754 & n40646 ;
  assign n40648 = ~n40645 & ~n40647 ;
  assign n40649 = ~\a[62]  & ~n7761 ;
  assign n40650 = ~n40648 & n40649 ;
  assign n40651 = ~n40644 & ~n40650 ;
  assign n40652 = ~n39931 & ~n40251 ;
  assign n40653 = \b[34]  & n21958 ;
  assign n40654 = \b[33]  & n21957 ;
  assign n40655 = ~n40653 & ~n40654 ;
  assign n40656 = n40247 & ~n40655 ;
  assign n40657 = ~n40652 & n40656 ;
  assign n40658 = n40247 & ~n40652 ;
  assign n40659 = n40655 & ~n40658 ;
  assign n40660 = ~n40657 & ~n40659 ;
  assign n40661 = \a[62]  & ~n40636 ;
  assign n40662 = ~n40634 & n40661 ;
  assign n40663 = n40642 & n40662 ;
  assign n40664 = ~n40660 & ~n40663 ;
  assign n40665 = ~n7761 & ~n40660 ;
  assign n40666 = ~n40648 & n40665 ;
  assign n40667 = ~n40664 & ~n40666 ;
  assign n40668 = n40651 & ~n40667 ;
  assign n40669 = ~n7761 & ~n40648 ;
  assign n40670 = \a[62]  & n40643 ;
  assign n40671 = ~n40669 & n40670 ;
  assign n40672 = n40651 & ~n40671 ;
  assign n40673 = n40660 & ~n40672 ;
  assign n40674 = ~n40668 & ~n40673 ;
  assign n40675 = n40633 & n40674 ;
  assign n40676 = ~n40633 & ~n40674 ;
  assign n40677 = ~n40675 & ~n40676 ;
  assign n40678 = n40632 & n40677 ;
  assign n40679 = ~n40632 & ~n40677 ;
  assign n40680 = ~n40678 & ~n40679 ;
  assign n40681 = n40609 & ~n40680 ;
  assign n40682 = ~n40609 & n40680 ;
  assign n40683 = ~n40681 & ~n40682 ;
  assign n40684 = ~n10406 & n37945 ;
  assign n40685 = ~n9929 & n37945 ;
  assign n40686 = ~n10402 & n40685 ;
  assign n40687 = ~n40684 & ~n40686 ;
  assign n40688 = ~n10409 & ~n40687 ;
  assign n40689 = \b[41]  & n17308 ;
  assign n40690 = n17305 & n40689 ;
  assign n40691 = ~\a[54]  & \b[42]  ;
  assign n40692 = n16647 & n40691 ;
  assign n40693 = ~n40690 & ~n40692 ;
  assign n40694 = \b[43]  & n16653 ;
  assign n40695 = \a[54]  & \b[42]  ;
  assign n40696 = n16644 & n40695 ;
  assign n40697 = \a[56]  & ~n40696 ;
  assign n40698 = ~n40694 & n40697 ;
  assign n40699 = n40693 & n40698 ;
  assign n40700 = ~n40688 & n40699 ;
  assign n40701 = ~n40694 & ~n40696 ;
  assign n40702 = n40693 & n40701 ;
  assign n40703 = ~\a[56]  & ~n40702 ;
  assign n40704 = ~\a[56]  & ~n10409 ;
  assign n40705 = ~n40687 & n40704 ;
  assign n40706 = ~n40703 & ~n40705 ;
  assign n40707 = ~n40700 & n40706 ;
  assign n40708 = n40683 & ~n40707 ;
  assign n40709 = ~n40683 & n40707 ;
  assign n40710 = ~n40708 & ~n40709 ;
  assign n40711 = ~n40606 & ~n40710 ;
  assign n40712 = n40606 & n40710 ;
  assign n40713 = ~n40711 & ~n40712 ;
  assign n40714 = n11906 & n14793 ;
  assign n40715 = ~n11903 & n40714 ;
  assign n40716 = n13483 & n14793 ;
  assign n40717 = ~n11902 & n40716 ;
  assign n40718 = \b[44]  & n15517 ;
  assign n40719 = n15514 & n40718 ;
  assign n40720 = ~\a[51]  & \b[45]  ;
  assign n40721 = n14785 & n40720 ;
  assign n40722 = ~n40719 & ~n40721 ;
  assign n40723 = \b[46]  & n14791 ;
  assign n40724 = \a[51]  & \b[45]  ;
  assign n40725 = n14782 & n40724 ;
  assign n40726 = \a[53]  & ~n40725 ;
  assign n40727 = ~n40723 & n40726 ;
  assign n40728 = n40722 & n40727 ;
  assign n40729 = ~n40717 & n40728 ;
  assign n40730 = ~n40715 & n40729 ;
  assign n40731 = ~n40723 & ~n40725 ;
  assign n40732 = n40722 & n40731 ;
  assign n40733 = ~n40717 & n40732 ;
  assign n40734 = ~n40715 & n40733 ;
  assign n40735 = ~\a[53]  & ~n40734 ;
  assign n40736 = ~n40730 & ~n40735 ;
  assign n40737 = ~n40713 & n40736 ;
  assign n40738 = n40713 & ~n40736 ;
  assign n40739 = ~n40737 & ~n40738 ;
  assign n40740 = ~n40604 & ~n40739 ;
  assign n40741 = n40604 & n40739 ;
  assign n40742 = ~n40740 & ~n40741 ;
  assign n40743 = n13125 & ~n13524 ;
  assign n40744 = ~n13522 & n40743 ;
  assign n40745 = \b[47]  & n13794 ;
  assign n40746 = n13792 & n40745 ;
  assign n40747 = ~\a[48]  & \b[48]  ;
  assign n40748 = n13117 & n40747 ;
  assign n40749 = ~n40746 & ~n40748 ;
  assign n40750 = \b[49]  & n13123 ;
  assign n40751 = \a[48]  & \b[48]  ;
  assign n40752 = n13786 & n40751 ;
  assign n40753 = \a[50]  & ~n40752 ;
  assign n40754 = ~n40750 & n40753 ;
  assign n40755 = n40749 & n40754 ;
  assign n40756 = ~n40744 & n40755 ;
  assign n40757 = ~n40750 & ~n40752 ;
  assign n40758 = n40749 & n40757 ;
  assign n40759 = ~n40744 & n40758 ;
  assign n40760 = ~\a[50]  & ~n40759 ;
  assign n40761 = ~n40756 & ~n40760 ;
  assign n40762 = n40742 & ~n40761 ;
  assign n40763 = ~n40742 & n40761 ;
  assign n40764 = ~n40762 & ~n40763 ;
  assign n40765 = n40383 & ~n40393 ;
  assign n40766 = n40388 & ~n40765 ;
  assign n40767 = ~n10988 & ~n14093 ;
  assign n40768 = ~n15201 & n40767 ;
  assign n40769 = ~n15197 & n40768 ;
  assign n40770 = ~n11569 & n40769 ;
  assign n40771 = n11572 & n15201 ;
  assign n40772 = ~n15198 & n40771 ;
  assign n40773 = ~n40770 & ~n40772 ;
  assign n40774 = \b[50]  & n12159 ;
  assign n40775 = n12156 & n40774 ;
  assign n40776 = ~\a[45]  & \b[51]  ;
  assign n40777 = n11564 & n40776 ;
  assign n40778 = ~n40775 & ~n40777 ;
  assign n40779 = \b[52]  & n11570 ;
  assign n40780 = \a[45]  & \b[51]  ;
  assign n40781 = n11561 & n40780 ;
  assign n40782 = \a[47]  & ~n40781 ;
  assign n40783 = ~n40779 & n40782 ;
  assign n40784 = n40778 & n40783 ;
  assign n40785 = n40773 & n40784 ;
  assign n40786 = ~n40779 & ~n40781 ;
  assign n40787 = n40778 & n40786 ;
  assign n40788 = n40773 & n40787 ;
  assign n40789 = ~\a[47]  & ~n40788 ;
  assign n40790 = ~n40785 & ~n40789 ;
  assign n40791 = ~n40766 & n40790 ;
  assign n40792 = ~n40764 & n40791 ;
  assign n40793 = n40766 & n40790 ;
  assign n40794 = n40764 & n40793 ;
  assign n40795 = ~n40792 & ~n40794 ;
  assign n40796 = n40766 & ~n40790 ;
  assign n40797 = ~n40764 & n40796 ;
  assign n40798 = ~n40766 & ~n40790 ;
  assign n40799 = n40764 & n40798 ;
  assign n40800 = ~n40797 & ~n40799 ;
  assign n40801 = n40795 & n40800 ;
  assign n40802 = n10082 & ~n16446 ;
  assign n40803 = ~n16444 & n40802 ;
  assign n40804 = \b[55]  & n10080 ;
  assign n40805 = \a[41]  & \b[54]  ;
  assign n40806 = n10679 & n40805 ;
  assign n40807 = ~\a[42]  & \b[54]  ;
  assign n40808 = n10074 & n40807 ;
  assign n40809 = ~n40806 & ~n40808 ;
  assign n40810 = ~n40804 & n40809 ;
  assign n40811 = \b[53]  & n10681 ;
  assign n40812 = n10678 & n40811 ;
  assign n40813 = \a[44]  & ~n40812 ;
  assign n40814 = n40810 & n40813 ;
  assign n40815 = ~n40803 & n40814 ;
  assign n40816 = n40810 & ~n40812 ;
  assign n40817 = ~n40803 & n40816 ;
  assign n40818 = ~\a[44]  & ~n40817 ;
  assign n40819 = ~n40815 & ~n40818 ;
  assign n40820 = n40422 & n40448 ;
  assign n40821 = n40417 & ~n40820 ;
  assign n40822 = n40819 & ~n40821 ;
  assign n40823 = n40801 & n40822 ;
  assign n40824 = n40819 & n40821 ;
  assign n40825 = ~n40801 & n40824 ;
  assign n40826 = ~n40823 & ~n40825 ;
  assign n40827 = ~n40819 & ~n40821 ;
  assign n40828 = ~n40801 & n40827 ;
  assign n40829 = ~n40819 & n40821 ;
  assign n40830 = n40801 & n40829 ;
  assign n40831 = ~n40828 & ~n40830 ;
  assign n40832 = n40826 & n40831 ;
  assign n40833 = n40458 & ~n40463 ;
  assign n40834 = n40453 & ~n40833 ;
  assign n40835 = n8759 & ~n19543 ;
  assign n40836 = ~n38598 & n40835 ;
  assign n40837 = \b[56]  & n9301 ;
  assign n40838 = n9298 & n40837 ;
  assign n40839 = ~\a[39]  & \b[57]  ;
  assign n40840 = n8751 & n40839 ;
  assign n40841 = ~n40838 & ~n40840 ;
  assign n40842 = \b[58]  & n8757 ;
  assign n40843 = \a[39]  & \b[57]  ;
  assign n40844 = n8748 & n40843 ;
  assign n40845 = \a[41]  & ~n40844 ;
  assign n40846 = ~n40842 & n40845 ;
  assign n40847 = n40841 & n40846 ;
  assign n40848 = ~n40836 & n40847 ;
  assign n40849 = ~n40842 & ~n40844 ;
  assign n40850 = n40841 & n40849 ;
  assign n40851 = ~n40836 & n40850 ;
  assign n40852 = ~\a[41]  & ~n40851 ;
  assign n40853 = ~n40848 & ~n40852 ;
  assign n40854 = ~n40834 & ~n40853 ;
  assign n40855 = ~n40832 & n40854 ;
  assign n40856 = n40834 & ~n40853 ;
  assign n40857 = n40832 & n40856 ;
  assign n40858 = ~n40855 & ~n40857 ;
  assign n40859 = n40834 & n40853 ;
  assign n40860 = ~n40832 & n40859 ;
  assign n40861 = ~n40834 & n40853 ;
  assign n40862 = n40832 & n40861 ;
  assign n40863 = ~n40860 & ~n40862 ;
  assign n40864 = n40858 & n40863 ;
  assign n40865 = n40487 & n40495 ;
  assign n40866 = n40492 & ~n40865 ;
  assign n40867 = n7534 & ~n20971 ;
  assign n40868 = ~n20969 & n40867 ;
  assign n40869 = \b[59]  & n7973 ;
  assign n40870 = n7970 & n40869 ;
  assign n40871 = ~\a[36]  & \b[60]  ;
  assign n40872 = n7526 & n40871 ;
  assign n40873 = ~n40870 & ~n40872 ;
  assign n40874 = \b[61]  & n7532 ;
  assign n40875 = \a[36]  & \b[60]  ;
  assign n40876 = n17801 & n40875 ;
  assign n40877 = \a[38]  & ~n40876 ;
  assign n40878 = ~n40874 & n40877 ;
  assign n40879 = n40873 & n40878 ;
  assign n40880 = ~n40868 & n40879 ;
  assign n40881 = ~n40874 & ~n40876 ;
  assign n40882 = n40873 & n40881 ;
  assign n40883 = ~n40868 & n40882 ;
  assign n40884 = ~\a[38]  & ~n40883 ;
  assign n40885 = ~n40880 & ~n40884 ;
  assign n40886 = n40866 & ~n40885 ;
  assign n40887 = ~n40864 & n40886 ;
  assign n40888 = ~n40866 & ~n40885 ;
  assign n40889 = n40864 & n40888 ;
  assign n40890 = ~n40887 & ~n40889 ;
  assign n40891 = ~n40866 & n40885 ;
  assign n40892 = ~n40864 & n40891 ;
  assign n40893 = n40866 & n40885 ;
  assign n40894 = n40864 & n40893 ;
  assign n40895 = ~n40892 & ~n40894 ;
  assign n40896 = n40890 & n40895 ;
  assign n40897 = n40602 & n40896 ;
  assign n40898 = ~n40602 & ~n40896 ;
  assign n40899 = ~n40897 & ~n40898 ;
  assign n40900 = n40578 & n40899 ;
  assign n40901 = ~n40578 & ~n40899 ;
  assign n40902 = ~n40900 & ~n40901 ;
  assign n40903 = ~n40576 & n40902 ;
  assign n40904 = ~n40568 & ~n40902 ;
  assign n40905 = ~n40572 & n40904 ;
  assign n40906 = ~n40903 & ~n40905 ;
  assign n40907 = ~n40568 & ~n40900 ;
  assign n40908 = ~n40572 & n40907 ;
  assign n40909 = ~n40599 & ~n40896 ;
  assign n40910 = ~n40601 & ~n40909 ;
  assign n40911 = n40864 & n40866 ;
  assign n40912 = n40885 & ~n40911 ;
  assign n40913 = ~n40864 & ~n40866 ;
  assign n40914 = ~n6306 & n39033 ;
  assign n40915 = ~n23171 & n40914 ;
  assign n40916 = ~n5952 & n40915 ;
  assign n40917 = \a[32]  & \a[34]  ;
  assign n40918 = \a[33]  & ~\a[35]  ;
  assign n40919 = n40917 & n40918 ;
  assign n40920 = ~\a[32]  & ~\a[34]  ;
  assign n40921 = ~\a[33]  & \a[35]  ;
  assign n40922 = n40920 & n40921 ;
  assign n40923 = ~n40919 & ~n40922 ;
  assign n40924 = \b[63]  & ~n40923 ;
  assign n40925 = \a[35]  & ~n40924 ;
  assign n40926 = ~n40916 & n40925 ;
  assign n40927 = ~\a[35]  & n40924 ;
  assign n40928 = ~\a[35]  & ~n5952 ;
  assign n40929 = n40915 & n40928 ;
  assign n40930 = ~n40927 & ~n40929 ;
  assign n40931 = ~n40926 & n40930 ;
  assign n40932 = ~n40913 & ~n40931 ;
  assign n40933 = ~n40912 & n40932 ;
  assign n40934 = ~n40912 & ~n40913 ;
  assign n40935 = n40931 & ~n40934 ;
  assign n40936 = ~n40933 & ~n40935 ;
  assign n40937 = n10082 & n17647 ;
  assign n40938 = ~n17644 & n40937 ;
  assign n40939 = n10082 & n19567 ;
  assign n40940 = ~n17643 & n40939 ;
  assign n40941 = \b[54]  & n10681 ;
  assign n40942 = n10678 & n40941 ;
  assign n40943 = \b[56]  & n10080 ;
  assign n40944 = \a[41]  & \b[55]  ;
  assign n40945 = n10679 & n40944 ;
  assign n40946 = ~\a[42]  & \b[55]  ;
  assign n40947 = n10074 & n40946 ;
  assign n40948 = ~n40945 & ~n40947 ;
  assign n40949 = ~n40943 & n40948 ;
  assign n40950 = ~n40942 & n40949 ;
  assign n40951 = ~n40940 & n40950 ;
  assign n40952 = ~n40938 & n40951 ;
  assign n40953 = ~\a[44]  & ~n40952 ;
  assign n40954 = \a[44]  & n40950 ;
  assign n40955 = ~n40940 & n40954 ;
  assign n40956 = ~n40938 & n40955 ;
  assign n40957 = ~n40953 & ~n40956 ;
  assign n40958 = ~n10889 & ~n16016 ;
  assign n40959 = ~n16652 & n40958 ;
  assign n40960 = n10886 & n40959 ;
  assign n40961 = n10889 & ~n16016 ;
  assign n40962 = ~n16652 & n40961 ;
  assign n40963 = ~n10886 & n40962 ;
  assign n40964 = ~n40960 & ~n40963 ;
  assign n40965 = \b[42]  & n17308 ;
  assign n40966 = n17305 & n40965 ;
  assign n40967 = ~\a[54]  & \b[43]  ;
  assign n40968 = n16647 & n40967 ;
  assign n40969 = ~n40966 & ~n40968 ;
  assign n40970 = \b[44]  & n16653 ;
  assign n40971 = \a[54]  & \b[43]  ;
  assign n40972 = n16644 & n40971 ;
  assign n40973 = \a[56]  & ~n40972 ;
  assign n40974 = ~n40970 & n40973 ;
  assign n40975 = n40969 & n40974 ;
  assign n40976 = n40964 & n40975 ;
  assign n40977 = ~n40970 & ~n40972 ;
  assign n40978 = n40969 & n40977 ;
  assign n40979 = n40964 & n40978 ;
  assign n40980 = ~\a[56]  & ~n40979 ;
  assign n40981 = ~n40976 & ~n40980 ;
  assign n40982 = n40632 & ~n40675 ;
  assign n40983 = ~n40676 & ~n40982 ;
  assign n40984 = ~n40659 & ~n40673 ;
  assign n40985 = \b[35]  & n21958 ;
  assign n40986 = \b[34]  & n21957 ;
  assign n40987 = ~n40985 & ~n40986 ;
  assign n40988 = ~n40655 & n40987 ;
  assign n40989 = n40655 & ~n40987 ;
  assign n40990 = ~n40988 & ~n40989 ;
  assign n40991 = ~n40984 & n40990 ;
  assign n40992 = n8175 & n20521 ;
  assign n40993 = ~n8172 & n40992 ;
  assign n40994 = n20521 & n25622 ;
  assign n40995 = ~n8171 & n40994 ;
  assign n40996 = \b[36]  & n21315 ;
  assign n40997 = n21312 & n40996 ;
  assign n40998 = ~\a[60]  & \b[37]  ;
  assign n40999 = n20513 & n40998 ;
  assign n41000 = ~n40997 & ~n40999 ;
  assign n41001 = \b[38]  & n20519 ;
  assign n41002 = \a[60]  & \b[37]  ;
  assign n41003 = n20510 & n41002 ;
  assign n41004 = \a[62]  & ~n41003 ;
  assign n41005 = ~n41001 & n41004 ;
  assign n41006 = n41000 & n41005 ;
  assign n41007 = ~n40995 & n41006 ;
  assign n41008 = ~n40993 & n41007 ;
  assign n41009 = ~n41001 & ~n41003 ;
  assign n41010 = n41000 & n41009 ;
  assign n41011 = ~n40995 & n41010 ;
  assign n41012 = ~n40993 & n41011 ;
  assign n41013 = ~\a[62]  & ~n41012 ;
  assign n41014 = ~n41008 & ~n41013 ;
  assign n41015 = ~n40657 & ~n40672 ;
  assign n41016 = ~n40659 & ~n40990 ;
  assign n41017 = ~n41015 & n41016 ;
  assign n41018 = ~n41014 & ~n41017 ;
  assign n41019 = ~n40991 & n41018 ;
  assign n41020 = n41014 & n41017 ;
  assign n41021 = n40990 & n41014 ;
  assign n41022 = ~n40984 & n41021 ;
  assign n41023 = ~n41020 & ~n41022 ;
  assign n41024 = ~n41019 & n41023 ;
  assign n41025 = ~n9479 & n18516 ;
  assign n41026 = ~n9043 & n18516 ;
  assign n41027 = ~n9475 & n41026 ;
  assign n41028 = ~n41025 & ~n41027 ;
  assign n41029 = ~n9482 & ~n41028 ;
  assign n41030 = \b[41]  & n18514 ;
  assign n41031 = \a[56]  & \b[40]  ;
  assign n41032 = n19181 & n41031 ;
  assign n41033 = ~\a[57]  & \b[40]  ;
  assign n41034 = n18508 & n41033 ;
  assign n41035 = ~n41032 & ~n41034 ;
  assign n41036 = ~n41030 & n41035 ;
  assign n41037 = \b[39]  & n19183 ;
  assign n41038 = n19180 & n41037 ;
  assign n41039 = \a[59]  & ~n41038 ;
  assign n41040 = n41036 & n41039 ;
  assign n41041 = ~n41029 & n41040 ;
  assign n41042 = n41036 & ~n41038 ;
  assign n41043 = ~\a[59]  & ~n41042 ;
  assign n41044 = ~\a[59]  & ~n9482 ;
  assign n41045 = ~n41028 & n41044 ;
  assign n41046 = ~n41043 & ~n41045 ;
  assign n41047 = ~n41041 & n41046 ;
  assign n41048 = ~n41024 & n41047 ;
  assign n41049 = ~n40983 & n41048 ;
  assign n41050 = ~n41024 & ~n41047 ;
  assign n41051 = n40983 & n41050 ;
  assign n41052 = ~n41049 & ~n41051 ;
  assign n41053 = ~n40983 & n41047 ;
  assign n41054 = ~n40676 & ~n41047 ;
  assign n41055 = ~n40982 & n41054 ;
  assign n41056 = n41024 & ~n41055 ;
  assign n41057 = ~n41053 & n41056 ;
  assign n41058 = n41052 & ~n41057 ;
  assign n41059 = n40981 & n41058 ;
  assign n41060 = ~n40981 & ~n41058 ;
  assign n41061 = ~n41059 & ~n41060 ;
  assign n41062 = ~n40681 & n40707 ;
  assign n41063 = ~n40682 & ~n41062 ;
  assign n41064 = ~n12435 & n14793 ;
  assign n41065 = ~n11905 & n14793 ;
  assign n41066 = ~n12431 & n41065 ;
  assign n41067 = ~n41064 & ~n41066 ;
  assign n41068 = ~n12438 & ~n41067 ;
  assign n41069 = \b[45]  & n15517 ;
  assign n41070 = n15514 & n41069 ;
  assign n41071 = ~\a[51]  & \b[46]  ;
  assign n41072 = n14785 & n41071 ;
  assign n41073 = ~n41070 & ~n41072 ;
  assign n41074 = \b[47]  & n14791 ;
  assign n41075 = \a[51]  & \b[46]  ;
  assign n41076 = n14782 & n41075 ;
  assign n41077 = \a[53]  & ~n41076 ;
  assign n41078 = ~n41074 & n41077 ;
  assign n41079 = n41073 & n41078 ;
  assign n41080 = ~n41068 & n41079 ;
  assign n41081 = ~n41074 & ~n41076 ;
  assign n41082 = n41073 & n41081 ;
  assign n41083 = ~\a[53]  & ~n41082 ;
  assign n41084 = ~\a[53]  & ~n12438 ;
  assign n41085 = ~n41067 & n41084 ;
  assign n41086 = ~n41083 & ~n41085 ;
  assign n41087 = ~n41080 & n41086 ;
  assign n41088 = ~n41063 & ~n41087 ;
  assign n41089 = ~n41061 & n41088 ;
  assign n41090 = n41063 & ~n41087 ;
  assign n41091 = n41061 & n41090 ;
  assign n41092 = ~n41089 & ~n41091 ;
  assign n41093 = ~n41063 & n41087 ;
  assign n41094 = n41061 & n41093 ;
  assign n41095 = n41063 & n41087 ;
  assign n41096 = ~n41061 & n41095 ;
  assign n41097 = ~n41094 & ~n41096 ;
  assign n41098 = n41092 & n41097 ;
  assign n41099 = ~n40712 & n40736 ;
  assign n41100 = ~n40711 & ~n41099 ;
  assign n41101 = ~n41098 & ~n41100 ;
  assign n41102 = n41098 & n41100 ;
  assign n41103 = ~n41101 & ~n41102 ;
  assign n41104 = ~n12606 & ~n13519 ;
  assign n41105 = ~n14052 & n41104 ;
  assign n41106 = ~n14048 & n41105 ;
  assign n41107 = ~n13122 & n41106 ;
  assign n41108 = n13125 & n14052 ;
  assign n41109 = ~n14049 & n41108 ;
  assign n41110 = ~n41107 & ~n41109 ;
  assign n41111 = \b[48]  & n13794 ;
  assign n41112 = n13792 & n41111 ;
  assign n41113 = ~\a[48]  & \b[49]  ;
  assign n41114 = n13117 & n41113 ;
  assign n41115 = ~n41112 & ~n41114 ;
  assign n41116 = \b[50]  & n13123 ;
  assign n41117 = \a[48]  & \b[49]  ;
  assign n41118 = n13786 & n41117 ;
  assign n41119 = \a[50]  & ~n41118 ;
  assign n41120 = ~n41116 & n41119 ;
  assign n41121 = n41115 & n41120 ;
  assign n41122 = n41110 & n41121 ;
  assign n41123 = ~n41116 & ~n41118 ;
  assign n41124 = n41115 & n41123 ;
  assign n41125 = n41110 & n41124 ;
  assign n41126 = ~\a[50]  & ~n41125 ;
  assign n41127 = ~n41122 & ~n41126 ;
  assign n41128 = ~n41103 & n41127 ;
  assign n41129 = n41103 & ~n41127 ;
  assign n41130 = ~n41128 & ~n41129 ;
  assign n41131 = n11572 & ~n15246 ;
  assign n41132 = ~n15244 & n41131 ;
  assign n41133 = \b[51]  & n12159 ;
  assign n41134 = n12156 & n41133 ;
  assign n41135 = ~\a[45]  & \b[52]  ;
  assign n41136 = n11564 & n41135 ;
  assign n41137 = ~n41134 & ~n41136 ;
  assign n41138 = \b[53]  & n11570 ;
  assign n41139 = \a[45]  & \b[52]  ;
  assign n41140 = n11561 & n41139 ;
  assign n41141 = \a[47]  & ~n41140 ;
  assign n41142 = ~n41138 & n41141 ;
  assign n41143 = n41137 & n41142 ;
  assign n41144 = ~n41132 & n41143 ;
  assign n41145 = ~n41138 & ~n41140 ;
  assign n41146 = n41137 & n41145 ;
  assign n41147 = ~n41132 & n41146 ;
  assign n41148 = ~\a[47]  & ~n41147 ;
  assign n41149 = ~n41144 & ~n41148 ;
  assign n41150 = ~n40741 & n40761 ;
  assign n41151 = ~n40740 & ~n41150 ;
  assign n41152 = n41149 & ~n41151 ;
  assign n41153 = n41130 & n41152 ;
  assign n41154 = n41149 & n41151 ;
  assign n41155 = ~n41130 & n41154 ;
  assign n41156 = ~n41153 & ~n41155 ;
  assign n41157 = ~n41149 & ~n41151 ;
  assign n41158 = ~n41130 & n41157 ;
  assign n41159 = ~n41149 & n41151 ;
  assign n41160 = n41130 & n41159 ;
  assign n41161 = ~n41158 & ~n41160 ;
  assign n41162 = n41156 & n41161 ;
  assign n41163 = ~n40764 & ~n40766 ;
  assign n41164 = n40764 & n40766 ;
  assign n41165 = n40790 & ~n41164 ;
  assign n41166 = ~n41163 & ~n41165 ;
  assign n41167 = ~n41162 & n41166 ;
  assign n41168 = n41162 & ~n41166 ;
  assign n41169 = ~n41167 & ~n41168 ;
  assign n41170 = ~n40957 & n41169 ;
  assign n41171 = n40957 & ~n41169 ;
  assign n41172 = ~n41170 & ~n41171 ;
  assign n41173 = ~n40801 & ~n40821 ;
  assign n41174 = n40801 & n40821 ;
  assign n41175 = n40819 & ~n41174 ;
  assign n41176 = ~n41173 & ~n41175 ;
  assign n41177 = n8759 & ~n19550 ;
  assign n41178 = ~n19548 & n41177 ;
  assign n41179 = \b[57]  & n9301 ;
  assign n41180 = n9298 & n41179 ;
  assign n41181 = ~\a[39]  & \b[58]  ;
  assign n41182 = n8751 & n41181 ;
  assign n41183 = ~n41180 & ~n41182 ;
  assign n41184 = \b[59]  & n8757 ;
  assign n41185 = \a[39]  & \b[58]  ;
  assign n41186 = n8748 & n41185 ;
  assign n41187 = \a[41]  & ~n41186 ;
  assign n41188 = ~n41184 & n41187 ;
  assign n41189 = n41183 & n41188 ;
  assign n41190 = ~n41178 & n41189 ;
  assign n41191 = ~n41184 & ~n41186 ;
  assign n41192 = n41183 & n41191 ;
  assign n41193 = ~n41178 & n41192 ;
  assign n41194 = ~\a[41]  & ~n41193 ;
  assign n41195 = ~n41190 & ~n41194 ;
  assign n41196 = n41176 & ~n41195 ;
  assign n41197 = ~n41172 & n41196 ;
  assign n41198 = ~n41176 & ~n41195 ;
  assign n41199 = n41172 & n41198 ;
  assign n41200 = ~n41197 & ~n41199 ;
  assign n41201 = ~n41176 & n41195 ;
  assign n41202 = ~n41172 & n41201 ;
  assign n41203 = n41176 & n41195 ;
  assign n41204 = n41172 & n41203 ;
  assign n41205 = ~n41202 & ~n41204 ;
  assign n41206 = n41200 & n41205 ;
  assign n41207 = n40832 & ~n40834 ;
  assign n41208 = ~n40832 & n40834 ;
  assign n41209 = n40853 & ~n41208 ;
  assign n41210 = ~n41207 & ~n41209 ;
  assign n41211 = n7534 & n21696 ;
  assign n41212 = ~n21693 & n41211 ;
  assign n41213 = ~n20966 & ~n21696 ;
  assign n41214 = n7534 & n41213 ;
  assign n41215 = ~n21692 & n41214 ;
  assign n41216 = \b[60]  & n7973 ;
  assign n41217 = n7970 & n41216 ;
  assign n41218 = ~\a[36]  & \b[61]  ;
  assign n41219 = n7526 & n41218 ;
  assign n41220 = ~n41217 & ~n41219 ;
  assign n41221 = \b[62]  & n7532 ;
  assign n41222 = \a[36]  & \b[61]  ;
  assign n41223 = n17801 & n41222 ;
  assign n41224 = \a[38]  & ~n41223 ;
  assign n41225 = ~n41221 & n41224 ;
  assign n41226 = n41220 & n41225 ;
  assign n41227 = ~n41215 & n41226 ;
  assign n41228 = ~n41212 & n41227 ;
  assign n41229 = ~n41221 & ~n41223 ;
  assign n41230 = n41220 & n41229 ;
  assign n41231 = ~n41215 & n41230 ;
  assign n41232 = ~n41212 & n41231 ;
  assign n41233 = ~\a[38]  & ~n41232 ;
  assign n41234 = ~n41228 & ~n41233 ;
  assign n41235 = ~n41210 & n41234 ;
  assign n41236 = ~n41206 & n41235 ;
  assign n41237 = n41210 & n41234 ;
  assign n41238 = n41206 & n41237 ;
  assign n41239 = ~n41236 & ~n41238 ;
  assign n41240 = ~n41210 & ~n41234 ;
  assign n41241 = n41206 & n41240 ;
  assign n41242 = n41210 & ~n41234 ;
  assign n41243 = ~n41206 & n41242 ;
  assign n41244 = ~n41241 & ~n41243 ;
  assign n41245 = n41239 & n41244 ;
  assign n41246 = n40936 & n41245 ;
  assign n41247 = ~n40936 & ~n41245 ;
  assign n41248 = ~n41246 & ~n41247 ;
  assign n41249 = n40910 & n41248 ;
  assign n41250 = ~n40910 & ~n41248 ;
  assign n41251 = ~n41249 & ~n41250 ;
  assign n41252 = ~n40901 & n41251 ;
  assign n41253 = ~n40908 & n41252 ;
  assign n41254 = ~n40901 & ~n40908 ;
  assign n41255 = ~n41251 & ~n41254 ;
  assign n41256 = ~n41253 & ~n41255 ;
  assign n41257 = ~n41249 & ~n41253 ;
  assign n41258 = ~n11397 & n37945 ;
  assign n41259 = ~n11395 & n41258 ;
  assign n41260 = \b[43]  & n17308 ;
  assign n41261 = n17305 & n41260 ;
  assign n41262 = ~\a[54]  & \b[44]  ;
  assign n41263 = n16647 & n41262 ;
  assign n41264 = ~n41261 & ~n41263 ;
  assign n41265 = \b[45]  & n16653 ;
  assign n41266 = \a[54]  & \b[44]  ;
  assign n41267 = n16644 & n41266 ;
  assign n41268 = \a[56]  & ~n41267 ;
  assign n41269 = ~n41265 & n41268 ;
  assign n41270 = n41264 & n41269 ;
  assign n41271 = ~n41259 & n41270 ;
  assign n41272 = ~n41265 & ~n41267 ;
  assign n41273 = n41264 & n41272 ;
  assign n41274 = ~n41259 & n41273 ;
  assign n41275 = ~\a[56]  & ~n41274 ;
  assign n41276 = ~n41271 & ~n41275 ;
  assign n41277 = n41024 & ~n41047 ;
  assign n41278 = ~n40983 & n41277 ;
  assign n41279 = ~n41049 & ~n41278 ;
  assign n41280 = n41024 & n41047 ;
  assign n41281 = n40983 & n41280 ;
  assign n41282 = ~n41051 & ~n41281 ;
  assign n41283 = n40981 & n41282 ;
  assign n41284 = n41279 & ~n41283 ;
  assign n41285 = ~n41019 & ~n41023 ;
  assign n41286 = ~n41019 & n41047 ;
  assign n41287 = ~n41285 & ~n41286 ;
  assign n41288 = ~n40659 & ~n40988 ;
  assign n41289 = ~n41015 & n41288 ;
  assign n41290 = ~n40989 & ~n41289 ;
  assign n41291 = ~\a[35]  & \b[34]  ;
  assign n41292 = n21957 & n41291 ;
  assign n41293 = ~\a[35]  & \b[35]  ;
  assign n41294 = n21958 & n41293 ;
  assign n41295 = ~n41292 & ~n41294 ;
  assign n41296 = \a[35]  & ~n40986 ;
  assign n41297 = ~n40985 & n41296 ;
  assign n41298 = n41295 & ~n41297 ;
  assign n41299 = \b[36]  & n21958 ;
  assign n41300 = \b[35]  & n21957 ;
  assign n41301 = ~n41299 & ~n41300 ;
  assign n41302 = ~n41298 & ~n41301 ;
  assign n41303 = n41298 & n41301 ;
  assign n41304 = ~n41302 & ~n41303 ;
  assign n41305 = ~n8599 & n20521 ;
  assign n41306 = ~n8174 & n20521 ;
  assign n41307 = ~n8595 & n41306 ;
  assign n41308 = ~n41305 & ~n41307 ;
  assign n41309 = ~n8602 & ~n41308 ;
  assign n41310 = \b[37]  & n21315 ;
  assign n41311 = n21312 & n41310 ;
  assign n41312 = ~\a[60]  & \b[38]  ;
  assign n41313 = n20513 & n41312 ;
  assign n41314 = ~n41311 & ~n41313 ;
  assign n41315 = \b[39]  & n20519 ;
  assign n41316 = \a[60]  & \b[38]  ;
  assign n41317 = n20510 & n41316 ;
  assign n41318 = \a[62]  & ~n41317 ;
  assign n41319 = ~n41315 & n41318 ;
  assign n41320 = n41314 & n41319 ;
  assign n41321 = ~n41309 & n41320 ;
  assign n41322 = ~n41315 & ~n41317 ;
  assign n41323 = n41314 & n41322 ;
  assign n41324 = ~\a[62]  & ~n41323 ;
  assign n41325 = ~\a[62]  & ~n8602 ;
  assign n41326 = ~n41308 & n41325 ;
  assign n41327 = ~n41324 & ~n41326 ;
  assign n41328 = ~n41321 & n41327 ;
  assign n41329 = ~n41304 & n41328 ;
  assign n41330 = n41290 & n41329 ;
  assign n41331 = n41304 & n41328 ;
  assign n41332 = ~n41290 & n41331 ;
  assign n41333 = ~n41330 & ~n41332 ;
  assign n41334 = ~n41290 & n41304 ;
  assign n41335 = ~n40989 & ~n41304 ;
  assign n41336 = ~n41289 & n41335 ;
  assign n41337 = ~n41328 & ~n41336 ;
  assign n41338 = ~n41334 & n41337 ;
  assign n41339 = n41333 & ~n41338 ;
  assign n41340 = ~n9930 & ~n17912 ;
  assign n41341 = ~n18513 & n41340 ;
  assign n41342 = n9927 & n41341 ;
  assign n41343 = n9930 & ~n17912 ;
  assign n41344 = ~n18513 & n41343 ;
  assign n41345 = ~n9927 & n41344 ;
  assign n41346 = ~n41342 & ~n41345 ;
  assign n41347 = \b[40]  & n19183 ;
  assign n41348 = n19180 & n41347 ;
  assign n41349 = \b[42]  & n18514 ;
  assign n41350 = \a[56]  & \b[41]  ;
  assign n41351 = n19181 & n41350 ;
  assign n41352 = ~\a[57]  & \b[41]  ;
  assign n41353 = n18508 & n41352 ;
  assign n41354 = ~n41351 & ~n41353 ;
  assign n41355 = ~n41349 & n41354 ;
  assign n41356 = ~n41348 & n41355 ;
  assign n41357 = n41346 & n41356 ;
  assign n41358 = ~\a[59]  & ~n41357 ;
  assign n41359 = \a[59]  & n41356 ;
  assign n41360 = n41346 & n41359 ;
  assign n41361 = ~n41358 & ~n41360 ;
  assign n41362 = n41339 & ~n41361 ;
  assign n41363 = ~n41339 & n41361 ;
  assign n41364 = ~n41362 & ~n41363 ;
  assign n41365 = n41287 & n41364 ;
  assign n41366 = ~n41287 & ~n41364 ;
  assign n41367 = ~n41365 & ~n41366 ;
  assign n41368 = ~n41284 & ~n41367 ;
  assign n41369 = n41276 & n41368 ;
  assign n41370 = ~n41284 & n41367 ;
  assign n41371 = ~n41276 & n41370 ;
  assign n41372 = ~n41369 & ~n41371 ;
  assign n41373 = n41276 & n41367 ;
  assign n41374 = n41284 & n41373 ;
  assign n41375 = n41284 & ~n41367 ;
  assign n41376 = ~n41276 & n41375 ;
  assign n41377 = ~n41374 & ~n41376 ;
  assign n41378 = n41372 & n41377 ;
  assign n41379 = ~n12478 & ~n14276 ;
  assign n41380 = ~n14790 & n41379 ;
  assign n41381 = n12475 & n41380 ;
  assign n41382 = n12478 & ~n14276 ;
  assign n41383 = ~n14790 & n41382 ;
  assign n41384 = ~n12475 & n41383 ;
  assign n41385 = ~n41381 & ~n41384 ;
  assign n41386 = \b[46]  & n15517 ;
  assign n41387 = n15514 & n41386 ;
  assign n41388 = ~\a[51]  & \b[47]  ;
  assign n41389 = n14785 & n41388 ;
  assign n41390 = ~n41387 & ~n41389 ;
  assign n41391 = \b[48]  & n14791 ;
  assign n41392 = \a[51]  & \b[47]  ;
  assign n41393 = n14782 & n41392 ;
  assign n41394 = \a[53]  & ~n41393 ;
  assign n41395 = ~n41391 & n41394 ;
  assign n41396 = n41390 & n41395 ;
  assign n41397 = n41385 & n41396 ;
  assign n41398 = ~n41391 & ~n41393 ;
  assign n41399 = n41390 & n41398 ;
  assign n41400 = n41385 & n41399 ;
  assign n41401 = ~\a[53]  & ~n41400 ;
  assign n41402 = ~n41397 & ~n41401 ;
  assign n41403 = n41378 & ~n41402 ;
  assign n41404 = ~n41378 & n41402 ;
  assign n41405 = ~n41403 & ~n41404 ;
  assign n41406 = n41061 & ~n41063 ;
  assign n41407 = ~n41061 & n41063 ;
  assign n41408 = n41087 & ~n41407 ;
  assign n41409 = ~n41406 & ~n41408 ;
  assign n41410 = n13125 & ~n14098 ;
  assign n41411 = ~n14096 & n41410 ;
  assign n41412 = \b[49]  & n13794 ;
  assign n41413 = n13792 & n41412 ;
  assign n41414 = ~\a[48]  & \b[50]  ;
  assign n41415 = n13117 & n41414 ;
  assign n41416 = ~n41413 & ~n41415 ;
  assign n41417 = \b[51]  & n13123 ;
  assign n41418 = \a[48]  & \b[50]  ;
  assign n41419 = n13786 & n41418 ;
  assign n41420 = \a[50]  & ~n41419 ;
  assign n41421 = ~n41417 & n41420 ;
  assign n41422 = n41416 & n41421 ;
  assign n41423 = ~n41411 & n41422 ;
  assign n41424 = ~n41417 & ~n41419 ;
  assign n41425 = n41416 & n41424 ;
  assign n41426 = ~n41411 & n41425 ;
  assign n41427 = ~\a[50]  & ~n41426 ;
  assign n41428 = ~n41423 & ~n41427 ;
  assign n41429 = ~n41409 & n41428 ;
  assign n41430 = ~n41405 & n41429 ;
  assign n41431 = n41409 & n41428 ;
  assign n41432 = n41405 & n41431 ;
  assign n41433 = ~n41430 & ~n41432 ;
  assign n41434 = ~n41409 & ~n41428 ;
  assign n41435 = n41405 & n41434 ;
  assign n41436 = n41409 & ~n41428 ;
  assign n41437 = ~n41405 & n41436 ;
  assign n41438 = ~n41435 & ~n41437 ;
  assign n41439 = n41433 & n41438 ;
  assign n41440 = ~n10988 & ~n15241 ;
  assign n41441 = ~n16398 & n41440 ;
  assign n41442 = ~n16404 & n41441 ;
  assign n41443 = ~n11569 & n41442 ;
  assign n41444 = n11572 & n16398 ;
  assign n41445 = n15241 & n41444 ;
  assign n41446 = n16400 & n41444 ;
  assign n41447 = ~n15239 & n41446 ;
  assign n41448 = ~n41445 & ~n41447 ;
  assign n41449 = \b[52]  & n12159 ;
  assign n41450 = n12156 & n41449 ;
  assign n41451 = ~\a[45]  & \b[53]  ;
  assign n41452 = n11564 & n41451 ;
  assign n41453 = ~n41450 & ~n41452 ;
  assign n41454 = \b[54]  & n11570 ;
  assign n41455 = \a[45]  & \b[53]  ;
  assign n41456 = n11561 & n41455 ;
  assign n41457 = \a[47]  & ~n41456 ;
  assign n41458 = ~n41454 & n41457 ;
  assign n41459 = n41453 & n41458 ;
  assign n41460 = n41448 & n41459 ;
  assign n41461 = ~n41443 & n41460 ;
  assign n41462 = ~n41454 & ~n41456 ;
  assign n41463 = n41453 & n41462 ;
  assign n41464 = n41448 & n41463 ;
  assign n41465 = ~n41443 & n41464 ;
  assign n41466 = ~\a[47]  & ~n41465 ;
  assign n41467 = ~n41461 & ~n41466 ;
  assign n41468 = ~n41102 & n41127 ;
  assign n41469 = n41101 & ~n41102 ;
  assign n41470 = ~n41468 & ~n41469 ;
  assign n41471 = ~n41467 & n41470 ;
  assign n41472 = ~n41439 & n41471 ;
  assign n41473 = ~n41467 & ~n41470 ;
  assign n41474 = n41439 & n41473 ;
  assign n41475 = ~n41472 & ~n41474 ;
  assign n41476 = n41467 & ~n41470 ;
  assign n41477 = ~n41439 & n41476 ;
  assign n41478 = n41467 & n41470 ;
  assign n41479 = n41439 & n41478 ;
  assign n41480 = ~n41477 & ~n41479 ;
  assign n41481 = n41475 & n41480 ;
  assign n41482 = ~n41130 & ~n41151 ;
  assign n41483 = n41130 & n41151 ;
  assign n41484 = n41149 & ~n41483 ;
  assign n41485 = ~n41482 & ~n41484 ;
  assign n41486 = n10082 & ~n17690 ;
  assign n41487 = ~n17688 & n41486 ;
  assign n41488 = \b[55]  & n10681 ;
  assign n41489 = n10678 & n41488 ;
  assign n41490 = \b[57]  & n10080 ;
  assign n41491 = \a[41]  & \b[56]  ;
  assign n41492 = n10679 & n41491 ;
  assign n41493 = ~\a[42]  & \b[56]  ;
  assign n41494 = n10074 & n41493 ;
  assign n41495 = ~n41492 & ~n41494 ;
  assign n41496 = ~n41490 & n41495 ;
  assign n41497 = ~n41489 & n41496 ;
  assign n41498 = ~\a[44]  & n41497 ;
  assign n41499 = ~n41487 & n41498 ;
  assign n41500 = ~n41487 & n41497 ;
  assign n41501 = \a[44]  & ~n41500 ;
  assign n41502 = ~n41499 & ~n41501 ;
  assign n41503 = n41485 & n41502 ;
  assign n41504 = ~n41481 & n41503 ;
  assign n41505 = ~n41485 & n41502 ;
  assign n41506 = n41481 & n41505 ;
  assign n41507 = ~n41504 & ~n41506 ;
  assign n41508 = ~n41485 & ~n41502 ;
  assign n41509 = ~n41481 & n41508 ;
  assign n41510 = n41485 & ~n41502 ;
  assign n41511 = n41481 & n41510 ;
  assign n41512 = ~n41509 & ~n41511 ;
  assign n41513 = n41507 & n41512 ;
  assign n41514 = n40957 & ~n41167 ;
  assign n41515 = ~n41167 & n41168 ;
  assign n41516 = ~n41514 & ~n41515 ;
  assign n41517 = n8759 & n20260 ;
  assign n41518 = ~n20257 & n41517 ;
  assign n41519 = n8759 & n40498 ;
  assign n41520 = ~n20256 & n41519 ;
  assign n41521 = \b[58]  & n9301 ;
  assign n41522 = n9298 & n41521 ;
  assign n41523 = ~\a[39]  & \b[59]  ;
  assign n41524 = n8751 & n41523 ;
  assign n41525 = ~n41522 & ~n41524 ;
  assign n41526 = \b[60]  & n8757 ;
  assign n41527 = \a[39]  & \b[59]  ;
  assign n41528 = n8748 & n41527 ;
  assign n41529 = \a[41]  & ~n41528 ;
  assign n41530 = ~n41526 & n41529 ;
  assign n41531 = n41525 & n41530 ;
  assign n41532 = ~n41520 & n41531 ;
  assign n41533 = ~n41518 & n41532 ;
  assign n41534 = ~n41526 & ~n41528 ;
  assign n41535 = n41525 & n41534 ;
  assign n41536 = ~n41520 & n41535 ;
  assign n41537 = ~n41518 & n41536 ;
  assign n41538 = ~\a[41]  & ~n41537 ;
  assign n41539 = ~n41533 & ~n41538 ;
  assign n41540 = n41516 & ~n41539 ;
  assign n41541 = ~n41513 & n41540 ;
  assign n41542 = ~n41516 & ~n41539 ;
  assign n41543 = n41513 & n41542 ;
  assign n41544 = ~n41541 & ~n41543 ;
  assign n41545 = ~n41516 & n41539 ;
  assign n41546 = ~n41513 & n41545 ;
  assign n41547 = n41516 & n41539 ;
  assign n41548 = n41513 & n41547 ;
  assign n41549 = ~n41546 & ~n41548 ;
  assign n41550 = n41544 & n41549 ;
  assign n41551 = ~n41172 & ~n41176 ;
  assign n41552 = n41172 & n41176 ;
  assign n41553 = n41195 & ~n41552 ;
  assign n41554 = ~n41551 & ~n41553 ;
  assign n41555 = ~n41550 & ~n41554 ;
  assign n41556 = n41550 & n41554 ;
  assign n41557 = ~n41555 & ~n41556 ;
  assign n41558 = n7534 & ~n22461 ;
  assign n41559 = ~n22459 & n41558 ;
  assign n41560 = \b[61]  & n7973 ;
  assign n41561 = n7970 & n41560 ;
  assign n41562 = ~\a[36]  & \b[62]  ;
  assign n41563 = n7526 & n41562 ;
  assign n41564 = ~n41561 & ~n41563 ;
  assign n41565 = \b[63]  & n7532 ;
  assign n41566 = \a[36]  & \b[62]  ;
  assign n41567 = n17801 & n41566 ;
  assign n41568 = \a[38]  & ~n41567 ;
  assign n41569 = ~n41565 & n41568 ;
  assign n41570 = n41564 & n41569 ;
  assign n41571 = ~n41559 & n41570 ;
  assign n41572 = ~n41565 & ~n41567 ;
  assign n41573 = n41564 & n41572 ;
  assign n41574 = ~n41559 & n41573 ;
  assign n41575 = ~\a[38]  & ~n41574 ;
  assign n41576 = ~n41571 & ~n41575 ;
  assign n41577 = n41557 & ~n41576 ;
  assign n41578 = ~n41557 & n41576 ;
  assign n41579 = ~n41577 & ~n41578 ;
  assign n41580 = ~n41206 & ~n41210 ;
  assign n41581 = n41206 & n41210 ;
  assign n41582 = n41234 & ~n41581 ;
  assign n41583 = ~n41580 & ~n41582 ;
  assign n41584 = ~n41579 & ~n41583 ;
  assign n41585 = n41579 & n41583 ;
  assign n41586 = ~n41584 & ~n41585 ;
  assign n41587 = ~n40933 & ~n41245 ;
  assign n41588 = ~n40935 & ~n41587 ;
  assign n41589 = n41586 & n41588 ;
  assign n41590 = ~n41586 & ~n41588 ;
  assign n41591 = ~n41589 & ~n41590 ;
  assign n41592 = ~n41257 & n41591 ;
  assign n41593 = ~n41249 & ~n41591 ;
  assign n41594 = ~n41253 & n41593 ;
  assign n41595 = ~n41592 & ~n41594 ;
  assign n41596 = ~n41249 & ~n41589 ;
  assign n41597 = ~n41253 & n41596 ;
  assign n41598 = ~n41577 & ~n41583 ;
  assign n41599 = ~n41578 & ~n41598 ;
  assign n41600 = n41544 & ~n41554 ;
  assign n41601 = n41549 & ~n41600 ;
  assign n41602 = n7534 & ~n22458 ;
  assign n41603 = ~n23173 & n41602 ;
  assign n41604 = \b[62]  & n7973 ;
  assign n41605 = n7970 & n41604 ;
  assign n41606 = \a[36]  & \b[63]  ;
  assign n41607 = n17801 & n41606 ;
  assign n41608 = ~\a[36]  & \b[63]  ;
  assign n41609 = n7526 & n41608 ;
  assign n41610 = \a[38]  & ~n41609 ;
  assign n41611 = ~n41607 & n41610 ;
  assign n41612 = ~n41605 & n41611 ;
  assign n41613 = ~n41603 & n41612 ;
  assign n41614 = ~n41607 & ~n41609 ;
  assign n41615 = ~n41605 & n41614 ;
  assign n41616 = ~n41603 & n41615 ;
  assign n41617 = ~\a[38]  & ~n41616 ;
  assign n41618 = ~n41613 & ~n41617 ;
  assign n41619 = ~n41601 & n41618 ;
  assign n41620 = n41549 & ~n41618 ;
  assign n41621 = ~n41600 & n41620 ;
  assign n41622 = ~n41403 & ~n41409 ;
  assign n41623 = ~n41404 & ~n41622 ;
  assign n41624 = ~n41276 & n41367 ;
  assign n41625 = n41276 & ~n41367 ;
  assign n41626 = ~n41624 & n41625 ;
  assign n41627 = ~n41284 & ~n41624 ;
  assign n41628 = ~n41626 & ~n41627 ;
  assign n41629 = ~n41287 & ~n41362 ;
  assign n41630 = ~n41363 & ~n41629 ;
  assign n41631 = n41328 & ~n41336 ;
  assign n41632 = ~n41334 & ~n41631 ;
  assign n41633 = ~n9044 & ~n19861 ;
  assign n41634 = ~n20518 & n41633 ;
  assign n41635 = n9041 & n41634 ;
  assign n41636 = n9044 & ~n19861 ;
  assign n41637 = ~n20518 & n41636 ;
  assign n41638 = ~n9041 & n41637 ;
  assign n41639 = ~n41635 & ~n41638 ;
  assign n41640 = \b[40]  & n20519 ;
  assign n41641 = \a[60]  & \b[39]  ;
  assign n41642 = n20510 & n41641 ;
  assign n41643 = ~n41640 & ~n41642 ;
  assign n41644 = \b[38]  & n21315 ;
  assign n41645 = n21312 & n41644 ;
  assign n41646 = ~\a[60]  & \b[39]  ;
  assign n41647 = n20513 & n41646 ;
  assign n41648 = ~n41645 & ~n41647 ;
  assign n41649 = n41643 & n41648 ;
  assign n41650 = n41639 & n41649 ;
  assign n41651 = n41295 & n41301 ;
  assign n41652 = n41295 & n41297 ;
  assign n41653 = ~n41651 & ~n41652 ;
  assign n41654 = \b[37]  & n21958 ;
  assign n41655 = \b[36]  & n21957 ;
  assign n41656 = ~n41654 & ~n41655 ;
  assign n41657 = ~\a[62]  & ~n41656 ;
  assign n41658 = n41653 & n41657 ;
  assign n41659 = ~\a[62]  & n41656 ;
  assign n41660 = ~n41653 & n41659 ;
  assign n41661 = ~n41658 & ~n41660 ;
  assign n41662 = ~n41650 & ~n41661 ;
  assign n41663 = \a[62]  & ~n41656 ;
  assign n41664 = n41653 & n41663 ;
  assign n41665 = \a[62]  & n41656 ;
  assign n41666 = ~n41653 & n41665 ;
  assign n41667 = ~n41664 & ~n41666 ;
  assign n41668 = n41649 & ~n41667 ;
  assign n41669 = n41639 & n41668 ;
  assign n41670 = ~n41662 & ~n41669 ;
  assign n41671 = ~\a[62]  & ~n41650 ;
  assign n41672 = n41653 & n41656 ;
  assign n41673 = ~n41653 & ~n41656 ;
  assign n41674 = ~n41672 & ~n41673 ;
  assign n41675 = \a[62]  & n41649 ;
  assign n41676 = n41639 & n41675 ;
  assign n41677 = ~n41674 & ~n41676 ;
  assign n41678 = ~n41671 & n41677 ;
  assign n41679 = n41670 & ~n41678 ;
  assign n41680 = ~n41632 & ~n41679 ;
  assign n41681 = n41632 & n41679 ;
  assign n41682 = ~n41680 & ~n41681 ;
  assign n41683 = ~n10406 & n18516 ;
  assign n41684 = ~n9929 & n18516 ;
  assign n41685 = ~n10402 & n41684 ;
  assign n41686 = ~n41683 & ~n41685 ;
  assign n41687 = ~n10409 & ~n41686 ;
  assign n41688 = \b[43]  & n18514 ;
  assign n41689 = \a[56]  & \b[42]  ;
  assign n41690 = n19181 & n41689 ;
  assign n41691 = ~\a[57]  & \b[42]  ;
  assign n41692 = n18508 & n41691 ;
  assign n41693 = ~n41690 & ~n41692 ;
  assign n41694 = ~n41688 & n41693 ;
  assign n41695 = \b[41]  & n19183 ;
  assign n41696 = n19180 & n41695 ;
  assign n41697 = \a[59]  & ~n41696 ;
  assign n41698 = n41694 & n41697 ;
  assign n41699 = ~n41687 & n41698 ;
  assign n41700 = n41694 & ~n41696 ;
  assign n41701 = ~\a[59]  & ~n41700 ;
  assign n41702 = ~\a[59]  & ~n10409 ;
  assign n41703 = ~n41686 & n41702 ;
  assign n41704 = ~n41701 & ~n41703 ;
  assign n41705 = ~n41699 & n41704 ;
  assign n41706 = n41682 & ~n41705 ;
  assign n41707 = ~n41682 & n41705 ;
  assign n41708 = ~n41706 & ~n41707 ;
  assign n41709 = ~n41630 & ~n41708 ;
  assign n41710 = n41630 & n41708 ;
  assign n41711 = ~n41709 & ~n41710 ;
  assign n41712 = n11906 & n16655 ;
  assign n41713 = ~n11903 & n41712 ;
  assign n41714 = n13483 & n37945 ;
  assign n41715 = ~n11902 & n41714 ;
  assign n41716 = \b[44]  & n17308 ;
  assign n41717 = n17305 & n41716 ;
  assign n41718 = ~\a[54]  & \b[45]  ;
  assign n41719 = n16647 & n41718 ;
  assign n41720 = ~n41717 & ~n41719 ;
  assign n41721 = \b[46]  & n16653 ;
  assign n41722 = \a[54]  & \b[45]  ;
  assign n41723 = n16644 & n41722 ;
  assign n41724 = \a[56]  & ~n41723 ;
  assign n41725 = ~n41721 & n41724 ;
  assign n41726 = n41720 & n41725 ;
  assign n41727 = ~n41715 & n41726 ;
  assign n41728 = ~n41713 & n41727 ;
  assign n41729 = ~n41721 & ~n41723 ;
  assign n41730 = n41720 & n41729 ;
  assign n41731 = ~n41715 & n41730 ;
  assign n41732 = ~n41713 & n41731 ;
  assign n41733 = ~\a[56]  & ~n41732 ;
  assign n41734 = ~n41728 & ~n41733 ;
  assign n41735 = ~n41711 & n41734 ;
  assign n41736 = n41711 & ~n41734 ;
  assign n41737 = ~n41735 & ~n41736 ;
  assign n41738 = ~n41628 & ~n41737 ;
  assign n41739 = n41628 & n41737 ;
  assign n41740 = ~n41738 & ~n41739 ;
  assign n41741 = ~n13524 & n14793 ;
  assign n41742 = ~n13522 & n41741 ;
  assign n41743 = \b[47]  & n15517 ;
  assign n41744 = n15514 & n41743 ;
  assign n41745 = ~\a[51]  & \b[48]  ;
  assign n41746 = n14785 & n41745 ;
  assign n41747 = ~n41744 & ~n41746 ;
  assign n41748 = \b[49]  & n14791 ;
  assign n41749 = \a[51]  & \b[48]  ;
  assign n41750 = n14782 & n41749 ;
  assign n41751 = \a[53]  & ~n41750 ;
  assign n41752 = ~n41748 & n41751 ;
  assign n41753 = n41747 & n41752 ;
  assign n41754 = ~n41742 & n41753 ;
  assign n41755 = ~n41748 & ~n41750 ;
  assign n41756 = n41747 & n41755 ;
  assign n41757 = ~n41742 & n41756 ;
  assign n41758 = ~\a[53]  & ~n41757 ;
  assign n41759 = ~n41754 & ~n41758 ;
  assign n41760 = n41740 & ~n41759 ;
  assign n41761 = ~n41740 & n41759 ;
  assign n41762 = ~n41760 & ~n41761 ;
  assign n41763 = ~n41623 & ~n41762 ;
  assign n41764 = n41623 & n41762 ;
  assign n41765 = ~n41763 & ~n41764 ;
  assign n41766 = ~n12606 & ~n14093 ;
  assign n41767 = ~n15201 & n41766 ;
  assign n41768 = ~n15197 & n41767 ;
  assign n41769 = ~n13122 & n41768 ;
  assign n41770 = n13125 & n15201 ;
  assign n41771 = ~n15198 & n41770 ;
  assign n41772 = ~n41769 & ~n41771 ;
  assign n41773 = \b[50]  & n13794 ;
  assign n41774 = n13792 & n41773 ;
  assign n41775 = ~\a[48]  & \b[51]  ;
  assign n41776 = n13117 & n41775 ;
  assign n41777 = ~n41774 & ~n41776 ;
  assign n41778 = \b[52]  & n13123 ;
  assign n41779 = \a[48]  & \b[51]  ;
  assign n41780 = n13786 & n41779 ;
  assign n41781 = \a[50]  & ~n41780 ;
  assign n41782 = ~n41778 & n41781 ;
  assign n41783 = n41777 & n41782 ;
  assign n41784 = n41772 & n41783 ;
  assign n41785 = ~n41778 & ~n41780 ;
  assign n41786 = n41777 & n41785 ;
  assign n41787 = n41772 & n41786 ;
  assign n41788 = ~\a[50]  & ~n41787 ;
  assign n41789 = ~n41784 & ~n41788 ;
  assign n41790 = ~n41765 & n41789 ;
  assign n41791 = n41765 & ~n41789 ;
  assign n41792 = ~n41790 & ~n41791 ;
  assign n41793 = n11572 & ~n16446 ;
  assign n41794 = ~n16444 & n41793 ;
  assign n41795 = \b[53]  & n12159 ;
  assign n41796 = n12156 & n41795 ;
  assign n41797 = ~\a[45]  & \b[54]  ;
  assign n41798 = n11564 & n41797 ;
  assign n41799 = ~n41796 & ~n41798 ;
  assign n41800 = \b[55]  & n11570 ;
  assign n41801 = \a[45]  & \b[54]  ;
  assign n41802 = n11561 & n41801 ;
  assign n41803 = \a[47]  & ~n41802 ;
  assign n41804 = ~n41800 & n41803 ;
  assign n41805 = n41799 & n41804 ;
  assign n41806 = ~n41794 & n41805 ;
  assign n41807 = ~n41800 & ~n41802 ;
  assign n41808 = n41799 & n41807 ;
  assign n41809 = ~n41794 & n41808 ;
  assign n41810 = ~\a[47]  & ~n41809 ;
  assign n41811 = ~n41806 & ~n41810 ;
  assign n41812 = n41438 & ~n41470 ;
  assign n41813 = n41433 & ~n41812 ;
  assign n41814 = n41811 & n41813 ;
  assign n41815 = ~n41792 & n41814 ;
  assign n41816 = n41811 & ~n41813 ;
  assign n41817 = n41792 & n41816 ;
  assign n41818 = ~n41815 & ~n41817 ;
  assign n41819 = ~n41811 & ~n41813 ;
  assign n41820 = ~n41792 & n41819 ;
  assign n41821 = ~n41811 & n41813 ;
  assign n41822 = n41792 & n41821 ;
  assign n41823 = ~n41820 & ~n41822 ;
  assign n41824 = n41818 & n41823 ;
  assign n41825 = n41475 & ~n41485 ;
  assign n41826 = n41480 & ~n41825 ;
  assign n41827 = n10082 & ~n19543 ;
  assign n41828 = ~n38598 & n41827 ;
  assign n41829 = \b[56]  & n10681 ;
  assign n41830 = n10678 & n41829 ;
  assign n41831 = \b[58]  & n10080 ;
  assign n41832 = \a[41]  & \b[57]  ;
  assign n41833 = n10679 & n41832 ;
  assign n41834 = ~\a[42]  & \b[57]  ;
  assign n41835 = n10074 & n41834 ;
  assign n41836 = ~n41833 & ~n41835 ;
  assign n41837 = ~n41831 & n41836 ;
  assign n41838 = ~n41830 & n41837 ;
  assign n41839 = ~n41828 & n41838 ;
  assign n41840 = ~\a[44]  & ~n41839 ;
  assign n41841 = \a[44]  & n41838 ;
  assign n41842 = ~n41828 & n41841 ;
  assign n41843 = ~n41840 & ~n41842 ;
  assign n41844 = ~n41826 & ~n41843 ;
  assign n41845 = ~n41824 & n41844 ;
  assign n41846 = n41826 & ~n41843 ;
  assign n41847 = n41824 & n41846 ;
  assign n41848 = ~n41845 & ~n41847 ;
  assign n41849 = n41826 & n41843 ;
  assign n41850 = ~n41824 & n41849 ;
  assign n41851 = ~n41826 & n41843 ;
  assign n41852 = n41824 & n41851 ;
  assign n41853 = ~n41850 & ~n41852 ;
  assign n41854 = n41848 & n41853 ;
  assign n41855 = n41507 & ~n41516 ;
  assign n41856 = n41512 & ~n41855 ;
  assign n41857 = n8759 & ~n20971 ;
  assign n41858 = ~n20969 & n41857 ;
  assign n41859 = \b[59]  & n9301 ;
  assign n41860 = n9298 & n41859 ;
  assign n41861 = ~\a[39]  & \b[60]  ;
  assign n41862 = n8751 & n41861 ;
  assign n41863 = ~n41860 & ~n41862 ;
  assign n41864 = \b[61]  & n8757 ;
  assign n41865 = \a[39]  & \b[60]  ;
  assign n41866 = n8748 & n41865 ;
  assign n41867 = \a[41]  & ~n41866 ;
  assign n41868 = ~n41864 & n41867 ;
  assign n41869 = n41863 & n41868 ;
  assign n41870 = ~n41858 & n41869 ;
  assign n41871 = ~n41864 & ~n41866 ;
  assign n41872 = n41863 & n41871 ;
  assign n41873 = ~n41858 & n41872 ;
  assign n41874 = ~\a[41]  & ~n41873 ;
  assign n41875 = ~n41870 & ~n41874 ;
  assign n41876 = n41856 & ~n41875 ;
  assign n41877 = ~n41854 & n41876 ;
  assign n41878 = ~n41856 & ~n41875 ;
  assign n41879 = n41854 & n41878 ;
  assign n41880 = ~n41877 & ~n41879 ;
  assign n41881 = ~n41856 & n41875 ;
  assign n41882 = ~n41854 & n41881 ;
  assign n41883 = n41856 & n41875 ;
  assign n41884 = n41854 & n41883 ;
  assign n41885 = ~n41882 & ~n41884 ;
  assign n41886 = n41880 & n41885 ;
  assign n41887 = ~n41621 & n41886 ;
  assign n41888 = ~n41619 & n41887 ;
  assign n41889 = ~n41619 & ~n41621 ;
  assign n41890 = ~n41886 & ~n41889 ;
  assign n41891 = ~n41888 & ~n41890 ;
  assign n41892 = ~n41599 & ~n41891 ;
  assign n41893 = n41599 & n41891 ;
  assign n41894 = ~n41892 & ~n41893 ;
  assign n41895 = ~n41590 & n41894 ;
  assign n41896 = ~n41597 & n41895 ;
  assign n41897 = ~n41590 & ~n41597 ;
  assign n41898 = ~n41894 & ~n41897 ;
  assign n41899 = ~n41896 & ~n41898 ;
  assign n41900 = ~n41893 & ~n41896 ;
  assign n41901 = ~n41621 & ~n41886 ;
  assign n41902 = ~n41619 & ~n41901 ;
  assign n41903 = n41854 & n41856 ;
  assign n41904 = n41875 & ~n41903 ;
  assign n41905 = ~n41854 & ~n41856 ;
  assign n41906 = n7534 & n39033 ;
  assign n41907 = ~n23171 & n41906 ;
  assign n41908 = \a[35]  & \a[37]  ;
  assign n41909 = \a[36]  & ~\a[38]  ;
  assign n41910 = n41908 & n41909 ;
  assign n41911 = ~\a[35]  & ~\a[37]  ;
  assign n41912 = ~\a[36]  & \a[38]  ;
  assign n41913 = n41911 & n41912 ;
  assign n41914 = ~n41910 & ~n41913 ;
  assign n41915 = \b[63]  & ~n41914 ;
  assign n41916 = \a[38]  & ~n41915 ;
  assign n41917 = ~n41907 & n41916 ;
  assign n41918 = ~n41907 & ~n41915 ;
  assign n41919 = ~\a[38]  & ~n41918 ;
  assign n41920 = ~n41917 & ~n41919 ;
  assign n41921 = ~n41905 & ~n41920 ;
  assign n41922 = ~n41904 & n41921 ;
  assign n41923 = ~n41904 & ~n41905 ;
  assign n41924 = n41920 & ~n41923 ;
  assign n41925 = ~n41922 & ~n41924 ;
  assign n41926 = ~n41792 & ~n41813 ;
  assign n41927 = n41792 & n41813 ;
  assign n41928 = n41811 & ~n41927 ;
  assign n41929 = ~n41926 & ~n41928 ;
  assign n41930 = ~n10889 & ~n17912 ;
  assign n41931 = ~n18513 & n41930 ;
  assign n41932 = n10886 & n41931 ;
  assign n41933 = n10889 & ~n17912 ;
  assign n41934 = ~n18513 & n41933 ;
  assign n41935 = ~n10886 & n41934 ;
  assign n41936 = ~n41932 & ~n41935 ;
  assign n41937 = \b[44]  & n18514 ;
  assign n41938 = \a[56]  & \b[43]  ;
  assign n41939 = n19181 & n41938 ;
  assign n41940 = ~\a[57]  & \b[43]  ;
  assign n41941 = n18508 & n41940 ;
  assign n41942 = ~n41939 & ~n41941 ;
  assign n41943 = ~n41937 & n41942 ;
  assign n41944 = \b[42]  & n19183 ;
  assign n41945 = n19180 & n41944 ;
  assign n41946 = \a[59]  & ~n41945 ;
  assign n41947 = n41943 & n41946 ;
  assign n41948 = n41936 & n41947 ;
  assign n41949 = n41943 & ~n41945 ;
  assign n41950 = n41936 & n41949 ;
  assign n41951 = ~\a[59]  & ~n41950 ;
  assign n41952 = ~n41948 & ~n41951 ;
  assign n41953 = ~n9479 & n20521 ;
  assign n41954 = ~n9043 & n20521 ;
  assign n41955 = ~n9475 & n41954 ;
  assign n41956 = ~n41953 & ~n41955 ;
  assign n41957 = ~n9482 & ~n41956 ;
  assign n41958 = \b[39]  & n21315 ;
  assign n41959 = n21312 & n41958 ;
  assign n41960 = ~\a[60]  & \b[40]  ;
  assign n41961 = n20513 & n41960 ;
  assign n41962 = ~n41959 & ~n41961 ;
  assign n41963 = \b[41]  & n20519 ;
  assign n41964 = \a[60]  & \b[40]  ;
  assign n41965 = n20510 & n41964 ;
  assign n41966 = \a[62]  & ~n41965 ;
  assign n41967 = ~n41963 & n41966 ;
  assign n41968 = n41962 & n41967 ;
  assign n41969 = ~n41957 & n41968 ;
  assign n41970 = ~n41963 & ~n41965 ;
  assign n41971 = n41962 & n41970 ;
  assign n41972 = ~\a[62]  & ~n41971 ;
  assign n41973 = ~\a[62]  & ~n9482 ;
  assign n41974 = ~n41956 & n41973 ;
  assign n41975 = ~n41972 & ~n41974 ;
  assign n41976 = ~n41969 & n41975 ;
  assign n41977 = ~n41669 & ~n41672 ;
  assign n41978 = ~n41662 & n41977 ;
  assign n41979 = \b[38]  & n21958 ;
  assign n41980 = \b[37]  & n21957 ;
  assign n41981 = ~n41979 & ~n41980 ;
  assign n41982 = n41656 & ~n41981 ;
  assign n41983 = ~n41656 & n41981 ;
  assign n41984 = ~n41982 & ~n41983 ;
  assign n41985 = n41978 & n41984 ;
  assign n41986 = ~n41978 & ~n41984 ;
  assign n41987 = ~n41985 & ~n41986 ;
  assign n41988 = ~n41976 & ~n41987 ;
  assign n41989 = n41976 & n41987 ;
  assign n41990 = ~n41988 & ~n41989 ;
  assign n41991 = n41952 & n41990 ;
  assign n41992 = ~n41952 & ~n41990 ;
  assign n41993 = ~n41991 & ~n41992 ;
  assign n41994 = ~n41681 & n41705 ;
  assign n41995 = ~n41680 & ~n41994 ;
  assign n41996 = n41993 & ~n41995 ;
  assign n41997 = ~n41993 & n41995 ;
  assign n41998 = ~n41996 & ~n41997 ;
  assign n41999 = ~n12438 & n16655 ;
  assign n42000 = ~n12436 & n41999 ;
  assign n42001 = \b[45]  & n17308 ;
  assign n42002 = n17305 & n42001 ;
  assign n42003 = ~\a[54]  & \b[46]  ;
  assign n42004 = n16647 & n42003 ;
  assign n42005 = ~n42002 & ~n42004 ;
  assign n42006 = \b[47]  & n16653 ;
  assign n42007 = \a[54]  & \b[46]  ;
  assign n42008 = n16644 & n42007 ;
  assign n42009 = \a[56]  & ~n42008 ;
  assign n42010 = ~n42006 & n42009 ;
  assign n42011 = n42005 & n42010 ;
  assign n42012 = ~n42000 & n42011 ;
  assign n42013 = ~n42006 & ~n42008 ;
  assign n42014 = n42005 & n42013 ;
  assign n42015 = ~n42000 & n42014 ;
  assign n42016 = ~\a[56]  & ~n42015 ;
  assign n42017 = ~n42012 & ~n42016 ;
  assign n42018 = ~n41998 & n42017 ;
  assign n42019 = n41998 & ~n42017 ;
  assign n42020 = ~n42018 & ~n42019 ;
  assign n42021 = ~n41710 & n41734 ;
  assign n42022 = ~n41709 & ~n42021 ;
  assign n42023 = ~n42020 & ~n42022 ;
  assign n42024 = n42020 & n42022 ;
  assign n42025 = ~n42023 & ~n42024 ;
  assign n42026 = ~n14052 & ~n14276 ;
  assign n42027 = ~n14790 & n42026 ;
  assign n42028 = n14049 & n42027 ;
  assign n42029 = n14052 & ~n14276 ;
  assign n42030 = ~n14790 & n42029 ;
  assign n42031 = ~n14049 & n42030 ;
  assign n42032 = ~n42028 & ~n42031 ;
  assign n42033 = \b[48]  & n15517 ;
  assign n42034 = n15514 & n42033 ;
  assign n42035 = ~\a[51]  & \b[49]  ;
  assign n42036 = n14785 & n42035 ;
  assign n42037 = ~n42034 & ~n42036 ;
  assign n42038 = \b[50]  & n14791 ;
  assign n42039 = \a[51]  & \b[49]  ;
  assign n42040 = n14782 & n42039 ;
  assign n42041 = \a[53]  & ~n42040 ;
  assign n42042 = ~n42038 & n42041 ;
  assign n42043 = n42037 & n42042 ;
  assign n42044 = n42032 & n42043 ;
  assign n42045 = ~n42038 & ~n42040 ;
  assign n42046 = n42037 & n42045 ;
  assign n42047 = n42032 & n42046 ;
  assign n42048 = ~\a[53]  & ~n42047 ;
  assign n42049 = ~n42044 & ~n42048 ;
  assign n42050 = ~n42025 & n42049 ;
  assign n42051 = n42025 & ~n42049 ;
  assign n42052 = ~n42050 & ~n42051 ;
  assign n42053 = n13125 & ~n15246 ;
  assign n42054 = ~n15244 & n42053 ;
  assign n42055 = \b[51]  & n13794 ;
  assign n42056 = n13792 & n42055 ;
  assign n42057 = ~\a[48]  & \b[52]  ;
  assign n42058 = n13117 & n42057 ;
  assign n42059 = ~n42056 & ~n42058 ;
  assign n42060 = \b[53]  & n13123 ;
  assign n42061 = \a[48]  & \b[52]  ;
  assign n42062 = n13786 & n42061 ;
  assign n42063 = \a[50]  & ~n42062 ;
  assign n42064 = ~n42060 & n42063 ;
  assign n42065 = n42059 & n42064 ;
  assign n42066 = ~n42054 & n42065 ;
  assign n42067 = ~n42060 & ~n42062 ;
  assign n42068 = n42059 & n42067 ;
  assign n42069 = ~n42054 & n42068 ;
  assign n42070 = ~\a[50]  & ~n42069 ;
  assign n42071 = ~n42066 & ~n42070 ;
  assign n42072 = ~n41739 & n41759 ;
  assign n42073 = ~n41738 & ~n42072 ;
  assign n42074 = n42071 & ~n42073 ;
  assign n42075 = n42052 & n42074 ;
  assign n42076 = n42071 & n42073 ;
  assign n42077 = ~n42052 & n42076 ;
  assign n42078 = ~n42075 & ~n42077 ;
  assign n42079 = ~n42071 & ~n42073 ;
  assign n42080 = ~n42052 & n42079 ;
  assign n42081 = ~n42071 & n42073 ;
  assign n42082 = n42052 & n42081 ;
  assign n42083 = ~n42080 & ~n42082 ;
  assign n42084 = n42078 & n42083 ;
  assign n42085 = ~n10988 & ~n16441 ;
  assign n42086 = ~n17647 & n42085 ;
  assign n42087 = ~n17643 & n42086 ;
  assign n42088 = ~n11569 & n42087 ;
  assign n42089 = n11572 & n17647 ;
  assign n42090 = ~n17644 & n42089 ;
  assign n42091 = ~n42088 & ~n42090 ;
  assign n42092 = \b[54]  & n12159 ;
  assign n42093 = n12156 & n42092 ;
  assign n42094 = ~\a[45]  & \b[55]  ;
  assign n42095 = n11564 & n42094 ;
  assign n42096 = ~n42093 & ~n42095 ;
  assign n42097 = \b[56]  & n11570 ;
  assign n42098 = \a[45]  & \b[55]  ;
  assign n42099 = n11561 & n42098 ;
  assign n42100 = \a[47]  & ~n42099 ;
  assign n42101 = ~n42097 & n42100 ;
  assign n42102 = n42096 & n42101 ;
  assign n42103 = n42091 & n42102 ;
  assign n42104 = ~n42097 & ~n42099 ;
  assign n42105 = n42096 & n42104 ;
  assign n42106 = n42091 & n42105 ;
  assign n42107 = ~\a[47]  & ~n42106 ;
  assign n42108 = ~n42103 & ~n42107 ;
  assign n42109 = ~n41764 & n41789 ;
  assign n42110 = ~n41763 & ~n42109 ;
  assign n42111 = ~n42108 & ~n42110 ;
  assign n42112 = ~n42084 & n42111 ;
  assign n42113 = ~n42108 & n42110 ;
  assign n42114 = n42084 & n42113 ;
  assign n42115 = ~n42112 & ~n42114 ;
  assign n42116 = n42108 & ~n42110 ;
  assign n42117 = n42084 & n42116 ;
  assign n42118 = n42108 & n42110 ;
  assign n42119 = ~n42084 & n42118 ;
  assign n42120 = ~n42117 & ~n42119 ;
  assign n42121 = n42115 & n42120 ;
  assign n42122 = n41929 & n42121 ;
  assign n42123 = ~n41929 & ~n42121 ;
  assign n42124 = ~n42122 & ~n42123 ;
  assign n42125 = n10082 & ~n19550 ;
  assign n42126 = ~n19548 & n42125 ;
  assign n42127 = \b[59]  & n10080 ;
  assign n42128 = \a[41]  & \b[58]  ;
  assign n42129 = n10679 & n42128 ;
  assign n42130 = ~\a[42]  & \b[58]  ;
  assign n42131 = n10074 & n42130 ;
  assign n42132 = ~n42129 & ~n42131 ;
  assign n42133 = ~n42127 & n42132 ;
  assign n42134 = \b[57]  & n10681 ;
  assign n42135 = n10678 & n42134 ;
  assign n42136 = \a[44]  & ~n42135 ;
  assign n42137 = n42133 & n42136 ;
  assign n42138 = ~n42126 & n42137 ;
  assign n42139 = n42133 & ~n42135 ;
  assign n42140 = ~n42126 & n42139 ;
  assign n42141 = ~\a[44]  & ~n42140 ;
  assign n42142 = ~n42138 & ~n42141 ;
  assign n42143 = n42124 & ~n42142 ;
  assign n42144 = ~n42124 & n42142 ;
  assign n42145 = ~n42143 & ~n42144 ;
  assign n42146 = n41824 & ~n41826 ;
  assign n42147 = ~n41824 & n41826 ;
  assign n42148 = n41843 & ~n42147 ;
  assign n42149 = ~n42146 & ~n42148 ;
  assign n42150 = ~n8272 & ~n20966 ;
  assign n42151 = ~n21696 & n42150 ;
  assign n42152 = ~n21692 & n42151 ;
  assign n42153 = ~n8756 & n42152 ;
  assign n42154 = n8759 & n21696 ;
  assign n42155 = ~n21693 & n42154 ;
  assign n42156 = ~n42153 & ~n42155 ;
  assign n42157 = \b[60]  & n9301 ;
  assign n42158 = n9298 & n42157 ;
  assign n42159 = ~\a[39]  & \b[61]  ;
  assign n42160 = n8751 & n42159 ;
  assign n42161 = ~n42158 & ~n42160 ;
  assign n42162 = \b[62]  & n8757 ;
  assign n42163 = \a[39]  & \b[61]  ;
  assign n42164 = n8748 & n42163 ;
  assign n42165 = \a[41]  & ~n42164 ;
  assign n42166 = ~n42162 & n42165 ;
  assign n42167 = n42161 & n42166 ;
  assign n42168 = n42156 & n42167 ;
  assign n42169 = ~n42162 & ~n42164 ;
  assign n42170 = n42161 & n42169 ;
  assign n42171 = n42156 & n42170 ;
  assign n42172 = ~\a[41]  & ~n42171 ;
  assign n42173 = ~n42168 & ~n42172 ;
  assign n42174 = ~n42149 & n42173 ;
  assign n42175 = ~n42145 & n42174 ;
  assign n42176 = n42149 & n42173 ;
  assign n42177 = n42145 & n42176 ;
  assign n42178 = ~n42175 & ~n42177 ;
  assign n42179 = ~n42149 & ~n42173 ;
  assign n42180 = n42145 & n42179 ;
  assign n42181 = n42149 & ~n42173 ;
  assign n42182 = ~n42145 & n42181 ;
  assign n42183 = ~n42180 & ~n42182 ;
  assign n42184 = n42178 & n42183 ;
  assign n42185 = n41925 & n42184 ;
  assign n42186 = ~n41925 & ~n42184 ;
  assign n42187 = ~n42185 & ~n42186 ;
  assign n42188 = n41902 & n42187 ;
  assign n42189 = ~n41902 & ~n42187 ;
  assign n42190 = ~n42188 & ~n42189 ;
  assign n42191 = ~n41900 & n42190 ;
  assign n42192 = ~n41893 & ~n42190 ;
  assign n42193 = ~n41896 & n42192 ;
  assign n42194 = ~n42191 & ~n42193 ;
  assign n42195 = ~n41893 & ~n42188 ;
  assign n42196 = ~n41896 & n42195 ;
  assign n42197 = ~n12478 & ~n16016 ;
  assign n42198 = ~n16652 & n42197 ;
  assign n42199 = n12475 & n42198 ;
  assign n42200 = n12478 & ~n16016 ;
  assign n42201 = ~n16652 & n42200 ;
  assign n42202 = ~n12475 & n42201 ;
  assign n42203 = ~n42199 & ~n42202 ;
  assign n42204 = \b[46]  & n17308 ;
  assign n42205 = n17305 & n42204 ;
  assign n42206 = ~\a[54]  & \b[47]  ;
  assign n42207 = n16647 & n42206 ;
  assign n42208 = ~n42205 & ~n42207 ;
  assign n42209 = \b[48]  & n16653 ;
  assign n42210 = \a[54]  & \b[47]  ;
  assign n42211 = n16644 & n42210 ;
  assign n42212 = \a[56]  & ~n42211 ;
  assign n42213 = ~n42209 & n42212 ;
  assign n42214 = n42208 & n42213 ;
  assign n42215 = n42203 & n42214 ;
  assign n42216 = ~n42209 & ~n42211 ;
  assign n42217 = n42208 & n42216 ;
  assign n42218 = n42203 & n42217 ;
  assign n42219 = ~\a[56]  & ~n42218 ;
  assign n42220 = ~n42215 & ~n42219 ;
  assign n42221 = ~n11397 & n18516 ;
  assign n42222 = ~n11395 & n42221 ;
  assign n42223 = \b[45]  & n18514 ;
  assign n42224 = \a[56]  & \b[44]  ;
  assign n42225 = n19181 & n42224 ;
  assign n42226 = ~\a[57]  & \b[44]  ;
  assign n42227 = n18508 & n42226 ;
  assign n42228 = ~n42225 & ~n42227 ;
  assign n42229 = ~n42223 & n42228 ;
  assign n42230 = \b[43]  & n19183 ;
  assign n42231 = n19180 & n42230 ;
  assign n42232 = \a[59]  & ~n42231 ;
  assign n42233 = n42229 & n42232 ;
  assign n42234 = ~n42222 & n42233 ;
  assign n42235 = n42229 & ~n42231 ;
  assign n42236 = ~n42222 & n42235 ;
  assign n42237 = ~\a[59]  & ~n42236 ;
  assign n42238 = ~n42234 & ~n42237 ;
  assign n42239 = ~n41672 & ~n41982 ;
  assign n42240 = ~n41669 & n42239 ;
  assign n42241 = ~n41662 & n42240 ;
  assign n42242 = ~\a[38]  & n41655 ;
  assign n42243 = ~\a[38]  & \b[37]  ;
  assign n42244 = n21958 & n42243 ;
  assign n42245 = ~n42242 & ~n42244 ;
  assign n42246 = \a[38]  & ~n41655 ;
  assign n42247 = ~n41654 & n42246 ;
  assign n42248 = n42245 & ~n42247 ;
  assign n42249 = \b[39]  & n21958 ;
  assign n42250 = \b[38]  & n21957 ;
  assign n42251 = ~n42249 & ~n42250 ;
  assign n42252 = ~n42248 & ~n42251 ;
  assign n42253 = n42248 & n42251 ;
  assign n42254 = ~n42252 & ~n42253 ;
  assign n42255 = ~n41983 & ~n42254 ;
  assign n42256 = ~n42241 & n42255 ;
  assign n42257 = ~n41983 & ~n42241 ;
  assign n42258 = n42254 & ~n42257 ;
  assign n42259 = ~n42256 & ~n42258 ;
  assign n42260 = ~n9930 & ~n19861 ;
  assign n42261 = ~n20518 & n42260 ;
  assign n42262 = n9927 & n42261 ;
  assign n42263 = n9930 & ~n19861 ;
  assign n42264 = ~n20518 & n42263 ;
  assign n42265 = ~n9927 & n42264 ;
  assign n42266 = ~n42262 & ~n42265 ;
  assign n42267 = \b[40]  & n21315 ;
  assign n42268 = n21312 & n42267 ;
  assign n42269 = ~\a[60]  & \b[41]  ;
  assign n42270 = n20513 & n42269 ;
  assign n42271 = ~n42268 & ~n42270 ;
  assign n42272 = \b[42]  & n20519 ;
  assign n42273 = \a[60]  & \b[41]  ;
  assign n42274 = n20510 & n42273 ;
  assign n42275 = \a[62]  & ~n42274 ;
  assign n42276 = ~n42272 & n42275 ;
  assign n42277 = n42271 & n42276 ;
  assign n42278 = n42266 & n42277 ;
  assign n42279 = ~n42272 & ~n42274 ;
  assign n42280 = n42271 & n42279 ;
  assign n42281 = n42266 & n42280 ;
  assign n42282 = ~\a[62]  & ~n42281 ;
  assign n42283 = ~n42278 & ~n42282 ;
  assign n42284 = n42259 & ~n42283 ;
  assign n42285 = ~n42259 & n42283 ;
  assign n42286 = ~n42284 & ~n42285 ;
  assign n42287 = ~n42238 & n42286 ;
  assign n42288 = n42238 & ~n42286 ;
  assign n42289 = n41952 & ~n41988 ;
  assign n42290 = ~n41989 & ~n42289 ;
  assign n42291 = ~n42288 & n42290 ;
  assign n42292 = ~n42287 & n42291 ;
  assign n42293 = n42288 & ~n42290 ;
  assign n42294 = n42287 & ~n42290 ;
  assign n42295 = ~n42293 & ~n42294 ;
  assign n42296 = ~n42292 & n42295 ;
  assign n42297 = ~n42220 & n42296 ;
  assign n42298 = n42220 & ~n42296 ;
  assign n42299 = ~n42297 & ~n42298 ;
  assign n42300 = ~n41997 & n42017 ;
  assign n42301 = ~n41996 & ~n42300 ;
  assign n42302 = ~n42299 & ~n42301 ;
  assign n42303 = n42299 & n42301 ;
  assign n42304 = ~n42302 & ~n42303 ;
  assign n42305 = ~n14098 & n14793 ;
  assign n42306 = ~n14096 & n42305 ;
  assign n42307 = \b[49]  & n15517 ;
  assign n42308 = n15514 & n42307 ;
  assign n42309 = ~\a[51]  & \b[50]  ;
  assign n42310 = n14785 & n42309 ;
  assign n42311 = ~n42308 & ~n42310 ;
  assign n42312 = \b[51]  & n14791 ;
  assign n42313 = \a[51]  & \b[50]  ;
  assign n42314 = n14782 & n42313 ;
  assign n42315 = \a[53]  & ~n42314 ;
  assign n42316 = ~n42312 & n42315 ;
  assign n42317 = n42311 & n42316 ;
  assign n42318 = ~n42306 & n42317 ;
  assign n42319 = ~n42312 & ~n42314 ;
  assign n42320 = n42311 & n42319 ;
  assign n42321 = ~n42306 & n42320 ;
  assign n42322 = ~\a[53]  & ~n42321 ;
  assign n42323 = ~n42318 & ~n42322 ;
  assign n42324 = ~n42304 & n42323 ;
  assign n42325 = n42304 & ~n42323 ;
  assign n42326 = ~n42324 & ~n42325 ;
  assign n42327 = ~n12606 & ~n15241 ;
  assign n42328 = ~n16398 & n42327 ;
  assign n42329 = ~n16404 & n42328 ;
  assign n42330 = ~n13122 & n42329 ;
  assign n42331 = n13125 & n16398 ;
  assign n42332 = n15241 & n42331 ;
  assign n42333 = n16400 & n42331 ;
  assign n42334 = ~n15239 & n42333 ;
  assign n42335 = ~n42332 & ~n42334 ;
  assign n42336 = \b[52]  & n13794 ;
  assign n42337 = n13792 & n42336 ;
  assign n42338 = ~\a[48]  & \b[53]  ;
  assign n42339 = n13117 & n42338 ;
  assign n42340 = ~n42337 & ~n42339 ;
  assign n42341 = \b[54]  & n13123 ;
  assign n42342 = \a[48]  & \b[53]  ;
  assign n42343 = n13786 & n42342 ;
  assign n42344 = \a[50]  & ~n42343 ;
  assign n42345 = ~n42341 & n42344 ;
  assign n42346 = n42340 & n42345 ;
  assign n42347 = n42335 & n42346 ;
  assign n42348 = ~n42330 & n42347 ;
  assign n42349 = ~n42341 & ~n42343 ;
  assign n42350 = n42340 & n42349 ;
  assign n42351 = n42335 & n42350 ;
  assign n42352 = ~n42330 & n42351 ;
  assign n42353 = ~\a[50]  & ~n42352 ;
  assign n42354 = ~n42348 & ~n42353 ;
  assign n42355 = ~n42024 & n42049 ;
  assign n42356 = n42023 & ~n42024 ;
  assign n42357 = ~n42355 & ~n42356 ;
  assign n42358 = ~n42354 & n42357 ;
  assign n42359 = ~n42326 & n42358 ;
  assign n42360 = ~n42354 & ~n42357 ;
  assign n42361 = n42326 & n42360 ;
  assign n42362 = ~n42359 & ~n42361 ;
  assign n42363 = n42354 & ~n42357 ;
  assign n42364 = ~n42326 & n42363 ;
  assign n42365 = n42354 & n42357 ;
  assign n42366 = n42326 & n42365 ;
  assign n42367 = ~n42364 & ~n42366 ;
  assign n42368 = n42362 & n42367 ;
  assign n42369 = ~n42052 & ~n42073 ;
  assign n42370 = n42052 & n42073 ;
  assign n42371 = n42071 & ~n42370 ;
  assign n42372 = ~n42369 & ~n42371 ;
  assign n42373 = n11572 & ~n17690 ;
  assign n42374 = ~n17688 & n42373 ;
  assign n42375 = \b[55]  & n12159 ;
  assign n42376 = n12156 & n42375 ;
  assign n42377 = ~\a[45]  & \b[56]  ;
  assign n42378 = n11564 & n42377 ;
  assign n42379 = ~n42376 & ~n42378 ;
  assign n42380 = \b[57]  & n11570 ;
  assign n42381 = \a[45]  & \b[56]  ;
  assign n42382 = n11561 & n42381 ;
  assign n42383 = \a[47]  & ~n42382 ;
  assign n42384 = ~n42380 & n42383 ;
  assign n42385 = n42379 & n42384 ;
  assign n42386 = ~n42374 & n42385 ;
  assign n42387 = ~n42380 & ~n42382 ;
  assign n42388 = n42379 & n42387 ;
  assign n42389 = ~n42374 & n42388 ;
  assign n42390 = ~\a[47]  & ~n42389 ;
  assign n42391 = ~n42386 & ~n42390 ;
  assign n42392 = n42372 & ~n42391 ;
  assign n42393 = ~n42368 & n42392 ;
  assign n42394 = ~n42372 & ~n42391 ;
  assign n42395 = n42368 & n42394 ;
  assign n42396 = ~n42393 & ~n42395 ;
  assign n42397 = ~n42372 & n42391 ;
  assign n42398 = ~n42368 & n42397 ;
  assign n42399 = n42372 & n42391 ;
  assign n42400 = n42368 & n42399 ;
  assign n42401 = ~n42398 & ~n42400 ;
  assign n42402 = n42396 & n42401 ;
  assign n42403 = ~n42084 & n42110 ;
  assign n42404 = n42115 & ~n42403 ;
  assign n42405 = n10082 & n20260 ;
  assign n42406 = ~n20257 & n42405 ;
  assign n42407 = n10082 & n40498 ;
  assign n42408 = ~n20256 & n42407 ;
  assign n42409 = \b[58]  & n10681 ;
  assign n42410 = n10678 & n42409 ;
  assign n42411 = \b[60]  & n10080 ;
  assign n42412 = \a[41]  & \b[59]  ;
  assign n42413 = n10679 & n42412 ;
  assign n42414 = ~\a[42]  & \b[59]  ;
  assign n42415 = n10074 & n42414 ;
  assign n42416 = ~n42413 & ~n42415 ;
  assign n42417 = ~n42411 & n42416 ;
  assign n42418 = ~n42410 & n42417 ;
  assign n42419 = ~n42408 & n42418 ;
  assign n42420 = ~n42406 & n42419 ;
  assign n42421 = ~\a[44]  & ~n42420 ;
  assign n42422 = \a[44]  & n42418 ;
  assign n42423 = ~n42408 & n42422 ;
  assign n42424 = ~n42406 & n42423 ;
  assign n42425 = ~n42421 & ~n42424 ;
  assign n42426 = ~n42404 & ~n42425 ;
  assign n42427 = ~n42402 & n42426 ;
  assign n42428 = n42404 & ~n42425 ;
  assign n42429 = n42402 & n42428 ;
  assign n42430 = ~n42427 & ~n42429 ;
  assign n42431 = n42404 & n42425 ;
  assign n42432 = ~n42402 & n42431 ;
  assign n42433 = ~n42404 & n42425 ;
  assign n42434 = n42402 & n42433 ;
  assign n42435 = ~n42432 & ~n42434 ;
  assign n42436 = n42430 & n42435 ;
  assign n42437 = ~n42122 & n42142 ;
  assign n42438 = ~n42123 & ~n42437 ;
  assign n42439 = n8759 & ~n22461 ;
  assign n42440 = ~n22459 & n42439 ;
  assign n42441 = \b[61]  & n9301 ;
  assign n42442 = n9298 & n42441 ;
  assign n42443 = ~\a[39]  & \b[62]  ;
  assign n42444 = n8751 & n42443 ;
  assign n42445 = ~n42442 & ~n42444 ;
  assign n42446 = \b[63]  & n8757 ;
  assign n42447 = \a[39]  & \b[62]  ;
  assign n42448 = n8748 & n42447 ;
  assign n42449 = \a[41]  & ~n42448 ;
  assign n42450 = ~n42446 & n42449 ;
  assign n42451 = n42445 & n42450 ;
  assign n42452 = ~n42440 & n42451 ;
  assign n42453 = ~n42446 & ~n42448 ;
  assign n42454 = n42445 & n42453 ;
  assign n42455 = ~n42440 & n42454 ;
  assign n42456 = ~\a[41]  & ~n42455 ;
  assign n42457 = ~n42452 & ~n42456 ;
  assign n42458 = ~n42438 & ~n42457 ;
  assign n42459 = n42436 & n42458 ;
  assign n42460 = n42438 & ~n42457 ;
  assign n42461 = ~n42436 & n42460 ;
  assign n42462 = ~n42459 & ~n42461 ;
  assign n42463 = ~n42438 & n42457 ;
  assign n42464 = ~n42436 & n42463 ;
  assign n42465 = n42438 & n42457 ;
  assign n42466 = n42436 & n42465 ;
  assign n42467 = ~n42464 & ~n42466 ;
  assign n42468 = n42462 & n42467 ;
  assign n42469 = ~n42145 & ~n42149 ;
  assign n42470 = n42145 & n42149 ;
  assign n42471 = n42173 & ~n42470 ;
  assign n42472 = ~n42469 & ~n42471 ;
  assign n42473 = ~n42468 & ~n42472 ;
  assign n42474 = n42468 & n42472 ;
  assign n42475 = ~n42473 & ~n42474 ;
  assign n42476 = ~n41922 & ~n42184 ;
  assign n42477 = ~n41924 & ~n42476 ;
  assign n42478 = n42475 & n42477 ;
  assign n42479 = ~n42475 & ~n42477 ;
  assign n42480 = ~n42478 & ~n42479 ;
  assign n42481 = ~n42189 & n42480 ;
  assign n42482 = ~n42196 & n42481 ;
  assign n42483 = ~n42189 & ~n42196 ;
  assign n42484 = ~n42480 & ~n42483 ;
  assign n42485 = ~n42482 & ~n42484 ;
  assign n42486 = n42462 & ~n42472 ;
  assign n42487 = n42467 & ~n42486 ;
  assign n42488 = n42430 & ~n42438 ;
  assign n42489 = \b[62]  & n9301 ;
  assign n42490 = n9298 & n42489 ;
  assign n42491 = ~\a[39]  & \b[63]  ;
  assign n42492 = n8751 & n42491 ;
  assign n42493 = \a[39]  & \b[63]  ;
  assign n42494 = n8748 & n42493 ;
  assign n42495 = ~n42492 & ~n42494 ;
  assign n42496 = ~n42490 & n42495 ;
  assign n42497 = ~\a[41]  & ~n42496 ;
  assign n42498 = n8759 & ~n22458 ;
  assign n42499 = ~\a[41]  & n42498 ;
  assign n42500 = ~n23173 & n42499 ;
  assign n42501 = ~n42497 & ~n42500 ;
  assign n42502 = ~n23173 & n42498 ;
  assign n42503 = \a[41]  & n42496 ;
  assign n42504 = ~n42502 & n42503 ;
  assign n42505 = n42501 & ~n42504 ;
  assign n42506 = n42435 & ~n42505 ;
  assign n42507 = ~n42488 & n42506 ;
  assign n42508 = n42435 & ~n42488 ;
  assign n42509 = n42505 & ~n42508 ;
  assign n42510 = ~n42507 & ~n42509 ;
  assign n42511 = n13125 & ~n16446 ;
  assign n42512 = ~n16444 & n42511 ;
  assign n42513 = \b[53]  & n13794 ;
  assign n42514 = n13792 & n42513 ;
  assign n42515 = ~\a[48]  & \b[54]  ;
  assign n42516 = n13117 & n42515 ;
  assign n42517 = ~n42514 & ~n42516 ;
  assign n42518 = \b[55]  & n13123 ;
  assign n42519 = \a[48]  & \b[54]  ;
  assign n42520 = n13786 & n42519 ;
  assign n42521 = \a[50]  & ~n42520 ;
  assign n42522 = ~n42518 & n42521 ;
  assign n42523 = n42517 & n42522 ;
  assign n42524 = ~n42512 & n42523 ;
  assign n42525 = ~n42518 & ~n42520 ;
  assign n42526 = n42517 & n42525 ;
  assign n42527 = ~n42512 & n42526 ;
  assign n42528 = ~\a[50]  & ~n42527 ;
  assign n42529 = ~n42524 & ~n42528 ;
  assign n42530 = ~n42325 & ~n42357 ;
  assign n42531 = ~n42324 & ~n42530 ;
  assign n42532 = ~n42297 & ~n42301 ;
  assign n42533 = ~n42298 & ~n42532 ;
  assign n42534 = ~n42287 & ~n42291 ;
  assign n42535 = \b[43]  & n20519 ;
  assign n42536 = \a[60]  & \b[42]  ;
  assign n42537 = n20510 & n42536 ;
  assign n42538 = ~n42535 & ~n42537 ;
  assign n42539 = \b[41]  & n21315 ;
  assign n42540 = n21312 & n42539 ;
  assign n42541 = ~\a[60]  & \b[42]  ;
  assign n42542 = n20513 & n42541 ;
  assign n42543 = ~n42540 & ~n42542 ;
  assign n42544 = n42538 & n42543 ;
  assign n42545 = n42245 & n42251 ;
  assign n42546 = ~n42247 & ~n42545 ;
  assign n42547 = \b[40]  & n21958 ;
  assign n42548 = \b[39]  & n21957 ;
  assign n42549 = ~n42547 & ~n42548 ;
  assign n42550 = ~n42546 & ~n42549 ;
  assign n42551 = ~n42247 & n42549 ;
  assign n42552 = ~n42545 & n42551 ;
  assign n42553 = ~\a[62]  & ~n42552 ;
  assign n42554 = ~n42550 & n42553 ;
  assign n42555 = ~n42544 & n42554 ;
  assign n42556 = ~n10406 & n20521 ;
  assign n42557 = ~n9929 & n20521 ;
  assign n42558 = ~n10402 & n42557 ;
  assign n42559 = ~n42556 & ~n42558 ;
  assign n42560 = ~n10409 & n42554 ;
  assign n42561 = ~n42559 & n42560 ;
  assign n42562 = ~n42555 & ~n42561 ;
  assign n42563 = ~n10409 & ~n42559 ;
  assign n42564 = \a[62]  & ~n42552 ;
  assign n42565 = ~n42550 & n42564 ;
  assign n42566 = n42544 & n42565 ;
  assign n42567 = ~n42563 & n42566 ;
  assign n42568 = n42562 & ~n42567 ;
  assign n42569 = ~\a[62]  & ~n42544 ;
  assign n42570 = ~\a[62]  & ~n10409 ;
  assign n42571 = ~n42559 & n42570 ;
  assign n42572 = ~n42569 & ~n42571 ;
  assign n42573 = ~n42550 & ~n42552 ;
  assign n42574 = \a[62]  & n42544 ;
  assign n42575 = ~n42563 & n42574 ;
  assign n42576 = ~n42573 & ~n42575 ;
  assign n42577 = n42572 & n42576 ;
  assign n42578 = n42568 & ~n42577 ;
  assign n42579 = ~n42256 & n42283 ;
  assign n42580 = ~n42258 & ~n42579 ;
  assign n42581 = n42578 & n42580 ;
  assign n42582 = ~n42578 & ~n42580 ;
  assign n42583 = ~n42581 & ~n42582 ;
  assign n42584 = n11906 & n18516 ;
  assign n42585 = ~n11903 & n42584 ;
  assign n42586 = n13483 & n18516 ;
  assign n42587 = ~n11902 & n42586 ;
  assign n42588 = \b[46]  & n18514 ;
  assign n42589 = \a[56]  & \b[45]  ;
  assign n42590 = n19181 & n42589 ;
  assign n42591 = ~\a[57]  & \b[45]  ;
  assign n42592 = n18508 & n42591 ;
  assign n42593 = ~n42590 & ~n42592 ;
  assign n42594 = ~n42588 & n42593 ;
  assign n42595 = \b[44]  & n19183 ;
  assign n42596 = n19180 & n42595 ;
  assign n42597 = \a[59]  & ~n42596 ;
  assign n42598 = n42594 & n42597 ;
  assign n42599 = ~n42587 & n42598 ;
  assign n42600 = ~n42585 & n42599 ;
  assign n42601 = n42594 & ~n42596 ;
  assign n42602 = ~n42587 & n42601 ;
  assign n42603 = ~n42585 & n42602 ;
  assign n42604 = ~\a[59]  & ~n42603 ;
  assign n42605 = ~n42600 & ~n42604 ;
  assign n42606 = n42583 & ~n42605 ;
  assign n42607 = ~n42583 & n42605 ;
  assign n42608 = ~n42606 & ~n42607 ;
  assign n42609 = n42534 & ~n42608 ;
  assign n42610 = ~n42534 & n42608 ;
  assign n42611 = ~n42609 & ~n42610 ;
  assign n42612 = ~n13524 & n37945 ;
  assign n42613 = ~n13522 & n42612 ;
  assign n42614 = \b[47]  & n17308 ;
  assign n42615 = n17305 & n42614 ;
  assign n42616 = ~\a[54]  & \b[48]  ;
  assign n42617 = n16647 & n42616 ;
  assign n42618 = ~n42615 & ~n42617 ;
  assign n42619 = \b[49]  & n16653 ;
  assign n42620 = \a[54]  & \b[48]  ;
  assign n42621 = n16644 & n42620 ;
  assign n42622 = \a[56]  & ~n42621 ;
  assign n42623 = ~n42619 & n42622 ;
  assign n42624 = n42618 & n42623 ;
  assign n42625 = ~n42613 & n42624 ;
  assign n42626 = ~n42619 & ~n42621 ;
  assign n42627 = n42618 & n42626 ;
  assign n42628 = ~n42613 & n42627 ;
  assign n42629 = ~\a[56]  & ~n42628 ;
  assign n42630 = ~n42625 & ~n42629 ;
  assign n42631 = ~n42611 & n42630 ;
  assign n42632 = n42611 & ~n42630 ;
  assign n42633 = ~n42631 & ~n42632 ;
  assign n42634 = ~n42533 & ~n42633 ;
  assign n42635 = n42533 & n42633 ;
  assign n42636 = ~n42634 & ~n42635 ;
  assign n42637 = ~n14276 & ~n15201 ;
  assign n42638 = ~n14790 & n42637 ;
  assign n42639 = n15198 & n42638 ;
  assign n42640 = ~n14276 & n15201 ;
  assign n42641 = ~n14790 & n42640 ;
  assign n42642 = ~n15198 & n42641 ;
  assign n42643 = ~n42639 & ~n42642 ;
  assign n42644 = \b[50]  & n15517 ;
  assign n42645 = n15514 & n42644 ;
  assign n42646 = ~\a[51]  & \b[51]  ;
  assign n42647 = n14785 & n42646 ;
  assign n42648 = ~n42645 & ~n42647 ;
  assign n42649 = \b[52]  & n14791 ;
  assign n42650 = \a[51]  & \b[51]  ;
  assign n42651 = n14782 & n42650 ;
  assign n42652 = \a[53]  & ~n42651 ;
  assign n42653 = ~n42649 & n42652 ;
  assign n42654 = n42648 & n42653 ;
  assign n42655 = n42643 & n42654 ;
  assign n42656 = ~n42649 & ~n42651 ;
  assign n42657 = n42648 & n42656 ;
  assign n42658 = n42643 & n42657 ;
  assign n42659 = ~\a[53]  & ~n42658 ;
  assign n42660 = ~n42655 & ~n42659 ;
  assign n42661 = n42636 & n42660 ;
  assign n42662 = ~n42636 & ~n42660 ;
  assign n42663 = ~n42661 & ~n42662 ;
  assign n42664 = n42531 & ~n42663 ;
  assign n42665 = ~n42531 & n42663 ;
  assign n42666 = ~n42664 & ~n42665 ;
  assign n42667 = n42529 & n42666 ;
  assign n42668 = ~n42529 & ~n42666 ;
  assign n42669 = ~n42667 & ~n42668 ;
  assign n42670 = n42362 & ~n42372 ;
  assign n42671 = n42367 & ~n42670 ;
  assign n42672 = n11572 & ~n19543 ;
  assign n42673 = ~n38598 & n42672 ;
  assign n42674 = \b[56]  & n12159 ;
  assign n42675 = n12156 & n42674 ;
  assign n42676 = ~\a[45]  & \b[57]  ;
  assign n42677 = n11564 & n42676 ;
  assign n42678 = ~n42675 & ~n42677 ;
  assign n42679 = \b[58]  & n11570 ;
  assign n42680 = \a[45]  & \b[57]  ;
  assign n42681 = n11561 & n42680 ;
  assign n42682 = \a[47]  & ~n42681 ;
  assign n42683 = ~n42679 & n42682 ;
  assign n42684 = n42678 & n42683 ;
  assign n42685 = ~n42673 & n42684 ;
  assign n42686 = ~n42679 & ~n42681 ;
  assign n42687 = n42678 & n42686 ;
  assign n42688 = ~n42673 & n42687 ;
  assign n42689 = ~\a[47]  & ~n42688 ;
  assign n42690 = ~n42685 & ~n42689 ;
  assign n42691 = ~n42671 & ~n42690 ;
  assign n42692 = ~n42669 & n42691 ;
  assign n42693 = n42671 & ~n42690 ;
  assign n42694 = n42669 & n42693 ;
  assign n42695 = ~n42692 & ~n42694 ;
  assign n42696 = n42671 & n42690 ;
  assign n42697 = ~n42669 & n42696 ;
  assign n42698 = ~n42671 & n42690 ;
  assign n42699 = n42669 & n42698 ;
  assign n42700 = ~n42697 & ~n42699 ;
  assign n42701 = n42695 & n42700 ;
  assign n42702 = n42396 & n42404 ;
  assign n42703 = n42401 & ~n42702 ;
  assign n42704 = n10082 & ~n20971 ;
  assign n42705 = ~n20969 & n42704 ;
  assign n42706 = \b[61]  & n10080 ;
  assign n42707 = \a[41]  & \b[60]  ;
  assign n42708 = n10679 & n42707 ;
  assign n42709 = ~\a[42]  & \b[60]  ;
  assign n42710 = n10074 & n42709 ;
  assign n42711 = ~n42708 & ~n42710 ;
  assign n42712 = ~n42706 & n42711 ;
  assign n42713 = \b[59]  & n10681 ;
  assign n42714 = n10678 & n42713 ;
  assign n42715 = \a[44]  & ~n42714 ;
  assign n42716 = n42712 & n42715 ;
  assign n42717 = ~n42705 & n42716 ;
  assign n42718 = n42712 & ~n42714 ;
  assign n42719 = ~n42705 & n42718 ;
  assign n42720 = ~\a[44]  & ~n42719 ;
  assign n42721 = ~n42717 & ~n42720 ;
  assign n42722 = n42703 & ~n42721 ;
  assign n42723 = ~n42701 & n42722 ;
  assign n42724 = ~n42703 & ~n42721 ;
  assign n42725 = n42701 & n42724 ;
  assign n42726 = ~n42723 & ~n42725 ;
  assign n42727 = ~n42703 & n42721 ;
  assign n42728 = ~n42701 & n42727 ;
  assign n42729 = n42703 & n42721 ;
  assign n42730 = n42701 & n42729 ;
  assign n42731 = ~n42728 & ~n42730 ;
  assign n42732 = n42726 & n42731 ;
  assign n42733 = n42510 & n42732 ;
  assign n42734 = ~n42510 & ~n42732 ;
  assign n42735 = ~n42733 & ~n42734 ;
  assign n42736 = ~n42487 & ~n42735 ;
  assign n42737 = n42487 & n42735 ;
  assign n42738 = ~n42736 & ~n42737 ;
  assign n42739 = n42478 & n42738 ;
  assign n42740 = n42481 & n42738 ;
  assign n42741 = ~n42196 & n42740 ;
  assign n42742 = ~n42739 & ~n42741 ;
  assign n42743 = ~n42478 & ~n42738 ;
  assign n42744 = ~n42482 & n42743 ;
  assign n42745 = n42742 & ~n42744 ;
  assign n42746 = ~n42737 & ~n42739 ;
  assign n42747 = ~n42741 & n42746 ;
  assign n42748 = ~n42507 & ~n42732 ;
  assign n42749 = ~n42509 & ~n42748 ;
  assign n42750 = n42701 & n42703 ;
  assign n42751 = n42721 & ~n42750 ;
  assign n42752 = ~n42701 & ~n42703 ;
  assign n42753 = ~n8756 & n39033 ;
  assign n42754 = ~n23171 & n42753 ;
  assign n42755 = ~n8272 & n42754 ;
  assign n42756 = \a[38]  & \a[40]  ;
  assign n42757 = \a[39]  & ~\a[41]  ;
  assign n42758 = n42756 & n42757 ;
  assign n42759 = ~\a[38]  & ~\a[40]  ;
  assign n42760 = ~\a[39]  & \a[41]  ;
  assign n42761 = n42759 & n42760 ;
  assign n42762 = ~n42758 & ~n42761 ;
  assign n42763 = \b[63]  & ~n42762 ;
  assign n42764 = \a[41]  & ~n42763 ;
  assign n42765 = ~n42755 & n42764 ;
  assign n42766 = ~\a[41]  & n42763 ;
  assign n42767 = ~\a[41]  & ~n8272 ;
  assign n42768 = n42754 & n42767 ;
  assign n42769 = ~n42766 & ~n42768 ;
  assign n42770 = ~n42765 & n42769 ;
  assign n42771 = ~n42752 & ~n42770 ;
  assign n42772 = ~n42751 & n42771 ;
  assign n42773 = ~n42751 & ~n42752 ;
  assign n42774 = n42770 & ~n42773 ;
  assign n42775 = ~n42772 & ~n42774 ;
  assign n42776 = n14793 & ~n15246 ;
  assign n42777 = ~n15244 & n42776 ;
  assign n42778 = \b[51]  & n15517 ;
  assign n42779 = n15514 & n42778 ;
  assign n42780 = ~\a[51]  & \b[52]  ;
  assign n42781 = n14785 & n42780 ;
  assign n42782 = ~n42779 & ~n42781 ;
  assign n42783 = \b[53]  & n14791 ;
  assign n42784 = \a[51]  & \b[52]  ;
  assign n42785 = n14782 & n42784 ;
  assign n42786 = \a[53]  & ~n42785 ;
  assign n42787 = ~n42783 & n42786 ;
  assign n42788 = n42782 & n42787 ;
  assign n42789 = ~n42777 & n42788 ;
  assign n42790 = ~n42783 & ~n42785 ;
  assign n42791 = n42782 & n42790 ;
  assign n42792 = ~n42777 & n42791 ;
  assign n42793 = ~\a[53]  & ~n42792 ;
  assign n42794 = ~n42789 & ~n42793 ;
  assign n42795 = ~n12435 & n18516 ;
  assign n42796 = ~n11905 & n18516 ;
  assign n42797 = ~n12431 & n42796 ;
  assign n42798 = ~n42795 & ~n42797 ;
  assign n42799 = ~n12438 & ~n42798 ;
  assign n42800 = \b[47]  & n18514 ;
  assign n42801 = \a[56]  & \b[46]  ;
  assign n42802 = n19181 & n42801 ;
  assign n42803 = ~\a[57]  & \b[46]  ;
  assign n42804 = n18508 & n42803 ;
  assign n42805 = ~n42802 & ~n42804 ;
  assign n42806 = ~n42800 & n42805 ;
  assign n42807 = \b[45]  & n19183 ;
  assign n42808 = n19180 & n42807 ;
  assign n42809 = \a[59]  & ~n42808 ;
  assign n42810 = n42806 & n42809 ;
  assign n42811 = ~n42799 & n42810 ;
  assign n42812 = n42806 & ~n42808 ;
  assign n42813 = ~\a[59]  & ~n42812 ;
  assign n42814 = ~\a[59]  & ~n12438 ;
  assign n42815 = ~n42798 & n42814 ;
  assign n42816 = ~n42813 & ~n42815 ;
  assign n42817 = ~n42811 & n42816 ;
  assign n42818 = ~n42552 & n42568 ;
  assign n42819 = \b[41]  & n21958 ;
  assign n42820 = \b[40]  & n21957 ;
  assign n42821 = ~n42819 & ~n42820 ;
  assign n42822 = n42549 & ~n42821 ;
  assign n42823 = ~n42549 & n42821 ;
  assign n42824 = ~n42822 & ~n42823 ;
  assign n42825 = ~n42818 & n42824 ;
  assign n42826 = ~n10889 & ~n19861 ;
  assign n42827 = ~n20518 & n42826 ;
  assign n42828 = n10886 & n42827 ;
  assign n42829 = n10889 & ~n19861 ;
  assign n42830 = ~n20518 & n42829 ;
  assign n42831 = ~n10886 & n42830 ;
  assign n42832 = ~n42828 & ~n42831 ;
  assign n42833 = \b[42]  & n21315 ;
  assign n42834 = n21312 & n42833 ;
  assign n42835 = ~\a[60]  & \b[43]  ;
  assign n42836 = n20513 & n42835 ;
  assign n42837 = ~n42834 & ~n42836 ;
  assign n42838 = \b[44]  & n20519 ;
  assign n42839 = \a[60]  & \b[43]  ;
  assign n42840 = n20510 & n42839 ;
  assign n42841 = \a[62]  & ~n42840 ;
  assign n42842 = ~n42838 & n42841 ;
  assign n42843 = n42837 & n42842 ;
  assign n42844 = n42832 & n42843 ;
  assign n42845 = ~n42838 & ~n42840 ;
  assign n42846 = n42837 & n42845 ;
  assign n42847 = n42832 & n42846 ;
  assign n42848 = ~\a[62]  & ~n42847 ;
  assign n42849 = ~n42844 & ~n42848 ;
  assign n42850 = ~n42552 & ~n42824 ;
  assign n42851 = n42568 & n42850 ;
  assign n42852 = ~n42849 & ~n42851 ;
  assign n42853 = ~n42825 & n42852 ;
  assign n42854 = ~n42825 & ~n42851 ;
  assign n42855 = n42849 & ~n42854 ;
  assign n42856 = ~n42853 & ~n42855 ;
  assign n42857 = ~n42581 & n42605 ;
  assign n42858 = ~n42582 & ~n42857 ;
  assign n42859 = ~n42856 & ~n42858 ;
  assign n42860 = n42817 & n42859 ;
  assign n42861 = n42856 & ~n42858 ;
  assign n42862 = ~n42817 & n42861 ;
  assign n42863 = ~n42860 & ~n42862 ;
  assign n42864 = ~n42817 & ~n42856 ;
  assign n42865 = n42858 & n42864 ;
  assign n42866 = n42856 & n42858 ;
  assign n42867 = n42817 & n42866 ;
  assign n42868 = ~n42865 & ~n42867 ;
  assign n42869 = n42863 & n42868 ;
  assign n42870 = n14052 & n16655 ;
  assign n42871 = ~n14049 & n42870 ;
  assign n42872 = n15779 & n37945 ;
  assign n42873 = ~n14048 & n42872 ;
  assign n42874 = \b[48]  & n17308 ;
  assign n42875 = n17305 & n42874 ;
  assign n42876 = ~\a[54]  & \b[49]  ;
  assign n42877 = n16647 & n42876 ;
  assign n42878 = ~n42875 & ~n42877 ;
  assign n42879 = \b[50]  & n16653 ;
  assign n42880 = \a[54]  & \b[49]  ;
  assign n42881 = n16644 & n42880 ;
  assign n42882 = \a[56]  & ~n42881 ;
  assign n42883 = ~n42879 & n42882 ;
  assign n42884 = n42878 & n42883 ;
  assign n42885 = ~n42873 & n42884 ;
  assign n42886 = ~n42871 & n42885 ;
  assign n42887 = ~n42879 & ~n42881 ;
  assign n42888 = n42878 & n42887 ;
  assign n42889 = ~n42873 & n42888 ;
  assign n42890 = ~n42871 & n42889 ;
  assign n42891 = ~\a[56]  & ~n42890 ;
  assign n42892 = ~n42886 & ~n42891 ;
  assign n42893 = ~n42869 & n42892 ;
  assign n42894 = n42869 & ~n42892 ;
  assign n42895 = ~n42893 & ~n42894 ;
  assign n42896 = ~n42610 & n42630 ;
  assign n42897 = ~n42609 & ~n42896 ;
  assign n42898 = n42895 & n42897 ;
  assign n42899 = ~n42895 & ~n42897 ;
  assign n42900 = ~n42898 & ~n42899 ;
  assign n42901 = n42794 & n42900 ;
  assign n42902 = ~n42794 & ~n42900 ;
  assign n42903 = ~n42901 & ~n42902 ;
  assign n42904 = ~n12606 & ~n16441 ;
  assign n42905 = ~n17647 & n42904 ;
  assign n42906 = ~n17643 & n42905 ;
  assign n42907 = ~n13122 & n42906 ;
  assign n42908 = n13125 & n17647 ;
  assign n42909 = ~n17644 & n42908 ;
  assign n42910 = ~n42907 & ~n42909 ;
  assign n42911 = \b[54]  & n13794 ;
  assign n42912 = n13792 & n42911 ;
  assign n42913 = ~\a[48]  & \b[55]  ;
  assign n42914 = n13117 & n42913 ;
  assign n42915 = ~n42912 & ~n42914 ;
  assign n42916 = \b[56]  & n13123 ;
  assign n42917 = \a[48]  & \b[55]  ;
  assign n42918 = n13786 & n42917 ;
  assign n42919 = \a[50]  & ~n42918 ;
  assign n42920 = ~n42916 & n42919 ;
  assign n42921 = n42915 & n42920 ;
  assign n42922 = n42910 & n42921 ;
  assign n42923 = ~n42916 & ~n42918 ;
  assign n42924 = n42915 & n42923 ;
  assign n42925 = n42910 & n42924 ;
  assign n42926 = ~\a[50]  & ~n42925 ;
  assign n42927 = ~n42922 & ~n42926 ;
  assign n42928 = ~n42635 & n42660 ;
  assign n42929 = ~n42634 & ~n42928 ;
  assign n42930 = ~n42927 & ~n42929 ;
  assign n42931 = ~n42903 & n42930 ;
  assign n42932 = ~n42927 & n42929 ;
  assign n42933 = n42903 & n42932 ;
  assign n42934 = ~n42931 & ~n42933 ;
  assign n42935 = n42927 & ~n42929 ;
  assign n42936 = n42903 & n42935 ;
  assign n42937 = n42927 & n42929 ;
  assign n42938 = ~n42903 & n42937 ;
  assign n42939 = ~n42936 & ~n42938 ;
  assign n42940 = n42934 & n42939 ;
  assign n42941 = n42529 & ~n42664 ;
  assign n42942 = ~n42665 & ~n42941 ;
  assign n42943 = n11572 & ~n19550 ;
  assign n42944 = ~n19548 & n42943 ;
  assign n42945 = \b[57]  & n12159 ;
  assign n42946 = n12156 & n42945 ;
  assign n42947 = ~\a[45]  & \b[58]  ;
  assign n42948 = n11564 & n42947 ;
  assign n42949 = ~n42946 & ~n42948 ;
  assign n42950 = \b[59]  & n11570 ;
  assign n42951 = \a[45]  & \b[58]  ;
  assign n42952 = n11561 & n42951 ;
  assign n42953 = \a[47]  & ~n42952 ;
  assign n42954 = ~n42950 & n42953 ;
  assign n42955 = n42949 & n42954 ;
  assign n42956 = ~n42944 & n42955 ;
  assign n42957 = ~n42950 & ~n42952 ;
  assign n42958 = n42949 & n42957 ;
  assign n42959 = ~n42944 & n42958 ;
  assign n42960 = ~\a[47]  & ~n42959 ;
  assign n42961 = ~n42956 & ~n42960 ;
  assign n42962 = n42942 & ~n42961 ;
  assign n42963 = ~n42940 & n42962 ;
  assign n42964 = ~n42942 & ~n42961 ;
  assign n42965 = n42940 & n42964 ;
  assign n42966 = ~n42963 & ~n42965 ;
  assign n42967 = ~n42942 & n42961 ;
  assign n42968 = ~n42940 & n42967 ;
  assign n42969 = n42942 & n42961 ;
  assign n42970 = n42940 & n42969 ;
  assign n42971 = ~n42968 & ~n42970 ;
  assign n42972 = n42966 & n42971 ;
  assign n42973 = n42669 & ~n42671 ;
  assign n42974 = ~n42669 & n42671 ;
  assign n42975 = n42690 & ~n42974 ;
  assign n42976 = ~n42973 & ~n42975 ;
  assign n42977 = ~n42972 & ~n42976 ;
  assign n42978 = n42972 & n42976 ;
  assign n42979 = ~n42977 & ~n42978 ;
  assign n42980 = n10082 & n21696 ;
  assign n42981 = ~n21693 & n42980 ;
  assign n42982 = n10082 & n41213 ;
  assign n42983 = ~n21692 & n42982 ;
  assign n42984 = \b[60]  & n10681 ;
  assign n42985 = n10678 & n42984 ;
  assign n42986 = \b[62]  & n10080 ;
  assign n42987 = \a[41]  & \b[61]  ;
  assign n42988 = n10679 & n42987 ;
  assign n42989 = ~\a[42]  & \b[61]  ;
  assign n42990 = n10074 & n42989 ;
  assign n42991 = ~n42988 & ~n42990 ;
  assign n42992 = ~n42986 & n42991 ;
  assign n42993 = ~n42985 & n42992 ;
  assign n42994 = ~n42983 & n42993 ;
  assign n42995 = ~n42981 & n42994 ;
  assign n42996 = ~\a[44]  & ~n42995 ;
  assign n42997 = \a[44]  & n42993 ;
  assign n42998 = ~n42983 & n42997 ;
  assign n42999 = ~n42981 & n42998 ;
  assign n43000 = ~n42996 & ~n42999 ;
  assign n43001 = ~n42979 & n43000 ;
  assign n43002 = n42979 & ~n43000 ;
  assign n43003 = ~n43001 & ~n43002 ;
  assign n43004 = n42775 & n43003 ;
  assign n43005 = ~n42775 & ~n43003 ;
  assign n43006 = ~n43004 & ~n43005 ;
  assign n43007 = n42749 & n43006 ;
  assign n43008 = ~n42749 & ~n43006 ;
  assign n43009 = ~n43007 & ~n43008 ;
  assign n43010 = n42747 & n43009 ;
  assign n43011 = ~n42747 & ~n43009 ;
  assign n43012 = ~n43010 & ~n43011 ;
  assign n43013 = ~n42737 & ~n43007 ;
  assign n43014 = ~n42739 & n43013 ;
  assign n43015 = ~n42741 & n43014 ;
  assign n43016 = n13125 & ~n17690 ;
  assign n43017 = ~n17688 & n43016 ;
  assign n43018 = \b[57]  & n13123 ;
  assign n43019 = \a[48]  & \b[56]  ;
  assign n43020 = n13786 & n43019 ;
  assign n43021 = ~n43018 & ~n43020 ;
  assign n43022 = \b[55]  & n13794 ;
  assign n43023 = n13792 & n43022 ;
  assign n43024 = ~\a[48]  & \b[56]  ;
  assign n43025 = n13117 & n43024 ;
  assign n43026 = ~n43023 & ~n43025 ;
  assign n43027 = n43021 & n43026 ;
  assign n43028 = ~n43017 & n43027 ;
  assign n43029 = ~\a[50]  & ~n43028 ;
  assign n43030 = \a[50]  & n43027 ;
  assign n43031 = ~n43017 & n43030 ;
  assign n43032 = ~n43029 & ~n43031 ;
  assign n43033 = n42794 & ~n42898 ;
  assign n43034 = ~n42899 & ~n43033 ;
  assign n43035 = ~n14098 & n37945 ;
  assign n43036 = ~n14096 & n43035 ;
  assign n43037 = \b[49]  & n17308 ;
  assign n43038 = n17305 & n43037 ;
  assign n43039 = ~\a[54]  & \b[50]  ;
  assign n43040 = n16647 & n43039 ;
  assign n43041 = ~n43038 & ~n43040 ;
  assign n43042 = \b[51]  & n16653 ;
  assign n43043 = \a[54]  & \b[50]  ;
  assign n43044 = n16644 & n43043 ;
  assign n43045 = \a[56]  & ~n43044 ;
  assign n43046 = ~n43042 & n43045 ;
  assign n43047 = n43041 & n43046 ;
  assign n43048 = ~n43036 & n43047 ;
  assign n43049 = ~n43042 & ~n43044 ;
  assign n43050 = n43041 & n43049 ;
  assign n43051 = ~n43036 & n43050 ;
  assign n43052 = ~\a[56]  & ~n43051 ;
  assign n43053 = ~n43048 & ~n43052 ;
  assign n43054 = ~n42817 & n42856 ;
  assign n43055 = ~n42858 & n43054 ;
  assign n43056 = n42817 & ~n42856 ;
  assign n43057 = ~n42858 & n43056 ;
  assign n43058 = ~n43055 & ~n43057 ;
  assign n43059 = n42868 & n42892 ;
  assign n43060 = n43058 & ~n43059 ;
  assign n43061 = n43053 & ~n43060 ;
  assign n43062 = ~n43053 & n43060 ;
  assign n43063 = ~n43061 & ~n43062 ;
  assign n43064 = n14793 & n38142 ;
  assign n43065 = ~n16404 & n43064 ;
  assign n43066 = n14793 & n16398 ;
  assign n43067 = n15241 & n43066 ;
  assign n43068 = n16400 & n43066 ;
  assign n43069 = ~n15239 & n43068 ;
  assign n43070 = ~n43067 & ~n43069 ;
  assign n43071 = ~n43065 & n43070 ;
  assign n43072 = \b[52]  & n15517 ;
  assign n43073 = n15514 & n43072 ;
  assign n43074 = ~\a[51]  & \b[53]  ;
  assign n43075 = n14785 & n43074 ;
  assign n43076 = ~n43073 & ~n43075 ;
  assign n43077 = \b[54]  & n14791 ;
  assign n43078 = \a[51]  & \b[53]  ;
  assign n43079 = n14782 & n43078 ;
  assign n43080 = \a[53]  & ~n43079 ;
  assign n43081 = ~n43077 & n43080 ;
  assign n43082 = n43076 & n43081 ;
  assign n43083 = n43071 & n43082 ;
  assign n43084 = ~n43077 & ~n43079 ;
  assign n43085 = n43076 & n43084 ;
  assign n43086 = n43071 & n43085 ;
  assign n43087 = ~\a[53]  & ~n43086 ;
  assign n43088 = ~n43083 & ~n43087 ;
  assign n43089 = n42825 & n42849 ;
  assign n43090 = n42849 & n42851 ;
  assign n43091 = ~n43089 & ~n43090 ;
  assign n43092 = n42817 & ~n42853 ;
  assign n43093 = n43091 & ~n43092 ;
  assign n43094 = ~n42552 & ~n42822 ;
  assign n43095 = n42568 & n43094 ;
  assign n43096 = ~n42823 & ~n43095 ;
  assign n43097 = \b[45]  & n20519 ;
  assign n43098 = \a[60]  & \b[44]  ;
  assign n43099 = n20510 & n43098 ;
  assign n43100 = ~n43097 & ~n43099 ;
  assign n43101 = \b[43]  & n21315 ;
  assign n43102 = n21312 & n43101 ;
  assign n43103 = ~\a[60]  & \b[44]  ;
  assign n43104 = n20513 & n43103 ;
  assign n43105 = ~n43102 & ~n43104 ;
  assign n43106 = n43100 & n43105 ;
  assign n43107 = ~\a[41]  & n42548 ;
  assign n43108 = ~\a[41]  & \b[40]  ;
  assign n43109 = n21958 & n43108 ;
  assign n43110 = ~n43107 & ~n43109 ;
  assign n43111 = \a[41]  & ~n42548 ;
  assign n43112 = ~n42547 & n43111 ;
  assign n43113 = n43110 & ~n43112 ;
  assign n43114 = \b[42]  & n21958 ;
  assign n43115 = \b[41]  & n21957 ;
  assign n43116 = ~n43114 & ~n43115 ;
  assign n43117 = ~\a[62]  & ~n43116 ;
  assign n43118 = ~n43113 & n43117 ;
  assign n43119 = ~\a[62]  & n43116 ;
  assign n43120 = n43113 & n43119 ;
  assign n43121 = ~n43118 & ~n43120 ;
  assign n43122 = ~n43106 & ~n43121 ;
  assign n43123 = ~n11394 & n20521 ;
  assign n43124 = ~n10888 & n20521 ;
  assign n43125 = ~n10892 & n43124 ;
  assign n43126 = ~n43123 & ~n43125 ;
  assign n43127 = ~n11397 & ~n43121 ;
  assign n43128 = ~n43126 & n43127 ;
  assign n43129 = ~n43122 & ~n43128 ;
  assign n43130 = ~n11397 & ~n43126 ;
  assign n43131 = \a[62]  & ~n43116 ;
  assign n43132 = ~n43113 & n43131 ;
  assign n43133 = \a[62]  & n43116 ;
  assign n43134 = n43113 & n43133 ;
  assign n43135 = ~n43132 & ~n43134 ;
  assign n43136 = n43106 & ~n43135 ;
  assign n43137 = ~n43130 & n43136 ;
  assign n43138 = n43129 & ~n43137 ;
  assign n43139 = ~\a[62]  & ~n43106 ;
  assign n43140 = ~\a[62]  & ~n11397 ;
  assign n43141 = ~n43126 & n43140 ;
  assign n43142 = ~n43139 & ~n43141 ;
  assign n43143 = ~n43113 & ~n43116 ;
  assign n43144 = n43113 & n43116 ;
  assign n43145 = ~n43143 & ~n43144 ;
  assign n43146 = \a[62]  & n43106 ;
  assign n43147 = ~n43130 & n43146 ;
  assign n43148 = n43145 & ~n43147 ;
  assign n43149 = n43142 & n43148 ;
  assign n43150 = n43138 & ~n43149 ;
  assign n43151 = ~n43096 & ~n43150 ;
  assign n43152 = n43096 & n43138 ;
  assign n43153 = ~n43149 & n43152 ;
  assign n43154 = ~n43151 & ~n43153 ;
  assign n43155 = ~n12478 & ~n17912 ;
  assign n43156 = ~n18513 & n43155 ;
  assign n43157 = n12475 & n43156 ;
  assign n43158 = n12478 & ~n17912 ;
  assign n43159 = ~n18513 & n43158 ;
  assign n43160 = ~n12475 & n43159 ;
  assign n43161 = ~n43157 & ~n43160 ;
  assign n43162 = \b[46]  & n19183 ;
  assign n43163 = n19180 & n43162 ;
  assign n43164 = \b[48]  & n18514 ;
  assign n43165 = \a[56]  & \b[47]  ;
  assign n43166 = n19181 & n43165 ;
  assign n43167 = ~\a[57]  & \b[47]  ;
  assign n43168 = n18508 & n43167 ;
  assign n43169 = ~n43166 & ~n43168 ;
  assign n43170 = ~n43164 & n43169 ;
  assign n43171 = ~n43163 & n43170 ;
  assign n43172 = n43161 & n43171 ;
  assign n43173 = ~\a[59]  & ~n43172 ;
  assign n43174 = \a[59]  & n43171 ;
  assign n43175 = n43161 & n43174 ;
  assign n43176 = ~n43173 & ~n43175 ;
  assign n43177 = n43154 & ~n43176 ;
  assign n43178 = ~n43154 & n43176 ;
  assign n43179 = ~n43177 & ~n43178 ;
  assign n43180 = n43093 & n43179 ;
  assign n43181 = ~n43093 & ~n43179 ;
  assign n43182 = ~n43180 & ~n43181 ;
  assign n43183 = n43088 & ~n43182 ;
  assign n43184 = ~n43063 & n43183 ;
  assign n43185 = n43088 & n43182 ;
  assign n43186 = n43063 & n43185 ;
  assign n43187 = ~n43184 & ~n43186 ;
  assign n43188 = ~n43088 & n43182 ;
  assign n43189 = ~n43063 & n43188 ;
  assign n43190 = ~n43088 & ~n43182 ;
  assign n43191 = n43063 & n43190 ;
  assign n43192 = ~n43189 & ~n43191 ;
  assign n43193 = n43187 & n43192 ;
  assign n43194 = n43034 & n43193 ;
  assign n43195 = ~n43034 & ~n43193 ;
  assign n43196 = ~n43194 & ~n43195 ;
  assign n43197 = n43032 & ~n43196 ;
  assign n43198 = ~n43032 & n43196 ;
  assign n43199 = ~n43197 & ~n43198 ;
  assign n43200 = ~n42903 & n42929 ;
  assign n43201 = n42934 & ~n43200 ;
  assign n43202 = ~n10988 & ~n19545 ;
  assign n43203 = ~n20260 & n43202 ;
  assign n43204 = ~n20256 & n43203 ;
  assign n43205 = ~n11569 & n43204 ;
  assign n43206 = n11572 & n20260 ;
  assign n43207 = ~n20257 & n43206 ;
  assign n43208 = ~n43205 & ~n43207 ;
  assign n43209 = \b[58]  & n12159 ;
  assign n43210 = n12156 & n43209 ;
  assign n43211 = ~\a[45]  & \b[59]  ;
  assign n43212 = n11564 & n43211 ;
  assign n43213 = ~n43210 & ~n43212 ;
  assign n43214 = \b[60]  & n11570 ;
  assign n43215 = \a[45]  & \b[59]  ;
  assign n43216 = n11561 & n43215 ;
  assign n43217 = \a[47]  & ~n43216 ;
  assign n43218 = ~n43214 & n43217 ;
  assign n43219 = n43213 & n43218 ;
  assign n43220 = n43208 & n43219 ;
  assign n43221 = ~n43214 & ~n43216 ;
  assign n43222 = n43213 & n43221 ;
  assign n43223 = n43208 & n43222 ;
  assign n43224 = ~\a[47]  & ~n43223 ;
  assign n43225 = ~n43220 & ~n43224 ;
  assign n43226 = ~n43201 & ~n43225 ;
  assign n43227 = ~n43199 & n43226 ;
  assign n43228 = n43201 & ~n43225 ;
  assign n43229 = n43199 & n43228 ;
  assign n43230 = ~n43227 & ~n43229 ;
  assign n43231 = n43201 & n43225 ;
  assign n43232 = ~n43199 & n43231 ;
  assign n43233 = ~n43201 & n43225 ;
  assign n43234 = n43199 & n43233 ;
  assign n43235 = ~n43232 & ~n43234 ;
  assign n43236 = n43230 & n43235 ;
  assign n43237 = ~n42940 & ~n42942 ;
  assign n43238 = n42940 & n42942 ;
  assign n43239 = n42961 & ~n43238 ;
  assign n43240 = ~n43237 & ~n43239 ;
  assign n43241 = n10082 & ~n22461 ;
  assign n43242 = ~n22459 & n43241 ;
  assign n43243 = \b[61]  & n10681 ;
  assign n43244 = n10678 & n43243 ;
  assign n43245 = \b[63]  & n10080 ;
  assign n43246 = \a[41]  & \b[62]  ;
  assign n43247 = n10679 & n43246 ;
  assign n43248 = ~\a[42]  & \b[62]  ;
  assign n43249 = n10074 & n43248 ;
  assign n43250 = ~n43247 & ~n43249 ;
  assign n43251 = ~n43245 & n43250 ;
  assign n43252 = ~n43244 & n43251 ;
  assign n43253 = ~\a[44]  & n43252 ;
  assign n43254 = ~n43242 & n43253 ;
  assign n43255 = ~n43242 & n43252 ;
  assign n43256 = \a[44]  & ~n43255 ;
  assign n43257 = ~n43254 & ~n43256 ;
  assign n43258 = ~n43240 & n43257 ;
  assign n43259 = n43236 & n43258 ;
  assign n43260 = n43240 & n43257 ;
  assign n43261 = ~n43236 & n43260 ;
  assign n43262 = ~n43259 & ~n43261 ;
  assign n43263 = ~n43240 & ~n43257 ;
  assign n43264 = ~n43236 & n43263 ;
  assign n43265 = n43240 & ~n43257 ;
  assign n43266 = n43236 & n43265 ;
  assign n43267 = ~n43264 & ~n43266 ;
  assign n43268 = n43262 & n43267 ;
  assign n43269 = ~n42978 & n43000 ;
  assign n43270 = ~n42977 & ~n43269 ;
  assign n43271 = ~n43268 & ~n43270 ;
  assign n43272 = n43268 & n43270 ;
  assign n43273 = ~n43271 & ~n43272 ;
  assign n43274 = ~n42772 & ~n43003 ;
  assign n43275 = ~n42774 & ~n43274 ;
  assign n43276 = n43273 & n43275 ;
  assign n43277 = ~n43273 & ~n43275 ;
  assign n43278 = ~n43276 & ~n43277 ;
  assign n43279 = ~n43008 & n43278 ;
  assign n43280 = ~n43015 & n43279 ;
  assign n43281 = ~n43008 & ~n43015 ;
  assign n43282 = ~n43278 & ~n43281 ;
  assign n43283 = ~n43280 & ~n43282 ;
  assign n43284 = n43262 & ~n43270 ;
  assign n43285 = n43267 & ~n43284 ;
  assign n43286 = n43230 & ~n43240 ;
  assign n43287 = n10082 & ~n22458 ;
  assign n43288 = ~n23173 & n43287 ;
  assign n43289 = \b[62]  & n10681 ;
  assign n43290 = n10678 & n43289 ;
  assign n43291 = \a[41]  & \b[63]  ;
  assign n43292 = n10679 & n43291 ;
  assign n43293 = ~\a[42]  & \b[63]  ;
  assign n43294 = n10074 & n43293 ;
  assign n43295 = ~n43292 & ~n43294 ;
  assign n43296 = ~n43290 & n43295 ;
  assign n43297 = ~\a[44]  & n43296 ;
  assign n43298 = ~n43288 & n43297 ;
  assign n43299 = ~n43288 & n43296 ;
  assign n43300 = \a[44]  & ~n43299 ;
  assign n43301 = ~n43298 & ~n43300 ;
  assign n43302 = n43235 & n43301 ;
  assign n43303 = ~n43286 & n43302 ;
  assign n43304 = n43235 & ~n43286 ;
  assign n43305 = ~n43301 & ~n43304 ;
  assign n43306 = ~n43303 & ~n43305 ;
  assign n43307 = n11572 & ~n20971 ;
  assign n43308 = ~n20969 & n43307 ;
  assign n43309 = \b[59]  & n12159 ;
  assign n43310 = n12156 & n43309 ;
  assign n43311 = ~\a[45]  & \b[60]  ;
  assign n43312 = n11564 & n43311 ;
  assign n43313 = ~n43310 & ~n43312 ;
  assign n43314 = \b[61]  & n11570 ;
  assign n43315 = \a[45]  & \b[60]  ;
  assign n43316 = n11561 & n43315 ;
  assign n43317 = \a[47]  & ~n43316 ;
  assign n43318 = ~n43314 & n43317 ;
  assign n43319 = n43313 & n43318 ;
  assign n43320 = ~n43308 & n43319 ;
  assign n43321 = ~n43314 & ~n43316 ;
  assign n43322 = n43313 & n43321 ;
  assign n43323 = ~n43308 & n43322 ;
  assign n43324 = ~\a[47]  & ~n43323 ;
  assign n43325 = ~n43320 & ~n43324 ;
  assign n43326 = ~n43198 & n43201 ;
  assign n43327 = ~n43197 & ~n43326 ;
  assign n43328 = n43053 & ~n43182 ;
  assign n43329 = ~n43060 & ~n43182 ;
  assign n43330 = ~n43061 & ~n43329 ;
  assign n43331 = ~n43328 & n43330 ;
  assign n43332 = ~n43093 & ~n43177 ;
  assign n43333 = ~n43178 & ~n43332 ;
  assign n43334 = ~n43096 & n43138 ;
  assign n43335 = n43106 & ~n43130 ;
  assign n43336 = \a[62]  & n43145 ;
  assign n43337 = ~n43335 & n43336 ;
  assign n43338 = ~\a[62]  & n43145 ;
  assign n43339 = n43335 & n43338 ;
  assign n43340 = ~n43337 & ~n43339 ;
  assign n43341 = ~n43334 & n43340 ;
  assign n43342 = n11906 & n20521 ;
  assign n43343 = ~n11903 & n43342 ;
  assign n43344 = n13483 & n20521 ;
  assign n43345 = ~n11902 & n43344 ;
  assign n43346 = \b[46]  & n20519 ;
  assign n43347 = \a[60]  & \b[45]  ;
  assign n43348 = n20510 & n43347 ;
  assign n43349 = ~n43346 & ~n43348 ;
  assign n43350 = \b[44]  & n21315 ;
  assign n43351 = n21312 & n43350 ;
  assign n43352 = ~\a[60]  & \b[45]  ;
  assign n43353 = n20513 & n43352 ;
  assign n43354 = ~n43351 & ~n43353 ;
  assign n43355 = n43349 & n43354 ;
  assign n43356 = ~n43345 & n43355 ;
  assign n43357 = ~n43343 & n43356 ;
  assign n43358 = n43110 & n43116 ;
  assign n43359 = ~n43112 & ~n43358 ;
  assign n43360 = \b[43]  & n21958 ;
  assign n43361 = \b[42]  & n21957 ;
  assign n43362 = ~n43360 & ~n43361 ;
  assign n43363 = ~n43359 & ~n43362 ;
  assign n43364 = ~n43112 & n43362 ;
  assign n43365 = ~n43358 & n43364 ;
  assign n43366 = ~\a[62]  & ~n43365 ;
  assign n43367 = ~n43363 & n43366 ;
  assign n43368 = ~n43357 & n43367 ;
  assign n43369 = \a[62]  & ~n43365 ;
  assign n43370 = ~n43363 & n43369 ;
  assign n43371 = n43355 & n43370 ;
  assign n43372 = ~n43345 & n43371 ;
  assign n43373 = ~n43343 & n43372 ;
  assign n43374 = ~n43368 & ~n43373 ;
  assign n43375 = ~\a[62]  & ~n43357 ;
  assign n43376 = ~n43363 & ~n43365 ;
  assign n43377 = \a[62]  & n43355 ;
  assign n43378 = ~n43345 & n43377 ;
  assign n43379 = ~n43343 & n43378 ;
  assign n43380 = ~n43376 & ~n43379 ;
  assign n43381 = ~n43375 & n43380 ;
  assign n43382 = n43374 & ~n43381 ;
  assign n43383 = n43341 & n43382 ;
  assign n43384 = ~n43341 & ~n43382 ;
  assign n43385 = ~n43383 & ~n43384 ;
  assign n43386 = ~n13521 & n18516 ;
  assign n43387 = ~n12477 & n18516 ;
  assign n43388 = ~n13517 & n43387 ;
  assign n43389 = ~n43386 & ~n43388 ;
  assign n43390 = ~n13524 & ~n43389 ;
  assign n43391 = \b[49]  & n18514 ;
  assign n43392 = \a[56]  & \b[48]  ;
  assign n43393 = n19181 & n43392 ;
  assign n43394 = ~\a[57]  & \b[48]  ;
  assign n43395 = n18508 & n43394 ;
  assign n43396 = ~n43393 & ~n43395 ;
  assign n43397 = ~n43391 & n43396 ;
  assign n43398 = \b[47]  & n19183 ;
  assign n43399 = n19180 & n43398 ;
  assign n43400 = \a[59]  & ~n43399 ;
  assign n43401 = n43397 & n43400 ;
  assign n43402 = ~n43390 & n43401 ;
  assign n43403 = n43397 & ~n43399 ;
  assign n43404 = ~\a[59]  & ~n43403 ;
  assign n43405 = ~\a[59]  & ~n13524 ;
  assign n43406 = ~n43389 & n43405 ;
  assign n43407 = ~n43404 & ~n43406 ;
  assign n43408 = ~n43402 & n43407 ;
  assign n43409 = n43385 & ~n43408 ;
  assign n43410 = ~n43385 & n43408 ;
  assign n43411 = ~n43409 & ~n43410 ;
  assign n43412 = ~n43333 & ~n43411 ;
  assign n43413 = n43333 & n43411 ;
  assign n43414 = ~n43412 & ~n43413 ;
  assign n43415 = ~n15201 & ~n16016 ;
  assign n43416 = ~n16652 & n43415 ;
  assign n43417 = n15198 & n43416 ;
  assign n43418 = n15201 & ~n16016 ;
  assign n43419 = ~n16652 & n43418 ;
  assign n43420 = ~n15198 & n43419 ;
  assign n43421 = ~n43417 & ~n43420 ;
  assign n43422 = \b[50]  & n17308 ;
  assign n43423 = n17305 & n43422 ;
  assign n43424 = ~\a[54]  & \b[51]  ;
  assign n43425 = n16647 & n43424 ;
  assign n43426 = ~n43423 & ~n43425 ;
  assign n43427 = \b[52]  & n16653 ;
  assign n43428 = \a[54]  & \b[51]  ;
  assign n43429 = n16644 & n43428 ;
  assign n43430 = \a[56]  & ~n43429 ;
  assign n43431 = ~n43427 & n43430 ;
  assign n43432 = n43426 & n43431 ;
  assign n43433 = n43421 & n43432 ;
  assign n43434 = ~n43427 & ~n43429 ;
  assign n43435 = n43426 & n43434 ;
  assign n43436 = n43421 & n43435 ;
  assign n43437 = ~\a[56]  & ~n43436 ;
  assign n43438 = ~n43433 & ~n43437 ;
  assign n43439 = ~n43414 & n43438 ;
  assign n43440 = n43414 & ~n43438 ;
  assign n43441 = ~n43439 & ~n43440 ;
  assign n43442 = ~n43331 & ~n43441 ;
  assign n43443 = n43331 & n43441 ;
  assign n43444 = ~n43442 & ~n43443 ;
  assign n43445 = n14793 & ~n16446 ;
  assign n43446 = ~n16444 & n43445 ;
  assign n43447 = \b[53]  & n15517 ;
  assign n43448 = n15514 & n43447 ;
  assign n43449 = ~\a[51]  & \b[54]  ;
  assign n43450 = n14785 & n43449 ;
  assign n43451 = ~n43448 & ~n43450 ;
  assign n43452 = \b[55]  & n14791 ;
  assign n43453 = \a[51]  & \b[54]  ;
  assign n43454 = n14782 & n43453 ;
  assign n43455 = \a[53]  & ~n43454 ;
  assign n43456 = ~n43452 & n43455 ;
  assign n43457 = n43451 & n43456 ;
  assign n43458 = ~n43446 & n43457 ;
  assign n43459 = ~n43452 & ~n43454 ;
  assign n43460 = n43451 & n43459 ;
  assign n43461 = ~n43446 & n43460 ;
  assign n43462 = ~\a[53]  & ~n43461 ;
  assign n43463 = ~n43458 & ~n43462 ;
  assign n43464 = n43444 & ~n43463 ;
  assign n43465 = ~n43444 & n43463 ;
  assign n43466 = ~n43464 & ~n43465 ;
  assign n43467 = n13125 & ~n19543 ;
  assign n43468 = ~n38598 & n43467 ;
  assign n43469 = \b[56]  & n13794 ;
  assign n43470 = n13792 & n43469 ;
  assign n43471 = ~\a[48]  & \b[57]  ;
  assign n43472 = n13117 & n43471 ;
  assign n43473 = ~n43470 & ~n43472 ;
  assign n43474 = \b[58]  & n13123 ;
  assign n43475 = \a[48]  & \b[57]  ;
  assign n43476 = n13786 & n43475 ;
  assign n43477 = \a[50]  & ~n43476 ;
  assign n43478 = ~n43474 & n43477 ;
  assign n43479 = n43473 & n43478 ;
  assign n43480 = ~n43468 & n43479 ;
  assign n43481 = ~n43474 & ~n43476 ;
  assign n43482 = n43473 & n43481 ;
  assign n43483 = ~n43468 & n43482 ;
  assign n43484 = ~\a[50]  & ~n43483 ;
  assign n43485 = ~n43480 & ~n43484 ;
  assign n43486 = ~n43034 & n43192 ;
  assign n43487 = n43187 & ~n43486 ;
  assign n43488 = n43485 & ~n43487 ;
  assign n43489 = ~n43466 & n43488 ;
  assign n43490 = n43485 & n43487 ;
  assign n43491 = n43466 & n43490 ;
  assign n43492 = ~n43489 & ~n43491 ;
  assign n43493 = ~n43485 & n43487 ;
  assign n43494 = ~n43466 & n43493 ;
  assign n43495 = ~n43485 & ~n43487 ;
  assign n43496 = n43466 & n43495 ;
  assign n43497 = ~n43494 & ~n43496 ;
  assign n43498 = n43492 & n43497 ;
  assign n43499 = n43327 & n43498 ;
  assign n43500 = ~n43327 & ~n43498 ;
  assign n43501 = ~n43499 & ~n43500 ;
  assign n43502 = n43325 & n43501 ;
  assign n43503 = ~n43325 & ~n43501 ;
  assign n43504 = ~n43502 & ~n43503 ;
  assign n43505 = n43306 & ~n43504 ;
  assign n43506 = ~n43306 & n43504 ;
  assign n43507 = ~n43505 & ~n43506 ;
  assign n43508 = ~n43285 & ~n43507 ;
  assign n43509 = n43285 & n43507 ;
  assign n43510 = ~n43508 & ~n43509 ;
  assign n43511 = n43276 & n43510 ;
  assign n43512 = n43279 & n43510 ;
  assign n43513 = ~n43015 & n43512 ;
  assign n43514 = ~n43511 & ~n43513 ;
  assign n43515 = ~n43276 & ~n43510 ;
  assign n43516 = ~n43280 & n43515 ;
  assign n43517 = n43514 & ~n43516 ;
  assign n43518 = ~n43509 & ~n43511 ;
  assign n43519 = ~n43513 & n43518 ;
  assign n43520 = n43325 & ~n43499 ;
  assign n43521 = ~n10079 & n39033 ;
  assign n43522 = ~n23171 & n43521 ;
  assign n43523 = ~n9646 & n43522 ;
  assign n43524 = \a[41]  & \a[43]  ;
  assign n43525 = \a[42]  & ~\a[44]  ;
  assign n43526 = n43524 & n43525 ;
  assign n43527 = ~\a[41]  & ~\a[43]  ;
  assign n43528 = ~\a[42]  & \a[44]  ;
  assign n43529 = n43527 & n43528 ;
  assign n43530 = ~n43526 & ~n43529 ;
  assign n43531 = \b[63]  & ~n43530 ;
  assign n43532 = \a[44]  & ~n43531 ;
  assign n43533 = ~n43523 & n43532 ;
  assign n43534 = ~\a[44]  & n43531 ;
  assign n43535 = ~\a[44]  & ~n9646 ;
  assign n43536 = n43522 & n43535 ;
  assign n43537 = ~n43534 & ~n43536 ;
  assign n43538 = ~n43533 & n43537 ;
  assign n43539 = ~n43500 & ~n43538 ;
  assign n43540 = ~n43520 & n43539 ;
  assign n43541 = n43500 & n43538 ;
  assign n43542 = n43325 & n43538 ;
  assign n43543 = ~n43499 & n43542 ;
  assign n43544 = ~n43541 & ~n43543 ;
  assign n43545 = ~n43540 & n43544 ;
  assign n43546 = n14793 & n17647 ;
  assign n43547 = ~n17644 & n43546 ;
  assign n43548 = n14793 & n19567 ;
  assign n43549 = ~n17643 & n43548 ;
  assign n43550 = \b[54]  & n15517 ;
  assign n43551 = n15514 & n43550 ;
  assign n43552 = ~\a[51]  & \b[55]  ;
  assign n43553 = n14785 & n43552 ;
  assign n43554 = ~n43551 & ~n43553 ;
  assign n43555 = \b[56]  & n14791 ;
  assign n43556 = \a[51]  & \b[55]  ;
  assign n43557 = n14782 & n43556 ;
  assign n43558 = \a[53]  & ~n43557 ;
  assign n43559 = ~n43555 & n43558 ;
  assign n43560 = n43554 & n43559 ;
  assign n43561 = ~n43549 & n43560 ;
  assign n43562 = ~n43547 & n43561 ;
  assign n43563 = ~n43555 & ~n43557 ;
  assign n43564 = n43554 & n43563 ;
  assign n43565 = ~n43549 & n43564 ;
  assign n43566 = ~n43547 & n43565 ;
  assign n43567 = ~\a[53]  & ~n43566 ;
  assign n43568 = ~n43562 & ~n43567 ;
  assign n43569 = ~n15246 & n37945 ;
  assign n43570 = ~n15244 & n43569 ;
  assign n43571 = \b[51]  & n17308 ;
  assign n43572 = n17305 & n43571 ;
  assign n43573 = ~\a[54]  & \b[52]  ;
  assign n43574 = n16647 & n43573 ;
  assign n43575 = ~n43572 & ~n43574 ;
  assign n43576 = \b[53]  & n16653 ;
  assign n43577 = \a[54]  & \b[52]  ;
  assign n43578 = n16644 & n43577 ;
  assign n43579 = \a[56]  & ~n43578 ;
  assign n43580 = ~n43576 & n43579 ;
  assign n43581 = n43575 & n43580 ;
  assign n43582 = ~n43570 & n43581 ;
  assign n43583 = ~n43576 & ~n43578 ;
  assign n43584 = n43575 & n43583 ;
  assign n43585 = ~n43570 & n43584 ;
  assign n43586 = ~\a[56]  & ~n43585 ;
  assign n43587 = ~n43582 & ~n43586 ;
  assign n43588 = n14052 & n18516 ;
  assign n43589 = ~n14049 & n43588 ;
  assign n43590 = n15779 & n18516 ;
  assign n43591 = ~n14048 & n43590 ;
  assign n43592 = \b[50]  & n18514 ;
  assign n43593 = \a[56]  & \b[49]  ;
  assign n43594 = n19181 & n43593 ;
  assign n43595 = ~\a[57]  & \b[49]  ;
  assign n43596 = n18508 & n43595 ;
  assign n43597 = ~n43594 & ~n43596 ;
  assign n43598 = ~n43592 & n43597 ;
  assign n43599 = \b[48]  & n19183 ;
  assign n43600 = n19180 & n43599 ;
  assign n43601 = \a[59]  & ~n43600 ;
  assign n43602 = n43598 & n43601 ;
  assign n43603 = ~n43591 & n43602 ;
  assign n43604 = ~n43589 & n43603 ;
  assign n43605 = n43598 & ~n43600 ;
  assign n43606 = ~n43591 & n43605 ;
  assign n43607 = ~n43589 & n43606 ;
  assign n43608 = ~\a[59]  & ~n43607 ;
  assign n43609 = ~n43604 & ~n43608 ;
  assign n43610 = \b[47]  & n20519 ;
  assign n43611 = \a[60]  & \b[46]  ;
  assign n43612 = n20510 & n43611 ;
  assign n43613 = ~n43610 & ~n43612 ;
  assign n43614 = \b[45]  & n21315 ;
  assign n43615 = n21312 & n43614 ;
  assign n43616 = ~\a[60]  & \b[46]  ;
  assign n43617 = n20513 & n43616 ;
  assign n43618 = ~n43615 & ~n43617 ;
  assign n43619 = n43613 & n43618 ;
  assign n43620 = ~\a[62]  & ~n43619 ;
  assign n43621 = ~n12435 & n20521 ;
  assign n43622 = ~n11905 & n20521 ;
  assign n43623 = ~n12431 & n43622 ;
  assign n43624 = ~n43621 & ~n43623 ;
  assign n43625 = ~\a[62]  & ~n12438 ;
  assign n43626 = ~n43624 & n43625 ;
  assign n43627 = ~n43620 & ~n43626 ;
  assign n43628 = \b[44]  & n21958 ;
  assign n43629 = \b[43]  & n21957 ;
  assign n43630 = ~n43628 & ~n43629 ;
  assign n43631 = n43362 & ~n43630 ;
  assign n43632 = ~n43362 & n43630 ;
  assign n43633 = ~n43631 & ~n43632 ;
  assign n43634 = ~n12438 & ~n43624 ;
  assign n43635 = \a[62]  & n43619 ;
  assign n43636 = ~n43634 & n43635 ;
  assign n43637 = ~n43633 & ~n43636 ;
  assign n43638 = n43627 & n43637 ;
  assign n43639 = ~n43365 & ~n43373 ;
  assign n43640 = ~n43368 & n43639 ;
  assign n43641 = ~\a[62]  & n43633 ;
  assign n43642 = ~n43619 & n43641 ;
  assign n43643 = ~n12438 & n43641 ;
  assign n43644 = ~n43624 & n43643 ;
  assign n43645 = ~n43642 & ~n43644 ;
  assign n43646 = \a[62]  & n43633 ;
  assign n43647 = n43619 & n43646 ;
  assign n43648 = ~n43634 & n43647 ;
  assign n43649 = n43645 & ~n43648 ;
  assign n43650 = ~n43640 & n43649 ;
  assign n43651 = ~n43638 & n43650 ;
  assign n43652 = n43640 & ~n43649 ;
  assign n43653 = n43627 & n43640 ;
  assign n43654 = n43637 & n43653 ;
  assign n43655 = ~n43652 & ~n43654 ;
  assign n43656 = ~n43651 & n43655 ;
  assign n43657 = n43609 & n43656 ;
  assign n43658 = ~n43609 & ~n43656 ;
  assign n43659 = ~n43657 & ~n43658 ;
  assign n43660 = ~n43383 & n43408 ;
  assign n43661 = ~n43384 & ~n43660 ;
  assign n43662 = ~n43659 & n43661 ;
  assign n43663 = n43659 & ~n43661 ;
  assign n43664 = ~n43662 & ~n43663 ;
  assign n43665 = n43587 & n43664 ;
  assign n43666 = ~n43587 & ~n43664 ;
  assign n43667 = ~n43665 & ~n43666 ;
  assign n43668 = ~n43413 & n43438 ;
  assign n43669 = ~n43412 & ~n43668 ;
  assign n43670 = ~n43667 & n43669 ;
  assign n43671 = n43667 & ~n43669 ;
  assign n43672 = ~n43670 & ~n43671 ;
  assign n43673 = ~n43568 & n43672 ;
  assign n43674 = n43568 & ~n43672 ;
  assign n43675 = ~n43673 & ~n43674 ;
  assign n43676 = ~n43443 & n43463 ;
  assign n43677 = ~n43442 & ~n43676 ;
  assign n43678 = n43675 & n43677 ;
  assign n43679 = ~n43675 & ~n43677 ;
  assign n43680 = ~n43678 & ~n43679 ;
  assign n43681 = n13125 & ~n19550 ;
  assign n43682 = ~n19548 & n43681 ;
  assign n43683 = \b[57]  & n13794 ;
  assign n43684 = n13792 & n43683 ;
  assign n43685 = ~\a[48]  & \b[58]  ;
  assign n43686 = n13117 & n43685 ;
  assign n43687 = ~n43684 & ~n43686 ;
  assign n43688 = \b[59]  & n13123 ;
  assign n43689 = \a[48]  & \b[58]  ;
  assign n43690 = n13786 & n43689 ;
  assign n43691 = \a[50]  & ~n43690 ;
  assign n43692 = ~n43688 & n43691 ;
  assign n43693 = n43687 & n43692 ;
  assign n43694 = ~n43682 & n43693 ;
  assign n43695 = ~n43688 & ~n43690 ;
  assign n43696 = n43687 & n43695 ;
  assign n43697 = ~n43682 & n43696 ;
  assign n43698 = ~\a[50]  & ~n43697 ;
  assign n43699 = ~n43694 & ~n43698 ;
  assign n43700 = n43680 & ~n43699 ;
  assign n43701 = ~n43680 & n43699 ;
  assign n43702 = ~n43700 & ~n43701 ;
  assign n43703 = ~n10988 & ~n20966 ;
  assign n43704 = ~n21696 & n43703 ;
  assign n43705 = ~n21692 & n43704 ;
  assign n43706 = ~n11569 & n43705 ;
  assign n43707 = n11572 & n21696 ;
  assign n43708 = ~n21693 & n43707 ;
  assign n43709 = ~n43706 & ~n43708 ;
  assign n43710 = \b[60]  & n12159 ;
  assign n43711 = n12156 & n43710 ;
  assign n43712 = ~\a[45]  & \b[61]  ;
  assign n43713 = n11564 & n43712 ;
  assign n43714 = ~n43711 & ~n43713 ;
  assign n43715 = \b[62]  & n11570 ;
  assign n43716 = \a[45]  & \b[61]  ;
  assign n43717 = n11561 & n43716 ;
  assign n43718 = \a[47]  & ~n43717 ;
  assign n43719 = ~n43715 & n43718 ;
  assign n43720 = n43714 & n43719 ;
  assign n43721 = n43709 & n43720 ;
  assign n43722 = ~n43715 & ~n43717 ;
  assign n43723 = n43714 & n43722 ;
  assign n43724 = n43709 & n43723 ;
  assign n43725 = ~\a[47]  & ~n43724 ;
  assign n43726 = ~n43721 & ~n43725 ;
  assign n43727 = n43466 & n43487 ;
  assign n43728 = n43497 & ~n43727 ;
  assign n43729 = n43726 & ~n43728 ;
  assign n43730 = ~n43702 & n43729 ;
  assign n43731 = n43726 & n43728 ;
  assign n43732 = n43702 & n43731 ;
  assign n43733 = ~n43730 & ~n43732 ;
  assign n43734 = ~n43726 & n43728 ;
  assign n43735 = ~n43702 & n43734 ;
  assign n43736 = ~n43726 & ~n43728 ;
  assign n43737 = n43702 & n43736 ;
  assign n43738 = ~n43735 & ~n43737 ;
  assign n43739 = n43733 & n43738 ;
  assign n43740 = n43545 & ~n43739 ;
  assign n43741 = ~n43545 & n43739 ;
  assign n43742 = ~n43740 & ~n43741 ;
  assign n43743 = ~n43303 & n43504 ;
  assign n43744 = ~n43305 & ~n43743 ;
  assign n43745 = n43742 & n43744 ;
  assign n43746 = ~n43742 & ~n43744 ;
  assign n43747 = ~n43745 & ~n43746 ;
  assign n43748 = n43519 & n43747 ;
  assign n43749 = ~n43519 & ~n43747 ;
  assign n43750 = ~n43748 & ~n43749 ;
  assign n43751 = ~n43509 & ~n43745 ;
  assign n43752 = ~n43511 & n43751 ;
  assign n43753 = ~n43513 & n43752 ;
  assign n43754 = ~n12606 & ~n19545 ;
  assign n43755 = ~n20260 & n43754 ;
  assign n43756 = ~n20256 & n43755 ;
  assign n43757 = ~n13122 & n43756 ;
  assign n43758 = n13125 & n20260 ;
  assign n43759 = ~n20257 & n43758 ;
  assign n43760 = ~n43757 & ~n43759 ;
  assign n43761 = \b[58]  & n13794 ;
  assign n43762 = n13792 & n43761 ;
  assign n43763 = ~\a[48]  & \b[59]  ;
  assign n43764 = n13117 & n43763 ;
  assign n43765 = ~n43762 & ~n43764 ;
  assign n43766 = \b[60]  & n13123 ;
  assign n43767 = \a[48]  & \b[59]  ;
  assign n43768 = n13786 & n43767 ;
  assign n43769 = \a[50]  & ~n43768 ;
  assign n43770 = ~n43766 & n43769 ;
  assign n43771 = n43765 & n43770 ;
  assign n43772 = n43760 & n43771 ;
  assign n43773 = ~n43766 & ~n43768 ;
  assign n43774 = n43765 & n43773 ;
  assign n43775 = n43760 & n43774 ;
  assign n43776 = ~\a[50]  & ~n43775 ;
  assign n43777 = ~n43772 & ~n43776 ;
  assign n43778 = n43587 & ~n43662 ;
  assign n43779 = ~n43663 & ~n43778 ;
  assign n43780 = ~n16404 & n38142 ;
  assign n43781 = n15241 & n16398 ;
  assign n43782 = n16398 & n16400 ;
  assign n43783 = ~n15239 & n43782 ;
  assign n43784 = ~n43781 & ~n43783 ;
  assign n43785 = ~n43780 & n43784 ;
  assign n43786 = n37945 & ~n43785 ;
  assign n43787 = \b[52]  & n17308 ;
  assign n43788 = n17305 & n43787 ;
  assign n43789 = ~\a[54]  & \b[53]  ;
  assign n43790 = n16647 & n43789 ;
  assign n43791 = ~n43788 & ~n43790 ;
  assign n43792 = \b[54]  & n16653 ;
  assign n43793 = \a[54]  & \b[53]  ;
  assign n43794 = n16644 & n43793 ;
  assign n43795 = \a[56]  & ~n43794 ;
  assign n43796 = ~n43792 & n43795 ;
  assign n43797 = n43791 & n43796 ;
  assign n43798 = ~n43786 & n43797 ;
  assign n43799 = ~n43792 & ~n43794 ;
  assign n43800 = n43791 & n43799 ;
  assign n43801 = ~n43786 & n43800 ;
  assign n43802 = ~\a[56]  & ~n43801 ;
  assign n43803 = ~n43798 & ~n43802 ;
  assign n43804 = n43609 & ~n43651 ;
  assign n43805 = n43655 & ~n43804 ;
  assign n43806 = ~n14098 & n18516 ;
  assign n43807 = ~n14096 & n43806 ;
  assign n43808 = \b[49]  & n19183 ;
  assign n43809 = n19180 & n43808 ;
  assign n43810 = \b[51]  & n18514 ;
  assign n43811 = \a[56]  & \b[50]  ;
  assign n43812 = n19181 & n43811 ;
  assign n43813 = ~\a[57]  & \b[50]  ;
  assign n43814 = n18508 & n43813 ;
  assign n43815 = ~n43812 & ~n43814 ;
  assign n43816 = ~n43810 & n43815 ;
  assign n43817 = ~n43809 & n43816 ;
  assign n43818 = ~\a[59]  & n43817 ;
  assign n43819 = ~n43807 & n43818 ;
  assign n43820 = ~n43807 & n43817 ;
  assign n43821 = \a[59]  & ~n43820 ;
  assign n43822 = ~n43819 & ~n43821 ;
  assign n43823 = ~n43631 & n43649 ;
  assign n43824 = ~\a[44]  & \b[44]  ;
  assign n43825 = n21957 & n43824 ;
  assign n43826 = ~\a[44]  & \b[45]  ;
  assign n43827 = n21958 & n43826 ;
  assign n43828 = ~n43825 & ~n43827 ;
  assign n43829 = \b[45]  & n21958 ;
  assign n43830 = \b[44]  & n21957 ;
  assign n43831 = \a[44]  & ~n43830 ;
  assign n43832 = ~n43829 & n43831 ;
  assign n43833 = n43828 & ~n43832 ;
  assign n43834 = ~n43362 & ~n43833 ;
  assign n43835 = n43362 & n43833 ;
  assign n43836 = ~n43834 & ~n43835 ;
  assign n43837 = ~n43823 & ~n43836 ;
  assign n43838 = ~n12478 & ~n19861 ;
  assign n43839 = ~n20518 & n43838 ;
  assign n43840 = n12475 & n43839 ;
  assign n43841 = n12478 & ~n19861 ;
  assign n43842 = ~n20518 & n43841 ;
  assign n43843 = ~n12475 & n43842 ;
  assign n43844 = ~n43840 & ~n43843 ;
  assign n43845 = \b[46]  & n21315 ;
  assign n43846 = n21312 & n43845 ;
  assign n43847 = ~\a[60]  & \b[47]  ;
  assign n43848 = n20513 & n43847 ;
  assign n43849 = ~n43846 & ~n43848 ;
  assign n43850 = \b[48]  & n20519 ;
  assign n43851 = \a[60]  & \b[47]  ;
  assign n43852 = n20510 & n43851 ;
  assign n43853 = \a[62]  & ~n43852 ;
  assign n43854 = ~n43850 & n43853 ;
  assign n43855 = n43849 & n43854 ;
  assign n43856 = n43844 & n43855 ;
  assign n43857 = ~n43850 & ~n43852 ;
  assign n43858 = n43849 & n43857 ;
  assign n43859 = n43844 & n43858 ;
  assign n43860 = ~\a[62]  & ~n43859 ;
  assign n43861 = ~n43856 & ~n43860 ;
  assign n43862 = ~n43631 & n43836 ;
  assign n43863 = n43649 & n43862 ;
  assign n43864 = ~n43861 & ~n43863 ;
  assign n43865 = ~n43837 & n43864 ;
  assign n43866 = ~n43837 & ~n43863 ;
  assign n43867 = n43861 & ~n43866 ;
  assign n43868 = ~n43865 & ~n43867 ;
  assign n43869 = n43822 & n43868 ;
  assign n43870 = ~n43822 & ~n43868 ;
  assign n43871 = ~n43869 & ~n43870 ;
  assign n43872 = n43805 & n43871 ;
  assign n43873 = ~n43805 & n43869 ;
  assign n43874 = ~n43805 & ~n43868 ;
  assign n43875 = ~n43822 & n43874 ;
  assign n43876 = ~n43873 & ~n43875 ;
  assign n43877 = ~n43872 & n43876 ;
  assign n43878 = n43803 & ~n43877 ;
  assign n43879 = ~n43803 & n43877 ;
  assign n43880 = ~n43878 & ~n43879 ;
  assign n43881 = n43779 & n43880 ;
  assign n43882 = ~n43779 & ~n43880 ;
  assign n43883 = ~n43881 & ~n43882 ;
  assign n43884 = n43568 & ~n43670 ;
  assign n43885 = ~n43670 & n43671 ;
  assign n43886 = ~n43884 & ~n43885 ;
  assign n43887 = n14793 & ~n17690 ;
  assign n43888 = ~n17688 & n43887 ;
  assign n43889 = \b[55]  & n15517 ;
  assign n43890 = n15514 & n43889 ;
  assign n43891 = ~\a[51]  & \b[56]  ;
  assign n43892 = n14785 & n43891 ;
  assign n43893 = ~n43890 & ~n43892 ;
  assign n43894 = \b[57]  & n14791 ;
  assign n43895 = \a[51]  & \b[56]  ;
  assign n43896 = n14782 & n43895 ;
  assign n43897 = \a[53]  & ~n43896 ;
  assign n43898 = ~n43894 & n43897 ;
  assign n43899 = n43893 & n43898 ;
  assign n43900 = ~n43888 & n43899 ;
  assign n43901 = ~n43894 & ~n43896 ;
  assign n43902 = n43893 & n43901 ;
  assign n43903 = ~n43888 & n43902 ;
  assign n43904 = ~\a[53]  & ~n43903 ;
  assign n43905 = ~n43900 & ~n43904 ;
  assign n43906 = n43886 & ~n43905 ;
  assign n43907 = ~n43883 & n43906 ;
  assign n43908 = n43886 & n43905 ;
  assign n43909 = n43883 & n43908 ;
  assign n43910 = ~n43907 & ~n43909 ;
  assign n43911 = ~n43886 & n43905 ;
  assign n43912 = ~n43883 & n43911 ;
  assign n43913 = ~n43886 & ~n43905 ;
  assign n43914 = n43883 & n43913 ;
  assign n43915 = ~n43912 & ~n43914 ;
  assign n43916 = n43910 & n43915 ;
  assign n43917 = n43777 & ~n43916 ;
  assign n43918 = ~n43777 & n43916 ;
  assign n43919 = ~n43917 & ~n43918 ;
  assign n43920 = ~n43678 & n43699 ;
  assign n43921 = ~n43679 & ~n43920 ;
  assign n43922 = n11572 & ~n22461 ;
  assign n43923 = ~n22459 & n43922 ;
  assign n43924 = \b[61]  & n12159 ;
  assign n43925 = n12156 & n43924 ;
  assign n43926 = ~\a[45]  & \b[62]  ;
  assign n43927 = n11564 & n43926 ;
  assign n43928 = ~n43925 & ~n43927 ;
  assign n43929 = \b[63]  & n11570 ;
  assign n43930 = \a[45]  & \b[62]  ;
  assign n43931 = n11561 & n43930 ;
  assign n43932 = \a[47]  & ~n43931 ;
  assign n43933 = ~n43929 & n43932 ;
  assign n43934 = n43928 & n43933 ;
  assign n43935 = ~n43923 & n43934 ;
  assign n43936 = ~n43929 & ~n43931 ;
  assign n43937 = n43928 & n43936 ;
  assign n43938 = ~n43923 & n43937 ;
  assign n43939 = ~\a[47]  & ~n43938 ;
  assign n43940 = ~n43935 & ~n43939 ;
  assign n43941 = ~n43921 & ~n43940 ;
  assign n43942 = n43919 & n43941 ;
  assign n43943 = n43921 & ~n43940 ;
  assign n43944 = ~n43919 & n43943 ;
  assign n43945 = ~n43942 & ~n43944 ;
  assign n43946 = ~n43921 & n43940 ;
  assign n43947 = ~n43919 & n43946 ;
  assign n43948 = n43921 & n43940 ;
  assign n43949 = n43919 & n43948 ;
  assign n43950 = ~n43947 & ~n43949 ;
  assign n43951 = n43945 & n43950 ;
  assign n43952 = ~n43702 & n43728 ;
  assign n43953 = n43702 & ~n43728 ;
  assign n43954 = n43726 & ~n43953 ;
  assign n43955 = ~n43952 & ~n43954 ;
  assign n43956 = ~n43951 & ~n43955 ;
  assign n43957 = n43951 & n43955 ;
  assign n43958 = ~n43956 & ~n43957 ;
  assign n43959 = ~n43540 & n43739 ;
  assign n43960 = n43544 & ~n43959 ;
  assign n43961 = n43958 & n43960 ;
  assign n43962 = ~n43958 & ~n43960 ;
  assign n43963 = ~n43961 & ~n43962 ;
  assign n43964 = ~n43746 & n43963 ;
  assign n43965 = ~n43753 & n43964 ;
  assign n43966 = ~n43746 & ~n43753 ;
  assign n43967 = ~n43963 & ~n43966 ;
  assign n43968 = ~n43965 & ~n43967 ;
  assign n43969 = n43945 & ~n43955 ;
  assign n43970 = n43950 & ~n43969 ;
  assign n43971 = ~n43918 & ~n43921 ;
  assign n43972 = \b[62]  & n12159 ;
  assign n43973 = n12156 & n43972 ;
  assign n43974 = ~\a[45]  & \b[63]  ;
  assign n43975 = n11564 & n43974 ;
  assign n43976 = \a[45]  & \b[63]  ;
  assign n43977 = n11561 & n43976 ;
  assign n43978 = ~n43975 & ~n43977 ;
  assign n43979 = ~n43973 & n43978 ;
  assign n43980 = ~\a[47]  & ~n43979 ;
  assign n43981 = n11572 & ~n22458 ;
  assign n43982 = ~\a[47]  & n43981 ;
  assign n43983 = ~n23173 & n43982 ;
  assign n43984 = ~n43980 & ~n43983 ;
  assign n43985 = ~n23173 & n43981 ;
  assign n43986 = \a[47]  & n43979 ;
  assign n43987 = ~n43985 & n43986 ;
  assign n43988 = n43984 & ~n43987 ;
  assign n43989 = ~n43917 & ~n43988 ;
  assign n43990 = ~n43971 & n43989 ;
  assign n43991 = n43917 & n43988 ;
  assign n43992 = ~n43921 & n43988 ;
  assign n43993 = ~n43918 & n43992 ;
  assign n43994 = ~n43991 & ~n43993 ;
  assign n43995 = ~n43990 & n43994 ;
  assign n43996 = n13125 & ~n20971 ;
  assign n43997 = ~n20969 & n43996 ;
  assign n43998 = \b[59]  & n13794 ;
  assign n43999 = n13792 & n43998 ;
  assign n44000 = ~\a[48]  & \b[60]  ;
  assign n44001 = n13117 & n44000 ;
  assign n44002 = ~n43999 & ~n44001 ;
  assign n44003 = \b[61]  & n13123 ;
  assign n44004 = \a[48]  & \b[60]  ;
  assign n44005 = n13786 & n44004 ;
  assign n44006 = \a[50]  & ~n44005 ;
  assign n44007 = ~n44003 & n44006 ;
  assign n44008 = n44002 & n44007 ;
  assign n44009 = ~n43997 & n44008 ;
  assign n44010 = ~n44003 & ~n44005 ;
  assign n44011 = n44002 & n44010 ;
  assign n44012 = ~n43997 & n44011 ;
  assign n44013 = ~\a[50]  & ~n44012 ;
  assign n44014 = ~n44009 & ~n44013 ;
  assign n44015 = ~n43883 & n43905 ;
  assign n44016 = n43883 & ~n43905 ;
  assign n44017 = ~n43886 & ~n44016 ;
  assign n44018 = ~n44015 & ~n44017 ;
  assign n44019 = n14793 & ~n19543 ;
  assign n44020 = ~n38598 & n44019 ;
  assign n44021 = \b[56]  & n15517 ;
  assign n44022 = n15514 & n44021 ;
  assign n44023 = ~\a[51]  & \b[57]  ;
  assign n44024 = n14785 & n44023 ;
  assign n44025 = ~n44022 & ~n44024 ;
  assign n44026 = \b[58]  & n14791 ;
  assign n44027 = \a[51]  & \b[57]  ;
  assign n44028 = n14782 & n44027 ;
  assign n44029 = \a[53]  & ~n44028 ;
  assign n44030 = ~n44026 & n44029 ;
  assign n44031 = n44025 & n44030 ;
  assign n44032 = ~n44020 & n44031 ;
  assign n44033 = ~n44026 & ~n44028 ;
  assign n44034 = n44025 & n44033 ;
  assign n44035 = ~n44020 & n44034 ;
  assign n44036 = ~\a[53]  & ~n44035 ;
  assign n44037 = ~n44032 & ~n44036 ;
  assign n44038 = ~n43779 & ~n43879 ;
  assign n44039 = ~n43878 & ~n44038 ;
  assign n44040 = ~n43869 & n43870 ;
  assign n44041 = ~n43805 & ~n43869 ;
  assign n44042 = ~n44040 & ~n44041 ;
  assign n44043 = ~n15201 & ~n17912 ;
  assign n44044 = ~n18513 & n44043 ;
  assign n44045 = n15198 & n44044 ;
  assign n44046 = n15201 & ~n17912 ;
  assign n44047 = ~n18513 & n44046 ;
  assign n44048 = ~n15198 & n44047 ;
  assign n44049 = ~n44045 & ~n44048 ;
  assign n44050 = \b[52]  & n18514 ;
  assign n44051 = \a[56]  & \b[51]  ;
  assign n44052 = n19181 & n44051 ;
  assign n44053 = ~\a[57]  & \b[51]  ;
  assign n44054 = n18508 & n44053 ;
  assign n44055 = ~n44052 & ~n44054 ;
  assign n44056 = ~n44050 & n44055 ;
  assign n44057 = \b[50]  & n19183 ;
  assign n44058 = n19180 & n44057 ;
  assign n44059 = \a[59]  & ~n44058 ;
  assign n44060 = n44056 & n44059 ;
  assign n44061 = n44049 & n44060 ;
  assign n44062 = n44056 & ~n44058 ;
  assign n44063 = n44049 & n44062 ;
  assign n44064 = ~\a[59]  & ~n44063 ;
  assign n44065 = ~n44061 & ~n44064 ;
  assign n44066 = ~n43837 & ~n43864 ;
  assign n44067 = \b[49]  & n20519 ;
  assign n44068 = \a[60]  & \b[48]  ;
  assign n44069 = n20510 & n44068 ;
  assign n44070 = ~n44067 & ~n44069 ;
  assign n44071 = \b[47]  & n21315 ;
  assign n44072 = n21312 & n44071 ;
  assign n44073 = ~\a[60]  & \b[48]  ;
  assign n44074 = n20513 & n44073 ;
  assign n44075 = ~n44072 & ~n44074 ;
  assign n44076 = n44070 & n44075 ;
  assign n44077 = ~\a[62]  & ~n44076 ;
  assign n44078 = ~n13521 & n20521 ;
  assign n44079 = ~n12477 & n20521 ;
  assign n44080 = ~n13517 & n44079 ;
  assign n44081 = ~n44078 & ~n44080 ;
  assign n44082 = ~\a[62]  & ~n13524 ;
  assign n44083 = ~n44081 & n44082 ;
  assign n44084 = ~n44077 & ~n44083 ;
  assign n44085 = ~n43362 & ~n43832 ;
  assign n44086 = \b[46]  & n21958 ;
  assign n44087 = \b[45]  & n21957 ;
  assign n44088 = ~n44086 & ~n44087 ;
  assign n44089 = n43828 & ~n44088 ;
  assign n44090 = ~n44085 & n44089 ;
  assign n44091 = n43828 & ~n44085 ;
  assign n44092 = n44088 & ~n44091 ;
  assign n44093 = ~n44090 & ~n44092 ;
  assign n44094 = \a[62]  & ~n44069 ;
  assign n44095 = ~n44067 & n44094 ;
  assign n44096 = n44075 & n44095 ;
  assign n44097 = ~n44093 & ~n44096 ;
  assign n44098 = ~n13524 & ~n44093 ;
  assign n44099 = ~n44081 & n44098 ;
  assign n44100 = ~n44097 & ~n44099 ;
  assign n44101 = n44084 & ~n44100 ;
  assign n44102 = ~n13524 & ~n44081 ;
  assign n44103 = \a[62]  & n44076 ;
  assign n44104 = ~n44102 & n44103 ;
  assign n44105 = n44084 & ~n44104 ;
  assign n44106 = n44093 & ~n44105 ;
  assign n44107 = ~n44101 & ~n44106 ;
  assign n44108 = ~n44066 & n44107 ;
  assign n44109 = n44066 & ~n44107 ;
  assign n44110 = ~n44108 & ~n44109 ;
  assign n44111 = n44065 & n44110 ;
  assign n44112 = ~n44065 & ~n44110 ;
  assign n44113 = ~n44111 & ~n44112 ;
  assign n44114 = n44042 & ~n44113 ;
  assign n44115 = ~n44042 & n44113 ;
  assign n44116 = ~n44114 & ~n44115 ;
  assign n44117 = ~n16446 & n37945 ;
  assign n44118 = ~n16444 & n44117 ;
  assign n44119 = \b[53]  & n17308 ;
  assign n44120 = n17305 & n44119 ;
  assign n44121 = ~\a[54]  & \b[54]  ;
  assign n44122 = n16647 & n44121 ;
  assign n44123 = ~n44120 & ~n44122 ;
  assign n44124 = \b[55]  & n16653 ;
  assign n44125 = \a[54]  & \b[54]  ;
  assign n44126 = n16644 & n44125 ;
  assign n44127 = \a[56]  & ~n44126 ;
  assign n44128 = ~n44124 & n44127 ;
  assign n44129 = n44123 & n44128 ;
  assign n44130 = ~n44118 & n44129 ;
  assign n44131 = ~n44124 & ~n44126 ;
  assign n44132 = n44123 & n44131 ;
  assign n44133 = ~n44118 & n44132 ;
  assign n44134 = ~\a[56]  & ~n44133 ;
  assign n44135 = ~n44130 & ~n44134 ;
  assign n44136 = n44116 & ~n44135 ;
  assign n44137 = ~n44116 & n44135 ;
  assign n44138 = ~n44136 & ~n44137 ;
  assign n44139 = n44039 & n44138 ;
  assign n44140 = ~n44039 & ~n44138 ;
  assign n44141 = ~n44139 & ~n44140 ;
  assign n44142 = n44037 & ~n44141 ;
  assign n44143 = ~n44037 & n44141 ;
  assign n44144 = ~n44142 & ~n44143 ;
  assign n44145 = n44018 & n44144 ;
  assign n44146 = ~n44018 & ~n44144 ;
  assign n44147 = ~n44145 & ~n44146 ;
  assign n44148 = n44014 & n44147 ;
  assign n44149 = ~n44014 & ~n44147 ;
  assign n44150 = ~n44148 & ~n44149 ;
  assign n44151 = n43995 & ~n44150 ;
  assign n44152 = ~n43995 & n44150 ;
  assign n44153 = ~n44151 & ~n44152 ;
  assign n44154 = ~n43970 & ~n44153 ;
  assign n44155 = n43970 & n44153 ;
  assign n44156 = ~n44154 & ~n44155 ;
  assign n44157 = n43961 & n44156 ;
  assign n44158 = ~n43746 & n44156 ;
  assign n44159 = n43963 & n44158 ;
  assign n44160 = ~n43753 & n44159 ;
  assign n44161 = ~n44157 & ~n44160 ;
  assign n44162 = ~n43961 & ~n44156 ;
  assign n44163 = ~n43965 & n44162 ;
  assign n44164 = n44161 & ~n44163 ;
  assign n44165 = n44014 & ~n44145 ;
  assign n44166 = \b[63]  & n11572 ;
  assign n44167 = ~n21694 & n44166 ;
  assign n44168 = ~n23171 & n44167 ;
  assign n44169 = \b[63]  & n12159 ;
  assign n44170 = n12156 & n44169 ;
  assign n44171 = \a[47]  & ~n44170 ;
  assign n44172 = ~n44168 & n44171 ;
  assign n44173 = ~n44168 & ~n44170 ;
  assign n44174 = ~\a[47]  & ~n44173 ;
  assign n44175 = ~n44172 & ~n44174 ;
  assign n44176 = ~n44146 & ~n44175 ;
  assign n44177 = ~n44165 & n44176 ;
  assign n44178 = n44146 & n44175 ;
  assign n44179 = n44014 & n44175 ;
  assign n44180 = ~n44145 & n44179 ;
  assign n44181 = ~n44178 & ~n44180 ;
  assign n44182 = ~n44177 & n44181 ;
  assign n44183 = n16655 & n17647 ;
  assign n44184 = ~n17644 & n44183 ;
  assign n44185 = n19567 & n37945 ;
  assign n44186 = ~n17643 & n44185 ;
  assign n44187 = \b[54]  & n17308 ;
  assign n44188 = n17305 & n44187 ;
  assign n44189 = ~\a[54]  & \b[55]  ;
  assign n44190 = n16647 & n44189 ;
  assign n44191 = ~n44188 & ~n44190 ;
  assign n44192 = \b[56]  & n16653 ;
  assign n44193 = \a[54]  & \b[55]  ;
  assign n44194 = n16644 & n44193 ;
  assign n44195 = \a[56]  & ~n44194 ;
  assign n44196 = ~n44192 & n44195 ;
  assign n44197 = n44191 & n44196 ;
  assign n44198 = ~n44186 & n44197 ;
  assign n44199 = ~n44184 & n44198 ;
  assign n44200 = ~n44192 & ~n44194 ;
  assign n44201 = n44191 & n44200 ;
  assign n44202 = ~n44186 & n44201 ;
  assign n44203 = ~n44184 & n44202 ;
  assign n44204 = ~\a[56]  & ~n44203 ;
  assign n44205 = ~n44199 & ~n44204 ;
  assign n44206 = n44065 & ~n44108 ;
  assign n44207 = ~n44109 & ~n44206 ;
  assign n44208 = ~n44092 & ~n44106 ;
  assign n44209 = \b[47]  & n21958 ;
  assign n44210 = \b[46]  & n21957 ;
  assign n44211 = ~n44209 & ~n44210 ;
  assign n44212 = n44088 & ~n44211 ;
  assign n44213 = ~n44088 & n44211 ;
  assign n44214 = ~n44212 & ~n44213 ;
  assign n44215 = ~n44208 & n44214 ;
  assign n44216 = n14052 & n20521 ;
  assign n44217 = ~n14049 & n44216 ;
  assign n44218 = n15779 & n20521 ;
  assign n44219 = ~n14048 & n44218 ;
  assign n44220 = \b[48]  & n21315 ;
  assign n44221 = n21312 & n44220 ;
  assign n44222 = ~\a[60]  & \b[49]  ;
  assign n44223 = n20513 & n44222 ;
  assign n44224 = ~n44221 & ~n44223 ;
  assign n44225 = \b[50]  & n20519 ;
  assign n44226 = \a[60]  & \b[49]  ;
  assign n44227 = n20510 & n44226 ;
  assign n44228 = \a[62]  & ~n44227 ;
  assign n44229 = ~n44225 & n44228 ;
  assign n44230 = n44224 & n44229 ;
  assign n44231 = ~n44219 & n44230 ;
  assign n44232 = ~n44217 & n44231 ;
  assign n44233 = ~n44225 & ~n44227 ;
  assign n44234 = n44224 & n44233 ;
  assign n44235 = ~n44219 & n44234 ;
  assign n44236 = ~n44217 & n44235 ;
  assign n44237 = ~\a[62]  & ~n44236 ;
  assign n44238 = ~n44232 & ~n44237 ;
  assign n44239 = ~n44090 & ~n44105 ;
  assign n44240 = ~n44092 & ~n44214 ;
  assign n44241 = ~n44239 & n44240 ;
  assign n44242 = ~n44238 & ~n44241 ;
  assign n44243 = ~n44215 & n44242 ;
  assign n44244 = ~n44214 & n44238 ;
  assign n44245 = n44208 & n44244 ;
  assign n44246 = n44214 & n44238 ;
  assign n44247 = ~n44208 & n44246 ;
  assign n44248 = ~n44245 & ~n44247 ;
  assign n44249 = ~n44243 & n44248 ;
  assign n44250 = ~n15246 & n18516 ;
  assign n44251 = ~n15244 & n44250 ;
  assign n44252 = \b[53]  & n18514 ;
  assign n44253 = \a[56]  & \b[52]  ;
  assign n44254 = n19181 & n44253 ;
  assign n44255 = ~\a[57]  & \b[52]  ;
  assign n44256 = n18508 & n44255 ;
  assign n44257 = ~n44254 & ~n44256 ;
  assign n44258 = ~n44252 & n44257 ;
  assign n44259 = \b[51]  & n19183 ;
  assign n44260 = n19180 & n44259 ;
  assign n44261 = \a[59]  & ~n44260 ;
  assign n44262 = n44258 & n44261 ;
  assign n44263 = ~n44251 & n44262 ;
  assign n44264 = n44258 & ~n44260 ;
  assign n44265 = ~n44251 & n44264 ;
  assign n44266 = ~\a[59]  & ~n44265 ;
  assign n44267 = ~n44263 & ~n44266 ;
  assign n44268 = ~n44249 & n44267 ;
  assign n44269 = ~n44207 & n44268 ;
  assign n44270 = ~n44249 & ~n44267 ;
  assign n44271 = n44207 & n44270 ;
  assign n44272 = ~n44269 & ~n44271 ;
  assign n44273 = n44249 & ~n44267 ;
  assign n44274 = ~n44207 & n44273 ;
  assign n44275 = n44249 & n44267 ;
  assign n44276 = n44207 & n44275 ;
  assign n44277 = ~n44274 & ~n44276 ;
  assign n44278 = n44272 & n44277 ;
  assign n44279 = n44205 & n44278 ;
  assign n44280 = ~n44205 & ~n44278 ;
  assign n44281 = ~n44279 & ~n44280 ;
  assign n44282 = ~n44114 & n44135 ;
  assign n44283 = ~n44115 & ~n44282 ;
  assign n44284 = ~n44281 & n44283 ;
  assign n44285 = n44281 & ~n44283 ;
  assign n44286 = ~n44284 & ~n44285 ;
  assign n44287 = n14793 & ~n19550 ;
  assign n44288 = ~n19548 & n44287 ;
  assign n44289 = \b[57]  & n15517 ;
  assign n44290 = n15514 & n44289 ;
  assign n44291 = ~\a[51]  & \b[58]  ;
  assign n44292 = n14785 & n44291 ;
  assign n44293 = ~n44290 & ~n44292 ;
  assign n44294 = \b[59]  & n14791 ;
  assign n44295 = \a[51]  & \b[58]  ;
  assign n44296 = n14782 & n44295 ;
  assign n44297 = \a[53]  & ~n44296 ;
  assign n44298 = ~n44294 & n44297 ;
  assign n44299 = n44293 & n44298 ;
  assign n44300 = ~n44288 & n44299 ;
  assign n44301 = ~n44294 & ~n44296 ;
  assign n44302 = n44293 & n44301 ;
  assign n44303 = ~n44288 & n44302 ;
  assign n44304 = ~\a[53]  & ~n44303 ;
  assign n44305 = ~n44300 & ~n44304 ;
  assign n44306 = n44286 & ~n44305 ;
  assign n44307 = ~n44286 & n44305 ;
  assign n44308 = ~n44306 & ~n44307 ;
  assign n44309 = ~n12606 & ~n20966 ;
  assign n44310 = ~n21696 & n44309 ;
  assign n44311 = ~n21692 & n44310 ;
  assign n44312 = ~n13122 & n44311 ;
  assign n44313 = n13125 & n21696 ;
  assign n44314 = ~n21693 & n44313 ;
  assign n44315 = ~n44312 & ~n44314 ;
  assign n44316 = \b[60]  & n13794 ;
  assign n44317 = n13792 & n44316 ;
  assign n44318 = ~\a[48]  & \b[61]  ;
  assign n44319 = n13117 & n44318 ;
  assign n44320 = ~n44317 & ~n44319 ;
  assign n44321 = \b[62]  & n13123 ;
  assign n44322 = \a[48]  & \b[61]  ;
  assign n44323 = n13786 & n44322 ;
  assign n44324 = \a[50]  & ~n44323 ;
  assign n44325 = ~n44321 & n44324 ;
  assign n44326 = n44320 & n44325 ;
  assign n44327 = n44315 & n44326 ;
  assign n44328 = ~n44321 & ~n44323 ;
  assign n44329 = n44320 & n44328 ;
  assign n44330 = n44315 & n44329 ;
  assign n44331 = ~\a[50]  & ~n44330 ;
  assign n44332 = ~n44327 & ~n44331 ;
  assign n44333 = n44037 & ~n44139 ;
  assign n44334 = ~n44139 & n44140 ;
  assign n44335 = ~n44333 & ~n44334 ;
  assign n44336 = n44332 & n44335 ;
  assign n44337 = ~n44308 & n44336 ;
  assign n44338 = n44332 & ~n44335 ;
  assign n44339 = n44308 & n44338 ;
  assign n44340 = ~n44337 & ~n44339 ;
  assign n44341 = ~n44332 & ~n44335 ;
  assign n44342 = ~n44308 & n44341 ;
  assign n44343 = ~n44332 & n44335 ;
  assign n44344 = n44308 & n44343 ;
  assign n44345 = ~n44342 & ~n44344 ;
  assign n44346 = n44340 & n44345 ;
  assign n44347 = n44182 & ~n44346 ;
  assign n44348 = ~n44182 & n44346 ;
  assign n44349 = ~n44347 & ~n44348 ;
  assign n44350 = ~n43990 & n44150 ;
  assign n44351 = n43994 & ~n44350 ;
  assign n44352 = ~n44349 & ~n44351 ;
  assign n44353 = n44349 & n44351 ;
  assign n44354 = ~n44352 & ~n44353 ;
  assign n44355 = ~n44155 & n44354 ;
  assign n44356 = ~n44157 & n44355 ;
  assign n44357 = ~n44160 & n44356 ;
  assign n44358 = ~n44155 & ~n44157 ;
  assign n44359 = ~n44160 & n44358 ;
  assign n44360 = ~n44354 & ~n44359 ;
  assign n44361 = ~n44357 & ~n44360 ;
  assign n44362 = ~n44155 & ~n44353 ;
  assign n44363 = ~n44157 & n44362 ;
  assign n44364 = ~n44160 & n44363 ;
  assign n44365 = ~n17690 & n37945 ;
  assign n44366 = ~n17688 & n44365 ;
  assign n44367 = \b[55]  & n17308 ;
  assign n44368 = n17305 & n44367 ;
  assign n44369 = ~\a[54]  & \b[56]  ;
  assign n44370 = n16647 & n44369 ;
  assign n44371 = ~n44368 & ~n44370 ;
  assign n44372 = \b[57]  & n16653 ;
  assign n44373 = \a[54]  & \b[56]  ;
  assign n44374 = n16644 & n44373 ;
  assign n44375 = \a[56]  & ~n44374 ;
  assign n44376 = ~n44372 & n44375 ;
  assign n44377 = n44371 & n44376 ;
  assign n44378 = ~n44366 & n44377 ;
  assign n44379 = ~n44372 & ~n44374 ;
  assign n44380 = n44371 & n44379 ;
  assign n44381 = ~n44366 & n44380 ;
  assign n44382 = ~\a[56]  & ~n44381 ;
  assign n44383 = ~n44378 & ~n44382 ;
  assign n44384 = ~n44269 & ~n44274 ;
  assign n44385 = ~n44271 & ~n44276 ;
  assign n44386 = n44205 & n44385 ;
  assign n44387 = n44384 & ~n44386 ;
  assign n44388 = n44383 & ~n44387 ;
  assign n44389 = ~n44383 & n44387 ;
  assign n44390 = ~n44388 & ~n44389 ;
  assign n44391 = n14793 & n20260 ;
  assign n44392 = ~n20257 & n44391 ;
  assign n44393 = n14793 & n40498 ;
  assign n44394 = ~n20256 & n44393 ;
  assign n44395 = \b[58]  & n15517 ;
  assign n44396 = n15514 & n44395 ;
  assign n44397 = ~\a[51]  & \b[59]  ;
  assign n44398 = n14785 & n44397 ;
  assign n44399 = ~n44396 & ~n44398 ;
  assign n44400 = \b[60]  & n14791 ;
  assign n44401 = \a[51]  & \b[59]  ;
  assign n44402 = n14782 & n44401 ;
  assign n44403 = \a[53]  & ~n44402 ;
  assign n44404 = ~n44400 & n44403 ;
  assign n44405 = n44399 & n44404 ;
  assign n44406 = ~n44394 & n44405 ;
  assign n44407 = ~n44392 & n44406 ;
  assign n44408 = ~n44400 & ~n44402 ;
  assign n44409 = n44399 & n44408 ;
  assign n44410 = ~n44394 & n44409 ;
  assign n44411 = ~n44392 & n44410 ;
  assign n44412 = ~\a[53]  & ~n44411 ;
  assign n44413 = ~n44407 & ~n44412 ;
  assign n44414 = ~n44243 & n44267 ;
  assign n44415 = n44248 & ~n44414 ;
  assign n44416 = ~n17912 & ~n18513 ;
  assign n44417 = ~n43785 & n44416 ;
  assign n44418 = \b[52]  & n19183 ;
  assign n44419 = n19180 & n44418 ;
  assign n44420 = \b[54]  & n18514 ;
  assign n44421 = \a[56]  & \b[53]  ;
  assign n44422 = n19181 & n44421 ;
  assign n44423 = ~\a[57]  & \b[53]  ;
  assign n44424 = n18508 & n44423 ;
  assign n44425 = ~n44422 & ~n44424 ;
  assign n44426 = ~n44420 & n44425 ;
  assign n44427 = ~n44419 & n44426 ;
  assign n44428 = ~n44417 & n44427 ;
  assign n44429 = ~\a[59]  & ~n44428 ;
  assign n44430 = \a[59]  & n44427 ;
  assign n44431 = ~n44417 & n44430 ;
  assign n44432 = ~n44429 & ~n44431 ;
  assign n44433 = ~n44092 & ~n44213 ;
  assign n44434 = ~n44239 & n44433 ;
  assign n44435 = ~n44212 & ~n44434 ;
  assign n44436 = ~n14098 & n20521 ;
  assign n44437 = ~n14096 & n44436 ;
  assign n44438 = \b[51]  & n20519 ;
  assign n44439 = \a[60]  & \b[50]  ;
  assign n44440 = n20510 & n44439 ;
  assign n44441 = ~n44438 & ~n44440 ;
  assign n44442 = \b[49]  & n21315 ;
  assign n44443 = n21312 & n44442 ;
  assign n44444 = ~\a[60]  & \b[50]  ;
  assign n44445 = n20513 & n44444 ;
  assign n44446 = ~n44443 & ~n44445 ;
  assign n44447 = n44441 & n44446 ;
  assign n44448 = ~n44437 & n44447 ;
  assign n44449 = ~\a[47]  & n44210 ;
  assign n44450 = ~\a[47]  & \b[47]  ;
  assign n44451 = n21958 & n44450 ;
  assign n44452 = ~n44449 & ~n44451 ;
  assign n44453 = \a[47]  & ~n44210 ;
  assign n44454 = ~n44209 & n44453 ;
  assign n44455 = n44452 & ~n44454 ;
  assign n44456 = \b[48]  & n21958 ;
  assign n44457 = \b[47]  & n21957 ;
  assign n44458 = ~n44456 & ~n44457 ;
  assign n44459 = ~\a[62]  & ~n44458 ;
  assign n44460 = ~n44455 & n44459 ;
  assign n44461 = ~\a[62]  & n44458 ;
  assign n44462 = n44455 & n44461 ;
  assign n44463 = ~n44460 & ~n44462 ;
  assign n44464 = ~n44448 & ~n44463 ;
  assign n44465 = \a[62]  & ~n44458 ;
  assign n44466 = ~n44455 & n44465 ;
  assign n44467 = \a[62]  & n44458 ;
  assign n44468 = n44455 & n44467 ;
  assign n44469 = ~n44466 & ~n44468 ;
  assign n44470 = n44447 & ~n44469 ;
  assign n44471 = ~n44437 & n44470 ;
  assign n44472 = ~n44464 & ~n44471 ;
  assign n44473 = ~\a[62]  & ~n44448 ;
  assign n44474 = ~n44455 & ~n44458 ;
  assign n44475 = n44455 & n44458 ;
  assign n44476 = ~n44474 & ~n44475 ;
  assign n44477 = \a[62]  & n44447 ;
  assign n44478 = ~n44437 & n44477 ;
  assign n44479 = n44476 & ~n44478 ;
  assign n44480 = ~n44473 & n44479 ;
  assign n44481 = n44472 & ~n44480 ;
  assign n44482 = n44435 & n44481 ;
  assign n44483 = ~n44435 & ~n44481 ;
  assign n44484 = ~n44482 & ~n44483 ;
  assign n44485 = n44432 & ~n44484 ;
  assign n44486 = ~n44432 & n44484 ;
  assign n44487 = ~n44485 & ~n44486 ;
  assign n44488 = n44415 & n44487 ;
  assign n44489 = ~n44415 & ~n44487 ;
  assign n44490 = ~n44488 & ~n44489 ;
  assign n44491 = n44413 & ~n44490 ;
  assign n44492 = ~n44390 & n44491 ;
  assign n44493 = n44413 & n44490 ;
  assign n44494 = n44390 & n44493 ;
  assign n44495 = ~n44492 & ~n44494 ;
  assign n44496 = ~n44413 & n44490 ;
  assign n44497 = ~n44390 & n44496 ;
  assign n44498 = ~n44413 & ~n44490 ;
  assign n44499 = n44390 & n44498 ;
  assign n44500 = ~n44497 & ~n44499 ;
  assign n44501 = n44495 & n44500 ;
  assign n44502 = ~n44284 & n44305 ;
  assign n44503 = ~n44285 & ~n44502 ;
  assign n44504 = n44501 & n44503 ;
  assign n44505 = ~n44501 & ~n44503 ;
  assign n44506 = ~n44504 & ~n44505 ;
  assign n44507 = n13125 & ~n22461 ;
  assign n44508 = ~n22459 & n44507 ;
  assign n44509 = \b[61]  & n13794 ;
  assign n44510 = n13792 & n44509 ;
  assign n44511 = ~\a[48]  & \b[62]  ;
  assign n44512 = n13117 & n44511 ;
  assign n44513 = ~n44510 & ~n44512 ;
  assign n44514 = \b[63]  & n13123 ;
  assign n44515 = \a[48]  & \b[62]  ;
  assign n44516 = n13786 & n44515 ;
  assign n44517 = \a[50]  & ~n44516 ;
  assign n44518 = ~n44514 & n44517 ;
  assign n44519 = n44513 & n44518 ;
  assign n44520 = ~n44508 & n44519 ;
  assign n44521 = ~n44514 & ~n44516 ;
  assign n44522 = n44513 & n44521 ;
  assign n44523 = ~n44508 & n44522 ;
  assign n44524 = ~\a[50]  & ~n44523 ;
  assign n44525 = ~n44520 & ~n44524 ;
  assign n44526 = n44506 & ~n44525 ;
  assign n44527 = ~n44506 & n44525 ;
  assign n44528 = ~n44526 & ~n44527 ;
  assign n44529 = ~n44308 & ~n44335 ;
  assign n44530 = n44308 & n44335 ;
  assign n44531 = n44332 & ~n44530 ;
  assign n44532 = ~n44529 & ~n44531 ;
  assign n44533 = ~n44528 & ~n44532 ;
  assign n44534 = n44528 & n44532 ;
  assign n44535 = ~n44533 & ~n44534 ;
  assign n44536 = ~n44177 & n44346 ;
  assign n44537 = n44181 & ~n44536 ;
  assign n44538 = ~n44535 & ~n44537 ;
  assign n44539 = n44535 & n44537 ;
  assign n44540 = ~n44538 & ~n44539 ;
  assign n44541 = ~n44352 & n44540 ;
  assign n44542 = ~n44364 & n44541 ;
  assign n44543 = ~n44352 & ~n44364 ;
  assign n44544 = ~n44540 & ~n44543 ;
  assign n44545 = ~n44542 & ~n44544 ;
  assign n44546 = ~n44526 & ~n44532 ;
  assign n44547 = ~n44527 & ~n44546 ;
  assign n44548 = n14793 & ~n20971 ;
  assign n44549 = ~n20969 & n44548 ;
  assign n44550 = \b[59]  & n15517 ;
  assign n44551 = n15514 & n44550 ;
  assign n44552 = ~\a[51]  & \b[60]  ;
  assign n44553 = n14785 & n44552 ;
  assign n44554 = ~n44551 & ~n44553 ;
  assign n44555 = \b[61]  & n14791 ;
  assign n44556 = \a[51]  & \b[60]  ;
  assign n44557 = n14782 & n44556 ;
  assign n44558 = \a[53]  & ~n44557 ;
  assign n44559 = ~n44555 & n44558 ;
  assign n44560 = n44554 & n44559 ;
  assign n44561 = ~n44549 & n44560 ;
  assign n44562 = ~n44555 & ~n44557 ;
  assign n44563 = n44554 & n44562 ;
  assign n44564 = ~n44549 & n44563 ;
  assign n44565 = ~\a[53]  & ~n44564 ;
  assign n44566 = ~n44561 & ~n44565 ;
  assign n44567 = n44383 & ~n44490 ;
  assign n44568 = ~n44387 & ~n44490 ;
  assign n44569 = ~n44388 & ~n44568 ;
  assign n44570 = ~n44567 & n44569 ;
  assign n44571 = n16655 & ~n19543 ;
  assign n44572 = ~n38598 & n44571 ;
  assign n44573 = \b[56]  & n17308 ;
  assign n44574 = n17305 & n44573 ;
  assign n44575 = ~\a[54]  & \b[57]  ;
  assign n44576 = n16647 & n44575 ;
  assign n44577 = ~n44574 & ~n44576 ;
  assign n44578 = \b[58]  & n16653 ;
  assign n44579 = \a[54]  & \b[57]  ;
  assign n44580 = n16644 & n44579 ;
  assign n44581 = \a[56]  & ~n44580 ;
  assign n44582 = ~n44578 & n44581 ;
  assign n44583 = n44577 & n44582 ;
  assign n44584 = ~n44572 & n44583 ;
  assign n44585 = ~n44578 & ~n44580 ;
  assign n44586 = n44577 & n44585 ;
  assign n44587 = ~n44572 & n44586 ;
  assign n44588 = ~\a[56]  & ~n44587 ;
  assign n44589 = ~n44584 & ~n44588 ;
  assign n44590 = ~n44415 & ~n44486 ;
  assign n44591 = ~n44485 & ~n44590 ;
  assign n44592 = ~n16446 & n18516 ;
  assign n44593 = ~n16444 & n44592 ;
  assign n44594 = \b[55]  & n18514 ;
  assign n44595 = \a[56]  & \b[54]  ;
  assign n44596 = n19181 & n44595 ;
  assign n44597 = ~\a[57]  & \b[54]  ;
  assign n44598 = n18508 & n44597 ;
  assign n44599 = ~n44596 & ~n44598 ;
  assign n44600 = ~n44594 & n44599 ;
  assign n44601 = \b[53]  & n19183 ;
  assign n44602 = n19180 & n44601 ;
  assign n44603 = \a[59]  & ~n44602 ;
  assign n44604 = n44600 & n44603 ;
  assign n44605 = ~n44593 & n44604 ;
  assign n44606 = n44600 & ~n44602 ;
  assign n44607 = ~n44593 & n44606 ;
  assign n44608 = ~\a[59]  & ~n44607 ;
  assign n44609 = ~n44605 & ~n44608 ;
  assign n44610 = ~n44435 & n44472 ;
  assign n44611 = \a[62]  & n44476 ;
  assign n44612 = ~n44448 & n44611 ;
  assign n44613 = ~\a[62]  & n44476 ;
  assign n44614 = n44448 & n44613 ;
  assign n44615 = ~n44612 & ~n44614 ;
  assign n44616 = ~n44610 & n44615 ;
  assign n44617 = ~n15201 & ~n19861 ;
  assign n44618 = ~n20518 & n44617 ;
  assign n44619 = n15198 & n44618 ;
  assign n44620 = n15201 & ~n19861 ;
  assign n44621 = ~n20518 & n44620 ;
  assign n44622 = ~n15198 & n44621 ;
  assign n44623 = ~n44619 & ~n44622 ;
  assign n44624 = \b[52]  & n20519 ;
  assign n44625 = \a[60]  & \b[51]  ;
  assign n44626 = n20510 & n44625 ;
  assign n44627 = ~n44624 & ~n44626 ;
  assign n44628 = \b[50]  & n21315 ;
  assign n44629 = n21312 & n44628 ;
  assign n44630 = ~\a[60]  & \b[51]  ;
  assign n44631 = n20513 & n44630 ;
  assign n44632 = ~n44629 & ~n44631 ;
  assign n44633 = n44627 & n44632 ;
  assign n44634 = n44623 & n44633 ;
  assign n44635 = n44452 & n44458 ;
  assign n44636 = ~n44454 & ~n44635 ;
  assign n44637 = \b[49]  & n21958 ;
  assign n44638 = \b[48]  & n21957 ;
  assign n44639 = ~n44637 & ~n44638 ;
  assign n44640 = ~n44636 & ~n44639 ;
  assign n44641 = ~n44454 & n44639 ;
  assign n44642 = ~n44635 & n44641 ;
  assign n44643 = ~\a[62]  & ~n44642 ;
  assign n44644 = ~n44640 & n44643 ;
  assign n44645 = ~n44634 & n44644 ;
  assign n44646 = \a[62]  & ~n44642 ;
  assign n44647 = ~n44640 & n44646 ;
  assign n44648 = n44633 & n44647 ;
  assign n44649 = n44623 & n44648 ;
  assign n44650 = ~n44645 & ~n44649 ;
  assign n44651 = ~\a[62]  & ~n44634 ;
  assign n44652 = ~n44640 & ~n44642 ;
  assign n44653 = \a[62]  & n44633 ;
  assign n44654 = n44623 & n44653 ;
  assign n44655 = ~n44652 & ~n44654 ;
  assign n44656 = ~n44651 & n44655 ;
  assign n44657 = n44650 & ~n44656 ;
  assign n44658 = n44616 & n44657 ;
  assign n44659 = ~n44616 & ~n44657 ;
  assign n44660 = ~n44658 & ~n44659 ;
  assign n44661 = n44609 & n44660 ;
  assign n44662 = ~n44609 & ~n44660 ;
  assign n44663 = ~n44661 & ~n44662 ;
  assign n44664 = n44591 & ~n44663 ;
  assign n44665 = ~n44591 & n44663 ;
  assign n44666 = ~n44664 & ~n44665 ;
  assign n44667 = ~n44589 & n44666 ;
  assign n44668 = n44589 & ~n44666 ;
  assign n44669 = ~n44667 & ~n44668 ;
  assign n44670 = n44570 & n44669 ;
  assign n44671 = ~n44570 & ~n44669 ;
  assign n44672 = ~n44670 & ~n44671 ;
  assign n44673 = n44566 & n44672 ;
  assign n44674 = ~n44566 & ~n44672 ;
  assign n44675 = ~n44673 & ~n44674 ;
  assign n44676 = n44500 & ~n44503 ;
  assign n44677 = n44495 & ~n44676 ;
  assign n44678 = \b[62]  & n13794 ;
  assign n44679 = n13792 & n44678 ;
  assign n44680 = ~\a[48]  & \b[63]  ;
  assign n44681 = n13117 & n44680 ;
  assign n44682 = \a[48]  & \b[63]  ;
  assign n44683 = n13786 & n44682 ;
  assign n44684 = ~n44681 & ~n44683 ;
  assign n44685 = ~n44679 & n44684 ;
  assign n44686 = ~\a[50]  & ~n44685 ;
  assign n44687 = n13125 & ~n22458 ;
  assign n44688 = ~\a[50]  & n44687 ;
  assign n44689 = ~n23173 & n44688 ;
  assign n44690 = ~n44686 & ~n44689 ;
  assign n44691 = ~n23173 & n44687 ;
  assign n44692 = \a[50]  & n44685 ;
  assign n44693 = ~n44691 & n44692 ;
  assign n44694 = n44690 & ~n44693 ;
  assign n44695 = ~n44677 & ~n44694 ;
  assign n44696 = ~n44675 & n44695 ;
  assign n44697 = n44677 & ~n44694 ;
  assign n44698 = n44675 & n44697 ;
  assign n44699 = ~n44696 & ~n44698 ;
  assign n44700 = n44677 & n44694 ;
  assign n44701 = ~n44675 & n44700 ;
  assign n44702 = ~n44677 & n44694 ;
  assign n44703 = n44675 & n44702 ;
  assign n44704 = ~n44701 & ~n44703 ;
  assign n44705 = n44699 & n44704 ;
  assign n44706 = ~n44547 & ~n44705 ;
  assign n44707 = n44547 & n44705 ;
  assign n44708 = ~n44706 & ~n44707 ;
  assign n44709 = n44539 & n44708 ;
  assign n44710 = ~n44539 & ~n44708 ;
  assign n44711 = ~n44709 & ~n44710 ;
  assign n44712 = ~n44542 & n44711 ;
  assign n44713 = ~n44708 & ~n44709 ;
  assign n44714 = n44542 & n44713 ;
  assign n44715 = ~n44712 & ~n44714 ;
  assign n44716 = n44542 & n44708 ;
  assign n44717 = n44566 & ~n44670 ;
  assign n44718 = ~n13122 & n39033 ;
  assign n44719 = ~n23171 & n44718 ;
  assign n44720 = ~n12606 & n44719 ;
  assign n44721 = \a[47]  & \a[49]  ;
  assign n44722 = \a[48]  & ~\a[50]  ;
  assign n44723 = n44721 & n44722 ;
  assign n44724 = ~\a[47]  & ~\a[49]  ;
  assign n44725 = ~\a[48]  & \a[50]  ;
  assign n44726 = n44724 & n44725 ;
  assign n44727 = ~n44723 & ~n44726 ;
  assign n44728 = \b[63]  & ~n44727 ;
  assign n44729 = \a[50]  & ~n44728 ;
  assign n44730 = ~n44720 & n44729 ;
  assign n44731 = ~\a[50]  & n44728 ;
  assign n44732 = ~\a[50]  & ~n12606 ;
  assign n44733 = n44719 & n44732 ;
  assign n44734 = ~n44731 & ~n44733 ;
  assign n44735 = ~n44730 & n44734 ;
  assign n44736 = ~n44671 & ~n44735 ;
  assign n44737 = ~n44717 & n44736 ;
  assign n44738 = ~n44671 & ~n44717 ;
  assign n44739 = n44735 & ~n44738 ;
  assign n44740 = ~n44737 & ~n44739 ;
  assign n44741 = n44609 & ~n44658 ;
  assign n44742 = ~n44659 & ~n44741 ;
  assign n44743 = ~n44642 & ~n44649 ;
  assign n44744 = ~n44645 & n44743 ;
  assign n44745 = ~n15246 & n20521 ;
  assign n44746 = ~n15244 & n44745 ;
  assign n44747 = \b[53]  & n20519 ;
  assign n44748 = \a[60]  & \b[52]  ;
  assign n44749 = n20510 & n44748 ;
  assign n44750 = ~n44747 & ~n44749 ;
  assign n44751 = \b[51]  & n21315 ;
  assign n44752 = n21312 & n44751 ;
  assign n44753 = ~\a[60]  & \b[52]  ;
  assign n44754 = n20513 & n44753 ;
  assign n44755 = ~n44752 & ~n44754 ;
  assign n44756 = n44750 & n44755 ;
  assign n44757 = ~n44746 & n44756 ;
  assign n44758 = \b[50]  & n21958 ;
  assign n44759 = \b[49]  & n21957 ;
  assign n44760 = ~n44758 & ~n44759 ;
  assign n44761 = n44639 & ~n44760 ;
  assign n44762 = ~n44639 & n44760 ;
  assign n44763 = ~n44761 & ~n44762 ;
  assign n44764 = ~\a[62]  & n44763 ;
  assign n44765 = ~n44757 & n44764 ;
  assign n44766 = \a[62]  & n44763 ;
  assign n44767 = n44756 & n44766 ;
  assign n44768 = ~n44746 & n44767 ;
  assign n44769 = ~n44765 & ~n44768 ;
  assign n44770 = ~\a[62]  & ~n44757 ;
  assign n44771 = \a[62]  & n44756 ;
  assign n44772 = ~n44746 & n44771 ;
  assign n44773 = ~n44763 & ~n44772 ;
  assign n44774 = ~n44770 & n44773 ;
  assign n44775 = n44769 & ~n44774 ;
  assign n44776 = n44744 & ~n44775 ;
  assign n44777 = ~n44744 & n44775 ;
  assign n44778 = ~n44776 & ~n44777 ;
  assign n44779 = ~n17647 & ~n17912 ;
  assign n44780 = ~n18513 & n44779 ;
  assign n44781 = n17644 & n44780 ;
  assign n44782 = n17647 & ~n17912 ;
  assign n44783 = ~n18513 & n44782 ;
  assign n44784 = ~n17644 & n44783 ;
  assign n44785 = ~n44781 & ~n44784 ;
  assign n44786 = \b[56]  & n18514 ;
  assign n44787 = \a[56]  & \b[55]  ;
  assign n44788 = n19181 & n44787 ;
  assign n44789 = ~\a[57]  & \b[55]  ;
  assign n44790 = n18508 & n44789 ;
  assign n44791 = ~n44788 & ~n44790 ;
  assign n44792 = ~n44786 & n44791 ;
  assign n44793 = \b[54]  & n19183 ;
  assign n44794 = n19180 & n44793 ;
  assign n44795 = \a[59]  & ~n44794 ;
  assign n44796 = n44792 & n44795 ;
  assign n44797 = n44785 & n44796 ;
  assign n44798 = n44792 & ~n44794 ;
  assign n44799 = n44785 & n44798 ;
  assign n44800 = ~\a[59]  & ~n44799 ;
  assign n44801 = ~n44797 & ~n44800 ;
  assign n44802 = ~n44778 & n44801 ;
  assign n44803 = n44778 & ~n44801 ;
  assign n44804 = ~n44802 & ~n44803 ;
  assign n44805 = n44742 & n44804 ;
  assign n44806 = ~n44742 & ~n44804 ;
  assign n44807 = ~n44805 & ~n44806 ;
  assign n44808 = ~n19550 & n37945 ;
  assign n44809 = ~n19548 & n44808 ;
  assign n44810 = \b[57]  & n17308 ;
  assign n44811 = n17305 & n44810 ;
  assign n44812 = ~\a[54]  & \b[58]  ;
  assign n44813 = n16647 & n44812 ;
  assign n44814 = ~n44811 & ~n44813 ;
  assign n44815 = \b[59]  & n16653 ;
  assign n44816 = \a[54]  & \b[58]  ;
  assign n44817 = n16644 & n44816 ;
  assign n44818 = \a[56]  & ~n44817 ;
  assign n44819 = ~n44815 & n44818 ;
  assign n44820 = n44814 & n44819 ;
  assign n44821 = ~n44809 & n44820 ;
  assign n44822 = ~n44815 & ~n44817 ;
  assign n44823 = n44814 & n44822 ;
  assign n44824 = ~n44809 & n44823 ;
  assign n44825 = ~\a[56]  & ~n44824 ;
  assign n44826 = ~n44821 & ~n44825 ;
  assign n44827 = n44807 & ~n44826 ;
  assign n44828 = ~n44807 & n44826 ;
  assign n44829 = ~n44827 & ~n44828 ;
  assign n44830 = n44589 & ~n44664 ;
  assign n44831 = ~n44664 & n44665 ;
  assign n44832 = ~n44830 & ~n44831 ;
  assign n44833 = n14793 & n21696 ;
  assign n44834 = ~n21693 & n44833 ;
  assign n44835 = n14793 & n41213 ;
  assign n44836 = ~n21692 & n44835 ;
  assign n44837 = \b[60]  & n15517 ;
  assign n44838 = n15514 & n44837 ;
  assign n44839 = ~\a[51]  & \b[61]  ;
  assign n44840 = n14785 & n44839 ;
  assign n44841 = ~n44838 & ~n44840 ;
  assign n44842 = \b[62]  & n14791 ;
  assign n44843 = \a[51]  & \b[61]  ;
  assign n44844 = n14782 & n44843 ;
  assign n44845 = \a[53]  & ~n44844 ;
  assign n44846 = ~n44842 & n44845 ;
  assign n44847 = n44841 & n44846 ;
  assign n44848 = ~n44836 & n44847 ;
  assign n44849 = ~n44834 & n44848 ;
  assign n44850 = ~n44842 & ~n44844 ;
  assign n44851 = n44841 & n44850 ;
  assign n44852 = ~n44836 & n44851 ;
  assign n44853 = ~n44834 & n44852 ;
  assign n44854 = ~\a[53]  & ~n44853 ;
  assign n44855 = ~n44849 & ~n44854 ;
  assign n44856 = ~n44832 & n44855 ;
  assign n44857 = ~n44829 & n44856 ;
  assign n44858 = n44832 & n44855 ;
  assign n44859 = n44829 & n44858 ;
  assign n44860 = ~n44857 & ~n44859 ;
  assign n44861 = n44832 & ~n44855 ;
  assign n44862 = ~n44829 & n44861 ;
  assign n44863 = ~n44832 & ~n44855 ;
  assign n44864 = n44829 & n44863 ;
  assign n44865 = ~n44862 & ~n44864 ;
  assign n44866 = n44860 & n44865 ;
  assign n44867 = n44740 & n44866 ;
  assign n44868 = ~n44740 & ~n44866 ;
  assign n44869 = ~n44867 & ~n44868 ;
  assign n44870 = n44675 & ~n44677 ;
  assign n44871 = n44566 & n44694 ;
  assign n44872 = ~n44672 & n44871 ;
  assign n44873 = ~n44566 & n44694 ;
  assign n44874 = n44672 & n44873 ;
  assign n44875 = ~n44872 & ~n44874 ;
  assign n44876 = ~n44702 & n44875 ;
  assign n44877 = ~n44870 & n44876 ;
  assign n44878 = ~n44869 & ~n44877 ;
  assign n44879 = n44869 & n44877 ;
  assign n44880 = ~n44878 & ~n44879 ;
  assign n44881 = ~n44707 & n44880 ;
  assign n44882 = ~n44709 & n44881 ;
  assign n44883 = ~n44716 & n44882 ;
  assign n44884 = ~n44707 & ~n44709 ;
  assign n44885 = ~n44716 & n44884 ;
  assign n44886 = ~n44880 & ~n44885 ;
  assign n44887 = ~n44883 & ~n44886 ;
  assign n44888 = ~n44707 & ~n44879 ;
  assign n44889 = ~n44709 & n44888 ;
  assign n44890 = ~n44716 & n44889 ;
  assign n44891 = n16655 & n20260 ;
  assign n44892 = ~n20257 & n44891 ;
  assign n44893 = n37945 & n40498 ;
  assign n44894 = ~n20256 & n44893 ;
  assign n44895 = \b[58]  & n17308 ;
  assign n44896 = n17305 & n44895 ;
  assign n44897 = ~\a[54]  & \b[59]  ;
  assign n44898 = n16647 & n44897 ;
  assign n44899 = ~n44896 & ~n44898 ;
  assign n44900 = \b[60]  & n16653 ;
  assign n44901 = \a[54]  & \b[59]  ;
  assign n44902 = n16644 & n44901 ;
  assign n44903 = \a[56]  & ~n44902 ;
  assign n44904 = ~n44900 & n44903 ;
  assign n44905 = n44899 & n44904 ;
  assign n44906 = ~n44894 & n44905 ;
  assign n44907 = ~n44892 & n44906 ;
  assign n44908 = ~n44900 & ~n44902 ;
  assign n44909 = n44899 & n44908 ;
  assign n44910 = ~n44894 & n44909 ;
  assign n44911 = ~n44892 & n44910 ;
  assign n44912 = ~\a[56]  & ~n44911 ;
  assign n44913 = ~n44907 & ~n44912 ;
  assign n44914 = ~n44777 & n44801 ;
  assign n44915 = ~n44776 & ~n44914 ;
  assign n44916 = ~n17690 & n18516 ;
  assign n44917 = ~n17688 & n44916 ;
  assign n44918 = \b[55]  & n19183 ;
  assign n44919 = n19180 & n44918 ;
  assign n44920 = \b[57]  & n18514 ;
  assign n44921 = \a[56]  & \b[56]  ;
  assign n44922 = n19181 & n44921 ;
  assign n44923 = ~\a[57]  & \b[56]  ;
  assign n44924 = n18508 & n44923 ;
  assign n44925 = ~n44922 & ~n44924 ;
  assign n44926 = ~n44920 & n44925 ;
  assign n44927 = ~n44919 & n44926 ;
  assign n44928 = ~\a[59]  & n44927 ;
  assign n44929 = ~n44917 & n44928 ;
  assign n44930 = ~n44917 & n44927 ;
  assign n44931 = \a[59]  & ~n44930 ;
  assign n44932 = ~n44929 & ~n44931 ;
  assign n44933 = ~n44761 & ~n44768 ;
  assign n44934 = ~n44765 & n44933 ;
  assign n44935 = ~\a[50]  & \b[50]  ;
  assign n44936 = n21957 & n44935 ;
  assign n44937 = ~\a[50]  & \b[51]  ;
  assign n44938 = n21958 & n44937 ;
  assign n44939 = ~n44936 & ~n44938 ;
  assign n44940 = \b[51]  & n21958 ;
  assign n44941 = \b[50]  & n21957 ;
  assign n44942 = \a[50]  & ~n44941 ;
  assign n44943 = ~n44940 & n44942 ;
  assign n44944 = n44939 & ~n44943 ;
  assign n44945 = ~n44639 & ~n44944 ;
  assign n44946 = n44639 & n44944 ;
  assign n44947 = ~n44945 & ~n44946 ;
  assign n44948 = ~n44934 & ~n44947 ;
  assign n44949 = n20521 & ~n43785 ;
  assign n44950 = \b[52]  & n21315 ;
  assign n44951 = n21312 & n44950 ;
  assign n44952 = ~\a[60]  & \b[53]  ;
  assign n44953 = n20513 & n44952 ;
  assign n44954 = ~n44951 & ~n44953 ;
  assign n44955 = \b[54]  & n20519 ;
  assign n44956 = \a[60]  & \b[53]  ;
  assign n44957 = n20510 & n44956 ;
  assign n44958 = \a[62]  & ~n44957 ;
  assign n44959 = ~n44955 & n44958 ;
  assign n44960 = n44954 & n44959 ;
  assign n44961 = ~n44949 & n44960 ;
  assign n44962 = ~n44955 & ~n44957 ;
  assign n44963 = n44954 & n44962 ;
  assign n44964 = ~n44949 & n44963 ;
  assign n44965 = ~\a[62]  & ~n44964 ;
  assign n44966 = ~n44961 & ~n44965 ;
  assign n44967 = n44934 & n44947 ;
  assign n44968 = ~n44966 & ~n44967 ;
  assign n44969 = ~n44948 & n44968 ;
  assign n44970 = ~n44948 & ~n44967 ;
  assign n44971 = n44966 & ~n44970 ;
  assign n44972 = ~n44969 & ~n44971 ;
  assign n44973 = n44932 & n44972 ;
  assign n44974 = ~n44932 & ~n44972 ;
  assign n44975 = ~n44973 & ~n44974 ;
  assign n44976 = n44915 & n44975 ;
  assign n44977 = ~n44915 & n44973 ;
  assign n44978 = ~n44915 & n44974 ;
  assign n44979 = ~n44977 & ~n44978 ;
  assign n44980 = ~n44976 & n44979 ;
  assign n44981 = ~n44913 & n44980 ;
  assign n44982 = n44913 & ~n44980 ;
  assign n44983 = ~n44981 & ~n44982 ;
  assign n44984 = ~n44805 & n44826 ;
  assign n44985 = ~n44806 & ~n44984 ;
  assign n44986 = n44983 & n44985 ;
  assign n44987 = ~n44983 & ~n44985 ;
  assign n44988 = ~n44986 & ~n44987 ;
  assign n44989 = n14793 & ~n22461 ;
  assign n44990 = ~n22459 & n44989 ;
  assign n44991 = \b[61]  & n15517 ;
  assign n44992 = n15514 & n44991 ;
  assign n44993 = ~\a[51]  & \b[62]  ;
  assign n44994 = n14785 & n44993 ;
  assign n44995 = ~n44992 & ~n44994 ;
  assign n44996 = \b[63]  & n14791 ;
  assign n44997 = \a[51]  & \b[62]  ;
  assign n44998 = n14782 & n44997 ;
  assign n44999 = \a[53]  & ~n44998 ;
  assign n45000 = ~n44996 & n44999 ;
  assign n45001 = n44995 & n45000 ;
  assign n45002 = ~n44990 & n45001 ;
  assign n45003 = ~n44996 & ~n44998 ;
  assign n45004 = n44995 & n45003 ;
  assign n45005 = ~n44990 & n45004 ;
  assign n45006 = ~\a[53]  & ~n45005 ;
  assign n45007 = ~n45002 & ~n45006 ;
  assign n45008 = n44988 & ~n45007 ;
  assign n45009 = ~n44988 & n45007 ;
  assign n45010 = ~n45008 & ~n45009 ;
  assign n45011 = ~n44829 & ~n44832 ;
  assign n45012 = n44829 & n44832 ;
  assign n45013 = n44855 & ~n45012 ;
  assign n45014 = ~n45011 & ~n45013 ;
  assign n45015 = ~n45010 & ~n45014 ;
  assign n45016 = n45010 & n45014 ;
  assign n45017 = ~n45015 & ~n45016 ;
  assign n45018 = ~n44737 & ~n44866 ;
  assign n45019 = ~n44739 & ~n45018 ;
  assign n45020 = ~n45017 & ~n45019 ;
  assign n45021 = n45017 & n45019 ;
  assign n45022 = ~n45020 & ~n45021 ;
  assign n45023 = ~n44878 & n45022 ;
  assign n45024 = ~n44890 & n45023 ;
  assign n45025 = ~n44878 & ~n44890 ;
  assign n45026 = ~n45022 & ~n45025 ;
  assign n45027 = ~n45024 & ~n45026 ;
  assign n45028 = ~n45008 & ~n45014 ;
  assign n45029 = ~n45009 & ~n45028 ;
  assign n45030 = ~n44981 & ~n44985 ;
  assign n45031 = ~n44982 & ~n45030 ;
  assign n45032 = ~n20971 & n37945 ;
  assign n45033 = ~n20969 & n45032 ;
  assign n45034 = \b[59]  & n17308 ;
  assign n45035 = n17305 & n45034 ;
  assign n45036 = ~\a[54]  & \b[60]  ;
  assign n45037 = n16647 & n45036 ;
  assign n45038 = ~n45035 & ~n45037 ;
  assign n45039 = \b[61]  & n16653 ;
  assign n45040 = \a[54]  & \b[60]  ;
  assign n45041 = n16644 & n45040 ;
  assign n45042 = \a[56]  & ~n45041 ;
  assign n45043 = ~n45039 & n45042 ;
  assign n45044 = n45038 & n45043 ;
  assign n45045 = ~n45033 & n45044 ;
  assign n45046 = ~n45039 & ~n45041 ;
  assign n45047 = n45038 & n45046 ;
  assign n45048 = ~n45033 & n45047 ;
  assign n45049 = ~\a[56]  & ~n45048 ;
  assign n45050 = ~n45045 & ~n45049 ;
  assign n45051 = ~n44973 & n44974 ;
  assign n45052 = ~n44915 & ~n44973 ;
  assign n45053 = ~n45051 & ~n45052 ;
  assign n45054 = n18516 & ~n19543 ;
  assign n45055 = ~n38598 & n45054 ;
  assign n45056 = \b[58]  & n18514 ;
  assign n45057 = \a[56]  & \b[57]  ;
  assign n45058 = n19181 & n45057 ;
  assign n45059 = ~\a[57]  & \b[57]  ;
  assign n45060 = n18508 & n45059 ;
  assign n45061 = ~n45058 & ~n45060 ;
  assign n45062 = ~n45056 & n45061 ;
  assign n45063 = \b[56]  & n19183 ;
  assign n45064 = n19180 & n45063 ;
  assign n45065 = \a[59]  & ~n45064 ;
  assign n45066 = n45062 & n45065 ;
  assign n45067 = ~n45055 & n45066 ;
  assign n45068 = n45062 & ~n45064 ;
  assign n45069 = ~n45055 & n45068 ;
  assign n45070 = ~\a[59]  & ~n45069 ;
  assign n45071 = ~n45067 & ~n45070 ;
  assign n45072 = ~n44948 & ~n44968 ;
  assign n45073 = ~n16446 & n20521 ;
  assign n45074 = ~n16444 & n45073 ;
  assign n45075 = \b[55]  & n20519 ;
  assign n45076 = \a[60]  & \b[54]  ;
  assign n45077 = n20510 & n45076 ;
  assign n45078 = ~n45075 & ~n45077 ;
  assign n45079 = \b[53]  & n21315 ;
  assign n45080 = n21312 & n45079 ;
  assign n45081 = ~\a[60]  & \b[54]  ;
  assign n45082 = n20513 & n45081 ;
  assign n45083 = ~n45080 & ~n45082 ;
  assign n45084 = n45078 & n45083 ;
  assign n45085 = ~n45074 & n45084 ;
  assign n45086 = ~\a[62]  & ~n45085 ;
  assign n45087 = ~n44639 & ~n44943 ;
  assign n45088 = \b[52]  & n21958 ;
  assign n45089 = \b[51]  & n21957 ;
  assign n45090 = ~n45088 & ~n45089 ;
  assign n45091 = n44939 & ~n45090 ;
  assign n45092 = ~n45087 & n45091 ;
  assign n45093 = n44939 & ~n45087 ;
  assign n45094 = n45090 & ~n45093 ;
  assign n45095 = ~n45092 & ~n45094 ;
  assign n45096 = \a[62]  & n45084 ;
  assign n45097 = ~n45074 & n45096 ;
  assign n45098 = ~n45095 & ~n45097 ;
  assign n45099 = ~n45086 & n45098 ;
  assign n45100 = ~\a[62]  & n45095 ;
  assign n45101 = ~n45085 & n45100 ;
  assign n45102 = \a[62]  & ~n45092 ;
  assign n45103 = ~n45094 & n45102 ;
  assign n45104 = n45084 & n45103 ;
  assign n45105 = ~n45074 & n45104 ;
  assign n45106 = ~n45101 & ~n45105 ;
  assign n45107 = ~n45099 & n45106 ;
  assign n45108 = ~n45072 & n45107 ;
  assign n45109 = n45072 & ~n45107 ;
  assign n45110 = ~n45108 & ~n45109 ;
  assign n45111 = n45071 & n45110 ;
  assign n45112 = ~n45071 & ~n45110 ;
  assign n45113 = ~n45111 & ~n45112 ;
  assign n45114 = n45053 & ~n45113 ;
  assign n45115 = ~n45053 & n45113 ;
  assign n45116 = ~n45114 & ~n45115 ;
  assign n45117 = n45050 & n45116 ;
  assign n45118 = ~n45050 & ~n45116 ;
  assign n45119 = ~n45117 & ~n45118 ;
  assign n45120 = n45031 & ~n45119 ;
  assign n45121 = ~n45031 & n45119 ;
  assign n45122 = ~n45120 & ~n45121 ;
  assign n45123 = n14793 & ~n22458 ;
  assign n45124 = ~n23173 & n45123 ;
  assign n45125 = \b[62]  & n15517 ;
  assign n45126 = n15514 & n45125 ;
  assign n45127 = \a[51]  & \b[63]  ;
  assign n45128 = n14782 & n45127 ;
  assign n45129 = ~\a[51]  & \b[63]  ;
  assign n45130 = n14785 & n45129 ;
  assign n45131 = \a[53]  & ~n45130 ;
  assign n45132 = ~n45128 & n45131 ;
  assign n45133 = ~n45126 & n45132 ;
  assign n45134 = ~n45124 & n45133 ;
  assign n45135 = ~n45128 & ~n45130 ;
  assign n45136 = ~n45126 & n45135 ;
  assign n45137 = ~n45124 & n45136 ;
  assign n45138 = ~\a[53]  & ~n45137 ;
  assign n45139 = ~n45134 & ~n45138 ;
  assign n45140 = n45122 & ~n45139 ;
  assign n45141 = ~n45122 & n45139 ;
  assign n45142 = ~n45140 & ~n45141 ;
  assign n45143 = ~n45029 & ~n45142 ;
  assign n45144 = n45029 & n45142 ;
  assign n45145 = ~n45143 & ~n45144 ;
  assign n45146 = n45021 & n45145 ;
  assign n45147 = ~n45021 & ~n45145 ;
  assign n45148 = ~n45146 & ~n45147 ;
  assign n45149 = ~n45024 & n45148 ;
  assign n45150 = ~n45145 & ~n45146 ;
  assign n45151 = n45024 & n45150 ;
  assign n45152 = ~n45149 & ~n45151 ;
  assign n45153 = n45024 & n45145 ;
  assign n45154 = n45050 & ~n45114 ;
  assign n45155 = n14793 & n39033 ;
  assign n45156 = ~n23171 & n45155 ;
  assign n45157 = \a[50]  & \a[52]  ;
  assign n45158 = \a[51]  & ~\a[53]  ;
  assign n45159 = n45157 & n45158 ;
  assign n45160 = ~\a[50]  & ~\a[52]  ;
  assign n45161 = ~\a[51]  & \a[53]  ;
  assign n45162 = n45160 & n45161 ;
  assign n45163 = ~n45159 & ~n45162 ;
  assign n45164 = \b[63]  & ~n45163 ;
  assign n45165 = \a[53]  & ~n45164 ;
  assign n45166 = ~n45156 & n45165 ;
  assign n45167 = ~n45156 & ~n45164 ;
  assign n45168 = ~\a[53]  & ~n45167 ;
  assign n45169 = ~n45166 & ~n45168 ;
  assign n45170 = ~n45115 & ~n45169 ;
  assign n45171 = ~n45154 & n45170 ;
  assign n45172 = ~n45115 & ~n45154 ;
  assign n45173 = n45169 & ~n45172 ;
  assign n45174 = ~n45171 & ~n45173 ;
  assign n45175 = n45071 & ~n45108 ;
  assign n45176 = ~n45109 & ~n45175 ;
  assign n45177 = n18516 & ~n19550 ;
  assign n45178 = ~n19548 & n45177 ;
  assign n45179 = \b[59]  & n18514 ;
  assign n45180 = \a[56]  & \b[58]  ;
  assign n45181 = n19181 & n45180 ;
  assign n45182 = ~\a[57]  & \b[58]  ;
  assign n45183 = n18508 & n45182 ;
  assign n45184 = ~n45181 & ~n45183 ;
  assign n45185 = ~n45179 & n45184 ;
  assign n45186 = \b[57]  & n19183 ;
  assign n45187 = n19180 & n45186 ;
  assign n45188 = \a[59]  & ~n45187 ;
  assign n45189 = n45185 & n45188 ;
  assign n45190 = ~n45178 & n45189 ;
  assign n45191 = n45185 & ~n45187 ;
  assign n45192 = ~n45178 & n45191 ;
  assign n45193 = ~\a[59]  & ~n45192 ;
  assign n45194 = ~n45190 & ~n45193 ;
  assign n45195 = ~n45094 & ~n45105 ;
  assign n45196 = ~n45101 & n45195 ;
  assign n45197 = \b[53]  & n21958 ;
  assign n45198 = \b[52]  & n21957 ;
  assign n45199 = ~n45197 & ~n45198 ;
  assign n45200 = n45090 & ~n45199 ;
  assign n45201 = ~n45090 & n45199 ;
  assign n45202 = ~n45200 & ~n45201 ;
  assign n45203 = ~n45196 & n45202 ;
  assign n45204 = ~n17647 & ~n19861 ;
  assign n45205 = ~n20518 & n45204 ;
  assign n45206 = n17644 & n45205 ;
  assign n45207 = n17647 & ~n19861 ;
  assign n45208 = ~n20518 & n45207 ;
  assign n45209 = ~n17644 & n45208 ;
  assign n45210 = ~n45206 & ~n45209 ;
  assign n45211 = \b[54]  & n21315 ;
  assign n45212 = n21312 & n45211 ;
  assign n45213 = ~\a[60]  & \b[55]  ;
  assign n45214 = n20513 & n45213 ;
  assign n45215 = ~n45212 & ~n45214 ;
  assign n45216 = \b[56]  & n20519 ;
  assign n45217 = \a[60]  & \b[55]  ;
  assign n45218 = n20510 & n45217 ;
  assign n45219 = \a[62]  & ~n45218 ;
  assign n45220 = ~n45216 & n45219 ;
  assign n45221 = n45215 & n45220 ;
  assign n45222 = n45210 & n45221 ;
  assign n45223 = ~n45216 & ~n45218 ;
  assign n45224 = n45215 & n45223 ;
  assign n45225 = n45210 & n45224 ;
  assign n45226 = ~\a[62]  & ~n45225 ;
  assign n45227 = ~n45222 & ~n45226 ;
  assign n45228 = n45196 & ~n45202 ;
  assign n45229 = ~n45227 & ~n45228 ;
  assign n45230 = ~n45203 & n45229 ;
  assign n45231 = ~n45203 & ~n45228 ;
  assign n45232 = n45227 & ~n45231 ;
  assign n45233 = ~n45230 & ~n45232 ;
  assign n45234 = n45194 & ~n45233 ;
  assign n45235 = ~n45176 & n45234 ;
  assign n45236 = ~n45194 & n45233 ;
  assign n45237 = ~n45176 & n45236 ;
  assign n45238 = ~n45235 & ~n45237 ;
  assign n45239 = ~n45234 & ~n45236 ;
  assign n45240 = n45176 & n45239 ;
  assign n45241 = n45238 & ~n45240 ;
  assign n45242 = n16655 & n21696 ;
  assign n45243 = ~n21693 & n45242 ;
  assign n45244 = n37945 & n41213 ;
  assign n45245 = ~n21692 & n45244 ;
  assign n45246 = \b[60]  & n17308 ;
  assign n45247 = n17305 & n45246 ;
  assign n45248 = ~\a[54]  & \b[61]  ;
  assign n45249 = n16647 & n45248 ;
  assign n45250 = ~n45247 & ~n45249 ;
  assign n45251 = \b[62]  & n16653 ;
  assign n45252 = \a[54]  & \b[61]  ;
  assign n45253 = n16644 & n45252 ;
  assign n45254 = \a[56]  & ~n45253 ;
  assign n45255 = ~n45251 & n45254 ;
  assign n45256 = n45250 & n45255 ;
  assign n45257 = ~n45245 & n45256 ;
  assign n45258 = ~n45243 & n45257 ;
  assign n45259 = ~n45251 & ~n45253 ;
  assign n45260 = n45250 & n45259 ;
  assign n45261 = ~n45245 & n45260 ;
  assign n45262 = ~n45243 & n45261 ;
  assign n45263 = ~\a[56]  & ~n45262 ;
  assign n45264 = ~n45258 & ~n45263 ;
  assign n45265 = n45241 & ~n45264 ;
  assign n45266 = ~n45241 & n45264 ;
  assign n45267 = ~n45265 & ~n45266 ;
  assign n45268 = n45174 & n45267 ;
  assign n45269 = ~n45174 & ~n45267 ;
  assign n45270 = ~n45268 & ~n45269 ;
  assign n45271 = ~n45120 & n45139 ;
  assign n45272 = ~n45121 & ~n45271 ;
  assign n45273 = ~n45270 & ~n45272 ;
  assign n45274 = n45270 & n45272 ;
  assign n45275 = ~n45273 & ~n45274 ;
  assign n45276 = ~n45144 & n45275 ;
  assign n45277 = ~n45146 & n45276 ;
  assign n45278 = ~n45153 & n45277 ;
  assign n45279 = ~n45144 & ~n45146 ;
  assign n45280 = ~n45153 & n45279 ;
  assign n45281 = ~n45275 & ~n45280 ;
  assign n45282 = ~n45278 & ~n45281 ;
  assign n45283 = ~n45144 & ~n45274 ;
  assign n45284 = ~n45146 & n45283 ;
  assign n45285 = ~n45153 & n45284 ;
  assign n45286 = ~n22461 & n37945 ;
  assign n45287 = ~n22459 & n45286 ;
  assign n45288 = \b[61]  & n17308 ;
  assign n45289 = n17305 & n45288 ;
  assign n45290 = ~\a[54]  & \b[62]  ;
  assign n45291 = n16647 & n45290 ;
  assign n45292 = ~n45289 & ~n45291 ;
  assign n45293 = \b[63]  & n16653 ;
  assign n45294 = \a[54]  & \b[62]  ;
  assign n45295 = n16644 & n45294 ;
  assign n45296 = \a[56]  & ~n45295 ;
  assign n45297 = ~n45293 & n45296 ;
  assign n45298 = n45292 & n45297 ;
  assign n45299 = ~n45287 & n45298 ;
  assign n45300 = ~n45293 & ~n45295 ;
  assign n45301 = n45292 & n45300 ;
  assign n45302 = ~n45287 & n45301 ;
  assign n45303 = ~\a[56]  & ~n45302 ;
  assign n45304 = ~n45299 & ~n45303 ;
  assign n45305 = ~n45240 & n45264 ;
  assign n45306 = n45238 & ~n45305 ;
  assign n45307 = n45227 & n45228 ;
  assign n45308 = n45203 & n45227 ;
  assign n45309 = ~n45307 & ~n45308 ;
  assign n45310 = n45194 & ~n45230 ;
  assign n45311 = n45309 & ~n45310 ;
  assign n45312 = n18516 & n20260 ;
  assign n45313 = ~n20257 & n45312 ;
  assign n45314 = n18516 & n40498 ;
  assign n45315 = ~n20256 & n45314 ;
  assign n45316 = \b[58]  & n19183 ;
  assign n45317 = n19180 & n45316 ;
  assign n45318 = \b[60]  & n18514 ;
  assign n45319 = \a[56]  & \b[59]  ;
  assign n45320 = n19181 & n45319 ;
  assign n45321 = ~\a[57]  & \b[59]  ;
  assign n45322 = n18508 & n45321 ;
  assign n45323 = ~n45320 & ~n45322 ;
  assign n45324 = ~n45318 & n45323 ;
  assign n45325 = ~n45317 & n45324 ;
  assign n45326 = ~n45315 & n45325 ;
  assign n45327 = ~n45313 & n45326 ;
  assign n45328 = ~\a[59]  & ~n45327 ;
  assign n45329 = \a[59]  & n45325 ;
  assign n45330 = ~n45315 & n45329 ;
  assign n45331 = ~n45313 & n45330 ;
  assign n45332 = ~n45328 & ~n45331 ;
  assign n45333 = ~n45094 & ~n45201 ;
  assign n45334 = ~n45105 & n45333 ;
  assign n45335 = ~n45101 & n45334 ;
  assign n45336 = ~n45200 & ~n45335 ;
  assign n45337 = ~n17690 & n20521 ;
  assign n45338 = ~n17688 & n45337 ;
  assign n45339 = \b[57]  & n20519 ;
  assign n45340 = \a[60]  & \b[56]  ;
  assign n45341 = n20510 & n45340 ;
  assign n45342 = ~n45339 & ~n45341 ;
  assign n45343 = \b[55]  & n21315 ;
  assign n45344 = n21312 & n45343 ;
  assign n45345 = ~\a[60]  & \b[56]  ;
  assign n45346 = n20513 & n45345 ;
  assign n45347 = ~n45344 & ~n45346 ;
  assign n45348 = n45342 & n45347 ;
  assign n45349 = ~n45338 & n45348 ;
  assign n45350 = ~\a[53]  & n45198 ;
  assign n45351 = ~\a[53]  & \b[53]  ;
  assign n45352 = n21958 & n45351 ;
  assign n45353 = ~n45350 & ~n45352 ;
  assign n45354 = \a[53]  & ~n45198 ;
  assign n45355 = ~n45197 & n45354 ;
  assign n45356 = n45353 & ~n45355 ;
  assign n45357 = \b[54]  & n21958 ;
  assign n45358 = \b[53]  & n21957 ;
  assign n45359 = ~n45357 & ~n45358 ;
  assign n45360 = ~\a[62]  & ~n45359 ;
  assign n45361 = ~n45356 & n45360 ;
  assign n45362 = ~\a[62]  & n45359 ;
  assign n45363 = n45356 & n45362 ;
  assign n45364 = ~n45361 & ~n45363 ;
  assign n45365 = ~n45349 & ~n45364 ;
  assign n45366 = \a[62]  & ~n45359 ;
  assign n45367 = ~n45356 & n45366 ;
  assign n45368 = \a[62]  & n45359 ;
  assign n45369 = n45356 & n45368 ;
  assign n45370 = ~n45367 & ~n45369 ;
  assign n45371 = n45348 & ~n45370 ;
  assign n45372 = ~n45338 & n45371 ;
  assign n45373 = ~n45365 & ~n45372 ;
  assign n45374 = ~\a[62]  & ~n45349 ;
  assign n45375 = ~n45356 & ~n45359 ;
  assign n45376 = n45356 & n45359 ;
  assign n45377 = ~n45375 & ~n45376 ;
  assign n45378 = \a[62]  & n45348 ;
  assign n45379 = ~n45338 & n45378 ;
  assign n45380 = n45377 & ~n45379 ;
  assign n45381 = ~n45374 & n45380 ;
  assign n45382 = n45373 & ~n45381 ;
  assign n45383 = n45336 & n45382 ;
  assign n45384 = ~n45336 & ~n45382 ;
  assign n45385 = ~n45383 & ~n45384 ;
  assign n45386 = ~n45332 & n45385 ;
  assign n45387 = n45332 & ~n45385 ;
  assign n45388 = ~n45386 & ~n45387 ;
  assign n45389 = n45311 & n45388 ;
  assign n45390 = ~n45311 & ~n45388 ;
  assign n45391 = ~n45389 & ~n45390 ;
  assign n45392 = ~n45306 & n45391 ;
  assign n45393 = ~n45304 & n45392 ;
  assign n45394 = n45306 & n45391 ;
  assign n45395 = n45304 & n45394 ;
  assign n45396 = ~n45393 & ~n45395 ;
  assign n45397 = n45304 & ~n45306 ;
  assign n45398 = ~n45391 & n45397 ;
  assign n45399 = n45306 & ~n45391 ;
  assign n45400 = ~n45304 & n45399 ;
  assign n45401 = ~n45398 & ~n45400 ;
  assign n45402 = n45396 & n45401 ;
  assign n45403 = ~n45171 & ~n45267 ;
  assign n45404 = ~n45173 & ~n45403 ;
  assign n45405 = n45402 & n45404 ;
  assign n45406 = ~n45402 & ~n45404 ;
  assign n45407 = ~n45405 & ~n45406 ;
  assign n45408 = ~n45273 & n45407 ;
  assign n45409 = ~n45285 & n45408 ;
  assign n45410 = ~n45273 & ~n45285 ;
  assign n45411 = ~n45407 & ~n45410 ;
  assign n45412 = ~n45409 & ~n45411 ;
  assign n45413 = ~n45405 & ~n45409 ;
  assign n45414 = n45304 & ~n45391 ;
  assign n45415 = ~n45306 & ~n45391 ;
  assign n45416 = ~n45414 & ~n45415 ;
  assign n45417 = ~n45397 & n45416 ;
  assign n45418 = ~n45311 & ~n45386 ;
  assign n45419 = ~n45387 & ~n45418 ;
  assign n45420 = n18516 & ~n20971 ;
  assign n45421 = ~n20969 & n45420 ;
  assign n45422 = \b[61]  & n18514 ;
  assign n45423 = \a[56]  & \b[60]  ;
  assign n45424 = n19181 & n45423 ;
  assign n45425 = ~\a[57]  & \b[60]  ;
  assign n45426 = n18508 & n45425 ;
  assign n45427 = ~n45424 & ~n45426 ;
  assign n45428 = ~n45422 & n45427 ;
  assign n45429 = \b[59]  & n19183 ;
  assign n45430 = n19180 & n45429 ;
  assign n45431 = \a[59]  & ~n45430 ;
  assign n45432 = n45428 & n45431 ;
  assign n45433 = ~n45421 & n45432 ;
  assign n45434 = n45428 & ~n45430 ;
  assign n45435 = ~n45421 & n45434 ;
  assign n45436 = ~\a[59]  & ~n45435 ;
  assign n45437 = ~n45433 & ~n45436 ;
  assign n45438 = ~n45336 & n45373 ;
  assign n45439 = \a[62]  & n45377 ;
  assign n45440 = ~n45349 & n45439 ;
  assign n45441 = ~\a[62]  & n45377 ;
  assign n45442 = n45349 & n45441 ;
  assign n45443 = ~n45440 & ~n45442 ;
  assign n45444 = ~n45438 & n45443 ;
  assign n45445 = ~n18940 & ~n19861 ;
  assign n45446 = ~n20518 & n45445 ;
  assign n45447 = n18937 & n45446 ;
  assign n45448 = n18940 & ~n19861 ;
  assign n45449 = ~n20518 & n45448 ;
  assign n45450 = ~n18937 & n45449 ;
  assign n45451 = ~n45447 & ~n45450 ;
  assign n45452 = \b[58]  & n20519 ;
  assign n45453 = \a[60]  & \b[57]  ;
  assign n45454 = n20510 & n45453 ;
  assign n45455 = ~n45452 & ~n45454 ;
  assign n45456 = \b[56]  & n21315 ;
  assign n45457 = n21312 & n45456 ;
  assign n45458 = ~\a[60]  & \b[57]  ;
  assign n45459 = n20513 & n45458 ;
  assign n45460 = ~n45457 & ~n45459 ;
  assign n45461 = n45455 & n45460 ;
  assign n45462 = n45451 & n45461 ;
  assign n45463 = n45353 & n45359 ;
  assign n45464 = ~n45355 & ~n45463 ;
  assign n45465 = \b[55]  & n21958 ;
  assign n45466 = \b[54]  & n21957 ;
  assign n45467 = ~n45465 & ~n45466 ;
  assign n45468 = ~n45464 & ~n45467 ;
  assign n45469 = ~n45355 & n45467 ;
  assign n45470 = ~n45463 & n45469 ;
  assign n45471 = ~\a[62]  & ~n45470 ;
  assign n45472 = ~n45468 & n45471 ;
  assign n45473 = ~n45462 & n45472 ;
  assign n45474 = \a[62]  & ~n45470 ;
  assign n45475 = ~n45468 & n45474 ;
  assign n45476 = n45461 & n45475 ;
  assign n45477 = n45451 & n45476 ;
  assign n45478 = ~n45473 & ~n45477 ;
  assign n45479 = ~\a[62]  & ~n45462 ;
  assign n45480 = ~n45468 & ~n45470 ;
  assign n45481 = \a[62]  & n45461 ;
  assign n45482 = n45451 & n45481 ;
  assign n45483 = ~n45480 & ~n45482 ;
  assign n45484 = ~n45479 & n45483 ;
  assign n45485 = n45478 & ~n45484 ;
  assign n45486 = n45444 & n45485 ;
  assign n45487 = ~n45444 & ~n45485 ;
  assign n45488 = ~n45486 & ~n45487 ;
  assign n45489 = n45437 & n45488 ;
  assign n45490 = ~n45437 & ~n45488 ;
  assign n45491 = ~n45489 & ~n45490 ;
  assign n45492 = n45419 & ~n45491 ;
  assign n45493 = ~n45419 & n45491 ;
  assign n45494 = ~n45492 & ~n45493 ;
  assign n45495 = ~n22458 & n37945 ;
  assign n45496 = ~n23173 & n45495 ;
  assign n45497 = \b[62]  & n17308 ;
  assign n45498 = n17305 & n45497 ;
  assign n45499 = \a[54]  & \b[63]  ;
  assign n45500 = n16644 & n45499 ;
  assign n45501 = ~\a[54]  & \b[63]  ;
  assign n45502 = n16647 & n45501 ;
  assign n45503 = \a[56]  & ~n45502 ;
  assign n45504 = ~n45500 & n45503 ;
  assign n45505 = ~n45498 & n45504 ;
  assign n45506 = ~n45496 & n45505 ;
  assign n45507 = ~n45500 & ~n45502 ;
  assign n45508 = ~n45498 & n45507 ;
  assign n45509 = ~n45496 & n45508 ;
  assign n45510 = ~\a[56]  & ~n45509 ;
  assign n45511 = ~n45506 & ~n45510 ;
  assign n45512 = n45494 & ~n45511 ;
  assign n45513 = ~n45494 & n45511 ;
  assign n45514 = ~n45512 & ~n45513 ;
  assign n45515 = n45417 & n45514 ;
  assign n45516 = ~n45417 & ~n45514 ;
  assign n45517 = ~n45515 & ~n45516 ;
  assign n45518 = ~n45413 & n45517 ;
  assign n45519 = ~n45405 & ~n45517 ;
  assign n45520 = ~n45409 & n45519 ;
  assign n45521 = ~n45518 & ~n45520 ;
  assign n45522 = ~n45405 & ~n45515 ;
  assign n45523 = ~n45409 & n45522 ;
  assign n45524 = n45437 & ~n45486 ;
  assign n45525 = n37945 & n39033 ;
  assign n45526 = ~n23171 & n45525 ;
  assign n45527 = \a[53]  & \a[55]  ;
  assign n45528 = \a[54]  & ~\a[56]  ;
  assign n45529 = n45527 & n45528 ;
  assign n45530 = ~\a[53]  & ~\a[55]  ;
  assign n45531 = ~\a[54]  & \a[56]  ;
  assign n45532 = n45530 & n45531 ;
  assign n45533 = ~n45529 & ~n45532 ;
  assign n45534 = \b[63]  & ~n45533 ;
  assign n45535 = \a[56]  & ~n45534 ;
  assign n45536 = ~n45526 & n45535 ;
  assign n45537 = ~n45526 & ~n45534 ;
  assign n45538 = ~\a[56]  & ~n45537 ;
  assign n45539 = ~n45536 & ~n45538 ;
  assign n45540 = ~n45487 & ~n45539 ;
  assign n45541 = ~n45524 & n45540 ;
  assign n45542 = n45487 & n45539 ;
  assign n45543 = ~n45486 & n45539 ;
  assign n45544 = n45437 & n45543 ;
  assign n45545 = ~n45542 & ~n45544 ;
  assign n45546 = ~n45541 & n45545 ;
  assign n45547 = ~n45470 & ~n45477 ;
  assign n45548 = ~n45473 & n45547 ;
  assign n45549 = ~n19550 & n20521 ;
  assign n45550 = ~n19548 & n45549 ;
  assign n45551 = \b[59]  & n20519 ;
  assign n45552 = \a[60]  & \b[58]  ;
  assign n45553 = n20510 & n45552 ;
  assign n45554 = ~n45551 & ~n45553 ;
  assign n45555 = \b[57]  & n21315 ;
  assign n45556 = n21312 & n45555 ;
  assign n45557 = ~\a[60]  & \b[58]  ;
  assign n45558 = n20513 & n45557 ;
  assign n45559 = ~n45556 & ~n45558 ;
  assign n45560 = n45554 & n45559 ;
  assign n45561 = ~n45550 & n45560 ;
  assign n45562 = \b[56]  & n21958 ;
  assign n45563 = \b[55]  & n21957 ;
  assign n45564 = ~n45562 & ~n45563 ;
  assign n45565 = n45467 & ~n45564 ;
  assign n45566 = ~n45467 & n45564 ;
  assign n45567 = ~n45565 & ~n45566 ;
  assign n45568 = ~\a[62]  & n45567 ;
  assign n45569 = ~n45561 & n45568 ;
  assign n45570 = \a[62]  & n45567 ;
  assign n45571 = n45560 & n45570 ;
  assign n45572 = ~n45550 & n45571 ;
  assign n45573 = ~n45569 & ~n45572 ;
  assign n45574 = ~\a[62]  & ~n45561 ;
  assign n45575 = \a[62]  & n45560 ;
  assign n45576 = ~n45550 & n45575 ;
  assign n45577 = ~n45567 & ~n45576 ;
  assign n45578 = ~n45574 & n45577 ;
  assign n45579 = n45573 & ~n45578 ;
  assign n45580 = n45548 & ~n45579 ;
  assign n45581 = ~n45548 & n45579 ;
  assign n45582 = ~n45580 & ~n45581 ;
  assign n45583 = n18516 & n21696 ;
  assign n45584 = ~n21693 & n45583 ;
  assign n45585 = n18516 & n41213 ;
  assign n45586 = ~n21692 & n45585 ;
  assign n45587 = \b[62]  & n18514 ;
  assign n45588 = \a[56]  & \b[61]  ;
  assign n45589 = n19181 & n45588 ;
  assign n45590 = ~\a[57]  & \b[61]  ;
  assign n45591 = n18508 & n45590 ;
  assign n45592 = ~n45589 & ~n45591 ;
  assign n45593 = ~n45587 & n45592 ;
  assign n45594 = \b[60]  & n19183 ;
  assign n45595 = n19180 & n45594 ;
  assign n45596 = \a[59]  & ~n45595 ;
  assign n45597 = n45593 & n45596 ;
  assign n45598 = ~n45586 & n45597 ;
  assign n45599 = ~n45584 & n45598 ;
  assign n45600 = n45593 & ~n45595 ;
  assign n45601 = ~n45586 & n45600 ;
  assign n45602 = ~n45584 & n45601 ;
  assign n45603 = ~\a[59]  & ~n45602 ;
  assign n45604 = ~n45599 & ~n45603 ;
  assign n45605 = n45582 & ~n45604 ;
  assign n45606 = ~n45582 & n45604 ;
  assign n45607 = ~n45605 & ~n45606 ;
  assign n45608 = n45546 & n45607 ;
  assign n45609 = ~n45546 & ~n45607 ;
  assign n45610 = ~n45608 & ~n45609 ;
  assign n45611 = ~n45492 & n45511 ;
  assign n45612 = ~n45493 & ~n45611 ;
  assign n45613 = ~n45610 & ~n45612 ;
  assign n45614 = n45610 & n45612 ;
  assign n45615 = ~n45613 & ~n45614 ;
  assign n45616 = ~n45516 & n45615 ;
  assign n45617 = ~n45523 & n45616 ;
  assign n45618 = ~n45516 & ~n45523 ;
  assign n45619 = ~n45615 & ~n45618 ;
  assign n45620 = ~n45617 & ~n45619 ;
  assign n45621 = ~n45565 & ~n45572 ;
  assign n45622 = ~n45569 & n45621 ;
  assign n45623 = ~\a[56]  & \b[56]  ;
  assign n45624 = n21957 & n45623 ;
  assign n45625 = ~\a[56]  & \b[57]  ;
  assign n45626 = n21958 & n45625 ;
  assign n45627 = ~n45624 & ~n45626 ;
  assign n45628 = \b[57]  & n21958 ;
  assign n45629 = \b[56]  & n21957 ;
  assign n45630 = \a[56]  & ~n45629 ;
  assign n45631 = ~n45628 & n45630 ;
  assign n45632 = n45627 & ~n45631 ;
  assign n45633 = ~n45467 & ~n45632 ;
  assign n45634 = n45467 & n45632 ;
  assign n45635 = ~n45633 & ~n45634 ;
  assign n45636 = ~n45622 & ~n45635 ;
  assign n45637 = n45622 & n45635 ;
  assign n45638 = ~n19861 & ~n20260 ;
  assign n45639 = ~n20518 & n45638 ;
  assign n45640 = n20257 & n45639 ;
  assign n45641 = ~n19861 & n20260 ;
  assign n45642 = ~n20518 & n45641 ;
  assign n45643 = ~n20257 & n45642 ;
  assign n45644 = ~n45640 & ~n45643 ;
  assign n45645 = \b[58]  & n21315 ;
  assign n45646 = n21312 & n45645 ;
  assign n45647 = ~\a[60]  & \b[59]  ;
  assign n45648 = n20513 & n45647 ;
  assign n45649 = ~n45646 & ~n45648 ;
  assign n45650 = \b[60]  & n20519 ;
  assign n45651 = \a[60]  & \b[59]  ;
  assign n45652 = n20510 & n45651 ;
  assign n45653 = \a[62]  & ~n45652 ;
  assign n45654 = ~n45650 & n45653 ;
  assign n45655 = n45649 & n45654 ;
  assign n45656 = n45644 & n45655 ;
  assign n45657 = ~n45650 & ~n45652 ;
  assign n45658 = n45649 & n45657 ;
  assign n45659 = n45644 & n45658 ;
  assign n45660 = ~\a[62]  & ~n45659 ;
  assign n45661 = ~n45656 & ~n45660 ;
  assign n45662 = ~n45637 & ~n45661 ;
  assign n45663 = ~n45636 & n45662 ;
  assign n45664 = ~n45636 & ~n45637 ;
  assign n45665 = n45661 & ~n45664 ;
  assign n45666 = ~n45663 & ~n45665 ;
  assign n45667 = ~n45581 & n45604 ;
  assign n45668 = ~n45580 & ~n45667 ;
  assign n45669 = n18516 & ~n22461 ;
  assign n45670 = ~n22459 & n45669 ;
  assign n45671 = \b[61]  & n19183 ;
  assign n45672 = n19180 & n45671 ;
  assign n45673 = \b[63]  & n18514 ;
  assign n45674 = \a[56]  & \b[62]  ;
  assign n45675 = n19181 & n45674 ;
  assign n45676 = ~\a[57]  & \b[62]  ;
  assign n45677 = n18508 & n45676 ;
  assign n45678 = ~n45675 & ~n45677 ;
  assign n45679 = ~n45673 & n45678 ;
  assign n45680 = ~n45672 & n45679 ;
  assign n45681 = ~\a[59]  & n45680 ;
  assign n45682 = ~n45670 & n45681 ;
  assign n45683 = ~n45670 & n45680 ;
  assign n45684 = \a[59]  & ~n45683 ;
  assign n45685 = ~n45682 & ~n45684 ;
  assign n45686 = ~n45668 & ~n45685 ;
  assign n45687 = n45668 & n45685 ;
  assign n45688 = ~n45686 & ~n45687 ;
  assign n45689 = n45666 & n45688 ;
  assign n45690 = ~n45666 & n45685 ;
  assign n45691 = n45668 & n45690 ;
  assign n45692 = ~n45666 & ~n45668 ;
  assign n45693 = ~n45685 & n45692 ;
  assign n45694 = ~n45691 & ~n45693 ;
  assign n45695 = ~n45689 & n45694 ;
  assign n45696 = ~n45541 & ~n45607 ;
  assign n45697 = n45545 & ~n45696 ;
  assign n45698 = ~n45695 & ~n45697 ;
  assign n45699 = n45695 & n45697 ;
  assign n45700 = ~n45698 & ~n45699 ;
  assign n45701 = n45614 & n45700 ;
  assign n45702 = ~n45614 & ~n45700 ;
  assign n45703 = ~n45701 & ~n45702 ;
  assign n45704 = ~n45617 & n45703 ;
  assign n45705 = ~n45700 & ~n45701 ;
  assign n45706 = n45617 & n45705 ;
  assign n45707 = ~n45704 & ~n45706 ;
  assign n45708 = n45617 & n45700 ;
  assign n45709 = n45686 & ~n45687 ;
  assign n45710 = ~n45666 & ~n45687 ;
  assign n45711 = ~n45709 & ~n45710 ;
  assign n45712 = ~n45636 & ~n45662 ;
  assign n45713 = n20521 & ~n20971 ;
  assign n45714 = ~n20969 & n45713 ;
  assign n45715 = \b[61]  & n20519 ;
  assign n45716 = \a[60]  & \b[60]  ;
  assign n45717 = n20510 & n45716 ;
  assign n45718 = ~n45715 & ~n45717 ;
  assign n45719 = \b[59]  & n21315 ;
  assign n45720 = n21312 & n45719 ;
  assign n45721 = ~\a[60]  & \b[60]  ;
  assign n45722 = n20513 & n45721 ;
  assign n45723 = ~n45720 & ~n45722 ;
  assign n45724 = n45718 & n45723 ;
  assign n45725 = ~n45714 & n45724 ;
  assign n45726 = ~n45467 & ~n45631 ;
  assign n45727 = n45627 & ~n45726 ;
  assign n45728 = \b[58]  & n21958 ;
  assign n45729 = \b[57]  & n21957 ;
  assign n45730 = ~n45728 & ~n45729 ;
  assign n45731 = ~n45727 & n45730 ;
  assign n45732 = n45627 & ~n45730 ;
  assign n45733 = ~n45726 & n45732 ;
  assign n45734 = ~\a[62]  & ~n45733 ;
  assign n45735 = ~n45731 & n45734 ;
  assign n45736 = ~n45725 & n45735 ;
  assign n45737 = \a[62]  & ~n45733 ;
  assign n45738 = ~n45731 & n45737 ;
  assign n45739 = n45724 & n45738 ;
  assign n45740 = ~n45714 & n45739 ;
  assign n45741 = ~n45736 & ~n45740 ;
  assign n45742 = ~\a[62]  & ~n45725 ;
  assign n45743 = ~n45731 & ~n45733 ;
  assign n45744 = \a[62]  & n45724 ;
  assign n45745 = ~n45714 & n45744 ;
  assign n45746 = ~n45743 & ~n45745 ;
  assign n45747 = ~n45742 & n45746 ;
  assign n45748 = n45741 & ~n45747 ;
  assign n45749 = ~n45712 & n45748 ;
  assign n45750 = n45712 & ~n45748 ;
  assign n45751 = ~n45749 & ~n45750 ;
  assign n45752 = n18516 & ~n22458 ;
  assign n45753 = ~n23173 & n45752 ;
  assign n45754 = \b[62]  & n19183 ;
  assign n45755 = n19180 & n45754 ;
  assign n45756 = \a[56]  & \b[63]  ;
  assign n45757 = n19181 & n45756 ;
  assign n45758 = ~\a[57]  & \b[63]  ;
  assign n45759 = n18508 & n45758 ;
  assign n45760 = ~n45757 & ~n45759 ;
  assign n45761 = ~n45755 & n45760 ;
  assign n45762 = ~\a[59]  & n45761 ;
  assign n45763 = ~n45753 & n45762 ;
  assign n45764 = ~n45753 & n45761 ;
  assign n45765 = \a[59]  & ~n45764 ;
  assign n45766 = ~n45763 & ~n45765 ;
  assign n45767 = n45751 & n45766 ;
  assign n45768 = ~n45751 & ~n45766 ;
  assign n45769 = ~n45767 & ~n45768 ;
  assign n45770 = ~n45711 & ~n45769 ;
  assign n45771 = n45711 & n45769 ;
  assign n45772 = ~n45770 & ~n45771 ;
  assign n45773 = ~n45699 & n45772 ;
  assign n45774 = ~n45701 & n45773 ;
  assign n45775 = ~n45708 & n45774 ;
  assign n45776 = ~n45699 & ~n45701 ;
  assign n45777 = ~n45708 & n45776 ;
  assign n45778 = ~n45772 & ~n45777 ;
  assign n45779 = ~n45775 & ~n45778 ;
  assign n45780 = ~n45699 & ~n45771 ;
  assign n45781 = ~n45701 & n45780 ;
  assign n45782 = ~n45708 & n45781 ;
  assign n45783 = ~n45731 & ~n45740 ;
  assign n45784 = ~n45736 & n45783 ;
  assign n45785 = \b[59]  & n21958 ;
  assign n45786 = \b[58]  & n21957 ;
  assign n45787 = ~n45785 & ~n45786 ;
  assign n45788 = n45730 & ~n45787 ;
  assign n45789 = ~n45730 & n45787 ;
  assign n45790 = ~n45788 & ~n45789 ;
  assign n45791 = n45784 & n45790 ;
  assign n45792 = ~n45784 & ~n45790 ;
  assign n45793 = ~n45791 & ~n45792 ;
  assign n45794 = n20521 & n21696 ;
  assign n45795 = ~n21693 & n45794 ;
  assign n45796 = n20521 & n41213 ;
  assign n45797 = ~n21692 & n45796 ;
  assign n45798 = \b[60]  & n21315 ;
  assign n45799 = n21312 & n45798 ;
  assign n45800 = ~\a[60]  & \b[61]  ;
  assign n45801 = n20513 & n45800 ;
  assign n45802 = ~n45799 & ~n45801 ;
  assign n45803 = \b[62]  & n20519 ;
  assign n45804 = \a[60]  & \b[61]  ;
  assign n45805 = n20510 & n45804 ;
  assign n45806 = \a[62]  & ~n45805 ;
  assign n45807 = ~n45803 & n45806 ;
  assign n45808 = n45802 & n45807 ;
  assign n45809 = ~n45797 & n45808 ;
  assign n45810 = ~n45795 & n45809 ;
  assign n45811 = ~n45803 & ~n45805 ;
  assign n45812 = n45802 & n45811 ;
  assign n45813 = ~n45797 & n45812 ;
  assign n45814 = ~n45795 & n45813 ;
  assign n45815 = ~\a[62]  & ~n45814 ;
  assign n45816 = ~n45810 & ~n45815 ;
  assign n45817 = n18516 & n39033 ;
  assign n45818 = ~n23171 & n45817 ;
  assign n45819 = \a[56]  & \a[58]  ;
  assign n45820 = \a[57]  & ~\a[59]  ;
  assign n45821 = n45819 & n45820 ;
  assign n45822 = ~\a[56]  & ~\a[58]  ;
  assign n45823 = ~\a[57]  & \a[59]  ;
  assign n45824 = n45822 & n45823 ;
  assign n45825 = ~n45821 & ~n45824 ;
  assign n45826 = \b[63]  & ~n45825 ;
  assign n45827 = \a[59]  & ~n45826 ;
  assign n45828 = ~n45818 & n45827 ;
  assign n45829 = ~n45818 & ~n45826 ;
  assign n45830 = ~\a[59]  & ~n45829 ;
  assign n45831 = ~n45828 & ~n45830 ;
  assign n45832 = ~n45816 & ~n45831 ;
  assign n45833 = n45816 & n45831 ;
  assign n45834 = ~n45832 & ~n45833 ;
  assign n45835 = ~n45793 & n45834 ;
  assign n45836 = n45793 & ~n45834 ;
  assign n45837 = ~n45835 & ~n45836 ;
  assign n45838 = ~n45749 & ~n45766 ;
  assign n45839 = ~n45750 & ~n45838 ;
  assign n45840 = n45837 & n45839 ;
  assign n45841 = ~n45837 & ~n45839 ;
  assign n45842 = ~n45840 & ~n45841 ;
  assign n45843 = ~n45770 & n45842 ;
  assign n45844 = ~n45782 & n45843 ;
  assign n45845 = ~n45770 & ~n45782 ;
  assign n45846 = ~n45842 & ~n45845 ;
  assign n45847 = ~n45844 & ~n45846 ;
  assign n45848 = ~n45840 & ~n45844 ;
  assign n45849 = ~n45832 & ~n45835 ;
  assign n45850 = ~n45731 & ~n45789 ;
  assign n45851 = ~n45740 & n45850 ;
  assign n45852 = ~n45736 & n45851 ;
  assign n45853 = ~n45788 & ~n45852 ;
  assign n45854 = n20521 & ~n22461 ;
  assign n45855 = ~n22459 & n45854 ;
  assign n45856 = \b[63]  & n20519 ;
  assign n45857 = \a[60]  & \b[62]  ;
  assign n45858 = n20510 & n45857 ;
  assign n45859 = ~n45856 & ~n45858 ;
  assign n45860 = \b[61]  & n21315 ;
  assign n45861 = n21312 & n45860 ;
  assign n45862 = ~\a[60]  & \b[62]  ;
  assign n45863 = n20513 & n45862 ;
  assign n45864 = ~n45861 & ~n45863 ;
  assign n45865 = n45859 & n45864 ;
  assign n45866 = ~n45855 & n45865 ;
  assign n45867 = ~\a[59]  & n45786 ;
  assign n45868 = ~\a[59]  & \b[59]  ;
  assign n45869 = n21958 & n45868 ;
  assign n45870 = ~n45867 & ~n45869 ;
  assign n45871 = \a[59]  & ~n45786 ;
  assign n45872 = ~n45785 & n45871 ;
  assign n45873 = n45870 & ~n45872 ;
  assign n45874 = \b[60]  & n21958 ;
  assign n45875 = \b[59]  & n21957 ;
  assign n45876 = ~n45874 & ~n45875 ;
  assign n45877 = ~\a[62]  & ~n45876 ;
  assign n45878 = ~n45873 & n45877 ;
  assign n45879 = ~\a[62]  & n45876 ;
  assign n45880 = n45873 & n45879 ;
  assign n45881 = ~n45878 & ~n45880 ;
  assign n45882 = ~n45866 & ~n45881 ;
  assign n45883 = \a[62]  & ~n45876 ;
  assign n45884 = ~n45873 & n45883 ;
  assign n45885 = \a[62]  & n45876 ;
  assign n45886 = n45873 & n45885 ;
  assign n45887 = ~n45884 & ~n45886 ;
  assign n45888 = n45865 & ~n45887 ;
  assign n45889 = ~n45855 & n45888 ;
  assign n45890 = ~n45882 & ~n45889 ;
  assign n45891 = ~\a[62]  & ~n45866 ;
  assign n45892 = ~n45873 & ~n45876 ;
  assign n45893 = n45873 & n45876 ;
  assign n45894 = ~n45892 & ~n45893 ;
  assign n45895 = \a[62]  & n45865 ;
  assign n45896 = ~n45855 & n45895 ;
  assign n45897 = n45894 & ~n45896 ;
  assign n45898 = ~n45891 & n45897 ;
  assign n45899 = n45890 & ~n45898 ;
  assign n45900 = n45853 & n45899 ;
  assign n45901 = ~n45853 & ~n45899 ;
  assign n45902 = ~n45900 & ~n45901 ;
  assign n45903 = ~n45849 & n45902 ;
  assign n45904 = n45849 & ~n45902 ;
  assign n45905 = ~n45903 & ~n45904 ;
  assign n45906 = ~n45848 & n45905 ;
  assign n45907 = ~n45840 & ~n45905 ;
  assign n45908 = ~n45844 & n45907 ;
  assign n45909 = ~n45906 & ~n45908 ;
  assign n45910 = ~n45840 & ~n45903 ;
  assign n45911 = ~n45844 & n45910 ;
  assign n45912 = ~n45853 & n45890 ;
  assign n45913 = \a[62]  & n45894 ;
  assign n45914 = ~n45866 & n45913 ;
  assign n45915 = ~\a[62]  & n45894 ;
  assign n45916 = n45866 & n45915 ;
  assign n45917 = ~n45914 & ~n45916 ;
  assign n45918 = n20521 & ~n22458 ;
  assign n45919 = ~n23173 & n45918 ;
  assign n45920 = \b[62]  & n21315 ;
  assign n45921 = n21312 & n45920 ;
  assign n45922 = ~\a[60]  & \b[63]  ;
  assign n45923 = n20513 & n45922 ;
  assign n45924 = \a[60]  & \b[63]  ;
  assign n45925 = n20510 & n45924 ;
  assign n45926 = ~n45923 & ~n45925 ;
  assign n45927 = ~n45921 & n45926 ;
  assign n45928 = ~n45919 & n45927 ;
  assign n45929 = n45870 & n45876 ;
  assign n45930 = ~n45872 & ~n45929 ;
  assign n45931 = \b[61]  & n21958 ;
  assign n45932 = \b[60]  & n21957 ;
  assign n45933 = ~n45931 & ~n45932 ;
  assign n45934 = ~n45930 & ~n45933 ;
  assign n45935 = ~n45872 & n45933 ;
  assign n45936 = ~n45929 & n45935 ;
  assign n45937 = ~\a[62]  & ~n45936 ;
  assign n45938 = ~n45934 & n45937 ;
  assign n45939 = ~n45928 & n45938 ;
  assign n45940 = \a[62]  & ~n45936 ;
  assign n45941 = ~n45934 & n45940 ;
  assign n45942 = n45927 & n45941 ;
  assign n45943 = ~n45919 & n45942 ;
  assign n45944 = ~n45939 & ~n45943 ;
  assign n45945 = ~\a[62]  & ~n45928 ;
  assign n45946 = ~n45934 & ~n45936 ;
  assign n45947 = \a[62]  & n45927 ;
  assign n45948 = ~n45919 & n45947 ;
  assign n45949 = ~n45946 & ~n45948 ;
  assign n45950 = ~n45945 & n45949 ;
  assign n45951 = n45944 & ~n45950 ;
  assign n45952 = n45917 & n45951 ;
  assign n45953 = ~n45912 & n45952 ;
  assign n45954 = ~n45912 & n45917 ;
  assign n45955 = ~n45951 & ~n45954 ;
  assign n45956 = ~n45953 & ~n45955 ;
  assign n45957 = ~n45904 & n45956 ;
  assign n45958 = ~n45911 & n45957 ;
  assign n45959 = ~n45904 & ~n45911 ;
  assign n45960 = ~n45956 & ~n45959 ;
  assign n45961 = ~n45958 & ~n45960 ;
  assign n45962 = ~n45936 & ~n45943 ;
  assign n45963 = ~n45939 & n45962 ;
  assign n45964 = n20521 & n39033 ;
  assign n45965 = ~n23171 & n45964 ;
  assign n45966 = \a[59]  & \a[61]  ;
  assign n45967 = \a[60]  & ~\a[62]  ;
  assign n45968 = n45966 & n45967 ;
  assign n45969 = ~\a[59]  & ~\a[61]  ;
  assign n45970 = ~\a[60]  & \a[62]  ;
  assign n45971 = n45969 & n45970 ;
  assign n45972 = ~n45968 & ~n45971 ;
  assign n45973 = \b[63]  & ~n45972 ;
  assign n45974 = \b[62]  & n21958 ;
  assign n45975 = \b[61]  & n21957 ;
  assign n45976 = ~n45974 & ~n45975 ;
  assign n45977 = n45933 & ~n45976 ;
  assign n45978 = ~n45933 & n45976 ;
  assign n45979 = ~n45977 & ~n45978 ;
  assign n45980 = \a[62]  & n45979 ;
  assign n45981 = ~n45973 & n45980 ;
  assign n45982 = ~n45965 & n45981 ;
  assign n45983 = ~n45965 & ~n45973 ;
  assign n45984 = ~\a[62]  & n45979 ;
  assign n45985 = ~n45983 & n45984 ;
  assign n45986 = ~n45982 & ~n45985 ;
  assign n45987 = ~\a[62]  & ~n45973 ;
  assign n45988 = ~n45979 & n45987 ;
  assign n45989 = ~n45965 & n45988 ;
  assign n45990 = \a[62]  & ~n45979 ;
  assign n45991 = ~n45983 & n45990 ;
  assign n45992 = ~n45989 & ~n45991 ;
  assign n45993 = n45986 & n45992 ;
  assign n45994 = ~n45963 & n45993 ;
  assign n45995 = n45963 & ~n45993 ;
  assign n45996 = ~n45994 & ~n45995 ;
  assign n45997 = ~n45953 & n45996 ;
  assign n45998 = ~n45958 & n45997 ;
  assign n45999 = ~n45953 & ~n45958 ;
  assign n46000 = ~n45996 & ~n45999 ;
  assign n46001 = ~n45998 & ~n46000 ;
  assign n46002 = ~n45953 & ~n45994 ;
  assign n46003 = ~n45958 & n46002 ;
  assign n46004 = ~n45977 & ~n45982 ;
  assign n46005 = ~n45985 & n46004 ;
  assign n46006 = \a[63]  & \b[63]  ;
  assign n46007 = \a[62]  & ~\b[63]  ;
  assign n46008 = ~n46006 & ~n46007 ;
  assign n46009 = \b[62]  & n21957 ;
  assign n46010 = ~n46008 & ~n46009 ;
  assign n46011 = ~n45933 & ~n46010 ;
  assign n46012 = n45933 & n46010 ;
  assign n46013 = ~n46011 & ~n46012 ;
  assign n46014 = n46005 & n46013 ;
  assign n46015 = ~n46005 & ~n46013 ;
  assign n46016 = ~n46014 & ~n46015 ;
  assign n46017 = ~n45995 & ~n46016 ;
  assign n46018 = ~n46003 & n46017 ;
  assign n46019 = ~n45995 & ~n46003 ;
  assign n46020 = n46016 & ~n46019 ;
  assign n46021 = ~n46018 & ~n46020 ;
  assign n46022 = \a[62]  & n46006 ;
  assign n46023 = ~n46010 & n46022 ;
  assign n46024 = ~n45933 & n46023 ;
  assign n46025 = ~n46006 & n46007 ;
  assign n46026 = ~n46009 & n46025 ;
  assign n46027 = ~n45932 & ~n46006 ;
  assign n46028 = ~n45931 & n46027 ;
  assign n46029 = ~n46026 & ~n46028 ;
  assign n46030 = ~n46024 & n46029 ;
  assign n46031 = ~n46005 & n46013 ;
  assign n46032 = n46030 & ~n46031 ;
  assign n46033 = ~n46018 & n46032 ;
  assign n46034 = ~n46018 & ~n46031 ;
  assign n46035 = ~n46030 & ~n46034 ;
  assign n46036 = ~n46033 & ~n46035 ;
  assign \f[0]  = n129 ;
  assign \f[1]  = n149 ;
  assign \f[2]  = n169 ;
  assign \f[3]  = n209 ;
  assign \f[4]  = n265 ;
  assign \f[5]  = n316 ;
  assign \f[6]  = n373 ;
  assign \f[7]  = n449 ;
  assign \f[8]  = n528 ;
  assign \f[9]  = n609 ;
  assign \f[10]  = n718 ;
  assign \f[11]  = n821 ;
  assign \f[12]  = n940 ;
  assign \f[13]  = n1076 ;
  assign \f[14]  = n1220 ;
  assign \f[15]  = n1369 ;
  assign \f[16]  = n1543 ;
  assign \f[17]  = n1723 ;
  assign \f[18]  = n1903 ;
  assign \f[19]  = n2108 ;
  assign \f[20]  = n2325 ;
  assign \f[21]  = n2552 ;
  assign \f[22]  = n2799 ;
  assign \f[23]  = n3051 ;
  assign \f[24]  = n3315 ;
  assign \f[25]  = n3595 ;
  assign \f[26]  = n3874 ;
  assign \f[27]  = n4177 ;
  assign \f[28]  = n4489 ;
  assign \f[29]  = n4802 ;
  assign \f[30]  = n5135 ;
  assign \f[31]  = n5491 ;
  assign \f[32]  = n5842 ;
  assign \f[33]  = n6205 ;
  assign \f[34]  = n6597 ;
  assign \f[35]  = n6970 ;
  assign \f[36]  = n7367 ;
  assign \f[37]  = n7790 ;
  assign \f[38]  = n8205 ;
  assign \f[39]  = n8631 ;
  assign \f[40]  = n9076 ;
  assign \f[41]  = n9511 ;
  assign \f[42]  = n9962 ;
  assign \f[43]  = n10439 ;
  assign \f[44]  = n10919 ;
  assign \f[45]  = n11425 ;
  assign \f[46]  = n11939 ;
  assign \f[47]  = n12467 ;
  assign \f[48]  = n12994 ;
  assign \f[49]  = n13553 ;
  assign \f[50]  = n14085 ;
  assign \f[51]  = n14653 ;
  assign \f[52]  = n15233 ;
  assign \f[53]  = n15823 ;
  assign \f[54]  = n16435 ;
  assign \f[55]  = n17060 ;
  assign \f[56]  = n17677 ;
  assign \f[57]  = n18326 ;
  assign \f[58]  = n18970 ;
  assign \f[59]  = n19652 ;
  assign \f[60]  = n20332 ;
  assign \f[61]  = n21057 ;
  assign \f[62]  = n21775 ;
  assign \f[63]  = ~n22487 ;
  assign \f[64]  = n23236 ;
  assign \f[65]  = n23994 ;
  assign \f[66]  = ~n24727 ;
  assign \f[67]  = n25436 ;
  assign \f[68]  = n26094 ;
  assign \f[69]  = n26847 ;
  assign \f[70]  = n27506 ;
  assign \f[71]  = n28134 ;
  assign \f[72]  = n28804 ;
  assign \f[73]  = n29429 ;
  assign \f[74]  = n30024 ;
  assign \f[75]  = n30680 ;
  assign \f[76]  = n31261 ;
  assign \f[77]  = n31829 ;
  assign \f[78]  = n32406 ;
  assign \f[79]  = ~n32947 ;
  assign \f[80]  = n33494 ;
  assign \f[81]  = n34013 ;
  assign \f[82]  = n34510 ;
  assign \f[83]  = n35019 ;
  assign \f[84]  = n35527 ;
  assign \f[85]  = ~n36003 ;
  assign \f[86]  = ~n36479 ;
  assign \f[87]  = n36932 ;
  assign \f[88]  = n37381 ;
  assign \f[89]  = n37814 ;
  assign \f[90]  = n38236 ;
  assign \f[91]  = ~n38646 ;
  assign \f[92]  = n39062 ;
  assign \f[93]  = n39459 ;
  assign \f[94]  = n39822 ;
  assign \f[95]  = n40210 ;
  assign \f[96]  = n40575 ;
  assign \f[97]  = n40906 ;
  assign \f[98]  = n41256 ;
  assign \f[99]  = n41595 ;
  assign \f[100]  = n41899 ;
  assign \f[101]  = n42194 ;
  assign \f[102]  = n42485 ;
  assign \f[103]  = n42745 ;
  assign \f[104]  = ~n43012 ;
  assign \f[105]  = n43283 ;
  assign \f[106]  = n43517 ;
  assign \f[107]  = ~n43750 ;
  assign \f[108]  = n43968 ;
  assign \f[109]  = n44164 ;
  assign \f[110]  = ~n44361 ;
  assign \f[111]  = n44545 ;
  assign \f[112]  = ~n44715 ;
  assign \f[113]  = ~n44887 ;
  assign \f[114]  = n45027 ;
  assign \f[115]  = ~n45152 ;
  assign \f[116]  = ~n45282 ;
  assign \f[117]  = n45412 ;
  assign \f[118]  = n45521 ;
  assign \f[119]  = n45620 ;
  assign \f[120]  = ~n45707 ;
  assign \f[121]  = ~n45779 ;
  assign \f[122]  = n45847 ;
  assign \f[123]  = n45909 ;
  assign \f[124]  = n45961 ;
  assign \f[125]  = ~n46001 ;
  assign \f[126]  = n46021 ;
  assign \f[127]  = n46036 ;
endmodule
