module top( \totalcoeffs[0]  , \totalcoeffs[1]  , \totalcoeffs[2]  , \totalcoeffs[3]  , \totalcoeffs[4]  , \ctable[0]  , \ctable[1]  , \ctable[2]  , \trailingones[0]  , \trailingones[1]  , \coeff_token[0]  , \coeff_token[1]  , \coeff_token[2]  , \coeff_token[3]  , \coeff_token[4]  , \coeff_token[5]  , \ctoken_len[0]  , \ctoken_len[1]  , \ctoken_len[2]  , \ctoken_len[3]  , \ctoken_len[4]  );
  input \totalcoeffs[0]  ;
  input \totalcoeffs[1]  ;
  input \totalcoeffs[2]  ;
  input \totalcoeffs[3]  ;
  input \totalcoeffs[4]  ;
  input \ctable[0]  ;
  input \ctable[1]  ;
  input \ctable[2]  ;
  input \trailingones[0]  ;
  input \trailingones[1]  ;
  output \coeff_token[0]  ;
  output \coeff_token[1]  ;
  output \coeff_token[2]  ;
  output \coeff_token[3]  ;
  output \coeff_token[4]  ;
  output \coeff_token[5]  ;
  output \ctoken_len[0]  ;
  output \ctoken_len[1]  ;
  output \ctoken_len[2]  ;
  output \ctoken_len[3]  ;
  output \ctoken_len[4]  ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 ;
  assign n11 = ~\totalcoeffs[0]  & ~\totalcoeffs[1]  ;
  assign n12 = \totalcoeffs[2]  & ~\trailingones[1]  ;
  assign n13 = n11 & n12 ;
  assign n14 = ~\ctable[0]  & \ctable[2]  ;
  assign n15 = ~\totalcoeffs[3]  & \trailingones[0]  ;
  assign n16 = n14 & n15 ;
  assign n17 = n13 & n16 ;
  assign n18 = ~\ctable[2]  & ~\trailingones[0]  ;
  assign n19 = ~\totalcoeffs[0]  & \ctable[0]  ;
  assign n20 = ~\trailingones[1]  & n19 ;
  assign n21 = \totalcoeffs[0]  & ~\totalcoeffs[1]  ;
  assign n22 = n12 & ~n21 ;
  assign n23 = ~n20 & ~n22 ;
  assign n24 = ~\totalcoeffs[1]  & \trailingones[1]  ;
  assign n25 = ~\totalcoeffs[2]  & ~\totalcoeffs[3]  ;
  assign n26 = n24 & ~n25 ;
  assign n27 = \totalcoeffs[0]  & \totalcoeffs[3]  ;
  assign n28 = ~\totalcoeffs[1]  & n27 ;
  assign n29 = \totalcoeffs[1]  & ~\totalcoeffs[3]  ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = ~n26 & n30 ;
  assign n32 = n23 & n31 ;
  assign n33 = n18 & ~n32 ;
  assign n34 = ~\ctable[2]  & \trailingones[1]  ;
  assign n35 = \totalcoeffs[1]  & n34 ;
  assign n36 = \totalcoeffs[1]  & \trailingones[0]  ;
  assign n37 = n14 & n36 ;
  assign n38 = ~n35 & ~n37 ;
  assign n39 = \totalcoeffs[1]  & ~\ctable[2]  ;
  assign n40 = ~\ctable[0]  & ~\trailingones[1]  ;
  assign n41 = ~n39 & n40 ;
  assign n42 = n38 & ~n41 ;
  assign n43 = \totalcoeffs[0]  & ~\totalcoeffs[2]  ;
  assign n44 = ~\totalcoeffs[3]  & n43 ;
  assign n45 = ~n42 & n44 ;
  assign n46 = ~\totalcoeffs[0]  & \trailingones[1]  ;
  assign n47 = \totalcoeffs[1]  & ~n46 ;
  assign n48 = ~\totalcoeffs[3]  & ~\ctable[0]  ;
  assign n49 = ~n24 & n48 ;
  assign n50 = ~n47 & n49 ;
  assign n51 = \totalcoeffs[0]  & ~\trailingones[1]  ;
  assign n52 = ~\totalcoeffs[1]  & ~n51 ;
  assign n53 = \totalcoeffs[1]  & ~\trailingones[1]  ;
  assign n54 = ~\ctable[2]  & ~n53 ;
  assign n55 = ~n52 & n54 ;
  assign n56 = ~n50 & ~n55 ;
  assign n57 = ~\totalcoeffs[2]  & ~\trailingones[0]  ;
  assign n58 = ~n56 & n57 ;
  assign n59 = ~n45 & ~n58 ;
  assign n60 = ~n33 & n59 ;
  assign n61 = ~n17 & n60 ;
  assign n62 = ~\ctable[1]  & ~n61 ;
  assign n63 = ~n46 & ~n51 ;
  assign n64 = \totalcoeffs[1]  & \ctable[0]  ;
  assign n65 = \totalcoeffs[2]  & \totalcoeffs[3]  ;
  assign n66 = n64 & n65 ;
  assign n67 = n63 & n66 ;
  assign n68 = ~\totalcoeffs[0]  & ~\totalcoeffs[2]  ;
  assign n69 = n24 & n68 ;
  assign n70 = ~\ctable[0]  & ~n69 ;
  assign n71 = \totalcoeffs[3]  & \ctable[1]  ;
  assign n72 = ~n70 & n71 ;
  assign n73 = ~n67 & ~n72 ;
  assign n74 = ~\totalcoeffs[0]  & ~\totalcoeffs[3]  ;
  assign n75 = \totalcoeffs[2]  & \trailingones[1]  ;
  assign n76 = \ctable[1]  & n75 ;
  assign n77 = ~\totalcoeffs[2]  & \ctable[1]  ;
  assign n78 = n53 & n77 ;
  assign n79 = ~n76 & ~n78 ;
  assign n80 = n74 & ~n79 ;
  assign n81 = ~\totalcoeffs[2]  & ~n51 ;
  assign n82 = n29 & ~n46 ;
  assign n83 = n81 & ~n82 ;
  assign n84 = \ctable[0]  & \ctable[1]  ;
  assign n85 = ~\totalcoeffs[2]  & \ctable[0]  ;
  assign n86 = ~n51 & n85 ;
  assign n87 = ~n84 & ~n86 ;
  assign n88 = ~n83 & ~n87 ;
  assign n89 = ~n80 & ~n88 ;
  assign n90 = n73 & n89 ;
  assign n91 = \trailingones[0]  & ~n90 ;
  assign n92 = ~\totalcoeffs[1]  & ~\trailingones[1]  ;
  assign n93 = ~\trailingones[0]  & n92 ;
  assign n94 = ~\totalcoeffs[3]  & n68 ;
  assign n95 = n93 & n94 ;
  assign n96 = \ctable[0]  & ~n95 ;
  assign n97 = \totalcoeffs[3]  & n12 ;
  assign n98 = n21 & n97 ;
  assign n99 = ~\totalcoeffs[1]  & ~n46 ;
  assign n100 = \totalcoeffs[3]  & ~\trailingones[0]  ;
  assign n101 = ~n99 & n100 ;
  assign n102 = ~n98 & ~n101 ;
  assign n103 = \totalcoeffs[1]  & ~\trailingones[0]  ;
  assign n104 = \totalcoeffs[2]  & ~\totalcoeffs[3]  ;
  assign n105 = n24 & n104 ;
  assign n106 = ~n103 & ~n105 ;
  assign n107 = ~\totalcoeffs[0]  & ~n106 ;
  assign n108 = n102 & ~n107 ;
  assign n109 = ~\trailingones[0]  & n75 ;
  assign n110 = \totalcoeffs[3]  & ~n77 ;
  assign n111 = n93 & ~n110 ;
  assign n112 = ~n109 & ~n111 ;
  assign n113 = ~n95 & n112 ;
  assign n114 = n108 & n113 ;
  assign n115 = ~n96 & ~n114 ;
  assign n116 = ~n91 & ~n115 ;
  assign n117 = ~\ctable[2]  & ~n116 ;
  assign n118 = ~n62 & ~n117 ;
  assign n119 = ~\totalcoeffs[4]  & ~n118 ;
  assign n120 = ~\ctable[1]  & \trailingones[0]  ;
  assign n121 = \ctable[0]  & ~n120 ;
  assign n122 = \totalcoeffs[4]  & \trailingones[0]  ;
  assign n123 = ~\ctable[1]  & ~\trailingones[1]  ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = n121 & ~n124 ;
  assign n126 = \ctable[1]  & ~\trailingones[1]  ;
  assign n127 = \totalcoeffs[4]  & \trailingones[1]  ;
  assign n128 = ~n126 & ~n127 ;
  assign n129 = ~\trailingones[0]  & ~n84 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = ~n125 & ~n130 ;
  assign n132 = ~\totalcoeffs[1]  & ~\totalcoeffs[3]  ;
  assign n133 = ~\ctable[2]  & n68 ;
  assign n134 = n132 & n133 ;
  assign n135 = ~n131 & n134 ;
  assign n136 = ~n119 & ~n135 ;
  assign n137 = \totalcoeffs[1]  & \totalcoeffs[2]  ;
  assign n138 = \totalcoeffs[3]  & n137 ;
  assign n139 = \totalcoeffs[3]  & \ctable[0]  ;
  assign n140 = \totalcoeffs[2]  & \ctable[0]  ;
  assign n141 = ~n139 & ~n140 ;
  assign n142 = ~n138 & n141 ;
  assign n143 = \ctable[1]  & ~n142 ;
  assign n144 = ~\totalcoeffs[1]  & \totalcoeffs[3]  ;
  assign n145 = n57 & n144 ;
  assign n146 = ~n64 & ~n145 ;
  assign n147 = \totalcoeffs[0]  & \ctable[1]  ;
  assign n148 = ~n146 & n147 ;
  assign n149 = ~n143 & ~n148 ;
  assign n150 = \ctable[0]  & ~\trailingones[0]  ;
  assign n151 = n138 & n150 ;
  assign n152 = \trailingones[1]  & ~n151 ;
  assign n153 = n149 & n152 ;
  assign n154 = ~\totalcoeffs[4]  & ~n153 ;
  assign n155 = ~\totalcoeffs[1]  & ~\trailingones[0]  ;
  assign n156 = ~\totalcoeffs[2]  & ~n155 ;
  assign n157 = ~\totalcoeffs[1]  & \trailingones[0]  ;
  assign n158 = \ctable[1]  & n157 ;
  assign n159 = ~n156 & ~n158 ;
  assign n160 = \totalcoeffs[3]  & ~\ctable[0]  ;
  assign n161 = ~n159 & n160 ;
  assign n162 = \totalcoeffs[0]  & \totalcoeffs[1]  ;
  assign n163 = ~\totalcoeffs[1]  & ~\ctable[1]  ;
  assign n164 = ~n162 & ~n163 ;
  assign n165 = ~\totalcoeffs[0]  & \trailingones[0]  ;
  assign n166 = ~\totalcoeffs[2]  & ~\ctable[0]  ;
  assign n167 = ~n165 & n166 ;
  assign n168 = n164 & n167 ;
  assign n169 = ~\trailingones[1]  & ~n168 ;
  assign n170 = ~n161 & n169 ;
  assign n171 = ~\ctable[2]  & ~n170 ;
  assign n172 = ~\totalcoeffs[2]  & \trailingones[0]  ;
  assign n173 = \totalcoeffs[0]  & n172 ;
  assign n174 = \totalcoeffs[0]  & ~\ctable[0]  ;
  assign n175 = ~n19 & ~n174 ;
  assign n176 = ~n173 & n175 ;
  assign n177 = \totalcoeffs[1]  & ~n176 ;
  assign n178 = ~\totalcoeffs[1]  & \ctable[0]  ;
  assign n179 = n57 & n178 ;
  assign n180 = ~\ctable[0]  & \trailingones[0]  ;
  assign n181 = ~\totalcoeffs[3]  & ~\trailingones[0]  ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = n21 & n182 ;
  assign n184 = ~n179 & ~n183 ;
  assign n185 = \totalcoeffs[3]  & \trailingones[0]  ;
  assign n186 = ~\totalcoeffs[2]  & ~n185 ;
  assign n187 = ~\totalcoeffs[0]  & ~n186 ;
  assign n188 = n184 & ~n187 ;
  assign n189 = ~n177 & n188 ;
  assign n190 = ~\ctable[1]  & ~\ctable[2]  ;
  assign n191 = ~n189 & n190 ;
  assign n192 = ~n171 & ~n191 ;
  assign n193 = n154 & ~n192 ;
  assign n194 = n12 & n120 ;
  assign n195 = ~\totalcoeffs[1]  & ~n194 ;
  assign n196 = ~\totalcoeffs[0]  & \ctable[1]  ;
  assign n197 = ~\totalcoeffs[2]  & ~n196 ;
  assign n198 = ~\trailingones[1]  & n180 ;
  assign n199 = ~n197 & n198 ;
  assign n200 = ~\ctable[1]  & ~\trailingones[0]  ;
  assign n201 = ~\trailingones[1]  & n200 ;
  assign n202 = ~n194 & ~n201 ;
  assign n203 = ~n199 & n202 ;
  assign n204 = ~n195 & ~n203 ;
  assign n205 = ~n122 & ~n150 ;
  assign n206 = ~\ctable[1]  & ~n205 ;
  assign n207 = ~n127 & ~n206 ;
  assign n208 = ~\ctable[1]  & \trailingones[1]  ;
  assign n209 = ~\totalcoeffs[2]  & n11 ;
  assign n210 = ~n208 & n209 ;
  assign n211 = ~n207 & n210 ;
  assign n212 = ~\totalcoeffs[2]  & ~\trailingones[1]  ;
  assign n213 = ~\totalcoeffs[0]  & ~\trailingones[0]  ;
  assign n214 = n212 & n213 ;
  assign n215 = \totalcoeffs[0]  & \trailingones[0]  ;
  assign n216 = n75 & n215 ;
  assign n217 = ~n214 & ~n216 ;
  assign n218 = n178 & ~n217 ;
  assign n219 = ~n211 & ~n218 ;
  assign n220 = ~\trailingones[0]  & \trailingones[1]  ;
  assign n221 = n19 & n220 ;
  assign n222 = \ctable[1]  & \trailingones[1]  ;
  assign n223 = ~n180 & ~n222 ;
  assign n224 = \ctable[1]  & \trailingones[0]  ;
  assign n225 = \totalcoeffs[0]  & ~n224 ;
  assign n226 = ~n223 & n225 ;
  assign n227 = ~n221 & ~n226 ;
  assign n228 = \totalcoeffs[1]  & ~\totalcoeffs[2]  ;
  assign n229 = ~n227 & n228 ;
  assign n230 = ~\totalcoeffs[0]  & ~n223 ;
  assign n231 = ~\trailingones[0]  & ~\trailingones[1]  ;
  assign n232 = \trailingones[0]  & \trailingones[1]  ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = ~n150 & ~n208 ;
  assign n235 = ~n233 & n234 ;
  assign n236 = ~n230 & ~n235 ;
  assign n237 = ~\totalcoeffs[1]  & \totalcoeffs[2]  ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ~n229 & ~n238 ;
  assign n240 = n219 & n239 ;
  assign n241 = ~n204 & n240 ;
  assign n242 = \totalcoeffs[4]  & ~n210 ;
  assign n243 = \totalcoeffs[4]  & ~\trailingones[1]  ;
  assign n244 = ~n206 & n243 ;
  assign n245 = ~n242 & ~n244 ;
  assign n246 = ~\totalcoeffs[3]  & ~\ctable[2]  ;
  assign n247 = n245 & n246 ;
  assign n248 = ~n241 & n247 ;
  assign n249 = ~n193 & ~n248 ;
  assign n250 = n81 & ~n162 ;
  assign n251 = \totalcoeffs[2]  & ~n11 ;
  assign n252 = ~\trailingones[0]  & ~n251 ;
  assign n253 = ~n250 & n252 ;
  assign n254 = n53 & n172 ;
  assign n255 = ~n13 & ~n254 ;
  assign n256 = ~n253 & n255 ;
  assign n257 = ~\ctable[2]  & ~n13 ;
  assign n258 = ~\totalcoeffs[4]  & ~\ctable[1]  ;
  assign n259 = n48 & n258 ;
  assign n260 = ~n257 & n259 ;
  assign n261 = ~n256 & n260 ;
  assign n262 = n249 & ~n261 ;
  assign n263 = ~\totalcoeffs[2]  & \trailingones[1]  ;
  assign n264 = ~n36 & n77 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = ~\trailingones[0]  & n24 ;
  assign n267 = n265 & ~n266 ;
  assign n268 = \totalcoeffs[3]  & ~n267 ;
  assign n269 = \totalcoeffs[2]  & ~n120 ;
  assign n270 = \totalcoeffs[1]  & ~n269 ;
  assign n271 = \ctable[0]  & ~n186 ;
  assign n272 = ~n270 & n271 ;
  assign n273 = ~n268 & ~n272 ;
  assign n274 = \totalcoeffs[3]  & ~n172 ;
  assign n275 = \ctable[0]  & ~n274 ;
  assign n276 = \totalcoeffs[2]  & ~\ctable[0]  ;
  assign n277 = \totalcoeffs[3]  & ~n276 ;
  assign n278 = \trailingones[0]  & ~n277 ;
  assign n279 = ~n275 & ~n278 ;
  assign n280 = n53 & ~n279 ;
  assign n281 = \ctable[1]  & ~\trailingones[0]  ;
  assign n282 = ~\totalcoeffs[3]  & \trailingones[1]  ;
  assign n283 = \totalcoeffs[1]  & n282 ;
  assign n284 = n281 & n283 ;
  assign n285 = ~n29 & ~n220 ;
  assign n286 = ~\ctable[1]  & ~n282 ;
  assign n287 = ~n285 & n286 ;
  assign n288 = ~n284 & ~n287 ;
  assign n289 = ~\ctable[0]  & \ctable[1]  ;
  assign n290 = n132 & n289 ;
  assign n291 = n231 & n290 ;
  assign n292 = ~\totalcoeffs[4]  & ~n291 ;
  assign n293 = n288 & n292 ;
  assign n294 = ~n280 & n293 ;
  assign n295 = n273 & n294 ;
  assign n296 = ~\totalcoeffs[1]  & n25 ;
  assign n297 = \totalcoeffs[4]  & ~n296 ;
  assign n298 = ~n232 & ~n281 ;
  assign n299 = \totalcoeffs[4]  & ~\ctable[0]  ;
  assign n300 = ~n298 & n299 ;
  assign n301 = ~n297 & ~n300 ;
  assign n302 = ~\totalcoeffs[0]  & n301 ;
  assign n303 = ~n295 & n302 ;
  assign n304 = ~\ctable[2]  & n303 ;
  assign n305 = ~n25 & n157 ;
  assign n306 = \trailingones[1]  & n305 ;
  assign n307 = \ctable[0]  & ~n144 ;
  assign n308 = ~\totalcoeffs[2]  & n231 ;
  assign n309 = ~n307 & n308 ;
  assign n310 = ~n306 & ~n309 ;
  assign n311 = \totalcoeffs[0]  & ~\ctable[1]  ;
  assign n312 = ~n310 & n311 ;
  assign n313 = ~n155 & ~n233 ;
  assign n314 = \totalcoeffs[2]  & ~n313 ;
  assign n315 = \trailingones[1]  & n215 ;
  assign n316 = \ctable[0]  & ~n231 ;
  assign n317 = ~n315 & n316 ;
  assign n318 = ~\ctable[0]  & ~n75 ;
  assign n319 = \totalcoeffs[1]  & ~n318 ;
  assign n320 = ~n317 & n319 ;
  assign n321 = ~n314 & ~n320 ;
  assign n322 = ~\totalcoeffs[3]  & ~\ctable[1]  ;
  assign n323 = ~n321 & n322 ;
  assign n324 = ~n312 & ~n323 ;
  assign n325 = \trailingones[0]  & n53 ;
  assign n326 = ~n24 & n224 ;
  assign n327 = ~n325 & ~n326 ;
  assign n328 = \totalcoeffs[1]  & \trailingones[1]  ;
  assign n329 = ~n92 & ~n328 ;
  assign n330 = n181 & ~n329 ;
  assign n331 = n327 & ~n330 ;
  assign n332 = ~\totalcoeffs[2]  & ~n331 ;
  assign n333 = \totalcoeffs[2]  & \ctable[1]  ;
  assign n334 = n328 & n333 ;
  assign n335 = ~n158 & ~n334 ;
  assign n336 = \trailingones[0]  & ~n12 ;
  assign n337 = \totalcoeffs[2]  & n231 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = n335 & n338 ;
  assign n340 = \totalcoeffs[3]  & ~n339 ;
  assign n341 = ~n332 & ~n340 ;
  assign n342 = n174 & ~n341 ;
  assign n343 = n324 & ~n342 ;
  assign n344 = ~\totalcoeffs[4]  & ~\ctable[2]  ;
  assign n345 = ~n343 & n344 ;
  assign n346 = ~n304 & ~n345 ;
  assign n347 = \ctable[2]  & n232 ;
  assign n348 = \totalcoeffs[0]  & ~n347 ;
  assign n349 = n47 & ~n348 ;
  assign n350 = n51 & n155 ;
  assign n351 = ~n349 & ~n350 ;
  assign n352 = ~\ctable[0]  & ~\ctable[1]  ;
  assign n353 = ~\totalcoeffs[4]  & n25 ;
  assign n354 = n352 & n353 ;
  assign n355 = ~n351 & n354 ;
  assign n356 = n346 & ~n355 ;
  assign n357 = \totalcoeffs[3]  & ~\ctable[1]  ;
  assign n358 = ~\trailingones[0]  & n357 ;
  assign n359 = n231 & n289 ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = ~\totalcoeffs[1]  & ~n360 ;
  assign n362 = \totalcoeffs[2]  & n357 ;
  assign n363 = ~n25 & n289 ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = n24 & ~n364 ;
  assign n366 = ~n361 & ~n365 ;
  assign n367 = ~\trailingones[1]  & n36 ;
  assign n368 = n289 & n367 ;
  assign n369 = ~n40 & ~n200 ;
  assign n370 = ~\totalcoeffs[2]  & ~n369 ;
  assign n371 = \ctable[0]  & \trailingones[1]  ;
  assign n372 = ~\ctable[1]  & ~n371 ;
  assign n373 = \ctable[0]  & \trailingones[0]  ;
  assign n374 = ~n328 & ~n373 ;
  assign n375 = n372 & ~n374 ;
  assign n376 = ~n370 & ~n375 ;
  assign n377 = \totalcoeffs[3]  & ~n376 ;
  assign n378 = ~n368 & ~n377 ;
  assign n379 = n366 & n378 ;
  assign n380 = ~\totalcoeffs[4]  & ~n379 ;
  assign n381 = ~n231 & ~n371 ;
  assign n382 = \totalcoeffs[2]  & ~n381 ;
  assign n383 = ~\totalcoeffs[3]  & ~n281 ;
  assign n384 = ~n382 & n383 ;
  assign n385 = \totalcoeffs[1]  & ~n121 ;
  assign n386 = ~n384 & n385 ;
  assign n387 = ~\trailingones[1]  & n144 ;
  assign n388 = ~\totalcoeffs[0]  & ~n387 ;
  assign n389 = \totalcoeffs[1]  & ~n276 ;
  assign n390 = \ctable[1]  & ~n25 ;
  assign n391 = ~n389 & n390 ;
  assign n392 = n388 & ~n391 ;
  assign n393 = ~n386 & n392 ;
  assign n394 = \ctable[0]  & n57 ;
  assign n395 = ~\trailingones[1]  & n163 ;
  assign n396 = n394 & n395 ;
  assign n397 = ~\totalcoeffs[3]  & ~\trailingones[1]  ;
  assign n398 = n289 & n397 ;
  assign n399 = \totalcoeffs[0]  & ~n398 ;
  assign n400 = ~n396 & n399 ;
  assign n401 = ~\totalcoeffs[4]  & ~n400 ;
  assign n402 = \totalcoeffs[2]  & n182 ;
  assign n403 = ~\totalcoeffs[2]  & ~n373 ;
  assign n404 = ~\trailingones[1]  & ~n403 ;
  assign n405 = ~n402 & n404 ;
  assign n406 = ~\totalcoeffs[2]  & \totalcoeffs[3]  ;
  assign n407 = n85 & n220 ;
  assign n408 = ~n406 & ~n407 ;
  assign n409 = ~\ctable[1]  & ~n100 ;
  assign n410 = ~n160 & ~n409 ;
  assign n411 = n408 & ~n410 ;
  assign n412 = ~n405 & n411 ;
  assign n413 = \totalcoeffs[1]  & ~\totalcoeffs[4]  ;
  assign n414 = ~n412 & n413 ;
  assign n415 = ~n401 & ~n414 ;
  assign n416 = ~n393 & ~n415 ;
  assign n417 = ~n380 & ~n416 ;
  assign n418 = ~\totalcoeffs[3]  & \totalcoeffs[4]  ;
  assign n419 = n209 & n418 ;
  assign n420 = ~n84 & ~n352 ;
  assign n421 = ~\ctable[0]  & ~n232 ;
  assign n422 = ~n420 & ~n421 ;
  assign n423 = n419 & n422 ;
  assign n424 = n417 & ~n423 ;
  assign n425 = ~\ctable[2]  & ~n424 ;
  assign n426 = \totalcoeffs[2]  & ~\totalcoeffs[4]  ;
  assign n427 = ~n11 & n426 ;
  assign n428 = \totalcoeffs[3]  & ~\totalcoeffs[4]  ;
  assign n429 = ~n418 & ~n428 ;
  assign n430 = n209 & ~n429 ;
  assign n431 = ~n427 & ~n430 ;
  assign n432 = ~\ctable[2]  & n84 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = ~n209 & n428 ;
  assign n435 = ~n419 & ~n434 ;
  assign n436 = n432 & ~n435 ;
  assign n437 = ~\totalcoeffs[2]  & ~\ctable[2]  ;
  assign n438 = n11 & n437 ;
  assign n439 = n418 & n438 ;
  assign n440 = ~n432 & ~n439 ;
  assign n441 = n53 & n68 ;
  assign n442 = \ctable[2]  & ~\trailingones[1]  ;
  assign n443 = \trailingones[0]  & ~n442 ;
  assign n444 = ~\totalcoeffs[0]  & n237 ;
  assign n445 = ~n443 & n444 ;
  assign n446 = ~n441 & ~n445 ;
  assign n447 = n215 & n328 ;
  assign n448 = ~n231 & ~n447 ;
  assign n449 = ~\totalcoeffs[2]  & \ctable[2]  ;
  assign n450 = ~n448 & n449 ;
  assign n451 = n446 & ~n450 ;
  assign n452 = ~\ctable[1]  & n48 ;
  assign n453 = ~\totalcoeffs[4]  & n452 ;
  assign n454 = ~n451 & n453 ;
  assign n455 = ~n344 & ~n454 ;
  assign n456 = n440 & n455 ;
  assign n457 = ~\totalcoeffs[1]  & ~n231 ;
  assign n458 = ~n53 & n174 ;
  assign n459 = ~n457 & n458 ;
  assign n460 = ~\totalcoeffs[0]  & ~\ctable[1]  ;
  assign n461 = ~n155 & n460 ;
  assign n462 = ~n137 & ~n461 ;
  assign n463 = ~\ctable[0]  & n329 ;
  assign n464 = ~n462 & n463 ;
  assign n465 = ~n459 & ~n464 ;
  assign n466 = ~n174 & ~n213 ;
  assign n467 = n53 & n466 ;
  assign n468 = ~\totalcoeffs[0]  & \totalcoeffs[2]  ;
  assign n469 = n103 & ~n468 ;
  assign n470 = n77 & n215 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = \trailingones[1]  & ~n471 ;
  assign n473 = ~n467 & ~n472 ;
  assign n474 = n465 & n473 ;
  assign n475 = \totalcoeffs[3]  & ~n474 ;
  assign n476 = ~n451 & n452 ;
  assign n477 = ~\totalcoeffs[1]  & ~\ctable[0]  ;
  assign n478 = \totalcoeffs[2]  & ~n477 ;
  assign n479 = \totalcoeffs[0]  & n123 ;
  assign n480 = ~n478 & n479 ;
  assign n481 = n162 & n371 ;
  assign n482 = ~n40 & n468 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = ~n480 & n483 ;
  assign n485 = n15 & ~n484 ;
  assign n486 = n57 & n126 ;
  assign n487 = \totalcoeffs[2]  & \trailingones[0]  ;
  assign n488 = n222 & n487 ;
  assign n489 = ~n486 & ~n488 ;
  assign n490 = ~\totalcoeffs[3]  & ~n489 ;
  assign n491 = \trailingones[1]  & n468 ;
  assign n492 = ~n93 & ~n491 ;
  assign n493 = ~\totalcoeffs[3]  & \ctable[0]  ;
  assign n494 = ~n492 & n493 ;
  assign n495 = ~n490 & ~n494 ;
  assign n496 = ~n485 & n495 ;
  assign n497 = ~n476 & n496 ;
  assign n498 = ~n475 & n497 ;
  assign n499 = n63 & n85 ;
  assign n500 = ~\ctable[1]  & ~n276 ;
  assign n501 = n46 & ~n500 ;
  assign n502 = ~n499 & ~n501 ;
  assign n503 = ~\trailingones[0]  & ~n502 ;
  assign n504 = \totalcoeffs[2]  & ~n231 ;
  assign n505 = ~n315 & ~n504 ;
  assign n506 = \ctable[1]  & ~n505 ;
  assign n507 = \totalcoeffs[1]  & ~n506 ;
  assign n508 = ~n503 & n507 ;
  assign n509 = \trailingones[0]  & ~n174 ;
  assign n510 = n212 & ~n460 ;
  assign n511 = ~n509 & n510 ;
  assign n512 = n46 & n487 ;
  assign n513 = ~\totalcoeffs[1]  & ~n512 ;
  assign n514 = ~n511 & n513 ;
  assign n515 = ~n508 & ~n514 ;
  assign n516 = n440 & ~n515 ;
  assign n517 = n498 & n516 ;
  assign n518 = ~n456 & ~n517 ;
  assign n519 = ~\ctable[0]  & ~\ctable[2]  ;
  assign n520 = n418 & n519 ;
  assign n521 = n209 & n520 ;
  assign n522 = ~\ctable[1]  & n521 ;
  assign n523 = \totalcoeffs[4]  & ~n522 ;
  assign n524 = n196 & ~n233 ;
  assign n525 = ~\ctable[1]  & ~n232 ;
  assign n526 = n81 & n525 ;
  assign n527 = ~n524 & ~n526 ;
  assign n528 = \totalcoeffs[3]  & ~n527 ;
  assign n529 = ~\ctable[1]  & ~n181 ;
  assign n530 = n504 & ~n529 ;
  assign n531 = ~\totalcoeffs[0]  & n57 ;
  assign n532 = \ctable[1]  & n215 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = ~\trailingones[1]  & ~n533 ;
  assign n535 = ~n530 & ~n534 ;
  assign n536 = ~n528 & n535 ;
  assign n537 = ~\totalcoeffs[1]  & ~n536 ;
  assign n538 = n165 & n357 ;
  assign n539 = ~n281 & ~n538 ;
  assign n540 = \trailingones[1]  & ~n539 ;
  assign n541 = ~\trailingones[0]  & ~n222 ;
  assign n542 = \totalcoeffs[0]  & ~n357 ;
  assign n543 = ~n126 & ~n542 ;
  assign n544 = ~n541 & ~n543 ;
  assign n545 = ~n540 & ~n544 ;
  assign n546 = n228 & ~n545 ;
  assign n547 = n123 & n181 ;
  assign n548 = ~\totalcoeffs[3]  & n232 ;
  assign n549 = ~n547 & ~n548 ;
  assign n550 = ~n232 & n357 ;
  assign n551 = ~\ctable[1]  & n215 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = n549 & n552 ;
  assign n554 = ~\totalcoeffs[2]  & ~n547 ;
  assign n555 = \totalcoeffs[1]  & ~n554 ;
  assign n556 = ~n553 & n555 ;
  assign n557 = ~\trailingones[1]  & n77 ;
  assign n558 = n100 & n557 ;
  assign n559 = ~n556 & ~n558 ;
  assign n560 = ~n546 & n559 ;
  assign n561 = ~n537 & n560 ;
  assign n562 = n519 & ~n561 ;
  assign n563 = ~n12 & ~n139 ;
  assign n564 = ~n232 & ~n563 ;
  assign n565 = \totalcoeffs[2]  & ~n213 ;
  assign n566 = \totalcoeffs[1]  & ~n565 ;
  assign n567 = n564 & n566 ;
  assign n568 = ~n75 & ~n212 ;
  assign n569 = n215 & n568 ;
  assign n570 = \trailingones[0]  & ~\trailingones[1]  ;
  assign n571 = n19 & n570 ;
  assign n572 = n140 & n220 ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = ~n569 & n573 ;
  assign n575 = n29 & ~n574 ;
  assign n576 = ~n567 & ~n575 ;
  assign n577 = \trailingones[0]  & n371 ;
  assign n578 = n65 & n577 ;
  assign n579 = \totalcoeffs[1]  & ~n578 ;
  assign n580 = ~n65 & n233 ;
  assign n581 = ~\totalcoeffs[2]  & ~n27 ;
  assign n582 = \ctable[0]  & ~n581 ;
  assign n583 = ~n580 & n582 ;
  assign n584 = n27 & n337 ;
  assign n585 = ~n578 & ~n584 ;
  assign n586 = ~n583 & n585 ;
  assign n587 = ~n579 & ~n586 ;
  assign n588 = n576 & ~n587 ;
  assign n589 = n190 & ~n588 ;
  assign n590 = n233 & n468 ;
  assign n591 = n173 & n442 ;
  assign n592 = ~n590 & ~n591 ;
  assign n593 = n48 & n163 ;
  assign n594 = ~n592 & n593 ;
  assign n595 = ~n522 & ~n594 ;
  assign n596 = ~n589 & n595 ;
  assign n597 = ~n562 & n596 ;
  assign n598 = ~n523 & ~n597 ;
  assign n599 = n85 & n92 ;
  assign n600 = ~n283 & ~n599 ;
  assign n601 = ~\totalcoeffs[0]  & ~n600 ;
  assign n602 = ~n64 & ~n160 ;
  assign n603 = ~\totalcoeffs[2]  & ~n92 ;
  assign n604 = ~n282 & n603 ;
  assign n605 = n602 & n604 ;
  assign n606 = n329 & ~n477 ;
  assign n607 = n104 & ~n606 ;
  assign n608 = ~n605 & ~n607 ;
  assign n609 = ~n601 & n608 ;
  assign n610 = ~\trailingones[0]  & ~n609 ;
  assign n611 = ~\ctable[0]  & ~n165 ;
  assign n612 = ~\trailingones[1]  & ~n139 ;
  assign n613 = ~n611 & n612 ;
  assign n614 = n137 & n613 ;
  assign n615 = n21 & n48 ;
  assign n616 = ~\totalcoeffs[2]  & ~n74 ;
  assign n617 = n602 & n616 ;
  assign n618 = ~n615 & ~n617 ;
  assign n619 = n570 & ~n618 ;
  assign n620 = ~n614 & ~n619 ;
  assign n621 = ~n139 & ~n276 ;
  assign n622 = ~n274 & ~n621 ;
  assign n623 = n328 & n622 ;
  assign n624 = ~n19 & n172 ;
  assign n625 = \trailingones[1]  & n144 ;
  assign n626 = n624 & n625 ;
  assign n627 = ~n623 & ~n626 ;
  assign n628 = n620 & n627 ;
  assign n629 = ~n610 & n628 ;
  assign n630 = n190 & ~n629 ;
  assign n631 = \totalcoeffs[0]  & ~n457 ;
  assign n632 = ~\ctable[1]  & ~n103 ;
  assign n633 = ~n631 & n632 ;
  assign n634 = \ctable[1]  & ~n24 ;
  assign n635 = ~n53 & n165 ;
  assign n636 = n634 & ~n635 ;
  assign n637 = ~\totalcoeffs[2]  & ~n636 ;
  assign n638 = ~n633 & ~n637 ;
  assign n639 = ~\ctable[2]  & n160 ;
  assign n640 = n638 & n639 ;
  assign n641 = n328 & n531 ;
  assign n642 = n452 & n641 ;
  assign n643 = \trailingones[0]  & n68 ;
  assign n644 = ~n232 & ~n263 ;
  assign n645 = ~n643 & n644 ;
  assign n646 = \totalcoeffs[0]  & ~\trailingones[0]  ;
  assign n647 = \totalcoeffs[0]  & \totalcoeffs[2]  ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = \totalcoeffs[2]  & ~\trailingones[0]  ;
  assign n650 = ~\trailingones[1]  & n649 ;
  assign n651 = n648 & ~n650 ;
  assign n652 = n645 & n651 ;
  assign n653 = ~\totalcoeffs[1]  & n452 ;
  assign n654 = n652 & n653 ;
  assign n655 = ~n642 & ~n654 ;
  assign n656 = ~n640 & n655 ;
  assign n657 = ~n630 & n656 ;
  assign n658 = ~\totalcoeffs[4]  & ~n657 ;
  assign n659 = ~n521 & ~n658 ;
  assign n660 = ~n421 & n457 ;
  assign n661 = n104 & n660 ;
  assign n662 = n165 & ~n372 ;
  assign n663 = \totalcoeffs[3]  & ~n222 ;
  assign n664 = ~n662 & n663 ;
  assign n665 = ~n352 & n418 ;
  assign n666 = ~\totalcoeffs[1]  & ~\totalcoeffs[2]  ;
  assign n667 = ~n665 & n666 ;
  assign n668 = ~n664 & n667 ;
  assign n669 = ~n661 & ~n668 ;
  assign n670 = n174 & n362 ;
  assign n671 = ~\ctable[2]  & ~n670 ;
  assign n672 = ~n457 & ~n671 ;
  assign n673 = n669 & ~n672 ;
  assign n674 = ~\totalcoeffs[0]  & n224 ;
  assign n675 = n263 & n674 ;
  assign n676 = n40 & ~n165 ;
  assign n677 = n25 & ~n676 ;
  assign n678 = ~n675 & ~n677 ;
  assign n679 = n362 & n421 ;
  assign n680 = ~\totalcoeffs[3]  & \ctable[1]  ;
  assign n681 = n15 & n371 ;
  assign n682 = ~n680 & ~n681 ;
  assign n683 = ~n679 & n682 ;
  assign n684 = n678 & n683 ;
  assign n685 = \totalcoeffs[1]  & ~n684 ;
  assign n686 = \ctable[2]  & ~n104 ;
  assign n687 = ~n297 & ~n686 ;
  assign n688 = \totalcoeffs[0]  & \ctable[2]  ;
  assign n689 = n43 & n132 ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = ~\ctable[0]  & ~n104 ;
  assign n692 = \ctable[1]  & ~n691 ;
  assign n693 = n690 & ~n692 ;
  assign n694 = n687 & n693 ;
  assign n695 = ~n685 & n694 ;
  assign n696 = n673 & n695 ;
  assign n697 = \trailingones[0]  & ~n47 ;
  assign n698 = \totalcoeffs[2]  & n428 ;
  assign n699 = ~n52 & n698 ;
  assign n700 = ~n697 & n699 ;
  assign n701 = ~n419 & ~n700 ;
  assign n702 = ~\ctable[2]  & n352 ;
  assign n703 = ~n701 & n702 ;
  assign \coeff_token[0]  = ~n136 ;
  assign \coeff_token[1]  = ~n262 ;
  assign \coeff_token[2]  = ~n356 ;
  assign \coeff_token[3]  = n425 ;
  assign \coeff_token[4]  = n433 ;
  assign \coeff_token[5]  = n436 ;
  assign \ctoken_len[0]  = ~n518 ;
  assign \ctoken_len[1]  = ~n598 ;
  assign \ctoken_len[2]  = n659 ;
  assign \ctoken_len[3]  = n696 ;
  assign \ctoken_len[4]  = n703 ;
endmodule
