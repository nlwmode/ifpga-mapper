module top( \a0_pad  , a_pad , \b0_pad  , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , \l0_pad  , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \d0_pad  , \e0_pad  , \f0_pad  , \g0_pad  , \h0_pad  , \i0_pad  , \j0_pad  , \k0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  , \t0_pad  , \u0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input \l0_pad  ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \d0_pad  ;
  output \e0_pad  ;
  output \f0_pad  ;
  output \g0_pad  ;
  output \h0_pad  ;
  output \i0_pad  ;
  output \j0_pad  ;
  output \k0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  output \t0_pad  ;
  output \u0_pad  ;
  wire n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 ;
  assign n29 = ~\l0_pad  & ~u_pad ;
  assign n30 = ~i_pad & \l0_pad  ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = ~\l0_pad  & ~v_pad ;
  assign n33 = ~j_pad & \l0_pad  ;
  assign n34 = ~n32 & ~n33 ;
  assign n35 = ~\l0_pad  & ~w_pad ;
  assign n36 = ~k_pad & \l0_pad  ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = ~\l0_pad  & ~x_pad ;
  assign n39 = \l0_pad  & ~l_pad ;
  assign n40 = ~n38 & ~n39 ;
  assign n41 = ~\l0_pad  & ~y_pad ;
  assign n42 = \l0_pad  & ~m_pad ;
  assign n43 = ~n41 & ~n42 ;
  assign n44 = ~\l0_pad  & ~z_pad ;
  assign n45 = \l0_pad  & ~n_pad ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = ~\a0_pad  & ~\l0_pad  ;
  assign n48 = \l0_pad  & ~o_pad ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = ~\b0_pad  & ~\l0_pad  ;
  assign n51 = \l0_pad  & ~p_pad ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = ~q_pad & ~s_pad ;
  assign n54 = i_pad & n53 ;
  assign n55 = ~r_pad & ~u_pad ;
  assign n56 = q_pad & n55 ;
  assign n61 = ~n54 & ~n56 ;
  assign n57 = ~q_pad & s_pad ;
  assign n58 = a_pad & n57 ;
  assign n59 = q_pad & r_pad ;
  assign n60 = u_pad & n59 ;
  assign n62 = ~n58 & ~n60 ;
  assign n63 = n61 & n62 ;
  assign n67 = v_pad & ~n55 ;
  assign n66 = ~v_pad & n55 ;
  assign n68 = q_pad & ~n66 ;
  assign n69 = ~n67 & n68 ;
  assign n64 = ~j_pad & n53 ;
  assign n65 = ~b_pad & n57 ;
  assign n70 = ~n64 & ~n65 ;
  assign n71 = ~n69 & n70 ;
  assign n73 = c_pad & s_pad ;
  assign n72 = k_pad & ~s_pad ;
  assign n74 = ~q_pad & ~n72 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = w_pad & ~n66 ;
  assign n77 = ~v_pad & ~w_pad ;
  assign n78 = n55 & n77 ;
  assign n79 = q_pad & ~n78 ;
  assign n80 = ~n76 & n79 ;
  assign n81 = ~n75 & ~n80 ;
  assign n82 = ~x_pad & n78 ;
  assign n83 = x_pad & ~n78 ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = q_pad & ~n84 ;
  assign n87 = ~d_pad & s_pad ;
  assign n86 = ~l_pad & ~s_pad ;
  assign n88 = ~q_pad & ~n86 ;
  assign n89 = ~n87 & n88 ;
  assign n90 = ~n85 & ~n89 ;
  assign n92 = e_pad & s_pad ;
  assign n91 = m_pad & ~s_pad ;
  assign n93 = ~q_pad & ~n91 ;
  assign n94 = ~n92 & n93 ;
  assign n96 = ~y_pad & n82 ;
  assign n95 = y_pad & ~n82 ;
  assign n97 = q_pad & ~n95 ;
  assign n98 = ~n96 & n97 ;
  assign n99 = ~n94 & ~n98 ;
  assign n101 = f_pad & s_pad ;
  assign n100 = n_pad & ~s_pad ;
  assign n102 = ~q_pad & ~n100 ;
  assign n103 = ~n101 & n102 ;
  assign n104 = z_pad & ~n96 ;
  assign n105 = ~x_pad & ~y_pad ;
  assign n106 = ~z_pad & n105 ;
  assign n107 = n78 & n106 ;
  assign n108 = q_pad & ~n107 ;
  assign n109 = ~n104 & n108 ;
  assign n110 = ~n103 & ~n109 ;
  assign n111 = \a0_pad  & ~n107 ;
  assign n112 = ~\a0_pad  & n107 ;
  assign n113 = ~n111 & ~n112 ;
  assign n114 = q_pad & ~n113 ;
  assign n116 = ~g_pad & s_pad ;
  assign n115 = ~o_pad & ~s_pad ;
  assign n117 = ~q_pad & ~n115 ;
  assign n118 = ~n116 & n117 ;
  assign n119 = ~n114 & ~n118 ;
  assign n120 = ~\a0_pad  & \b0_pad  ;
  assign n121 = ~y_pad & ~z_pad ;
  assign n122 = n120 & n121 ;
  assign n123 = n82 & n122 ;
  assign n124 = ~\b0_pad  & ~n112 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = q_pad & ~n125 ;
  assign n128 = h_pad & s_pad ;
  assign n127 = p_pad & ~s_pad ;
  assign n129 = ~q_pad & ~n127 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = ~n126 & ~n130 ;
  assign n133 = ~\a0_pad  & u_pad ;
  assign n134 = n77 & n133 ;
  assign n135 = n106 & n134 ;
  assign n136 = ~n122 & n135 ;
  assign n137 = ~r_pad & ~n136 ;
  assign n132 = ~\l0_pad  & r_pad ;
  assign n138 = q_pad & ~n132 ;
  assign n139 = ~n137 & n138 ;
  assign \d0_pad  = ~n31 ;
  assign \e0_pad  = ~n34 ;
  assign \f0_pad  = ~n37 ;
  assign \g0_pad  = ~n40 ;
  assign \h0_pad  = ~n43 ;
  assign \i0_pad  = ~n46 ;
  assign \j0_pad  = ~n49 ;
  assign \k0_pad  = ~n52 ;
  assign \m0_pad  = ~n63 ;
  assign \n0_pad  = n71 ;
  assign \o0_pad  = n81 ;
  assign \p0_pad  = ~n90 ;
  assign \q0_pad  = n99 ;
  assign \r0_pad  = n110 ;
  assign \s0_pad  = ~n119 ;
  assign \t0_pad  = n131 ;
  assign \u0_pad  = n139 ;
endmodule
