module top( \CarrierSense_Tx2_reg/NET0131  , \Collision_Tx1_reg/NET0131  , \Collision_Tx2_reg/NET0131  , \RstTxPauseRq_reg/NET0131  , \RxAbortRst_reg/NET0131  , \RxAbort_latch_reg/NET0131  , \RxAbort_wb_reg/NET0131  , \RxEnSync_reg/NET0131  , \TPauseRq_reg/NET0131  , \TxPauseRq_sync2_reg/NET0131  , \TxPauseRq_sync3_reg/NET0131  , \WillSendControlFrame_sync2_reg/NET0131  , \WillSendControlFrame_sync3_reg/NET0131  , \WillTransmit_q2_reg/P0001  , \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  , \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  , \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  , \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  , \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  , \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  , \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131  , \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131  , \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131  , \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131  , \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  , \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  , \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  , \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131  , \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131  , \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131  , \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131  , \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131  , \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131  , \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131  , \ethreg1_IPGR1_0_DataOut_reg[0]/NET0131  , \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131  , \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131  , \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131  , \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131  , \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131  , \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131  , \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131  , \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131  , \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131  , \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131  , \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131  , \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131  , \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131  , \ethreg1_IPGT_0_DataOut_reg[0]/NET0131  , \ethreg1_IPGT_0_DataOut_reg[1]/NET0131  , \ethreg1_IPGT_0_DataOut_reg[2]/NET0131  , \ethreg1_IPGT_0_DataOut_reg[3]/NET0131  , \ethreg1_IPGT_0_DataOut_reg[4]/NET0131  , \ethreg1_IPGT_0_DataOut_reg[5]/NET0131  , \ethreg1_IPGT_0_DataOut_reg[6]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  , \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  , \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  , \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  , \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  , \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  , \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  , \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131  , \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131  , \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131  , \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131  , \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131  , \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131  , \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131  , \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131  , \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131  , \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131  , \ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131  , \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131  , \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  , \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  , \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131  , \ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131  , \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131  , \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131  , \ethreg1_MODER_0_DataOut_reg[0]/NET0131  , \ethreg1_MODER_0_DataOut_reg[1]/NET0131  , \ethreg1_MODER_0_DataOut_reg[2]/NET0131  , \ethreg1_MODER_0_DataOut_reg[3]/NET0131  , \ethreg1_MODER_0_DataOut_reg[4]/NET0131  , \ethreg1_MODER_0_DataOut_reg[5]/NET0131  , \ethreg1_MODER_0_DataOut_reg[6]/NET0131  , \ethreg1_MODER_0_DataOut_reg[7]/NET0131  , \ethreg1_MODER_1_DataOut_reg[0]/NET0131  , \ethreg1_MODER_1_DataOut_reg[1]/NET0131  , \ethreg1_MODER_1_DataOut_reg[2]/NET0131  , \ethreg1_MODER_1_DataOut_reg[3]/NET0131  , \ethreg1_MODER_1_DataOut_reg[4]/NET0131  , \ethreg1_MODER_1_DataOut_reg[5]/NET0131  , \ethreg1_MODER_1_DataOut_reg[6]/NET0131  , \ethreg1_MODER_1_DataOut_reg[7]/NET0131  , \ethreg1_MODER_2_DataOut_reg[0]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  , \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  , \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  , \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  , \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131  , \ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131  , \ethreg1_ResetRxCIrq_sync2_reg/NET0131  , \ethreg1_ResetRxCIrq_sync3_reg/NET0131  , \ethreg1_ResetTxCIrq_sync2_reg/NET0131  , \ethreg1_SetRxCIrq_reg/NET0131  , \ethreg1_SetRxCIrq_rxclk_reg/NET0131  , \ethreg1_SetRxCIrq_sync2_reg/NET0131  , \ethreg1_SetRxCIrq_sync3_reg/NET0131  , \ethreg1_SetTxCIrq_reg/NET0131  , \ethreg1_SetTxCIrq_sync2_reg/NET0131  , \ethreg1_SetTxCIrq_sync3_reg/NET0131  , \ethreg1_SetTxCIrq_txclk_reg/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131  , \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131  , \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131  , \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131  , \ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131  , \ethreg1_irq_busy_reg/NET0131  , \ethreg1_irq_rxb_reg/NET0131  , \ethreg1_irq_rxc_reg/NET0131  , \ethreg1_irq_rxe_reg/NET0131  , \ethreg1_irq_txb_reg/NET0131  , \ethreg1_irq_txc_reg/NET0131  , \ethreg1_irq_txe_reg/NET0131  , m_wb_ack_i_pad , \m_wb_adr_o[10]_pad  , \m_wb_adr_o[11]_pad  , \m_wb_adr_o[12]_pad  , \m_wb_adr_o[13]_pad  , \m_wb_adr_o[14]_pad  , \m_wb_adr_o[15]_pad  , \m_wb_adr_o[16]_pad  , \m_wb_adr_o[17]_pad  , \m_wb_adr_o[18]_pad  , \m_wb_adr_o[19]_pad  , \m_wb_adr_o[20]_pad  , \m_wb_adr_o[21]_pad  , \m_wb_adr_o[22]_pad  , \m_wb_adr_o[23]_pad  , \m_wb_adr_o[24]_pad  , \m_wb_adr_o[25]_pad  , \m_wb_adr_o[26]_pad  , \m_wb_adr_o[27]_pad  , \m_wb_adr_o[28]_pad  , \m_wb_adr_o[29]_pad  , \m_wb_adr_o[2]_pad  , \m_wb_adr_o[30]_pad  , \m_wb_adr_o[31]_pad  , \m_wb_adr_o[3]_pad  , \m_wb_adr_o[4]_pad  , \m_wb_adr_o[5]_pad  , \m_wb_adr_o[6]_pad  , \m_wb_adr_o[7]_pad  , \m_wb_adr_o[8]_pad  , \m_wb_adr_o[9]_pad  , \m_wb_dat_i[10]_pad  , \m_wb_dat_i[11]_pad  , \m_wb_dat_i[12]_pad  , \m_wb_dat_i[13]_pad  , \m_wb_dat_i[14]_pad  , \m_wb_dat_i[15]_pad  , \m_wb_dat_i[16]_pad  , \m_wb_dat_i[17]_pad  , \m_wb_dat_i[18]_pad  , \m_wb_dat_i[19]_pad  , \m_wb_dat_i[1]_pad  , \m_wb_dat_i[20]_pad  , \m_wb_dat_i[22]_pad  , \m_wb_dat_i[23]_pad  , \m_wb_dat_i[24]_pad  , \m_wb_dat_i[25]_pad  , \m_wb_dat_i[26]_pad  , \m_wb_dat_i[27]_pad  , \m_wb_dat_i[28]_pad  , \m_wb_dat_i[29]_pad  , \m_wb_dat_i[2]_pad  , \m_wb_dat_i[30]_pad  , \m_wb_dat_i[31]_pad  , \m_wb_dat_i[3]_pad  , \m_wb_dat_i[4]_pad  , \m_wb_dat_i[5]_pad  , \m_wb_dat_i[6]_pad  , \m_wb_dat_i[7]_pad  , \m_wb_dat_i[8]_pad  , m_wb_err_i_pad , \m_wb_sel_o[0]_pad  , \m_wb_sel_o[1]_pad  , \m_wb_sel_o[2]_pad  , \m_wb_sel_o[3]_pad  , m_wb_stb_o_pad , m_wb_we_o_pad , \maccontrol1_MuxedAbort_reg/NET0131  , \maccontrol1_MuxedDone_reg/NET0131  , \maccontrol1_TxAbortInLatched_reg/NET0131  , \maccontrol1_TxDoneInLatched_reg/NET0131  , \maccontrol1_TxUsedDataOutDetected_reg/NET0131  , \maccontrol1_receivecontrol1_AddressOK_reg/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131  , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131  , \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  , \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  , \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  , \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  , \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  , \maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131  , \maccontrol1_receivecontrol1_Divider2_reg/NET0131  , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131  , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131  , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131  , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131  , \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131  , \maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131  , \maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  , \maccontrol1_receivecontrol1_Pause_reg/NET0131  , \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  , \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131  , \maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131  , \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  , \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131  , \maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131  , \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  , \maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131  , \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131  , \maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131  , \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  , \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  , \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  , \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  , \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  , \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131  , \maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131  , \maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001  , \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131  , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131  , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  , \maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131  , \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131  , \maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001  , \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  , \maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131  , \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131  , \macstatus1_CarrierSenseLost_reg/NET0131  , \macstatus1_DeferLatched_reg/NET0131  , \macstatus1_DribbleNibble_reg/NET0131  , \macstatus1_InvalidSymbol_reg/NET0131  , \macstatus1_LatchedCrcError_reg/NET0131  , \macstatus1_LatchedMRxErr_reg/NET0131  , \macstatus1_LateCollLatched_reg/P0002  , \macstatus1_LoadRxStatus_reg/NET0131  , \macstatus1_ReceiveEnd_reg/NET0131  , \macstatus1_ReceivedPacketTooBig_reg/NET0131  , \macstatus1_RetryCntLatched_reg[0]/P0002  , \macstatus1_RetryCntLatched_reg[1]/P0002  , \macstatus1_RetryCntLatched_reg[2]/P0002  , \macstatus1_RetryCntLatched_reg[3]/P0002  , \macstatus1_RetryLimit_reg/P0002  , \macstatus1_RxColWindow_reg/NET0131  , \macstatus1_RxLateCollision_reg/NET0131  , \macstatus1_ShortFrame_reg/NET0131  , mcoll_pad_i_pad , md_pad_i_pad , mdc_pad_o_pad , \miim1_BitCounter_reg[0]/NET0131  , \miim1_BitCounter_reg[1]/NET0131  , \miim1_BitCounter_reg[2]/NET0131  , \miim1_BitCounter_reg[3]/NET0131  , \miim1_BitCounter_reg[4]/NET0131  , \miim1_BitCounter_reg[5]/NET0131  , \miim1_BitCounter_reg[6]/NET0131  , \miim1_EndBusy_reg/NET0131  , \miim1_InProgress_q1_reg/NET0131  , \miim1_InProgress_q2_reg/NET0131  , \miim1_InProgress_q3_reg/NET0131  , \miim1_InProgress_reg/NET0131  , \miim1_LatchByte0_d_reg/NET0131  , \miim1_LatchByte1_d_reg/NET0131  , \miim1_LatchByte_reg[0]/NET0131  , \miim1_LatchByte_reg[1]/NET0131  , \miim1_Nvalid_reg/NET0131  , \miim1_RStatStart_q1_reg/NET0131  , \miim1_RStatStart_q2_reg/NET0131  , \miim1_RStatStart_reg/NET0131  , \miim1_RStat_q2_reg/NET0131  , \miim1_RStat_q3_reg/NET0131  , \miim1_ScanStat_q2_reg/NET0131  , \miim1_SyncStatMdcEn_reg/NET0131  , \miim1_WCtrlDataStart_q1_reg/NET0131  , \miim1_WCtrlDataStart_q2_reg/NET0131  , \miim1_WCtrlDataStart_q_reg/NET0131  , \miim1_WCtrlDataStart_reg/NET0131  , \miim1_WCtrlData_q2_reg/NET0131  , \miim1_WCtrlData_q3_reg/NET0131  , \miim1_WriteOp_reg/NET0131  , \miim1_clkgen_Counter_reg[0]/NET0131  , \miim1_clkgen_Counter_reg[1]/NET0131  , \miim1_clkgen_Counter_reg[2]/NET0131  , \miim1_clkgen_Counter_reg[3]/NET0131  , \miim1_clkgen_Counter_reg[4]/NET0131  , \miim1_clkgen_Counter_reg[5]/NET0131  , \miim1_clkgen_Counter_reg[6]/NET0131  , \miim1_outctrl_Mdo_2d_reg/NET0131  , \miim1_shftrg_LinkFail_reg/NET0131  , \miim1_shftrg_ShiftReg_reg[0]/NET0131  , \miim1_shftrg_ShiftReg_reg[1]/NET0131  , \miim1_shftrg_ShiftReg_reg[2]/NET0131  , \miim1_shftrg_ShiftReg_reg[3]/NET0131  , \miim1_shftrg_ShiftReg_reg[4]/NET0131  , \miim1_shftrg_ShiftReg_reg[5]/NET0131  , \miim1_shftrg_ShiftReg_reg[6]/NET0131  , \miim1_shftrg_ShiftReg_reg[7]/NET0131  , \mrxd_pad_i[0]_pad  , \mrxd_pad_i[1]_pad  , \mrxd_pad_i[2]_pad  , \mrxd_pad_i[3]_pad  , mrxdv_pad_i_pad , mrxerr_pad_i_pad , \mtxd_pad_o[0]_pad  , \mtxd_pad_o[1]_pad  , \mtxd_pad_o[2]_pad  , \mtxd_pad_o[3]_pad  , mtxen_pad_o_pad , mtxerr_pad_o_pad , \rxethmac1_Broadcast_reg/NET0131  , \rxethmac1_CrcHashGood_reg/P0001  , \rxethmac1_CrcHash_reg[0]/P0001  , \rxethmac1_CrcHash_reg[1]/P0001  , \rxethmac1_CrcHash_reg[2]/P0001  , \rxethmac1_CrcHash_reg[3]/P0001  , \rxethmac1_CrcHash_reg[4]/P0001  , \rxethmac1_CrcHash_reg[5]/P0001  , \rxethmac1_DelayData_reg/NET0131  , \rxethmac1_LatchedByte_reg[0]/NET0131  , \rxethmac1_LatchedByte_reg[1]/NET0131  , \rxethmac1_LatchedByte_reg[2]/NET0131  , \rxethmac1_LatchedByte_reg[3]/NET0131  , \rxethmac1_LatchedByte_reg[4]/NET0131  , \rxethmac1_LatchedByte_reg[5]/NET0131  , \rxethmac1_LatchedByte_reg[6]/NET0131  , \rxethmac1_LatchedByte_reg[7]/NET0131  , \rxethmac1_Multicast_reg/NET0131  , \rxethmac1_RxData_d_reg[0]/NET0131  , \rxethmac1_RxData_d_reg[1]/NET0131  , \rxethmac1_RxData_d_reg[2]/NET0131  , \rxethmac1_RxData_d_reg[3]/NET0131  , \rxethmac1_RxData_d_reg[4]/NET0131  , \rxethmac1_RxData_d_reg[5]/NET0131  , \rxethmac1_RxData_d_reg[6]/NET0131  , \rxethmac1_RxData_d_reg[7]/NET0131  , \rxethmac1_RxData_reg[0]/NET0131  , \rxethmac1_RxData_reg[1]/NET0131  , \rxethmac1_RxData_reg[2]/NET0131  , \rxethmac1_RxData_reg[3]/NET0131  , \rxethmac1_RxData_reg[4]/NET0131  , \rxethmac1_RxData_reg[5]/NET0131  , \rxethmac1_RxData_reg[6]/NET0131  , \rxethmac1_RxData_reg[7]/NET0131  , \rxethmac1_RxEndFrm_d_reg/NET0131  , \rxethmac1_RxEndFrm_reg/NET0131  , \rxethmac1_RxStartFrm_reg/NET0131  , \rxethmac1_RxValid_reg/NET0131  , \rxethmac1_crcrx_Crc_reg[0]/NET0131  , \rxethmac1_crcrx_Crc_reg[10]/NET0131  , \rxethmac1_crcrx_Crc_reg[11]/NET0131  , \rxethmac1_crcrx_Crc_reg[12]/NET0131  , \rxethmac1_crcrx_Crc_reg[13]/NET0131  , \rxethmac1_crcrx_Crc_reg[14]/NET0131  , \rxethmac1_crcrx_Crc_reg[15]/NET0131  , \rxethmac1_crcrx_Crc_reg[16]/NET0131  , \rxethmac1_crcrx_Crc_reg[17]/NET0131  , \rxethmac1_crcrx_Crc_reg[18]/NET0131  , \rxethmac1_crcrx_Crc_reg[19]/NET0131  , \rxethmac1_crcrx_Crc_reg[1]/NET0131  , \rxethmac1_crcrx_Crc_reg[20]/NET0131  , \rxethmac1_crcrx_Crc_reg[21]/NET0131  , \rxethmac1_crcrx_Crc_reg[22]/NET0131  , \rxethmac1_crcrx_Crc_reg[23]/NET0131  , \rxethmac1_crcrx_Crc_reg[24]/NET0131  , \rxethmac1_crcrx_Crc_reg[25]/NET0131  , \rxethmac1_crcrx_Crc_reg[26]/NET0131  , \rxethmac1_crcrx_Crc_reg[27]/NET0131  , \rxethmac1_crcrx_Crc_reg[28]/NET0131  , \rxethmac1_crcrx_Crc_reg[29]/NET0131  , \rxethmac1_crcrx_Crc_reg[2]/NET0131  , \rxethmac1_crcrx_Crc_reg[30]/NET0131  , \rxethmac1_crcrx_Crc_reg[31]/NET0131  , \rxethmac1_crcrx_Crc_reg[3]/NET0131  , \rxethmac1_crcrx_Crc_reg[4]/NET0131  , \rxethmac1_crcrx_Crc_reg[5]/NET0131  , \rxethmac1_crcrx_Crc_reg[6]/NET0131  , \rxethmac1_crcrx_Crc_reg[7]/NET0131  , \rxethmac1_crcrx_Crc_reg[8]/NET0131  , \rxethmac1_crcrx_Crc_reg[9]/NET0131  , \rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131  , \rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131  , \rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131  , \rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  , \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  , \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  , \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  , \rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  , \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  , \rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131  , \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  , \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  , \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131  , \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131  , \rxethmac1_rxstatem1_StateData0_reg/NET0131  , \rxethmac1_rxstatem1_StateData1_reg/NET0131  , \rxethmac1_rxstatem1_StateDrop_reg/NET0131  , \rxethmac1_rxstatem1_StateIdle_reg/NET0131  , \rxethmac1_rxstatem1_StatePreamble_reg/NET0131  , \rxethmac1_rxstatem1_StateSFD_reg/NET0131  , \txethmac1_ColWindow_reg/NET0131  , \txethmac1_PacketFinished_q_reg/NET0131  , \txethmac1_RetryCnt_reg[0]/NET0131  , \txethmac1_RetryCnt_reg[1]/NET0131  , \txethmac1_RetryCnt_reg[2]/NET0131  , \txethmac1_RetryCnt_reg[3]/NET0131  , \txethmac1_StatusLatch_reg/NET0131  , \txethmac1_StopExcessiveDeferOccured_reg/NET0131  , \txethmac1_TxAbort_reg/NET0131  , \txethmac1_TxDone_reg/NET0131  , \txethmac1_TxRetry_reg/NET0131  , \txethmac1_TxUsedData_reg/NET0131  , \txethmac1_random1_RandomLatched_reg[0]/NET0131  , \txethmac1_random1_RandomLatched_reg[1]/NET0131  , \txethmac1_random1_RandomLatched_reg[2]/NET0131  , \txethmac1_random1_RandomLatched_reg[3]/NET0131  , \txethmac1_random1_RandomLatched_reg[4]/NET0131  , \txethmac1_random1_RandomLatched_reg[5]/NET0131  , \txethmac1_random1_RandomLatched_reg[6]/NET0131  , \txethmac1_random1_RandomLatched_reg[7]/NET0131  , \txethmac1_random1_RandomLatched_reg[8]/NET0131  , \txethmac1_random1_RandomLatched_reg[9]/NET0131  , \txethmac1_random1_x_reg[1]/NET0131  , \txethmac1_random1_x_reg[2]/NET0131  , \txethmac1_random1_x_reg[3]/NET0131  , \txethmac1_random1_x_reg[4]/NET0131  , \txethmac1_random1_x_reg[5]/NET0131  , \txethmac1_random1_x_reg[6]/NET0131  , \txethmac1_random1_x_reg[7]/NET0131  , \txethmac1_random1_x_reg[8]/NET0131  , \txethmac1_random1_x_reg[9]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  , \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  , \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  , \txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131  , \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[14]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[15]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  , \txethmac1_txcounters1_NibCnt_reg[9]/NET0131  , \txethmac1_txcrc_Crc_reg[0]/NET0131  , \txethmac1_txcrc_Crc_reg[10]/NET0131  , \txethmac1_txcrc_Crc_reg[11]/NET0131  , \txethmac1_txcrc_Crc_reg[12]/NET0131  , \txethmac1_txcrc_Crc_reg[13]/NET0131  , \txethmac1_txcrc_Crc_reg[14]/NET0131  , \txethmac1_txcrc_Crc_reg[15]/NET0131  , \txethmac1_txcrc_Crc_reg[16]/NET0131  , \txethmac1_txcrc_Crc_reg[17]/NET0131  , \txethmac1_txcrc_Crc_reg[18]/NET0131  , \txethmac1_txcrc_Crc_reg[19]/NET0131  , \txethmac1_txcrc_Crc_reg[1]/NET0131  , \txethmac1_txcrc_Crc_reg[20]/NET0131  , \txethmac1_txcrc_Crc_reg[21]/NET0131  , \txethmac1_txcrc_Crc_reg[22]/NET0131  , \txethmac1_txcrc_Crc_reg[23]/NET0131  , \txethmac1_txcrc_Crc_reg[24]/NET0131  , \txethmac1_txcrc_Crc_reg[25]/NET0131  , \txethmac1_txcrc_Crc_reg[26]/NET0131  , \txethmac1_txcrc_Crc_reg[27]/NET0131  , \txethmac1_txcrc_Crc_reg[28]/NET0131  , \txethmac1_txcrc_Crc_reg[29]/NET0131  , \txethmac1_txcrc_Crc_reg[2]/NET0131  , \txethmac1_txcrc_Crc_reg[30]/NET0131  , \txethmac1_txcrc_Crc_reg[31]/NET0131  , \txethmac1_txcrc_Crc_reg[3]/NET0131  , \txethmac1_txcrc_Crc_reg[4]/NET0131  , \txethmac1_txcrc_Crc_reg[5]/NET0131  , \txethmac1_txcrc_Crc_reg[6]/NET0131  , \txethmac1_txcrc_Crc_reg[7]/NET0131  , \txethmac1_txcrc_Crc_reg[8]/NET0131  , \txethmac1_txcrc_Crc_reg[9]/NET0131  , \txethmac1_txstatem1_Rule1_reg/NET0131  , \txethmac1_txstatem1_StateBackOff_reg/NET0131  , \txethmac1_txstatem1_StateData_reg[0]/NET0131  , \txethmac1_txstatem1_StateData_reg[1]/NET0131  , \txethmac1_txstatem1_StateDefer_reg/NET0131  , \txethmac1_txstatem1_StateFCS_reg/NET0131  , \txethmac1_txstatem1_StateIPG_reg/NET0131  , \txethmac1_txstatem1_StateIdle_reg/NET0131  , \txethmac1_txstatem1_StateJam_q_reg/NET0131  , \txethmac1_txstatem1_StateJam_reg/NET0131  , \txethmac1_txstatem1_StatePAD_reg/NET0131  , \txethmac1_txstatem1_StatePreamble_reg/NET0131  , wb_ack_o_pad , \wb_adr_i[10]_pad  , \wb_adr_i[11]_pad  , \wb_adr_i[2]_pad  , \wb_adr_i[3]_pad  , \wb_adr_i[4]_pad  , \wb_adr_i[5]_pad  , \wb_adr_i[6]_pad  , \wb_adr_i[7]_pad  , \wb_adr_i[8]_pad  , \wb_adr_i[9]_pad  , wb_cyc_i_pad , \wb_dat_i[0]_pad  , \wb_dat_i[10]_pad  , \wb_dat_i[11]_pad  , \wb_dat_i[12]_pad  , \wb_dat_i[13]_pad  , \wb_dat_i[14]_pad  , \wb_dat_i[15]_pad  , \wb_dat_i[16]_pad  , \wb_dat_i[17]_pad  , \wb_dat_i[18]_pad  , \wb_dat_i[19]_pad  , \wb_dat_i[1]_pad  , \wb_dat_i[20]_pad  , \wb_dat_i[21]_pad  , \wb_dat_i[22]_pad  , \wb_dat_i[23]_pad  , \wb_dat_i[24]_pad  , \wb_dat_i[25]_pad  , \wb_dat_i[26]_pad  , \wb_dat_i[27]_pad  , \wb_dat_i[28]_pad  , \wb_dat_i[29]_pad  , \wb_dat_i[2]_pad  , \wb_dat_i[30]_pad  , \wb_dat_i[31]_pad  , \wb_dat_i[3]_pad  , \wb_dat_i[4]_pad  , \wb_dat_i[5]_pad  , \wb_dat_i[6]_pad  , \wb_dat_i[7]_pad  , \wb_dat_i[8]_pad  , \wb_dat_i[9]_pad  , wb_err_o_pad , wb_rst_i_pad , \wb_sel_i[0]_pad  , \wb_sel_i[1]_pad  , \wb_sel_i[2]_pad  , \wb_sel_i[3]_pad  , wb_stb_i_pad , wb_we_i_pad , \wishbone_BDRead_reg/NET0131  , \wishbone_BDWrite_reg[0]/NET0131  , \wishbone_BDWrite_reg[1]/NET0131  , \wishbone_BDWrite_reg[2]/NET0131  , \wishbone_BDWrite_reg[3]/NET0131  , \wishbone_BlockReadTxDataFromMemory_reg/NET0131  , \wishbone_BlockingIncrementTxPointer_reg/NET0131  , \wishbone_BlockingTxBDRead_reg/NET0131  , \wishbone_BlockingTxStatusWrite_reg/NET0131  , \wishbone_BlockingTxStatusWrite_sync2_reg/NET0131  , \wishbone_BlockingTxStatusWrite_sync3_reg/NET0131  , \wishbone_Busy_IRQ_rck_reg/NET0131  , \wishbone_Busy_IRQ_sync2_reg/P0001  , \wishbone_Busy_IRQ_sync3_reg/P0001  , \wishbone_Busy_IRQ_syncb2_reg/P0001  , \wishbone_Flop_reg/NET0131  , \wishbone_IncrTxPointer_reg/NET0131  , \wishbone_LastByteIn_reg/NET0131  , \wishbone_LastWord_reg/NET0131  , \wishbone_LatchValidBytes_q_reg/NET0131  , \wishbone_LatchValidBytes_reg/NET0131  , \wishbone_LatchedRxLength_reg[0]/NET0131  , \wishbone_LatchedRxLength_reg[10]/NET0131  , \wishbone_LatchedRxLength_reg[11]/NET0131  , \wishbone_LatchedRxLength_reg[12]/NET0131  , \wishbone_LatchedRxLength_reg[13]/NET0131  , \wishbone_LatchedRxLength_reg[14]/NET0131  , \wishbone_LatchedRxLength_reg[15]/NET0131  , \wishbone_LatchedRxLength_reg[1]/NET0131  , \wishbone_LatchedRxLength_reg[2]/NET0131  , \wishbone_LatchedRxLength_reg[3]/NET0131  , \wishbone_LatchedRxLength_reg[4]/NET0131  , \wishbone_LatchedRxLength_reg[5]/NET0131  , \wishbone_LatchedRxLength_reg[6]/NET0131  , \wishbone_LatchedRxLength_reg[7]/NET0131  , \wishbone_LatchedRxLength_reg[8]/NET0131  , \wishbone_LatchedRxLength_reg[9]/NET0131  , \wishbone_LatchedRxStartFrm_reg/NET0131  , \wishbone_LatchedTxLength_reg[0]/NET0131  , \wishbone_LatchedTxLength_reg[10]/NET0131  , \wishbone_LatchedTxLength_reg[11]/NET0131  , \wishbone_LatchedTxLength_reg[12]/NET0131  , \wishbone_LatchedTxLength_reg[13]/NET0131  , \wishbone_LatchedTxLength_reg[14]/NET0131  , \wishbone_LatchedTxLength_reg[15]/NET0131  , \wishbone_LatchedTxLength_reg[1]/NET0131  , \wishbone_LatchedTxLength_reg[2]/NET0131  , \wishbone_LatchedTxLength_reg[3]/NET0131  , \wishbone_LatchedTxLength_reg[4]/NET0131  , \wishbone_LatchedTxLength_reg[5]/NET0131  , \wishbone_LatchedTxLength_reg[6]/NET0131  , \wishbone_LatchedTxLength_reg[7]/NET0131  , \wishbone_LatchedTxLength_reg[8]/NET0131  , \wishbone_LatchedTxLength_reg[9]/NET0131  , \wishbone_MasterWbRX_reg/NET0131  , \wishbone_MasterWbTX_reg/NET0131  , \wishbone_ReadTxDataFromFifo_sync2_reg/NET0131  , \wishbone_ReadTxDataFromFifo_sync3_reg/NET0131  , \wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131  , \wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131  , \wishbone_ReadTxDataFromFifo_tck_reg/NET0131  , \wishbone_ReadTxDataFromMemory_reg/NET0131  , \wishbone_RxAbortLatched_reg/NET0131  , \wishbone_RxAbortSync2_reg/NET0131  , \wishbone_RxAbortSync3_reg/NET0131  , \wishbone_RxAbortSync4_reg/NET0131  , \wishbone_RxAbortSyncb2_reg/NET0131  , \wishbone_RxBDAddress_reg[1]/NET0131  , \wishbone_RxBDAddress_reg[2]/NET0131  , \wishbone_RxBDAddress_reg[3]/NET0131  , \wishbone_RxBDAddress_reg[4]/NET0131  , \wishbone_RxBDAddress_reg[5]/NET0131  , \wishbone_RxBDAddress_reg[6]/NET0131  , \wishbone_RxBDAddress_reg[7]/NET0131  , \wishbone_RxBDRead_reg/NET0131  , \wishbone_RxBDReady_reg/NET0131  , \wishbone_RxB_IRQ_reg/NET0131  , \wishbone_RxByteCnt_reg[0]/NET0131  , \wishbone_RxByteCnt_reg[1]/NET0131  , \wishbone_RxDataLatched1_reg[10]/NET0131  , \wishbone_RxDataLatched1_reg[11]/NET0131  , \wishbone_RxDataLatched1_reg[12]/NET0131  , \wishbone_RxDataLatched1_reg[13]/NET0131  , \wishbone_RxDataLatched1_reg[14]/NET0131  , \wishbone_RxDataLatched1_reg[15]/NET0131  , \wishbone_RxDataLatched1_reg[16]/NET0131  , \wishbone_RxDataLatched1_reg[17]/NET0131  , \wishbone_RxDataLatched1_reg[18]/NET0131  , \wishbone_RxDataLatched1_reg[19]/NET0131  , \wishbone_RxDataLatched1_reg[20]/NET0131  , \wishbone_RxDataLatched1_reg[21]/NET0131  , \wishbone_RxDataLatched1_reg[22]/NET0131  , \wishbone_RxDataLatched1_reg[23]/NET0131  , \wishbone_RxDataLatched1_reg[24]/NET0131  , \wishbone_RxDataLatched1_reg[25]/NET0131  , \wishbone_RxDataLatched1_reg[26]/NET0131  , \wishbone_RxDataLatched1_reg[27]/NET0131  , \wishbone_RxDataLatched1_reg[28]/NET0131  , \wishbone_RxDataLatched1_reg[29]/NET0131  , \wishbone_RxDataLatched1_reg[30]/NET0131  , \wishbone_RxDataLatched1_reg[31]/NET0131  , \wishbone_RxDataLatched1_reg[8]/NET0131  , \wishbone_RxDataLatched1_reg[9]/NET0131  , \wishbone_RxDataLatched2_reg[0]/NET0131  , \wishbone_RxDataLatched2_reg[10]/NET0131  , \wishbone_RxDataLatched2_reg[11]/NET0131  , \wishbone_RxDataLatched2_reg[12]/NET0131  , \wishbone_RxDataLatched2_reg[13]/NET0131  , \wishbone_RxDataLatched2_reg[14]/NET0131  , \wishbone_RxDataLatched2_reg[15]/NET0131  , \wishbone_RxDataLatched2_reg[16]/NET0131  , \wishbone_RxDataLatched2_reg[17]/NET0131  , \wishbone_RxDataLatched2_reg[18]/NET0131  , \wishbone_RxDataLatched2_reg[19]/NET0131  , \wishbone_RxDataLatched2_reg[1]/NET0131  , \wishbone_RxDataLatched2_reg[20]/NET0131  , \wishbone_RxDataLatched2_reg[21]/NET0131  , \wishbone_RxDataLatched2_reg[22]/NET0131  , \wishbone_RxDataLatched2_reg[23]/NET0131  , \wishbone_RxDataLatched2_reg[24]/NET0131  , \wishbone_RxDataLatched2_reg[25]/NET0131  , \wishbone_RxDataLatched2_reg[26]/NET0131  , \wishbone_RxDataLatched2_reg[27]/NET0131  , \wishbone_RxDataLatched2_reg[28]/NET0131  , \wishbone_RxDataLatched2_reg[29]/NET0131  , \wishbone_RxDataLatched2_reg[2]/NET0131  , \wishbone_RxDataLatched2_reg[30]/NET0131  , \wishbone_RxDataLatched2_reg[31]/NET0131  , \wishbone_RxDataLatched2_reg[3]/NET0131  , \wishbone_RxDataLatched2_reg[4]/NET0131  , \wishbone_RxDataLatched2_reg[5]/NET0131  , \wishbone_RxDataLatched2_reg[6]/NET0131  , \wishbone_RxDataLatched2_reg[7]/NET0131  , \wishbone_RxDataLatched2_reg[8]/NET0131  , \wishbone_RxDataLatched2_reg[9]/NET0131  , \wishbone_RxE_IRQ_reg/NET0131  , \wishbone_RxEn_needed_reg/NET0131  , \wishbone_RxEn_q_reg/NET0131  , \wishbone_RxEn_reg/NET0131  , \wishbone_RxEnableWindow_reg/NET0131  , \wishbone_RxOverrun_reg/NET0131  , \wishbone_RxPointerLSB_rst_reg[0]/NET0131  , \wishbone_RxPointerLSB_rst_reg[1]/NET0131  , \wishbone_RxPointerMSB_reg[10]/NET0131  , \wishbone_RxPointerMSB_reg[11]/NET0131  , \wishbone_RxPointerMSB_reg[12]/NET0131  , \wishbone_RxPointerMSB_reg[13]/NET0131  , \wishbone_RxPointerMSB_reg[14]/NET0131  , \wishbone_RxPointerMSB_reg[15]/NET0131  , \wishbone_RxPointerMSB_reg[16]/NET0131  , \wishbone_RxPointerMSB_reg[17]/NET0131  , \wishbone_RxPointerMSB_reg[18]/NET0131  , \wishbone_RxPointerMSB_reg[19]/NET0131  , \wishbone_RxPointerMSB_reg[20]/NET0131  , \wishbone_RxPointerMSB_reg[21]/NET0131  , \wishbone_RxPointerMSB_reg[22]/NET0131  , \wishbone_RxPointerMSB_reg[23]/NET0131  , \wishbone_RxPointerMSB_reg[24]/NET0131  , \wishbone_RxPointerMSB_reg[25]/NET0131  , \wishbone_RxPointerMSB_reg[26]/NET0131  , \wishbone_RxPointerMSB_reg[27]/NET0131  , \wishbone_RxPointerMSB_reg[28]/NET0131  , \wishbone_RxPointerMSB_reg[29]/NET0131  , \wishbone_RxPointerMSB_reg[2]/NET0131  , \wishbone_RxPointerMSB_reg[30]/NET0131  , \wishbone_RxPointerMSB_reg[31]/NET0131  , \wishbone_RxPointerMSB_reg[3]/NET0131  , \wishbone_RxPointerMSB_reg[4]/NET0131  , \wishbone_RxPointerMSB_reg[5]/NET0131  , \wishbone_RxPointerMSB_reg[6]/NET0131  , \wishbone_RxPointerMSB_reg[7]/NET0131  , \wishbone_RxPointerMSB_reg[8]/NET0131  , \wishbone_RxPointerMSB_reg[9]/NET0131  , \wishbone_RxPointerRead_reg/NET0131  , \wishbone_RxReady_reg/NET0131  , \wishbone_RxStatusInLatched_reg[0]/NET0131  , \wishbone_RxStatusInLatched_reg[1]/NET0131  , \wishbone_RxStatusInLatched_reg[2]/NET0131  , \wishbone_RxStatusInLatched_reg[3]/NET0131  , \wishbone_RxStatusInLatched_reg[4]/NET0131  , \wishbone_RxStatusInLatched_reg[5]/NET0131  , \wishbone_RxStatusInLatched_reg[6]/NET0131  , \wishbone_RxStatusInLatched_reg[7]/NET0131  , \wishbone_RxStatusInLatched_reg[8]/NET0131  , \wishbone_RxStatusWriteLatched_reg/NET0131  , \wishbone_RxStatusWriteLatched_sync2_reg/NET0131  , \wishbone_RxStatusWriteLatched_syncb2_reg/NET0131  , \wishbone_RxStatus_reg[13]/NET0131  , \wishbone_RxStatus_reg[14]/NET0131  , \wishbone_RxValidBytes_reg[0]/NET0131  , \wishbone_RxValidBytes_reg[1]/NET0131  , \wishbone_ShiftEndedSync1_reg/NET0131  , \wishbone_ShiftEndedSync2_reg/NET0131  , \wishbone_ShiftEndedSync3_reg/NET0131  , \wishbone_ShiftEndedSync_c1_reg/NET0131  , \wishbone_ShiftEndedSync_c2_reg/NET0131  , \wishbone_ShiftEnded_rck_reg/NET0131  , \wishbone_ShiftEnded_reg/NET0131  , \wishbone_ShiftWillEnd_reg/NET0131  , \wishbone_StartOccured_reg/NET0131  , \wishbone_SyncRxStartFrm_q2_reg/NET0131  , \wishbone_SyncRxStartFrm_q_reg/NET0131  , \wishbone_TxAbortPacketBlocked_reg/NET0131  , \wishbone_TxAbortPacket_NotCleared_reg/NET0131  , \wishbone_TxAbortPacket_reg/NET0131  , \wishbone_TxAbort_q_reg/NET0131  , \wishbone_TxAbort_wb_q_reg/NET0131  , \wishbone_TxAbort_wb_reg/NET0131  , \wishbone_TxBDAddress_reg[1]/NET0131  , \wishbone_TxBDAddress_reg[2]/NET0131  , \wishbone_TxBDAddress_reg[3]/NET0131  , \wishbone_TxBDAddress_reg[4]/NET0131  , \wishbone_TxBDAddress_reg[5]/NET0131  , \wishbone_TxBDAddress_reg[6]/NET0131  , \wishbone_TxBDAddress_reg[7]/NET0131  , \wishbone_TxBDRead_reg/NET0131  , \wishbone_TxBDReady_reg/NET0131  , \wishbone_TxB_IRQ_reg/NET0131  , \wishbone_TxByteCnt_reg[0]/NET0131  , \wishbone_TxByteCnt_reg[1]/NET0131  , \wishbone_TxDataLatched_reg[0]/NET0131  , \wishbone_TxDataLatched_reg[10]/NET0131  , \wishbone_TxDataLatched_reg[11]/NET0131  , \wishbone_TxDataLatched_reg[12]/NET0131  , \wishbone_TxDataLatched_reg[13]/NET0131  , \wishbone_TxDataLatched_reg[14]/NET0131  , \wishbone_TxDataLatched_reg[15]/NET0131  , \wishbone_TxDataLatched_reg[16]/NET0131  , \wishbone_TxDataLatched_reg[17]/NET0131  , \wishbone_TxDataLatched_reg[18]/NET0131  , \wishbone_TxDataLatched_reg[19]/NET0131  , \wishbone_TxDataLatched_reg[1]/NET0131  , \wishbone_TxDataLatched_reg[20]/NET0131  , \wishbone_TxDataLatched_reg[21]/NET0131  , \wishbone_TxDataLatched_reg[22]/NET0131  , \wishbone_TxDataLatched_reg[23]/NET0131  , \wishbone_TxDataLatched_reg[24]/NET0131  , \wishbone_TxDataLatched_reg[25]/NET0131  , \wishbone_TxDataLatched_reg[26]/NET0131  , \wishbone_TxDataLatched_reg[27]/NET0131  , \wishbone_TxDataLatched_reg[28]/NET0131  , \wishbone_TxDataLatched_reg[29]/NET0131  , \wishbone_TxDataLatched_reg[2]/NET0131  , \wishbone_TxDataLatched_reg[30]/NET0131  , \wishbone_TxDataLatched_reg[31]/NET0131  , \wishbone_TxDataLatched_reg[3]/NET0131  , \wishbone_TxDataLatched_reg[4]/NET0131  , \wishbone_TxDataLatched_reg[5]/NET0131  , \wishbone_TxDataLatched_reg[6]/NET0131  , \wishbone_TxDataLatched_reg[7]/NET0131  , \wishbone_TxDataLatched_reg[8]/NET0131  , \wishbone_TxDataLatched_reg[9]/NET0131  , \wishbone_TxData_reg[0]/NET0131  , \wishbone_TxData_reg[1]/NET0131  , \wishbone_TxData_reg[2]/NET0131  , \wishbone_TxData_reg[3]/NET0131  , \wishbone_TxData_reg[4]/NET0131  , \wishbone_TxData_reg[5]/NET0131  , \wishbone_TxData_reg[6]/NET0131  , \wishbone_TxData_reg[7]/NET0131  , \wishbone_TxDonePacketBlocked_reg/NET0131  , \wishbone_TxDonePacket_NotCleared_reg/NET0131  , \wishbone_TxDonePacket_reg/NET0131  , \wishbone_TxDone_wb_q_reg/NET0131  , \wishbone_TxDone_wb_reg/NET0131  , \wishbone_TxE_IRQ_reg/NET0131  , \wishbone_TxEn_needed_reg/NET0131  , \wishbone_TxEn_q_reg/NET0131  , \wishbone_TxEn_reg/NET0131  , \wishbone_TxEndFrm_reg/NET0131  , \wishbone_TxEndFrm_wb_reg/NET0131  , \wishbone_TxLength_reg[0]/NET0131  , \wishbone_TxLength_reg[10]/NET0131  , \wishbone_TxLength_reg[11]/NET0131  , \wishbone_TxLength_reg[12]/NET0131  , \wishbone_TxLength_reg[13]/NET0131  , \wishbone_TxLength_reg[14]/NET0131  , \wishbone_TxLength_reg[15]/NET0131  , \wishbone_TxLength_reg[1]/NET0131  , \wishbone_TxLength_reg[2]/NET0131  , \wishbone_TxLength_reg[3]/NET0131  , \wishbone_TxLength_reg[4]/NET0131  , \wishbone_TxLength_reg[5]/NET0131  , \wishbone_TxLength_reg[6]/NET0131  , \wishbone_TxLength_reg[7]/NET0131  , \wishbone_TxLength_reg[8]/NET0131  , \wishbone_TxLength_reg[9]/NET0131  , \wishbone_TxPointerLSB_reg[0]/NET0131  , \wishbone_TxPointerLSB_reg[1]/NET0131  , \wishbone_TxPointerLSB_rst_reg[0]/NET0131  , \wishbone_TxPointerLSB_rst_reg[1]/NET0131  , \wishbone_TxPointerMSB_reg[10]/NET0131  , \wishbone_TxPointerMSB_reg[11]/NET0131  , \wishbone_TxPointerMSB_reg[12]/NET0131  , \wishbone_TxPointerMSB_reg[13]/NET0131  , \wishbone_TxPointerMSB_reg[14]/NET0131  , \wishbone_TxPointerMSB_reg[15]/NET0131  , \wishbone_TxPointerMSB_reg[16]/NET0131  , \wishbone_TxPointerMSB_reg[17]/NET0131  , \wishbone_TxPointerMSB_reg[18]/NET0131  , \wishbone_TxPointerMSB_reg[19]/NET0131  , \wishbone_TxPointerMSB_reg[20]/NET0131  , \wishbone_TxPointerMSB_reg[21]/NET0131  , \wishbone_TxPointerMSB_reg[22]/NET0131  , \wishbone_TxPointerMSB_reg[23]/NET0131  , \wishbone_TxPointerMSB_reg[24]/NET0131  , \wishbone_TxPointerMSB_reg[25]/NET0131  , \wishbone_TxPointerMSB_reg[26]/NET0131  , \wishbone_TxPointerMSB_reg[27]/NET0131  , \wishbone_TxPointerMSB_reg[28]/NET0131  , \wishbone_TxPointerMSB_reg[29]/NET0131  , \wishbone_TxPointerMSB_reg[2]/NET0131  , \wishbone_TxPointerMSB_reg[30]/NET0131  , \wishbone_TxPointerMSB_reg[31]/NET0131  , \wishbone_TxPointerMSB_reg[3]/NET0131  , \wishbone_TxPointerMSB_reg[4]/NET0131  , \wishbone_TxPointerMSB_reg[5]/NET0131  , \wishbone_TxPointerMSB_reg[6]/NET0131  , \wishbone_TxPointerMSB_reg[7]/NET0131  , \wishbone_TxPointerMSB_reg[8]/NET0131  , \wishbone_TxPointerMSB_reg[9]/NET0131  , \wishbone_TxPointerRead_reg/NET0131  , \wishbone_TxRetryPacketBlocked_reg/NET0131  , \wishbone_TxRetryPacket_NotCleared_reg/NET0131  , \wishbone_TxRetryPacket_reg/NET0131  , \wishbone_TxRetry_q_reg/NET0131  , \wishbone_TxRetry_wb_q_reg/NET0131  , \wishbone_TxRetry_wb_reg/NET0131  , \wishbone_TxStartFrm_reg/NET0131  , \wishbone_TxStartFrm_sync2_reg/NET0131  , \wishbone_TxStartFrm_syncb2_reg/NET0131  , \wishbone_TxStartFrm_wb_reg/NET0131  , \wishbone_TxStatus_reg[11]/NET0131  , \wishbone_TxStatus_reg[12]/NET0131  , \wishbone_TxStatus_reg[13]/NET0131  , \wishbone_TxStatus_reg[14]/NET0131  , \wishbone_TxUnderRun_reg/NET0131  , \wishbone_TxUnderRun_sync1_reg/NET0131  , \wishbone_TxUnderRun_wb_reg/NET0131  , \wishbone_TxUsedData_q_reg/NET0131  , \wishbone_TxValidBytesLatched_reg[0]/NET0131  , \wishbone_TxValidBytesLatched_reg[1]/NET0131  , \wishbone_WB_ACK_O_reg/P0001  , \wishbone_WbEn_q_reg/NET0131  , \wishbone_WbEn_reg/NET0131  , \wishbone_WriteRxDataToFifoSync2_reg/NET0131  , \wishbone_WriteRxDataToFifoSync3_reg/NET0131  , \wishbone_WriteRxDataToFifo_reg/NET0131  , \wishbone_bd_ram_mem0_reg[0][0]/P0001  , \wishbone_bd_ram_mem0_reg[0][1]/P0001  , \wishbone_bd_ram_mem0_reg[0][2]/P0001  , \wishbone_bd_ram_mem0_reg[0][3]/P0001  , \wishbone_bd_ram_mem0_reg[0][4]/P0001  , \wishbone_bd_ram_mem0_reg[0][5]/P0001  , \wishbone_bd_ram_mem0_reg[0][6]/P0001  , \wishbone_bd_ram_mem0_reg[0][7]/P0001  , \wishbone_bd_ram_mem0_reg[100][0]/P0001  , \wishbone_bd_ram_mem0_reg[100][1]/P0001  , \wishbone_bd_ram_mem0_reg[100][2]/P0001  , \wishbone_bd_ram_mem0_reg[100][3]/P0001  , \wishbone_bd_ram_mem0_reg[100][4]/P0001  , \wishbone_bd_ram_mem0_reg[100][5]/P0001  , \wishbone_bd_ram_mem0_reg[100][6]/P0001  , \wishbone_bd_ram_mem0_reg[100][7]/P0001  , \wishbone_bd_ram_mem0_reg[101][0]/P0001  , \wishbone_bd_ram_mem0_reg[101][1]/P0001  , \wishbone_bd_ram_mem0_reg[101][2]/P0001  , \wishbone_bd_ram_mem0_reg[101][3]/P0001  , \wishbone_bd_ram_mem0_reg[101][4]/P0001  , \wishbone_bd_ram_mem0_reg[101][5]/P0001  , \wishbone_bd_ram_mem0_reg[101][6]/P0001  , \wishbone_bd_ram_mem0_reg[101][7]/P0001  , \wishbone_bd_ram_mem0_reg[102][0]/P0001  , \wishbone_bd_ram_mem0_reg[102][1]/P0001  , \wishbone_bd_ram_mem0_reg[102][2]/P0001  , \wishbone_bd_ram_mem0_reg[102][3]/P0001  , \wishbone_bd_ram_mem0_reg[102][4]/P0001  , \wishbone_bd_ram_mem0_reg[102][5]/P0001  , \wishbone_bd_ram_mem0_reg[102][6]/P0001  , \wishbone_bd_ram_mem0_reg[102][7]/P0001  , \wishbone_bd_ram_mem0_reg[103][0]/P0001  , \wishbone_bd_ram_mem0_reg[103][1]/P0001  , \wishbone_bd_ram_mem0_reg[103][2]/P0001  , \wishbone_bd_ram_mem0_reg[103][3]/P0001  , \wishbone_bd_ram_mem0_reg[103][4]/P0001  , \wishbone_bd_ram_mem0_reg[103][5]/P0001  , \wishbone_bd_ram_mem0_reg[103][6]/P0001  , \wishbone_bd_ram_mem0_reg[103][7]/P0001  , \wishbone_bd_ram_mem0_reg[104][0]/P0001  , \wishbone_bd_ram_mem0_reg[104][1]/P0001  , \wishbone_bd_ram_mem0_reg[104][2]/P0001  , \wishbone_bd_ram_mem0_reg[104][3]/P0001  , \wishbone_bd_ram_mem0_reg[104][4]/P0001  , \wishbone_bd_ram_mem0_reg[104][5]/P0001  , \wishbone_bd_ram_mem0_reg[104][6]/P0001  , \wishbone_bd_ram_mem0_reg[104][7]/P0001  , \wishbone_bd_ram_mem0_reg[105][0]/P0001  , \wishbone_bd_ram_mem0_reg[105][1]/P0001  , \wishbone_bd_ram_mem0_reg[105][2]/P0001  , \wishbone_bd_ram_mem0_reg[105][3]/P0001  , \wishbone_bd_ram_mem0_reg[105][4]/P0001  , \wishbone_bd_ram_mem0_reg[105][5]/P0001  , \wishbone_bd_ram_mem0_reg[105][6]/P0001  , \wishbone_bd_ram_mem0_reg[105][7]/P0001  , \wishbone_bd_ram_mem0_reg[106][0]/P0001  , \wishbone_bd_ram_mem0_reg[106][1]/P0001  , \wishbone_bd_ram_mem0_reg[106][2]/P0001  , \wishbone_bd_ram_mem0_reg[106][3]/P0001  , \wishbone_bd_ram_mem0_reg[106][4]/P0001  , \wishbone_bd_ram_mem0_reg[106][5]/P0001  , \wishbone_bd_ram_mem0_reg[106][6]/P0001  , \wishbone_bd_ram_mem0_reg[106][7]/P0001  , \wishbone_bd_ram_mem0_reg[107][0]/P0001  , \wishbone_bd_ram_mem0_reg[107][1]/P0001  , \wishbone_bd_ram_mem0_reg[107][2]/P0001  , \wishbone_bd_ram_mem0_reg[107][3]/P0001  , \wishbone_bd_ram_mem0_reg[107][4]/P0001  , \wishbone_bd_ram_mem0_reg[107][5]/P0001  , \wishbone_bd_ram_mem0_reg[107][6]/P0001  , \wishbone_bd_ram_mem0_reg[107][7]/P0001  , \wishbone_bd_ram_mem0_reg[108][0]/P0001  , \wishbone_bd_ram_mem0_reg[108][1]/P0001  , \wishbone_bd_ram_mem0_reg[108][2]/P0001  , \wishbone_bd_ram_mem0_reg[108][3]/P0001  , \wishbone_bd_ram_mem0_reg[108][4]/P0001  , \wishbone_bd_ram_mem0_reg[108][5]/P0001  , \wishbone_bd_ram_mem0_reg[108][6]/P0001  , \wishbone_bd_ram_mem0_reg[108][7]/P0001  , \wishbone_bd_ram_mem0_reg[109][0]/P0001  , \wishbone_bd_ram_mem0_reg[109][1]/P0001  , \wishbone_bd_ram_mem0_reg[109][2]/P0001  , \wishbone_bd_ram_mem0_reg[109][3]/P0001  , \wishbone_bd_ram_mem0_reg[109][4]/P0001  , \wishbone_bd_ram_mem0_reg[109][5]/P0001  , \wishbone_bd_ram_mem0_reg[109][6]/P0001  , \wishbone_bd_ram_mem0_reg[109][7]/P0001  , \wishbone_bd_ram_mem0_reg[10][0]/P0001  , \wishbone_bd_ram_mem0_reg[10][1]/P0001  , \wishbone_bd_ram_mem0_reg[10][2]/P0001  , \wishbone_bd_ram_mem0_reg[10][3]/P0001  , \wishbone_bd_ram_mem0_reg[10][4]/P0001  , \wishbone_bd_ram_mem0_reg[10][5]/P0001  , \wishbone_bd_ram_mem0_reg[10][6]/P0001  , \wishbone_bd_ram_mem0_reg[10][7]/P0001  , \wishbone_bd_ram_mem0_reg[110][0]/P0001  , \wishbone_bd_ram_mem0_reg[110][1]/P0001  , \wishbone_bd_ram_mem0_reg[110][2]/P0001  , \wishbone_bd_ram_mem0_reg[110][3]/P0001  , \wishbone_bd_ram_mem0_reg[110][4]/P0001  , \wishbone_bd_ram_mem0_reg[110][5]/P0001  , \wishbone_bd_ram_mem0_reg[110][6]/P0001  , \wishbone_bd_ram_mem0_reg[110][7]/P0001  , \wishbone_bd_ram_mem0_reg[111][0]/P0001  , \wishbone_bd_ram_mem0_reg[111][1]/P0001  , \wishbone_bd_ram_mem0_reg[111][2]/P0001  , \wishbone_bd_ram_mem0_reg[111][3]/P0001  , \wishbone_bd_ram_mem0_reg[111][4]/P0001  , \wishbone_bd_ram_mem0_reg[111][5]/P0001  , \wishbone_bd_ram_mem0_reg[111][6]/P0001  , \wishbone_bd_ram_mem0_reg[111][7]/P0001  , \wishbone_bd_ram_mem0_reg[112][0]/P0001  , \wishbone_bd_ram_mem0_reg[112][1]/P0001  , \wishbone_bd_ram_mem0_reg[112][2]/P0001  , \wishbone_bd_ram_mem0_reg[112][3]/P0001  , \wishbone_bd_ram_mem0_reg[112][4]/P0001  , \wishbone_bd_ram_mem0_reg[112][5]/P0001  , \wishbone_bd_ram_mem0_reg[112][6]/P0001  , \wishbone_bd_ram_mem0_reg[112][7]/P0001  , \wishbone_bd_ram_mem0_reg[113][0]/P0001  , \wishbone_bd_ram_mem0_reg[113][1]/P0001  , \wishbone_bd_ram_mem0_reg[113][2]/P0001  , \wishbone_bd_ram_mem0_reg[113][3]/P0001  , \wishbone_bd_ram_mem0_reg[113][4]/P0001  , \wishbone_bd_ram_mem0_reg[113][5]/P0001  , \wishbone_bd_ram_mem0_reg[113][6]/P0001  , \wishbone_bd_ram_mem0_reg[113][7]/P0001  , \wishbone_bd_ram_mem0_reg[114][0]/P0001  , \wishbone_bd_ram_mem0_reg[114][1]/P0001  , \wishbone_bd_ram_mem0_reg[114][2]/P0001  , \wishbone_bd_ram_mem0_reg[114][3]/P0001  , \wishbone_bd_ram_mem0_reg[114][4]/P0001  , \wishbone_bd_ram_mem0_reg[114][5]/P0001  , \wishbone_bd_ram_mem0_reg[114][6]/P0001  , \wishbone_bd_ram_mem0_reg[114][7]/P0001  , \wishbone_bd_ram_mem0_reg[115][0]/P0001  , \wishbone_bd_ram_mem0_reg[115][1]/P0001  , \wishbone_bd_ram_mem0_reg[115][2]/P0001  , \wishbone_bd_ram_mem0_reg[115][3]/P0001  , \wishbone_bd_ram_mem0_reg[115][4]/P0001  , \wishbone_bd_ram_mem0_reg[115][5]/P0001  , \wishbone_bd_ram_mem0_reg[115][6]/P0001  , \wishbone_bd_ram_mem0_reg[115][7]/P0001  , \wishbone_bd_ram_mem0_reg[116][0]/P0001  , \wishbone_bd_ram_mem0_reg[116][1]/P0001  , \wishbone_bd_ram_mem0_reg[116][2]/P0001  , \wishbone_bd_ram_mem0_reg[116][3]/P0001  , \wishbone_bd_ram_mem0_reg[116][4]/P0001  , \wishbone_bd_ram_mem0_reg[116][5]/P0001  , \wishbone_bd_ram_mem0_reg[116][6]/P0001  , \wishbone_bd_ram_mem0_reg[116][7]/P0001  , \wishbone_bd_ram_mem0_reg[117][0]/P0001  , \wishbone_bd_ram_mem0_reg[117][1]/P0001  , \wishbone_bd_ram_mem0_reg[117][2]/P0001  , \wishbone_bd_ram_mem0_reg[117][3]/P0001  , \wishbone_bd_ram_mem0_reg[117][4]/P0001  , \wishbone_bd_ram_mem0_reg[117][5]/P0001  , \wishbone_bd_ram_mem0_reg[117][6]/P0001  , \wishbone_bd_ram_mem0_reg[117][7]/P0001  , \wishbone_bd_ram_mem0_reg[118][0]/P0001  , \wishbone_bd_ram_mem0_reg[118][1]/P0001  , \wishbone_bd_ram_mem0_reg[118][2]/P0001  , \wishbone_bd_ram_mem0_reg[118][3]/P0001  , \wishbone_bd_ram_mem0_reg[118][4]/P0001  , \wishbone_bd_ram_mem0_reg[118][5]/P0001  , \wishbone_bd_ram_mem0_reg[118][6]/P0001  , \wishbone_bd_ram_mem0_reg[118][7]/P0001  , \wishbone_bd_ram_mem0_reg[119][0]/P0001  , \wishbone_bd_ram_mem0_reg[119][1]/P0001  , \wishbone_bd_ram_mem0_reg[119][2]/P0001  , \wishbone_bd_ram_mem0_reg[119][3]/P0001  , \wishbone_bd_ram_mem0_reg[119][4]/P0001  , \wishbone_bd_ram_mem0_reg[119][5]/P0001  , \wishbone_bd_ram_mem0_reg[119][6]/P0001  , \wishbone_bd_ram_mem0_reg[119][7]/P0001  , \wishbone_bd_ram_mem0_reg[11][0]/P0001  , \wishbone_bd_ram_mem0_reg[11][1]/P0001  , \wishbone_bd_ram_mem0_reg[11][2]/P0001  , \wishbone_bd_ram_mem0_reg[11][3]/P0001  , \wishbone_bd_ram_mem0_reg[11][4]/P0001  , \wishbone_bd_ram_mem0_reg[11][5]/P0001  , \wishbone_bd_ram_mem0_reg[11][6]/P0001  , \wishbone_bd_ram_mem0_reg[11][7]/P0001  , \wishbone_bd_ram_mem0_reg[120][0]/P0001  , \wishbone_bd_ram_mem0_reg[120][1]/P0001  , \wishbone_bd_ram_mem0_reg[120][2]/P0001  , \wishbone_bd_ram_mem0_reg[120][3]/P0001  , \wishbone_bd_ram_mem0_reg[120][4]/P0001  , \wishbone_bd_ram_mem0_reg[120][5]/P0001  , \wishbone_bd_ram_mem0_reg[120][6]/P0001  , \wishbone_bd_ram_mem0_reg[120][7]/P0001  , \wishbone_bd_ram_mem0_reg[121][0]/P0001  , \wishbone_bd_ram_mem0_reg[121][1]/P0001  , \wishbone_bd_ram_mem0_reg[121][2]/P0001  , \wishbone_bd_ram_mem0_reg[121][3]/P0001  , \wishbone_bd_ram_mem0_reg[121][4]/P0001  , \wishbone_bd_ram_mem0_reg[121][5]/P0001  , \wishbone_bd_ram_mem0_reg[121][6]/P0001  , \wishbone_bd_ram_mem0_reg[121][7]/P0001  , \wishbone_bd_ram_mem0_reg[122][0]/P0001  , \wishbone_bd_ram_mem0_reg[122][1]/P0001  , \wishbone_bd_ram_mem0_reg[122][2]/P0001  , \wishbone_bd_ram_mem0_reg[122][3]/P0001  , \wishbone_bd_ram_mem0_reg[122][4]/P0001  , \wishbone_bd_ram_mem0_reg[122][5]/P0001  , \wishbone_bd_ram_mem0_reg[122][6]/P0001  , \wishbone_bd_ram_mem0_reg[122][7]/P0001  , \wishbone_bd_ram_mem0_reg[123][0]/P0001  , \wishbone_bd_ram_mem0_reg[123][1]/P0001  , \wishbone_bd_ram_mem0_reg[123][2]/P0001  , \wishbone_bd_ram_mem0_reg[123][3]/P0001  , \wishbone_bd_ram_mem0_reg[123][4]/P0001  , \wishbone_bd_ram_mem0_reg[123][5]/P0001  , \wishbone_bd_ram_mem0_reg[123][6]/P0001  , \wishbone_bd_ram_mem0_reg[123][7]/P0001  , \wishbone_bd_ram_mem0_reg[124][0]/P0001  , \wishbone_bd_ram_mem0_reg[124][1]/P0001  , \wishbone_bd_ram_mem0_reg[124][2]/P0001  , \wishbone_bd_ram_mem0_reg[124][3]/P0001  , \wishbone_bd_ram_mem0_reg[124][4]/P0001  , \wishbone_bd_ram_mem0_reg[124][5]/P0001  , \wishbone_bd_ram_mem0_reg[124][6]/P0001  , \wishbone_bd_ram_mem0_reg[124][7]/P0001  , \wishbone_bd_ram_mem0_reg[125][0]/P0001  , \wishbone_bd_ram_mem0_reg[125][1]/P0001  , \wishbone_bd_ram_mem0_reg[125][2]/P0001  , \wishbone_bd_ram_mem0_reg[125][3]/P0001  , \wishbone_bd_ram_mem0_reg[125][4]/P0001  , \wishbone_bd_ram_mem0_reg[125][5]/P0001  , \wishbone_bd_ram_mem0_reg[125][6]/P0001  , \wishbone_bd_ram_mem0_reg[125][7]/P0001  , \wishbone_bd_ram_mem0_reg[126][0]/P0001  , \wishbone_bd_ram_mem0_reg[126][1]/P0001  , \wishbone_bd_ram_mem0_reg[126][2]/P0001  , \wishbone_bd_ram_mem0_reg[126][3]/P0001  , \wishbone_bd_ram_mem0_reg[126][4]/P0001  , \wishbone_bd_ram_mem0_reg[126][5]/P0001  , \wishbone_bd_ram_mem0_reg[126][6]/P0001  , \wishbone_bd_ram_mem0_reg[126][7]/P0001  , \wishbone_bd_ram_mem0_reg[127][0]/P0001  , \wishbone_bd_ram_mem0_reg[127][1]/P0001  , \wishbone_bd_ram_mem0_reg[127][2]/P0001  , \wishbone_bd_ram_mem0_reg[127][3]/P0001  , \wishbone_bd_ram_mem0_reg[127][4]/P0001  , \wishbone_bd_ram_mem0_reg[127][5]/P0001  , \wishbone_bd_ram_mem0_reg[127][6]/P0001  , \wishbone_bd_ram_mem0_reg[127][7]/P0001  , \wishbone_bd_ram_mem0_reg[128][0]/P0001  , \wishbone_bd_ram_mem0_reg[128][1]/P0001  , \wishbone_bd_ram_mem0_reg[128][2]/P0001  , \wishbone_bd_ram_mem0_reg[128][3]/P0001  , \wishbone_bd_ram_mem0_reg[128][4]/P0001  , \wishbone_bd_ram_mem0_reg[128][5]/P0001  , \wishbone_bd_ram_mem0_reg[128][6]/P0001  , \wishbone_bd_ram_mem0_reg[128][7]/P0001  , \wishbone_bd_ram_mem0_reg[129][0]/P0001  , \wishbone_bd_ram_mem0_reg[129][1]/P0001  , \wishbone_bd_ram_mem0_reg[129][2]/P0001  , \wishbone_bd_ram_mem0_reg[129][3]/P0001  , \wishbone_bd_ram_mem0_reg[129][4]/P0001  , \wishbone_bd_ram_mem0_reg[129][5]/P0001  , \wishbone_bd_ram_mem0_reg[129][6]/P0001  , \wishbone_bd_ram_mem0_reg[129][7]/P0001  , \wishbone_bd_ram_mem0_reg[12][0]/P0001  , \wishbone_bd_ram_mem0_reg[12][1]/P0001  , \wishbone_bd_ram_mem0_reg[12][2]/P0001  , \wishbone_bd_ram_mem0_reg[12][3]/P0001  , \wishbone_bd_ram_mem0_reg[12][4]/P0001  , \wishbone_bd_ram_mem0_reg[12][5]/P0001  , \wishbone_bd_ram_mem0_reg[12][6]/P0001  , \wishbone_bd_ram_mem0_reg[12][7]/P0001  , \wishbone_bd_ram_mem0_reg[130][0]/P0001  , \wishbone_bd_ram_mem0_reg[130][1]/P0001  , \wishbone_bd_ram_mem0_reg[130][2]/P0001  , \wishbone_bd_ram_mem0_reg[130][3]/P0001  , \wishbone_bd_ram_mem0_reg[130][4]/P0001  , \wishbone_bd_ram_mem0_reg[130][5]/P0001  , \wishbone_bd_ram_mem0_reg[130][6]/P0001  , \wishbone_bd_ram_mem0_reg[130][7]/P0001  , \wishbone_bd_ram_mem0_reg[131][0]/P0001  , \wishbone_bd_ram_mem0_reg[131][1]/P0001  , \wishbone_bd_ram_mem0_reg[131][2]/P0001  , \wishbone_bd_ram_mem0_reg[131][3]/P0001  , \wishbone_bd_ram_mem0_reg[131][4]/P0001  , \wishbone_bd_ram_mem0_reg[131][5]/P0001  , \wishbone_bd_ram_mem0_reg[131][6]/P0001  , \wishbone_bd_ram_mem0_reg[131][7]/P0001  , \wishbone_bd_ram_mem0_reg[132][0]/P0001  , \wishbone_bd_ram_mem0_reg[132][1]/P0001  , \wishbone_bd_ram_mem0_reg[132][2]/P0001  , \wishbone_bd_ram_mem0_reg[132][3]/P0001  , \wishbone_bd_ram_mem0_reg[132][4]/P0001  , \wishbone_bd_ram_mem0_reg[132][5]/P0001  , \wishbone_bd_ram_mem0_reg[132][6]/P0001  , \wishbone_bd_ram_mem0_reg[132][7]/P0001  , \wishbone_bd_ram_mem0_reg[133][0]/P0001  , \wishbone_bd_ram_mem0_reg[133][1]/P0001  , \wishbone_bd_ram_mem0_reg[133][2]/P0001  , \wishbone_bd_ram_mem0_reg[133][3]/P0001  , \wishbone_bd_ram_mem0_reg[133][4]/P0001  , \wishbone_bd_ram_mem0_reg[133][5]/P0001  , \wishbone_bd_ram_mem0_reg[133][6]/P0001  , \wishbone_bd_ram_mem0_reg[133][7]/P0001  , \wishbone_bd_ram_mem0_reg[134][0]/P0001  , \wishbone_bd_ram_mem0_reg[134][1]/P0001  , \wishbone_bd_ram_mem0_reg[134][2]/P0001  , \wishbone_bd_ram_mem0_reg[134][3]/P0001  , \wishbone_bd_ram_mem0_reg[134][4]/P0001  , \wishbone_bd_ram_mem0_reg[134][5]/P0001  , \wishbone_bd_ram_mem0_reg[134][6]/P0001  , \wishbone_bd_ram_mem0_reg[134][7]/P0001  , \wishbone_bd_ram_mem0_reg[135][0]/P0001  , \wishbone_bd_ram_mem0_reg[135][1]/P0001  , \wishbone_bd_ram_mem0_reg[135][2]/P0001  , \wishbone_bd_ram_mem0_reg[135][3]/P0001  , \wishbone_bd_ram_mem0_reg[135][4]/P0001  , \wishbone_bd_ram_mem0_reg[135][5]/P0001  , \wishbone_bd_ram_mem0_reg[135][6]/P0001  , \wishbone_bd_ram_mem0_reg[135][7]/P0001  , \wishbone_bd_ram_mem0_reg[136][0]/P0001  , \wishbone_bd_ram_mem0_reg[136][1]/P0001  , \wishbone_bd_ram_mem0_reg[136][2]/P0001  , \wishbone_bd_ram_mem0_reg[136][3]/P0001  , \wishbone_bd_ram_mem0_reg[136][4]/P0001  , \wishbone_bd_ram_mem0_reg[136][5]/P0001  , \wishbone_bd_ram_mem0_reg[136][6]/P0001  , \wishbone_bd_ram_mem0_reg[136][7]/P0001  , \wishbone_bd_ram_mem0_reg[137][0]/P0001  , \wishbone_bd_ram_mem0_reg[137][1]/P0001  , \wishbone_bd_ram_mem0_reg[137][2]/P0001  , \wishbone_bd_ram_mem0_reg[137][3]/P0001  , \wishbone_bd_ram_mem0_reg[137][4]/P0001  , \wishbone_bd_ram_mem0_reg[137][5]/P0001  , \wishbone_bd_ram_mem0_reg[137][6]/P0001  , \wishbone_bd_ram_mem0_reg[137][7]/P0001  , \wishbone_bd_ram_mem0_reg[138][0]/P0001  , \wishbone_bd_ram_mem0_reg[138][1]/P0001  , \wishbone_bd_ram_mem0_reg[138][2]/P0001  , \wishbone_bd_ram_mem0_reg[138][3]/P0001  , \wishbone_bd_ram_mem0_reg[138][4]/P0001  , \wishbone_bd_ram_mem0_reg[138][5]/P0001  , \wishbone_bd_ram_mem0_reg[138][6]/P0001  , \wishbone_bd_ram_mem0_reg[138][7]/P0001  , \wishbone_bd_ram_mem0_reg[139][0]/P0001  , \wishbone_bd_ram_mem0_reg[139][1]/P0001  , \wishbone_bd_ram_mem0_reg[139][2]/P0001  , \wishbone_bd_ram_mem0_reg[139][3]/P0001  , \wishbone_bd_ram_mem0_reg[139][4]/P0001  , \wishbone_bd_ram_mem0_reg[139][5]/P0001  , \wishbone_bd_ram_mem0_reg[139][6]/P0001  , \wishbone_bd_ram_mem0_reg[139][7]/P0001  , \wishbone_bd_ram_mem0_reg[13][0]/P0001  , \wishbone_bd_ram_mem0_reg[13][1]/P0001  , \wishbone_bd_ram_mem0_reg[13][2]/P0001  , \wishbone_bd_ram_mem0_reg[13][3]/P0001  , \wishbone_bd_ram_mem0_reg[13][4]/P0001  , \wishbone_bd_ram_mem0_reg[13][5]/P0001  , \wishbone_bd_ram_mem0_reg[13][6]/P0001  , \wishbone_bd_ram_mem0_reg[13][7]/P0001  , \wishbone_bd_ram_mem0_reg[140][0]/P0001  , \wishbone_bd_ram_mem0_reg[140][1]/P0001  , \wishbone_bd_ram_mem0_reg[140][2]/P0001  , \wishbone_bd_ram_mem0_reg[140][3]/P0001  , \wishbone_bd_ram_mem0_reg[140][4]/P0001  , \wishbone_bd_ram_mem0_reg[140][5]/P0001  , \wishbone_bd_ram_mem0_reg[140][6]/P0001  , \wishbone_bd_ram_mem0_reg[140][7]/P0001  , \wishbone_bd_ram_mem0_reg[141][0]/P0001  , \wishbone_bd_ram_mem0_reg[141][1]/P0001  , \wishbone_bd_ram_mem0_reg[141][2]/P0001  , \wishbone_bd_ram_mem0_reg[141][3]/P0001  , \wishbone_bd_ram_mem0_reg[141][4]/P0001  , \wishbone_bd_ram_mem0_reg[141][5]/P0001  , \wishbone_bd_ram_mem0_reg[141][6]/P0001  , \wishbone_bd_ram_mem0_reg[141][7]/P0001  , \wishbone_bd_ram_mem0_reg[142][0]/P0001  , \wishbone_bd_ram_mem0_reg[142][1]/P0001  , \wishbone_bd_ram_mem0_reg[142][2]/P0001  , \wishbone_bd_ram_mem0_reg[142][3]/P0001  , \wishbone_bd_ram_mem0_reg[142][4]/P0001  , \wishbone_bd_ram_mem0_reg[142][5]/P0001  , \wishbone_bd_ram_mem0_reg[142][6]/P0001  , \wishbone_bd_ram_mem0_reg[142][7]/P0001  , \wishbone_bd_ram_mem0_reg[143][0]/P0001  , \wishbone_bd_ram_mem0_reg[143][1]/P0001  , \wishbone_bd_ram_mem0_reg[143][2]/P0001  , \wishbone_bd_ram_mem0_reg[143][3]/P0001  , \wishbone_bd_ram_mem0_reg[143][4]/P0001  , \wishbone_bd_ram_mem0_reg[143][5]/P0001  , \wishbone_bd_ram_mem0_reg[143][6]/P0001  , \wishbone_bd_ram_mem0_reg[143][7]/P0001  , \wishbone_bd_ram_mem0_reg[144][0]/P0001  , \wishbone_bd_ram_mem0_reg[144][1]/P0001  , \wishbone_bd_ram_mem0_reg[144][2]/P0001  , \wishbone_bd_ram_mem0_reg[144][3]/P0001  , \wishbone_bd_ram_mem0_reg[144][4]/P0001  , \wishbone_bd_ram_mem0_reg[144][5]/P0001  , \wishbone_bd_ram_mem0_reg[144][6]/P0001  , \wishbone_bd_ram_mem0_reg[144][7]/P0001  , \wishbone_bd_ram_mem0_reg[145][0]/P0001  , \wishbone_bd_ram_mem0_reg[145][1]/P0001  , \wishbone_bd_ram_mem0_reg[145][2]/P0001  , \wishbone_bd_ram_mem0_reg[145][3]/P0001  , \wishbone_bd_ram_mem0_reg[145][4]/P0001  , \wishbone_bd_ram_mem0_reg[145][5]/P0001  , \wishbone_bd_ram_mem0_reg[145][6]/P0001  , \wishbone_bd_ram_mem0_reg[145][7]/P0001  , \wishbone_bd_ram_mem0_reg[146][0]/P0001  , \wishbone_bd_ram_mem0_reg[146][1]/P0001  , \wishbone_bd_ram_mem0_reg[146][2]/P0001  , \wishbone_bd_ram_mem0_reg[146][3]/P0001  , \wishbone_bd_ram_mem0_reg[146][4]/P0001  , \wishbone_bd_ram_mem0_reg[146][5]/P0001  , \wishbone_bd_ram_mem0_reg[146][6]/P0001  , \wishbone_bd_ram_mem0_reg[146][7]/P0001  , \wishbone_bd_ram_mem0_reg[147][0]/P0001  , \wishbone_bd_ram_mem0_reg[147][1]/P0001  , \wishbone_bd_ram_mem0_reg[147][2]/P0001  , \wishbone_bd_ram_mem0_reg[147][3]/P0001  , \wishbone_bd_ram_mem0_reg[147][4]/P0001  , \wishbone_bd_ram_mem0_reg[147][5]/P0001  , \wishbone_bd_ram_mem0_reg[147][6]/P0001  , \wishbone_bd_ram_mem0_reg[147][7]/P0001  , \wishbone_bd_ram_mem0_reg[148][0]/P0001  , \wishbone_bd_ram_mem0_reg[148][1]/P0001  , \wishbone_bd_ram_mem0_reg[148][2]/P0001  , \wishbone_bd_ram_mem0_reg[148][3]/P0001  , \wishbone_bd_ram_mem0_reg[148][4]/P0001  , \wishbone_bd_ram_mem0_reg[148][5]/P0001  , \wishbone_bd_ram_mem0_reg[148][6]/P0001  , \wishbone_bd_ram_mem0_reg[148][7]/P0001  , \wishbone_bd_ram_mem0_reg[149][0]/P0001  , \wishbone_bd_ram_mem0_reg[149][1]/P0001  , \wishbone_bd_ram_mem0_reg[149][2]/P0001  , \wishbone_bd_ram_mem0_reg[149][3]/P0001  , \wishbone_bd_ram_mem0_reg[149][4]/P0001  , \wishbone_bd_ram_mem0_reg[149][5]/P0001  , \wishbone_bd_ram_mem0_reg[149][6]/P0001  , \wishbone_bd_ram_mem0_reg[149][7]/P0001  , \wishbone_bd_ram_mem0_reg[14][0]/P0001  , \wishbone_bd_ram_mem0_reg[14][1]/P0001  , \wishbone_bd_ram_mem0_reg[14][2]/P0001  , \wishbone_bd_ram_mem0_reg[14][3]/P0001  , \wishbone_bd_ram_mem0_reg[14][4]/P0001  , \wishbone_bd_ram_mem0_reg[14][5]/P0001  , \wishbone_bd_ram_mem0_reg[14][6]/P0001  , \wishbone_bd_ram_mem0_reg[14][7]/P0001  , \wishbone_bd_ram_mem0_reg[150][0]/P0001  , \wishbone_bd_ram_mem0_reg[150][1]/P0001  , \wishbone_bd_ram_mem0_reg[150][2]/P0001  , \wishbone_bd_ram_mem0_reg[150][3]/P0001  , \wishbone_bd_ram_mem0_reg[150][4]/P0001  , \wishbone_bd_ram_mem0_reg[150][5]/P0001  , \wishbone_bd_ram_mem0_reg[150][6]/P0001  , \wishbone_bd_ram_mem0_reg[150][7]/P0001  , \wishbone_bd_ram_mem0_reg[151][0]/P0001  , \wishbone_bd_ram_mem0_reg[151][1]/P0001  , \wishbone_bd_ram_mem0_reg[151][2]/P0001  , \wishbone_bd_ram_mem0_reg[151][3]/P0001  , \wishbone_bd_ram_mem0_reg[151][4]/P0001  , \wishbone_bd_ram_mem0_reg[151][5]/P0001  , \wishbone_bd_ram_mem0_reg[151][6]/P0001  , \wishbone_bd_ram_mem0_reg[151][7]/P0001  , \wishbone_bd_ram_mem0_reg[152][0]/P0001  , \wishbone_bd_ram_mem0_reg[152][1]/P0001  , \wishbone_bd_ram_mem0_reg[152][2]/P0001  , \wishbone_bd_ram_mem0_reg[152][3]/P0001  , \wishbone_bd_ram_mem0_reg[152][4]/P0001  , \wishbone_bd_ram_mem0_reg[152][5]/P0001  , \wishbone_bd_ram_mem0_reg[152][6]/P0001  , \wishbone_bd_ram_mem0_reg[152][7]/P0001  , \wishbone_bd_ram_mem0_reg[153][0]/P0001  , \wishbone_bd_ram_mem0_reg[153][1]/P0001  , \wishbone_bd_ram_mem0_reg[153][2]/P0001  , \wishbone_bd_ram_mem0_reg[153][3]/P0001  , \wishbone_bd_ram_mem0_reg[153][4]/P0001  , \wishbone_bd_ram_mem0_reg[153][5]/P0001  , \wishbone_bd_ram_mem0_reg[153][6]/P0001  , \wishbone_bd_ram_mem0_reg[153][7]/P0001  , \wishbone_bd_ram_mem0_reg[154][0]/P0001  , \wishbone_bd_ram_mem0_reg[154][1]/P0001  , \wishbone_bd_ram_mem0_reg[154][2]/P0001  , \wishbone_bd_ram_mem0_reg[154][3]/P0001  , \wishbone_bd_ram_mem0_reg[154][4]/P0001  , \wishbone_bd_ram_mem0_reg[154][5]/P0001  , \wishbone_bd_ram_mem0_reg[154][6]/P0001  , \wishbone_bd_ram_mem0_reg[154][7]/P0001  , \wishbone_bd_ram_mem0_reg[155][0]/P0001  , \wishbone_bd_ram_mem0_reg[155][1]/P0001  , \wishbone_bd_ram_mem0_reg[155][2]/P0001  , \wishbone_bd_ram_mem0_reg[155][3]/P0001  , \wishbone_bd_ram_mem0_reg[155][4]/P0001  , \wishbone_bd_ram_mem0_reg[155][5]/P0001  , \wishbone_bd_ram_mem0_reg[155][6]/P0001  , \wishbone_bd_ram_mem0_reg[155][7]/P0001  , \wishbone_bd_ram_mem0_reg[156][0]/P0001  , \wishbone_bd_ram_mem0_reg[156][1]/P0001  , \wishbone_bd_ram_mem0_reg[156][2]/P0001  , \wishbone_bd_ram_mem0_reg[156][3]/P0001  , \wishbone_bd_ram_mem0_reg[156][4]/P0001  , \wishbone_bd_ram_mem0_reg[156][5]/P0001  , \wishbone_bd_ram_mem0_reg[156][6]/P0001  , \wishbone_bd_ram_mem0_reg[156][7]/P0001  , \wishbone_bd_ram_mem0_reg[157][0]/P0001  , \wishbone_bd_ram_mem0_reg[157][1]/P0001  , \wishbone_bd_ram_mem0_reg[157][2]/P0001  , \wishbone_bd_ram_mem0_reg[157][3]/P0001  , \wishbone_bd_ram_mem0_reg[157][4]/P0001  , \wishbone_bd_ram_mem0_reg[157][5]/P0001  , \wishbone_bd_ram_mem0_reg[157][6]/P0001  , \wishbone_bd_ram_mem0_reg[157][7]/P0001  , \wishbone_bd_ram_mem0_reg[158][0]/P0001  , \wishbone_bd_ram_mem0_reg[158][1]/P0001  , \wishbone_bd_ram_mem0_reg[158][2]/P0001  , \wishbone_bd_ram_mem0_reg[158][3]/P0001  , \wishbone_bd_ram_mem0_reg[158][4]/P0001  , \wishbone_bd_ram_mem0_reg[158][5]/P0001  , \wishbone_bd_ram_mem0_reg[158][6]/P0001  , \wishbone_bd_ram_mem0_reg[158][7]/P0001  , \wishbone_bd_ram_mem0_reg[159][0]/P0001  , \wishbone_bd_ram_mem0_reg[159][1]/P0001  , \wishbone_bd_ram_mem0_reg[159][2]/P0001  , \wishbone_bd_ram_mem0_reg[159][3]/P0001  , \wishbone_bd_ram_mem0_reg[159][4]/P0001  , \wishbone_bd_ram_mem0_reg[159][5]/P0001  , \wishbone_bd_ram_mem0_reg[159][6]/P0001  , \wishbone_bd_ram_mem0_reg[159][7]/P0001  , \wishbone_bd_ram_mem0_reg[15][0]/P0001  , \wishbone_bd_ram_mem0_reg[15][1]/P0001  , \wishbone_bd_ram_mem0_reg[15][2]/P0001  , \wishbone_bd_ram_mem0_reg[15][3]/P0001  , \wishbone_bd_ram_mem0_reg[15][4]/P0001  , \wishbone_bd_ram_mem0_reg[15][5]/P0001  , \wishbone_bd_ram_mem0_reg[15][6]/P0001  , \wishbone_bd_ram_mem0_reg[15][7]/P0001  , \wishbone_bd_ram_mem0_reg[160][0]/P0001  , \wishbone_bd_ram_mem0_reg[160][1]/P0001  , \wishbone_bd_ram_mem0_reg[160][2]/P0001  , \wishbone_bd_ram_mem0_reg[160][3]/P0001  , \wishbone_bd_ram_mem0_reg[160][4]/P0001  , \wishbone_bd_ram_mem0_reg[160][5]/P0001  , \wishbone_bd_ram_mem0_reg[160][6]/P0001  , \wishbone_bd_ram_mem0_reg[160][7]/P0001  , \wishbone_bd_ram_mem0_reg[161][0]/P0001  , \wishbone_bd_ram_mem0_reg[161][1]/P0001  , \wishbone_bd_ram_mem0_reg[161][2]/P0001  , \wishbone_bd_ram_mem0_reg[161][3]/P0001  , \wishbone_bd_ram_mem0_reg[161][4]/P0001  , \wishbone_bd_ram_mem0_reg[161][5]/P0001  , \wishbone_bd_ram_mem0_reg[161][6]/P0001  , \wishbone_bd_ram_mem0_reg[161][7]/P0001  , \wishbone_bd_ram_mem0_reg[162][0]/P0001  , \wishbone_bd_ram_mem0_reg[162][1]/P0001  , \wishbone_bd_ram_mem0_reg[162][2]/P0001  , \wishbone_bd_ram_mem0_reg[162][3]/P0001  , \wishbone_bd_ram_mem0_reg[162][4]/P0001  , \wishbone_bd_ram_mem0_reg[162][5]/P0001  , \wishbone_bd_ram_mem0_reg[162][6]/P0001  , \wishbone_bd_ram_mem0_reg[162][7]/P0001  , \wishbone_bd_ram_mem0_reg[163][0]/P0001  , \wishbone_bd_ram_mem0_reg[163][1]/P0001  , \wishbone_bd_ram_mem0_reg[163][2]/P0001  , \wishbone_bd_ram_mem0_reg[163][3]/P0001  , \wishbone_bd_ram_mem0_reg[163][4]/P0001  , \wishbone_bd_ram_mem0_reg[163][5]/P0001  , \wishbone_bd_ram_mem0_reg[163][6]/P0001  , \wishbone_bd_ram_mem0_reg[163][7]/P0001  , \wishbone_bd_ram_mem0_reg[164][0]/P0001  , \wishbone_bd_ram_mem0_reg[164][1]/P0001  , \wishbone_bd_ram_mem0_reg[164][2]/P0001  , \wishbone_bd_ram_mem0_reg[164][3]/P0001  , \wishbone_bd_ram_mem0_reg[164][4]/P0001  , \wishbone_bd_ram_mem0_reg[164][5]/P0001  , \wishbone_bd_ram_mem0_reg[164][6]/P0001  , \wishbone_bd_ram_mem0_reg[164][7]/P0001  , \wishbone_bd_ram_mem0_reg[165][0]/P0001  , \wishbone_bd_ram_mem0_reg[165][1]/P0001  , \wishbone_bd_ram_mem0_reg[165][2]/P0001  , \wishbone_bd_ram_mem0_reg[165][3]/P0001  , \wishbone_bd_ram_mem0_reg[165][4]/P0001  , \wishbone_bd_ram_mem0_reg[165][5]/P0001  , \wishbone_bd_ram_mem0_reg[165][6]/P0001  , \wishbone_bd_ram_mem0_reg[165][7]/P0001  , \wishbone_bd_ram_mem0_reg[166][0]/P0001  , \wishbone_bd_ram_mem0_reg[166][1]/P0001  , \wishbone_bd_ram_mem0_reg[166][2]/P0001  , \wishbone_bd_ram_mem0_reg[166][3]/P0001  , \wishbone_bd_ram_mem0_reg[166][4]/P0001  , \wishbone_bd_ram_mem0_reg[166][5]/P0001  , \wishbone_bd_ram_mem0_reg[166][6]/P0001  , \wishbone_bd_ram_mem0_reg[166][7]/P0001  , \wishbone_bd_ram_mem0_reg[167][0]/P0001  , \wishbone_bd_ram_mem0_reg[167][1]/P0001  , \wishbone_bd_ram_mem0_reg[167][2]/P0001  , \wishbone_bd_ram_mem0_reg[167][3]/P0001  , \wishbone_bd_ram_mem0_reg[167][4]/P0001  , \wishbone_bd_ram_mem0_reg[167][5]/P0001  , \wishbone_bd_ram_mem0_reg[167][6]/P0001  , \wishbone_bd_ram_mem0_reg[167][7]/P0001  , \wishbone_bd_ram_mem0_reg[168][0]/P0001  , \wishbone_bd_ram_mem0_reg[168][1]/P0001  , \wishbone_bd_ram_mem0_reg[168][2]/P0001  , \wishbone_bd_ram_mem0_reg[168][3]/P0001  , \wishbone_bd_ram_mem0_reg[168][4]/P0001  , \wishbone_bd_ram_mem0_reg[168][5]/P0001  , \wishbone_bd_ram_mem0_reg[168][6]/P0001  , \wishbone_bd_ram_mem0_reg[168][7]/P0001  , \wishbone_bd_ram_mem0_reg[169][0]/P0001  , \wishbone_bd_ram_mem0_reg[169][1]/P0001  , \wishbone_bd_ram_mem0_reg[169][2]/P0001  , \wishbone_bd_ram_mem0_reg[169][3]/P0001  , \wishbone_bd_ram_mem0_reg[169][4]/P0001  , \wishbone_bd_ram_mem0_reg[169][5]/P0001  , \wishbone_bd_ram_mem0_reg[169][6]/P0001  , \wishbone_bd_ram_mem0_reg[169][7]/P0001  , \wishbone_bd_ram_mem0_reg[16][0]/P0001  , \wishbone_bd_ram_mem0_reg[16][1]/P0001  , \wishbone_bd_ram_mem0_reg[16][2]/P0001  , \wishbone_bd_ram_mem0_reg[16][3]/P0001  , \wishbone_bd_ram_mem0_reg[16][4]/P0001  , \wishbone_bd_ram_mem0_reg[16][5]/P0001  , \wishbone_bd_ram_mem0_reg[16][6]/P0001  , \wishbone_bd_ram_mem0_reg[16][7]/P0001  , \wishbone_bd_ram_mem0_reg[170][0]/P0001  , \wishbone_bd_ram_mem0_reg[170][1]/P0001  , \wishbone_bd_ram_mem0_reg[170][2]/P0001  , \wishbone_bd_ram_mem0_reg[170][3]/P0001  , \wishbone_bd_ram_mem0_reg[170][4]/P0001  , \wishbone_bd_ram_mem0_reg[170][5]/P0001  , \wishbone_bd_ram_mem0_reg[170][6]/P0001  , \wishbone_bd_ram_mem0_reg[170][7]/P0001  , \wishbone_bd_ram_mem0_reg[171][0]/P0001  , \wishbone_bd_ram_mem0_reg[171][1]/P0001  , \wishbone_bd_ram_mem0_reg[171][2]/P0001  , \wishbone_bd_ram_mem0_reg[171][3]/P0001  , \wishbone_bd_ram_mem0_reg[171][4]/P0001  , \wishbone_bd_ram_mem0_reg[171][5]/P0001  , \wishbone_bd_ram_mem0_reg[171][6]/P0001  , \wishbone_bd_ram_mem0_reg[171][7]/P0001  , \wishbone_bd_ram_mem0_reg[172][0]/P0001  , \wishbone_bd_ram_mem0_reg[172][1]/P0001  , \wishbone_bd_ram_mem0_reg[172][2]/P0001  , \wishbone_bd_ram_mem0_reg[172][3]/P0001  , \wishbone_bd_ram_mem0_reg[172][4]/P0001  , \wishbone_bd_ram_mem0_reg[172][5]/P0001  , \wishbone_bd_ram_mem0_reg[172][6]/P0001  , \wishbone_bd_ram_mem0_reg[172][7]/P0001  , \wishbone_bd_ram_mem0_reg[173][0]/P0001  , \wishbone_bd_ram_mem0_reg[173][1]/P0001  , \wishbone_bd_ram_mem0_reg[173][2]/P0001  , \wishbone_bd_ram_mem0_reg[173][3]/P0001  , \wishbone_bd_ram_mem0_reg[173][4]/P0001  , \wishbone_bd_ram_mem0_reg[173][5]/P0001  , \wishbone_bd_ram_mem0_reg[173][6]/P0001  , \wishbone_bd_ram_mem0_reg[173][7]/P0001  , \wishbone_bd_ram_mem0_reg[174][0]/P0001  , \wishbone_bd_ram_mem0_reg[174][1]/P0001  , \wishbone_bd_ram_mem0_reg[174][2]/P0001  , \wishbone_bd_ram_mem0_reg[174][3]/P0001  , \wishbone_bd_ram_mem0_reg[174][4]/P0001  , \wishbone_bd_ram_mem0_reg[174][5]/P0001  , \wishbone_bd_ram_mem0_reg[174][6]/P0001  , \wishbone_bd_ram_mem0_reg[174][7]/P0001  , \wishbone_bd_ram_mem0_reg[175][0]/P0001  , \wishbone_bd_ram_mem0_reg[175][1]/P0001  , \wishbone_bd_ram_mem0_reg[175][2]/P0001  , \wishbone_bd_ram_mem0_reg[175][3]/P0001  , \wishbone_bd_ram_mem0_reg[175][4]/P0001  , \wishbone_bd_ram_mem0_reg[175][5]/P0001  , \wishbone_bd_ram_mem0_reg[175][6]/P0001  , \wishbone_bd_ram_mem0_reg[175][7]/P0001  , \wishbone_bd_ram_mem0_reg[176][0]/P0001  , \wishbone_bd_ram_mem0_reg[176][1]/P0001  , \wishbone_bd_ram_mem0_reg[176][2]/P0001  , \wishbone_bd_ram_mem0_reg[176][3]/P0001  , \wishbone_bd_ram_mem0_reg[176][4]/P0001  , \wishbone_bd_ram_mem0_reg[176][5]/P0001  , \wishbone_bd_ram_mem0_reg[176][6]/P0001  , \wishbone_bd_ram_mem0_reg[176][7]/P0001  , \wishbone_bd_ram_mem0_reg[177][0]/P0001  , \wishbone_bd_ram_mem0_reg[177][1]/P0001  , \wishbone_bd_ram_mem0_reg[177][2]/P0001  , \wishbone_bd_ram_mem0_reg[177][3]/P0001  , \wishbone_bd_ram_mem0_reg[177][4]/P0001  , \wishbone_bd_ram_mem0_reg[177][5]/P0001  , \wishbone_bd_ram_mem0_reg[177][6]/P0001  , \wishbone_bd_ram_mem0_reg[177][7]/P0001  , \wishbone_bd_ram_mem0_reg[178][0]/P0001  , \wishbone_bd_ram_mem0_reg[178][1]/P0001  , \wishbone_bd_ram_mem0_reg[178][2]/P0001  , \wishbone_bd_ram_mem0_reg[178][3]/P0001  , \wishbone_bd_ram_mem0_reg[178][4]/P0001  , \wishbone_bd_ram_mem0_reg[178][5]/P0001  , \wishbone_bd_ram_mem0_reg[178][6]/P0001  , \wishbone_bd_ram_mem0_reg[178][7]/P0001  , \wishbone_bd_ram_mem0_reg[179][0]/P0001  , \wishbone_bd_ram_mem0_reg[179][1]/P0001  , \wishbone_bd_ram_mem0_reg[179][2]/P0001  , \wishbone_bd_ram_mem0_reg[179][3]/P0001  , \wishbone_bd_ram_mem0_reg[179][4]/P0001  , \wishbone_bd_ram_mem0_reg[179][5]/P0001  , \wishbone_bd_ram_mem0_reg[179][6]/P0001  , \wishbone_bd_ram_mem0_reg[179][7]/P0001  , \wishbone_bd_ram_mem0_reg[17][0]/P0001  , \wishbone_bd_ram_mem0_reg[17][1]/P0001  , \wishbone_bd_ram_mem0_reg[17][2]/P0001  , \wishbone_bd_ram_mem0_reg[17][3]/P0001  , \wishbone_bd_ram_mem0_reg[17][4]/P0001  , \wishbone_bd_ram_mem0_reg[17][5]/P0001  , \wishbone_bd_ram_mem0_reg[17][6]/P0001  , \wishbone_bd_ram_mem0_reg[17][7]/P0001  , \wishbone_bd_ram_mem0_reg[180][0]/P0001  , \wishbone_bd_ram_mem0_reg[180][1]/P0001  , \wishbone_bd_ram_mem0_reg[180][2]/P0001  , \wishbone_bd_ram_mem0_reg[180][3]/P0001  , \wishbone_bd_ram_mem0_reg[180][4]/P0001  , \wishbone_bd_ram_mem0_reg[180][5]/P0001  , \wishbone_bd_ram_mem0_reg[180][6]/P0001  , \wishbone_bd_ram_mem0_reg[180][7]/P0001  , \wishbone_bd_ram_mem0_reg[181][0]/P0001  , \wishbone_bd_ram_mem0_reg[181][1]/P0001  , \wishbone_bd_ram_mem0_reg[181][2]/P0001  , \wishbone_bd_ram_mem0_reg[181][3]/P0001  , \wishbone_bd_ram_mem0_reg[181][4]/P0001  , \wishbone_bd_ram_mem0_reg[181][5]/P0001  , \wishbone_bd_ram_mem0_reg[181][6]/P0001  , \wishbone_bd_ram_mem0_reg[181][7]/P0001  , \wishbone_bd_ram_mem0_reg[182][0]/P0001  , \wishbone_bd_ram_mem0_reg[182][1]/P0001  , \wishbone_bd_ram_mem0_reg[182][2]/P0001  , \wishbone_bd_ram_mem0_reg[182][3]/P0001  , \wishbone_bd_ram_mem0_reg[182][4]/P0001  , \wishbone_bd_ram_mem0_reg[182][5]/P0001  , \wishbone_bd_ram_mem0_reg[182][6]/P0001  , \wishbone_bd_ram_mem0_reg[182][7]/P0001  , \wishbone_bd_ram_mem0_reg[183][0]/P0001  , \wishbone_bd_ram_mem0_reg[183][1]/P0001  , \wishbone_bd_ram_mem0_reg[183][2]/P0001  , \wishbone_bd_ram_mem0_reg[183][3]/P0001  , \wishbone_bd_ram_mem0_reg[183][4]/P0001  , \wishbone_bd_ram_mem0_reg[183][5]/P0001  , \wishbone_bd_ram_mem0_reg[183][6]/P0001  , \wishbone_bd_ram_mem0_reg[183][7]/P0001  , \wishbone_bd_ram_mem0_reg[184][0]/P0001  , \wishbone_bd_ram_mem0_reg[184][1]/P0001  , \wishbone_bd_ram_mem0_reg[184][2]/P0001  , \wishbone_bd_ram_mem0_reg[184][3]/P0001  , \wishbone_bd_ram_mem0_reg[184][4]/P0001  , \wishbone_bd_ram_mem0_reg[184][5]/P0001  , \wishbone_bd_ram_mem0_reg[184][6]/P0001  , \wishbone_bd_ram_mem0_reg[184][7]/P0001  , \wishbone_bd_ram_mem0_reg[185][0]/P0001  , \wishbone_bd_ram_mem0_reg[185][1]/P0001  , \wishbone_bd_ram_mem0_reg[185][2]/P0001  , \wishbone_bd_ram_mem0_reg[185][3]/P0001  , \wishbone_bd_ram_mem0_reg[185][4]/P0001  , \wishbone_bd_ram_mem0_reg[185][5]/P0001  , \wishbone_bd_ram_mem0_reg[185][6]/P0001  , \wishbone_bd_ram_mem0_reg[185][7]/P0001  , \wishbone_bd_ram_mem0_reg[186][0]/P0001  , \wishbone_bd_ram_mem0_reg[186][1]/P0001  , \wishbone_bd_ram_mem0_reg[186][2]/P0001  , \wishbone_bd_ram_mem0_reg[186][3]/P0001  , \wishbone_bd_ram_mem0_reg[186][4]/P0001  , \wishbone_bd_ram_mem0_reg[186][5]/P0001  , \wishbone_bd_ram_mem0_reg[186][6]/P0001  , \wishbone_bd_ram_mem0_reg[186][7]/P0001  , \wishbone_bd_ram_mem0_reg[187][0]/P0001  , \wishbone_bd_ram_mem0_reg[187][1]/P0001  , \wishbone_bd_ram_mem0_reg[187][2]/P0001  , \wishbone_bd_ram_mem0_reg[187][3]/P0001  , \wishbone_bd_ram_mem0_reg[187][4]/P0001  , \wishbone_bd_ram_mem0_reg[187][5]/P0001  , \wishbone_bd_ram_mem0_reg[187][6]/P0001  , \wishbone_bd_ram_mem0_reg[187][7]/P0001  , \wishbone_bd_ram_mem0_reg[188][0]/P0001  , \wishbone_bd_ram_mem0_reg[188][1]/P0001  , \wishbone_bd_ram_mem0_reg[188][2]/P0001  , \wishbone_bd_ram_mem0_reg[188][3]/P0001  , \wishbone_bd_ram_mem0_reg[188][4]/P0001  , \wishbone_bd_ram_mem0_reg[188][5]/P0001  , \wishbone_bd_ram_mem0_reg[188][6]/P0001  , \wishbone_bd_ram_mem0_reg[188][7]/P0001  , \wishbone_bd_ram_mem0_reg[189][0]/P0001  , \wishbone_bd_ram_mem0_reg[189][1]/P0001  , \wishbone_bd_ram_mem0_reg[189][2]/P0001  , \wishbone_bd_ram_mem0_reg[189][3]/P0001  , \wishbone_bd_ram_mem0_reg[189][4]/P0001  , \wishbone_bd_ram_mem0_reg[189][5]/P0001  , \wishbone_bd_ram_mem0_reg[189][6]/P0001  , \wishbone_bd_ram_mem0_reg[189][7]/P0001  , \wishbone_bd_ram_mem0_reg[18][0]/P0001  , \wishbone_bd_ram_mem0_reg[18][1]/P0001  , \wishbone_bd_ram_mem0_reg[18][2]/P0001  , \wishbone_bd_ram_mem0_reg[18][3]/P0001  , \wishbone_bd_ram_mem0_reg[18][4]/P0001  , \wishbone_bd_ram_mem0_reg[18][5]/P0001  , \wishbone_bd_ram_mem0_reg[18][6]/P0001  , \wishbone_bd_ram_mem0_reg[18][7]/P0001  , \wishbone_bd_ram_mem0_reg[190][0]/P0001  , \wishbone_bd_ram_mem0_reg[190][1]/P0001  , \wishbone_bd_ram_mem0_reg[190][2]/P0001  , \wishbone_bd_ram_mem0_reg[190][3]/P0001  , \wishbone_bd_ram_mem0_reg[190][4]/P0001  , \wishbone_bd_ram_mem0_reg[190][5]/P0001  , \wishbone_bd_ram_mem0_reg[190][6]/P0001  , \wishbone_bd_ram_mem0_reg[190][7]/P0001  , \wishbone_bd_ram_mem0_reg[191][0]/P0001  , \wishbone_bd_ram_mem0_reg[191][1]/P0001  , \wishbone_bd_ram_mem0_reg[191][2]/P0001  , \wishbone_bd_ram_mem0_reg[191][3]/P0001  , \wishbone_bd_ram_mem0_reg[191][4]/P0001  , \wishbone_bd_ram_mem0_reg[191][5]/P0001  , \wishbone_bd_ram_mem0_reg[191][6]/P0001  , \wishbone_bd_ram_mem0_reg[191][7]/P0001  , \wishbone_bd_ram_mem0_reg[192][0]/P0001  , \wishbone_bd_ram_mem0_reg[192][1]/P0001  , \wishbone_bd_ram_mem0_reg[192][2]/P0001  , \wishbone_bd_ram_mem0_reg[192][3]/P0001  , \wishbone_bd_ram_mem0_reg[192][4]/P0001  , \wishbone_bd_ram_mem0_reg[192][5]/P0001  , \wishbone_bd_ram_mem0_reg[192][6]/P0001  , \wishbone_bd_ram_mem0_reg[192][7]/P0001  , \wishbone_bd_ram_mem0_reg[193][0]/P0001  , \wishbone_bd_ram_mem0_reg[193][1]/P0001  , \wishbone_bd_ram_mem0_reg[193][2]/P0001  , \wishbone_bd_ram_mem0_reg[193][3]/P0001  , \wishbone_bd_ram_mem0_reg[193][4]/P0001  , \wishbone_bd_ram_mem0_reg[193][5]/P0001  , \wishbone_bd_ram_mem0_reg[193][6]/P0001  , \wishbone_bd_ram_mem0_reg[193][7]/P0001  , \wishbone_bd_ram_mem0_reg[194][0]/P0001  , \wishbone_bd_ram_mem0_reg[194][1]/P0001  , \wishbone_bd_ram_mem0_reg[194][2]/P0001  , \wishbone_bd_ram_mem0_reg[194][3]/P0001  , \wishbone_bd_ram_mem0_reg[194][4]/P0001  , \wishbone_bd_ram_mem0_reg[194][5]/P0001  , \wishbone_bd_ram_mem0_reg[194][6]/P0001  , \wishbone_bd_ram_mem0_reg[194][7]/P0001  , \wishbone_bd_ram_mem0_reg[195][0]/P0001  , \wishbone_bd_ram_mem0_reg[195][1]/P0001  , \wishbone_bd_ram_mem0_reg[195][2]/P0001  , \wishbone_bd_ram_mem0_reg[195][3]/P0001  , \wishbone_bd_ram_mem0_reg[195][4]/P0001  , \wishbone_bd_ram_mem0_reg[195][5]/P0001  , \wishbone_bd_ram_mem0_reg[195][6]/P0001  , \wishbone_bd_ram_mem0_reg[195][7]/P0001  , \wishbone_bd_ram_mem0_reg[196][0]/P0001  , \wishbone_bd_ram_mem0_reg[196][1]/P0001  , \wishbone_bd_ram_mem0_reg[196][2]/P0001  , \wishbone_bd_ram_mem0_reg[196][3]/P0001  , \wishbone_bd_ram_mem0_reg[196][4]/P0001  , \wishbone_bd_ram_mem0_reg[196][5]/P0001  , \wishbone_bd_ram_mem0_reg[196][6]/P0001  , \wishbone_bd_ram_mem0_reg[196][7]/P0001  , \wishbone_bd_ram_mem0_reg[197][0]/P0001  , \wishbone_bd_ram_mem0_reg[197][1]/P0001  , \wishbone_bd_ram_mem0_reg[197][2]/P0001  , \wishbone_bd_ram_mem0_reg[197][3]/P0001  , \wishbone_bd_ram_mem0_reg[197][4]/P0001  , \wishbone_bd_ram_mem0_reg[197][5]/P0001  , \wishbone_bd_ram_mem0_reg[197][6]/P0001  , \wishbone_bd_ram_mem0_reg[197][7]/P0001  , \wishbone_bd_ram_mem0_reg[198][0]/P0001  , \wishbone_bd_ram_mem0_reg[198][1]/P0001  , \wishbone_bd_ram_mem0_reg[198][2]/P0001  , \wishbone_bd_ram_mem0_reg[198][3]/P0001  , \wishbone_bd_ram_mem0_reg[198][4]/P0001  , \wishbone_bd_ram_mem0_reg[198][5]/P0001  , \wishbone_bd_ram_mem0_reg[198][6]/P0001  , \wishbone_bd_ram_mem0_reg[198][7]/P0001  , \wishbone_bd_ram_mem0_reg[199][0]/P0001  , \wishbone_bd_ram_mem0_reg[199][1]/P0001  , \wishbone_bd_ram_mem0_reg[199][2]/P0001  , \wishbone_bd_ram_mem0_reg[199][3]/P0001  , \wishbone_bd_ram_mem0_reg[199][4]/P0001  , \wishbone_bd_ram_mem0_reg[199][5]/P0001  , \wishbone_bd_ram_mem0_reg[199][6]/P0001  , \wishbone_bd_ram_mem0_reg[199][7]/P0001  , \wishbone_bd_ram_mem0_reg[19][0]/P0001  , \wishbone_bd_ram_mem0_reg[19][1]/P0001  , \wishbone_bd_ram_mem0_reg[19][2]/P0001  , \wishbone_bd_ram_mem0_reg[19][3]/P0001  , \wishbone_bd_ram_mem0_reg[19][4]/P0001  , \wishbone_bd_ram_mem0_reg[19][5]/P0001  , \wishbone_bd_ram_mem0_reg[19][6]/P0001  , \wishbone_bd_ram_mem0_reg[19][7]/P0001  , \wishbone_bd_ram_mem0_reg[1][0]/P0001  , \wishbone_bd_ram_mem0_reg[1][1]/P0001  , \wishbone_bd_ram_mem0_reg[1][2]/P0001  , \wishbone_bd_ram_mem0_reg[1][3]/P0001  , \wishbone_bd_ram_mem0_reg[1][4]/P0001  , \wishbone_bd_ram_mem0_reg[1][5]/P0001  , \wishbone_bd_ram_mem0_reg[1][6]/P0001  , \wishbone_bd_ram_mem0_reg[1][7]/P0001  , \wishbone_bd_ram_mem0_reg[200][0]/P0001  , \wishbone_bd_ram_mem0_reg[200][1]/P0001  , \wishbone_bd_ram_mem0_reg[200][2]/P0001  , \wishbone_bd_ram_mem0_reg[200][3]/P0001  , \wishbone_bd_ram_mem0_reg[200][4]/P0001  , \wishbone_bd_ram_mem0_reg[200][5]/P0001  , \wishbone_bd_ram_mem0_reg[200][6]/P0001  , \wishbone_bd_ram_mem0_reg[200][7]/P0001  , \wishbone_bd_ram_mem0_reg[201][0]/P0001  , \wishbone_bd_ram_mem0_reg[201][1]/P0001  , \wishbone_bd_ram_mem0_reg[201][2]/P0001  , \wishbone_bd_ram_mem0_reg[201][3]/P0001  , \wishbone_bd_ram_mem0_reg[201][4]/P0001  , \wishbone_bd_ram_mem0_reg[201][5]/P0001  , \wishbone_bd_ram_mem0_reg[201][6]/P0001  , \wishbone_bd_ram_mem0_reg[201][7]/P0001  , \wishbone_bd_ram_mem0_reg[202][0]/P0001  , \wishbone_bd_ram_mem0_reg[202][1]/P0001  , \wishbone_bd_ram_mem0_reg[202][2]/P0001  , \wishbone_bd_ram_mem0_reg[202][3]/P0001  , \wishbone_bd_ram_mem0_reg[202][4]/P0001  , \wishbone_bd_ram_mem0_reg[202][5]/P0001  , \wishbone_bd_ram_mem0_reg[202][6]/P0001  , \wishbone_bd_ram_mem0_reg[202][7]/P0001  , \wishbone_bd_ram_mem0_reg[203][0]/P0001  , \wishbone_bd_ram_mem0_reg[203][1]/P0001  , \wishbone_bd_ram_mem0_reg[203][2]/P0001  , \wishbone_bd_ram_mem0_reg[203][3]/P0001  , \wishbone_bd_ram_mem0_reg[203][4]/P0001  , \wishbone_bd_ram_mem0_reg[203][5]/P0001  , \wishbone_bd_ram_mem0_reg[203][6]/P0001  , \wishbone_bd_ram_mem0_reg[203][7]/P0001  , \wishbone_bd_ram_mem0_reg[204][0]/P0001  , \wishbone_bd_ram_mem0_reg[204][1]/P0001  , \wishbone_bd_ram_mem0_reg[204][2]/P0001  , \wishbone_bd_ram_mem0_reg[204][3]/P0001  , \wishbone_bd_ram_mem0_reg[204][4]/P0001  , \wishbone_bd_ram_mem0_reg[204][5]/P0001  , \wishbone_bd_ram_mem0_reg[204][6]/P0001  , \wishbone_bd_ram_mem0_reg[204][7]/P0001  , \wishbone_bd_ram_mem0_reg[205][0]/P0001  , \wishbone_bd_ram_mem0_reg[205][1]/P0001  , \wishbone_bd_ram_mem0_reg[205][2]/P0001  , \wishbone_bd_ram_mem0_reg[205][3]/P0001  , \wishbone_bd_ram_mem0_reg[205][4]/P0001  , \wishbone_bd_ram_mem0_reg[205][5]/P0001  , \wishbone_bd_ram_mem0_reg[205][6]/P0001  , \wishbone_bd_ram_mem0_reg[205][7]/P0001  , \wishbone_bd_ram_mem0_reg[206][0]/P0001  , \wishbone_bd_ram_mem0_reg[206][1]/P0001  , \wishbone_bd_ram_mem0_reg[206][2]/P0001  , \wishbone_bd_ram_mem0_reg[206][3]/P0001  , \wishbone_bd_ram_mem0_reg[206][4]/P0001  , \wishbone_bd_ram_mem0_reg[206][5]/P0001  , \wishbone_bd_ram_mem0_reg[206][6]/P0001  , \wishbone_bd_ram_mem0_reg[206][7]/P0001  , \wishbone_bd_ram_mem0_reg[207][0]/P0001  , \wishbone_bd_ram_mem0_reg[207][1]/P0001  , \wishbone_bd_ram_mem0_reg[207][2]/P0001  , \wishbone_bd_ram_mem0_reg[207][3]/P0001  , \wishbone_bd_ram_mem0_reg[207][4]/P0001  , \wishbone_bd_ram_mem0_reg[207][5]/P0001  , \wishbone_bd_ram_mem0_reg[207][6]/P0001  , \wishbone_bd_ram_mem0_reg[207][7]/P0001  , \wishbone_bd_ram_mem0_reg[208][0]/P0001  , \wishbone_bd_ram_mem0_reg[208][1]/P0001  , \wishbone_bd_ram_mem0_reg[208][2]/P0001  , \wishbone_bd_ram_mem0_reg[208][3]/P0001  , \wishbone_bd_ram_mem0_reg[208][4]/P0001  , \wishbone_bd_ram_mem0_reg[208][5]/P0001  , \wishbone_bd_ram_mem0_reg[208][6]/P0001  , \wishbone_bd_ram_mem0_reg[208][7]/P0001  , \wishbone_bd_ram_mem0_reg[209][0]/P0001  , \wishbone_bd_ram_mem0_reg[209][1]/P0001  , \wishbone_bd_ram_mem0_reg[209][2]/P0001  , \wishbone_bd_ram_mem0_reg[209][3]/P0001  , \wishbone_bd_ram_mem0_reg[209][4]/P0001  , \wishbone_bd_ram_mem0_reg[209][5]/P0001  , \wishbone_bd_ram_mem0_reg[209][6]/P0001  , \wishbone_bd_ram_mem0_reg[209][7]/P0001  , \wishbone_bd_ram_mem0_reg[20][0]/P0001  , \wishbone_bd_ram_mem0_reg[20][1]/P0001  , \wishbone_bd_ram_mem0_reg[20][2]/P0001  , \wishbone_bd_ram_mem0_reg[20][3]/P0001  , \wishbone_bd_ram_mem0_reg[20][4]/P0001  , \wishbone_bd_ram_mem0_reg[20][5]/P0001  , \wishbone_bd_ram_mem0_reg[20][6]/P0001  , \wishbone_bd_ram_mem0_reg[20][7]/P0001  , \wishbone_bd_ram_mem0_reg[210][0]/P0001  , \wishbone_bd_ram_mem0_reg[210][1]/P0001  , \wishbone_bd_ram_mem0_reg[210][2]/P0001  , \wishbone_bd_ram_mem0_reg[210][3]/P0001  , \wishbone_bd_ram_mem0_reg[210][4]/P0001  , \wishbone_bd_ram_mem0_reg[210][5]/P0001  , \wishbone_bd_ram_mem0_reg[210][6]/P0001  , \wishbone_bd_ram_mem0_reg[210][7]/P0001  , \wishbone_bd_ram_mem0_reg[211][0]/P0001  , \wishbone_bd_ram_mem0_reg[211][1]/P0001  , \wishbone_bd_ram_mem0_reg[211][2]/P0001  , \wishbone_bd_ram_mem0_reg[211][3]/P0001  , \wishbone_bd_ram_mem0_reg[211][4]/P0001  , \wishbone_bd_ram_mem0_reg[211][5]/P0001  , \wishbone_bd_ram_mem0_reg[211][6]/P0001  , \wishbone_bd_ram_mem0_reg[211][7]/P0001  , \wishbone_bd_ram_mem0_reg[212][0]/P0001  , \wishbone_bd_ram_mem0_reg[212][1]/P0001  , \wishbone_bd_ram_mem0_reg[212][2]/P0001  , \wishbone_bd_ram_mem0_reg[212][3]/P0001  , \wishbone_bd_ram_mem0_reg[212][4]/P0001  , \wishbone_bd_ram_mem0_reg[212][5]/P0001  , \wishbone_bd_ram_mem0_reg[212][6]/P0001  , \wishbone_bd_ram_mem0_reg[212][7]/P0001  , \wishbone_bd_ram_mem0_reg[213][0]/P0001  , \wishbone_bd_ram_mem0_reg[213][1]/P0001  , \wishbone_bd_ram_mem0_reg[213][2]/P0001  , \wishbone_bd_ram_mem0_reg[213][3]/P0001  , \wishbone_bd_ram_mem0_reg[213][4]/P0001  , \wishbone_bd_ram_mem0_reg[213][5]/P0001  , \wishbone_bd_ram_mem0_reg[213][6]/P0001  , \wishbone_bd_ram_mem0_reg[213][7]/P0001  , \wishbone_bd_ram_mem0_reg[214][0]/P0001  , \wishbone_bd_ram_mem0_reg[214][1]/P0001  , \wishbone_bd_ram_mem0_reg[214][2]/P0001  , \wishbone_bd_ram_mem0_reg[214][3]/P0001  , \wishbone_bd_ram_mem0_reg[214][4]/P0001  , \wishbone_bd_ram_mem0_reg[214][5]/P0001  , \wishbone_bd_ram_mem0_reg[214][6]/P0001  , \wishbone_bd_ram_mem0_reg[214][7]/P0001  , \wishbone_bd_ram_mem0_reg[215][0]/P0001  , \wishbone_bd_ram_mem0_reg[215][1]/P0001  , \wishbone_bd_ram_mem0_reg[215][2]/P0001  , \wishbone_bd_ram_mem0_reg[215][3]/P0001  , \wishbone_bd_ram_mem0_reg[215][4]/P0001  , \wishbone_bd_ram_mem0_reg[215][5]/P0001  , \wishbone_bd_ram_mem0_reg[215][6]/P0001  , \wishbone_bd_ram_mem0_reg[215][7]/P0001  , \wishbone_bd_ram_mem0_reg[216][0]/P0001  , \wishbone_bd_ram_mem0_reg[216][1]/P0001  , \wishbone_bd_ram_mem0_reg[216][2]/P0001  , \wishbone_bd_ram_mem0_reg[216][3]/P0001  , \wishbone_bd_ram_mem0_reg[216][4]/P0001  , \wishbone_bd_ram_mem0_reg[216][5]/P0001  , \wishbone_bd_ram_mem0_reg[216][6]/P0001  , \wishbone_bd_ram_mem0_reg[216][7]/P0001  , \wishbone_bd_ram_mem0_reg[217][0]/P0001  , \wishbone_bd_ram_mem0_reg[217][1]/P0001  , \wishbone_bd_ram_mem0_reg[217][2]/P0001  , \wishbone_bd_ram_mem0_reg[217][3]/P0001  , \wishbone_bd_ram_mem0_reg[217][4]/P0001  , \wishbone_bd_ram_mem0_reg[217][5]/P0001  , \wishbone_bd_ram_mem0_reg[217][6]/P0001  , \wishbone_bd_ram_mem0_reg[217][7]/P0001  , \wishbone_bd_ram_mem0_reg[218][0]/P0001  , \wishbone_bd_ram_mem0_reg[218][1]/P0001  , \wishbone_bd_ram_mem0_reg[218][2]/P0001  , \wishbone_bd_ram_mem0_reg[218][3]/P0001  , \wishbone_bd_ram_mem0_reg[218][4]/P0001  , \wishbone_bd_ram_mem0_reg[218][5]/P0001  , \wishbone_bd_ram_mem0_reg[218][6]/P0001  , \wishbone_bd_ram_mem0_reg[218][7]/P0001  , \wishbone_bd_ram_mem0_reg[219][0]/P0001  , \wishbone_bd_ram_mem0_reg[219][1]/P0001  , \wishbone_bd_ram_mem0_reg[219][2]/P0001  , \wishbone_bd_ram_mem0_reg[219][3]/P0001  , \wishbone_bd_ram_mem0_reg[219][4]/P0001  , \wishbone_bd_ram_mem0_reg[219][5]/P0001  , \wishbone_bd_ram_mem0_reg[219][6]/P0001  , \wishbone_bd_ram_mem0_reg[219][7]/P0001  , \wishbone_bd_ram_mem0_reg[21][0]/P0001  , \wishbone_bd_ram_mem0_reg[21][1]/P0001  , \wishbone_bd_ram_mem0_reg[21][2]/P0001  , \wishbone_bd_ram_mem0_reg[21][3]/P0001  , \wishbone_bd_ram_mem0_reg[21][4]/P0001  , \wishbone_bd_ram_mem0_reg[21][5]/P0001  , \wishbone_bd_ram_mem0_reg[21][6]/P0001  , \wishbone_bd_ram_mem0_reg[21][7]/P0001  , \wishbone_bd_ram_mem0_reg[220][0]/P0001  , \wishbone_bd_ram_mem0_reg[220][1]/P0001  , \wishbone_bd_ram_mem0_reg[220][2]/P0001  , \wishbone_bd_ram_mem0_reg[220][3]/P0001  , \wishbone_bd_ram_mem0_reg[220][4]/P0001  , \wishbone_bd_ram_mem0_reg[220][5]/P0001  , \wishbone_bd_ram_mem0_reg[220][6]/P0001  , \wishbone_bd_ram_mem0_reg[220][7]/P0001  , \wishbone_bd_ram_mem0_reg[221][0]/P0001  , \wishbone_bd_ram_mem0_reg[221][1]/P0001  , \wishbone_bd_ram_mem0_reg[221][2]/P0001  , \wishbone_bd_ram_mem0_reg[221][3]/P0001  , \wishbone_bd_ram_mem0_reg[221][4]/P0001  , \wishbone_bd_ram_mem0_reg[221][5]/P0001  , \wishbone_bd_ram_mem0_reg[221][6]/P0001  , \wishbone_bd_ram_mem0_reg[221][7]/P0001  , \wishbone_bd_ram_mem0_reg[222][0]/P0001  , \wishbone_bd_ram_mem0_reg[222][1]/P0001  , \wishbone_bd_ram_mem0_reg[222][2]/P0001  , \wishbone_bd_ram_mem0_reg[222][3]/P0001  , \wishbone_bd_ram_mem0_reg[222][4]/P0001  , \wishbone_bd_ram_mem0_reg[222][5]/P0001  , \wishbone_bd_ram_mem0_reg[222][6]/P0001  , \wishbone_bd_ram_mem0_reg[222][7]/P0001  , \wishbone_bd_ram_mem0_reg[223][0]/P0001  , \wishbone_bd_ram_mem0_reg[223][1]/P0001  , \wishbone_bd_ram_mem0_reg[223][2]/P0001  , \wishbone_bd_ram_mem0_reg[223][3]/P0001  , \wishbone_bd_ram_mem0_reg[223][4]/P0001  , \wishbone_bd_ram_mem0_reg[223][5]/P0001  , \wishbone_bd_ram_mem0_reg[223][6]/P0001  , \wishbone_bd_ram_mem0_reg[223][7]/P0001  , \wishbone_bd_ram_mem0_reg[224][0]/P0001  , \wishbone_bd_ram_mem0_reg[224][1]/P0001  , \wishbone_bd_ram_mem0_reg[224][2]/P0001  , \wishbone_bd_ram_mem0_reg[224][3]/P0001  , \wishbone_bd_ram_mem0_reg[224][4]/P0001  , \wishbone_bd_ram_mem0_reg[224][5]/P0001  , \wishbone_bd_ram_mem0_reg[224][6]/P0001  , \wishbone_bd_ram_mem0_reg[224][7]/P0001  , \wishbone_bd_ram_mem0_reg[225][0]/P0001  , \wishbone_bd_ram_mem0_reg[225][1]/P0001  , \wishbone_bd_ram_mem0_reg[225][2]/P0001  , \wishbone_bd_ram_mem0_reg[225][3]/P0001  , \wishbone_bd_ram_mem0_reg[225][4]/P0001  , \wishbone_bd_ram_mem0_reg[225][5]/P0001  , \wishbone_bd_ram_mem0_reg[225][6]/P0001  , \wishbone_bd_ram_mem0_reg[225][7]/P0001  , \wishbone_bd_ram_mem0_reg[226][0]/P0001  , \wishbone_bd_ram_mem0_reg[226][1]/P0001  , \wishbone_bd_ram_mem0_reg[226][2]/P0001  , \wishbone_bd_ram_mem0_reg[226][3]/P0001  , \wishbone_bd_ram_mem0_reg[226][4]/P0001  , \wishbone_bd_ram_mem0_reg[226][5]/P0001  , \wishbone_bd_ram_mem0_reg[226][6]/P0001  , \wishbone_bd_ram_mem0_reg[226][7]/P0001  , \wishbone_bd_ram_mem0_reg[227][0]/P0001  , \wishbone_bd_ram_mem0_reg[227][1]/P0001  , \wishbone_bd_ram_mem0_reg[227][2]/P0001  , \wishbone_bd_ram_mem0_reg[227][3]/P0001  , \wishbone_bd_ram_mem0_reg[227][4]/P0001  , \wishbone_bd_ram_mem0_reg[227][5]/P0001  , \wishbone_bd_ram_mem0_reg[227][6]/P0001  , \wishbone_bd_ram_mem0_reg[227][7]/P0001  , \wishbone_bd_ram_mem0_reg[228][0]/P0001  , \wishbone_bd_ram_mem0_reg[228][1]/P0001  , \wishbone_bd_ram_mem0_reg[228][2]/P0001  , \wishbone_bd_ram_mem0_reg[228][3]/P0001  , \wishbone_bd_ram_mem0_reg[228][4]/P0001  , \wishbone_bd_ram_mem0_reg[228][5]/P0001  , \wishbone_bd_ram_mem0_reg[228][6]/P0001  , \wishbone_bd_ram_mem0_reg[228][7]/P0001  , \wishbone_bd_ram_mem0_reg[229][0]/P0001  , \wishbone_bd_ram_mem0_reg[229][1]/P0001  , \wishbone_bd_ram_mem0_reg[229][2]/P0001  , \wishbone_bd_ram_mem0_reg[229][3]/P0001  , \wishbone_bd_ram_mem0_reg[229][4]/P0001  , \wishbone_bd_ram_mem0_reg[229][5]/P0001  , \wishbone_bd_ram_mem0_reg[229][6]/P0001  , \wishbone_bd_ram_mem0_reg[229][7]/P0001  , \wishbone_bd_ram_mem0_reg[22][0]/P0001  , \wishbone_bd_ram_mem0_reg[22][1]/P0001  , \wishbone_bd_ram_mem0_reg[22][2]/P0001  , \wishbone_bd_ram_mem0_reg[22][3]/P0001  , \wishbone_bd_ram_mem0_reg[22][4]/P0001  , \wishbone_bd_ram_mem0_reg[22][5]/P0001  , \wishbone_bd_ram_mem0_reg[22][6]/P0001  , \wishbone_bd_ram_mem0_reg[22][7]/P0001  , \wishbone_bd_ram_mem0_reg[230][0]/P0001  , \wishbone_bd_ram_mem0_reg[230][1]/P0001  , \wishbone_bd_ram_mem0_reg[230][2]/P0001  , \wishbone_bd_ram_mem0_reg[230][3]/P0001  , \wishbone_bd_ram_mem0_reg[230][4]/P0001  , \wishbone_bd_ram_mem0_reg[230][5]/P0001  , \wishbone_bd_ram_mem0_reg[230][6]/P0001  , \wishbone_bd_ram_mem0_reg[230][7]/P0001  , \wishbone_bd_ram_mem0_reg[231][0]/P0001  , \wishbone_bd_ram_mem0_reg[231][1]/P0001  , \wishbone_bd_ram_mem0_reg[231][2]/P0001  , \wishbone_bd_ram_mem0_reg[231][3]/P0001  , \wishbone_bd_ram_mem0_reg[231][4]/P0001  , \wishbone_bd_ram_mem0_reg[231][5]/P0001  , \wishbone_bd_ram_mem0_reg[231][6]/P0001  , \wishbone_bd_ram_mem0_reg[231][7]/P0001  , \wishbone_bd_ram_mem0_reg[232][0]/P0001  , \wishbone_bd_ram_mem0_reg[232][1]/P0001  , \wishbone_bd_ram_mem0_reg[232][2]/P0001  , \wishbone_bd_ram_mem0_reg[232][3]/P0001  , \wishbone_bd_ram_mem0_reg[232][4]/P0001  , \wishbone_bd_ram_mem0_reg[232][5]/P0001  , \wishbone_bd_ram_mem0_reg[232][6]/P0001  , \wishbone_bd_ram_mem0_reg[232][7]/P0001  , \wishbone_bd_ram_mem0_reg[233][0]/P0001  , \wishbone_bd_ram_mem0_reg[233][1]/P0001  , \wishbone_bd_ram_mem0_reg[233][2]/P0001  , \wishbone_bd_ram_mem0_reg[233][3]/P0001  , \wishbone_bd_ram_mem0_reg[233][4]/P0001  , \wishbone_bd_ram_mem0_reg[233][5]/P0001  , \wishbone_bd_ram_mem0_reg[233][6]/P0001  , \wishbone_bd_ram_mem0_reg[233][7]/P0001  , \wishbone_bd_ram_mem0_reg[234][0]/P0001  , \wishbone_bd_ram_mem0_reg[234][1]/P0001  , \wishbone_bd_ram_mem0_reg[234][2]/P0001  , \wishbone_bd_ram_mem0_reg[234][3]/P0001  , \wishbone_bd_ram_mem0_reg[234][4]/P0001  , \wishbone_bd_ram_mem0_reg[234][5]/P0001  , \wishbone_bd_ram_mem0_reg[234][6]/P0001  , \wishbone_bd_ram_mem0_reg[234][7]/P0001  , \wishbone_bd_ram_mem0_reg[235][0]/P0001  , \wishbone_bd_ram_mem0_reg[235][1]/P0001  , \wishbone_bd_ram_mem0_reg[235][2]/P0001  , \wishbone_bd_ram_mem0_reg[235][3]/P0001  , \wishbone_bd_ram_mem0_reg[235][4]/P0001  , \wishbone_bd_ram_mem0_reg[235][5]/P0001  , \wishbone_bd_ram_mem0_reg[235][6]/P0001  , \wishbone_bd_ram_mem0_reg[235][7]/P0001  , \wishbone_bd_ram_mem0_reg[236][0]/P0001  , \wishbone_bd_ram_mem0_reg[236][1]/P0001  , \wishbone_bd_ram_mem0_reg[236][2]/P0001  , \wishbone_bd_ram_mem0_reg[236][3]/P0001  , \wishbone_bd_ram_mem0_reg[236][4]/P0001  , \wishbone_bd_ram_mem0_reg[236][5]/P0001  , \wishbone_bd_ram_mem0_reg[236][6]/P0001  , \wishbone_bd_ram_mem0_reg[236][7]/P0001  , \wishbone_bd_ram_mem0_reg[237][0]/P0001  , \wishbone_bd_ram_mem0_reg[237][1]/P0001  , \wishbone_bd_ram_mem0_reg[237][2]/P0001  , \wishbone_bd_ram_mem0_reg[237][3]/P0001  , \wishbone_bd_ram_mem0_reg[237][4]/P0001  , \wishbone_bd_ram_mem0_reg[237][5]/P0001  , \wishbone_bd_ram_mem0_reg[237][6]/P0001  , \wishbone_bd_ram_mem0_reg[237][7]/P0001  , \wishbone_bd_ram_mem0_reg[238][0]/P0001  , \wishbone_bd_ram_mem0_reg[238][1]/P0001  , \wishbone_bd_ram_mem0_reg[238][2]/P0001  , \wishbone_bd_ram_mem0_reg[238][3]/P0001  , \wishbone_bd_ram_mem0_reg[238][4]/P0001  , \wishbone_bd_ram_mem0_reg[238][5]/P0001  , \wishbone_bd_ram_mem0_reg[238][6]/P0001  , \wishbone_bd_ram_mem0_reg[238][7]/P0001  , \wishbone_bd_ram_mem0_reg[239][0]/P0001  , \wishbone_bd_ram_mem0_reg[239][1]/P0001  , \wishbone_bd_ram_mem0_reg[239][2]/P0001  , \wishbone_bd_ram_mem0_reg[239][3]/P0001  , \wishbone_bd_ram_mem0_reg[239][4]/P0001  , \wishbone_bd_ram_mem0_reg[239][5]/P0001  , \wishbone_bd_ram_mem0_reg[239][6]/P0001  , \wishbone_bd_ram_mem0_reg[239][7]/P0001  , \wishbone_bd_ram_mem0_reg[23][0]/P0001  , \wishbone_bd_ram_mem0_reg[23][1]/P0001  , \wishbone_bd_ram_mem0_reg[23][2]/P0001  , \wishbone_bd_ram_mem0_reg[23][3]/P0001  , \wishbone_bd_ram_mem0_reg[23][4]/P0001  , \wishbone_bd_ram_mem0_reg[23][5]/P0001  , \wishbone_bd_ram_mem0_reg[23][6]/P0001  , \wishbone_bd_ram_mem0_reg[23][7]/P0001  , \wishbone_bd_ram_mem0_reg[240][0]/P0001  , \wishbone_bd_ram_mem0_reg[240][1]/P0001  , \wishbone_bd_ram_mem0_reg[240][2]/P0001  , \wishbone_bd_ram_mem0_reg[240][3]/P0001  , \wishbone_bd_ram_mem0_reg[240][4]/P0001  , \wishbone_bd_ram_mem0_reg[240][5]/P0001  , \wishbone_bd_ram_mem0_reg[240][6]/P0001  , \wishbone_bd_ram_mem0_reg[240][7]/P0001  , \wishbone_bd_ram_mem0_reg[241][0]/P0001  , \wishbone_bd_ram_mem0_reg[241][1]/P0001  , \wishbone_bd_ram_mem0_reg[241][2]/P0001  , \wishbone_bd_ram_mem0_reg[241][3]/P0001  , \wishbone_bd_ram_mem0_reg[241][4]/P0001  , \wishbone_bd_ram_mem0_reg[241][5]/P0001  , \wishbone_bd_ram_mem0_reg[241][6]/P0001  , \wishbone_bd_ram_mem0_reg[241][7]/P0001  , \wishbone_bd_ram_mem0_reg[242][0]/P0001  , \wishbone_bd_ram_mem0_reg[242][1]/P0001  , \wishbone_bd_ram_mem0_reg[242][2]/P0001  , \wishbone_bd_ram_mem0_reg[242][3]/P0001  , \wishbone_bd_ram_mem0_reg[242][4]/P0001  , \wishbone_bd_ram_mem0_reg[242][5]/P0001  , \wishbone_bd_ram_mem0_reg[242][6]/P0001  , \wishbone_bd_ram_mem0_reg[242][7]/P0001  , \wishbone_bd_ram_mem0_reg[243][0]/P0001  , \wishbone_bd_ram_mem0_reg[243][1]/P0001  , \wishbone_bd_ram_mem0_reg[243][2]/P0001  , \wishbone_bd_ram_mem0_reg[243][3]/P0001  , \wishbone_bd_ram_mem0_reg[243][4]/P0001  , \wishbone_bd_ram_mem0_reg[243][5]/P0001  , \wishbone_bd_ram_mem0_reg[243][6]/P0001  , \wishbone_bd_ram_mem0_reg[243][7]/P0001  , \wishbone_bd_ram_mem0_reg[244][0]/P0001  , \wishbone_bd_ram_mem0_reg[244][1]/P0001  , \wishbone_bd_ram_mem0_reg[244][2]/P0001  , \wishbone_bd_ram_mem0_reg[244][3]/P0001  , \wishbone_bd_ram_mem0_reg[244][4]/P0001  , \wishbone_bd_ram_mem0_reg[244][5]/P0001  , \wishbone_bd_ram_mem0_reg[244][6]/P0001  , \wishbone_bd_ram_mem0_reg[244][7]/P0001  , \wishbone_bd_ram_mem0_reg[245][0]/P0001  , \wishbone_bd_ram_mem0_reg[245][1]/P0001  , \wishbone_bd_ram_mem0_reg[245][2]/P0001  , \wishbone_bd_ram_mem0_reg[245][3]/P0001  , \wishbone_bd_ram_mem0_reg[245][4]/P0001  , \wishbone_bd_ram_mem0_reg[245][5]/P0001  , \wishbone_bd_ram_mem0_reg[245][6]/P0001  , \wishbone_bd_ram_mem0_reg[245][7]/P0001  , \wishbone_bd_ram_mem0_reg[246][0]/P0001  , \wishbone_bd_ram_mem0_reg[246][1]/P0001  , \wishbone_bd_ram_mem0_reg[246][2]/P0001  , \wishbone_bd_ram_mem0_reg[246][3]/P0001  , \wishbone_bd_ram_mem0_reg[246][4]/P0001  , \wishbone_bd_ram_mem0_reg[246][5]/P0001  , \wishbone_bd_ram_mem0_reg[246][6]/P0001  , \wishbone_bd_ram_mem0_reg[246][7]/P0001  , \wishbone_bd_ram_mem0_reg[247][0]/P0001  , \wishbone_bd_ram_mem0_reg[247][1]/P0001  , \wishbone_bd_ram_mem0_reg[247][2]/P0001  , \wishbone_bd_ram_mem0_reg[247][3]/P0001  , \wishbone_bd_ram_mem0_reg[247][4]/P0001  , \wishbone_bd_ram_mem0_reg[247][5]/P0001  , \wishbone_bd_ram_mem0_reg[247][6]/P0001  , \wishbone_bd_ram_mem0_reg[247][7]/P0001  , \wishbone_bd_ram_mem0_reg[248][0]/P0001  , \wishbone_bd_ram_mem0_reg[248][1]/P0001  , \wishbone_bd_ram_mem0_reg[248][2]/P0001  , \wishbone_bd_ram_mem0_reg[248][3]/P0001  , \wishbone_bd_ram_mem0_reg[248][4]/P0001  , \wishbone_bd_ram_mem0_reg[248][5]/P0001  , \wishbone_bd_ram_mem0_reg[248][6]/P0001  , \wishbone_bd_ram_mem0_reg[248][7]/P0001  , \wishbone_bd_ram_mem0_reg[249][0]/P0001  , \wishbone_bd_ram_mem0_reg[249][1]/P0001  , \wishbone_bd_ram_mem0_reg[249][2]/P0001  , \wishbone_bd_ram_mem0_reg[249][3]/P0001  , \wishbone_bd_ram_mem0_reg[249][4]/P0001  , \wishbone_bd_ram_mem0_reg[249][5]/P0001  , \wishbone_bd_ram_mem0_reg[249][6]/P0001  , \wishbone_bd_ram_mem0_reg[249][7]/P0001  , \wishbone_bd_ram_mem0_reg[24][0]/P0001  , \wishbone_bd_ram_mem0_reg[24][1]/P0001  , \wishbone_bd_ram_mem0_reg[24][2]/P0001  , \wishbone_bd_ram_mem0_reg[24][3]/P0001  , \wishbone_bd_ram_mem0_reg[24][4]/P0001  , \wishbone_bd_ram_mem0_reg[24][5]/P0001  , \wishbone_bd_ram_mem0_reg[24][6]/P0001  , \wishbone_bd_ram_mem0_reg[24][7]/P0001  , \wishbone_bd_ram_mem0_reg[250][0]/P0001  , \wishbone_bd_ram_mem0_reg[250][1]/P0001  , \wishbone_bd_ram_mem0_reg[250][2]/P0001  , \wishbone_bd_ram_mem0_reg[250][3]/P0001  , \wishbone_bd_ram_mem0_reg[250][4]/P0001  , \wishbone_bd_ram_mem0_reg[250][5]/P0001  , \wishbone_bd_ram_mem0_reg[250][6]/P0001  , \wishbone_bd_ram_mem0_reg[250][7]/P0001  , \wishbone_bd_ram_mem0_reg[251][0]/P0001  , \wishbone_bd_ram_mem0_reg[251][1]/P0001  , \wishbone_bd_ram_mem0_reg[251][2]/P0001  , \wishbone_bd_ram_mem0_reg[251][3]/P0001  , \wishbone_bd_ram_mem0_reg[251][4]/P0001  , \wishbone_bd_ram_mem0_reg[251][5]/P0001  , \wishbone_bd_ram_mem0_reg[251][6]/P0001  , \wishbone_bd_ram_mem0_reg[251][7]/P0001  , \wishbone_bd_ram_mem0_reg[252][0]/P0001  , \wishbone_bd_ram_mem0_reg[252][1]/P0001  , \wishbone_bd_ram_mem0_reg[252][2]/P0001  , \wishbone_bd_ram_mem0_reg[252][3]/P0001  , \wishbone_bd_ram_mem0_reg[252][4]/P0001  , \wishbone_bd_ram_mem0_reg[252][5]/P0001  , \wishbone_bd_ram_mem0_reg[252][6]/P0001  , \wishbone_bd_ram_mem0_reg[252][7]/P0001  , \wishbone_bd_ram_mem0_reg[253][0]/P0001  , \wishbone_bd_ram_mem0_reg[253][1]/P0001  , \wishbone_bd_ram_mem0_reg[253][2]/P0001  , \wishbone_bd_ram_mem0_reg[253][3]/P0001  , \wishbone_bd_ram_mem0_reg[253][4]/P0001  , \wishbone_bd_ram_mem0_reg[253][5]/P0001  , \wishbone_bd_ram_mem0_reg[253][6]/P0001  , \wishbone_bd_ram_mem0_reg[253][7]/P0001  , \wishbone_bd_ram_mem0_reg[254][0]/P0001  , \wishbone_bd_ram_mem0_reg[254][1]/P0001  , \wishbone_bd_ram_mem0_reg[254][2]/P0001  , \wishbone_bd_ram_mem0_reg[254][3]/P0001  , \wishbone_bd_ram_mem0_reg[254][4]/P0001  , \wishbone_bd_ram_mem0_reg[254][5]/P0001  , \wishbone_bd_ram_mem0_reg[254][6]/P0001  , \wishbone_bd_ram_mem0_reg[254][7]/P0001  , \wishbone_bd_ram_mem0_reg[255][0]/P0001  , \wishbone_bd_ram_mem0_reg[255][1]/P0001  , \wishbone_bd_ram_mem0_reg[255][2]/P0001  , \wishbone_bd_ram_mem0_reg[255][3]/P0001  , \wishbone_bd_ram_mem0_reg[255][4]/P0001  , \wishbone_bd_ram_mem0_reg[255][5]/P0001  , \wishbone_bd_ram_mem0_reg[255][6]/P0001  , \wishbone_bd_ram_mem0_reg[255][7]/P0001  , \wishbone_bd_ram_mem0_reg[25][0]/P0001  , \wishbone_bd_ram_mem0_reg[25][1]/P0001  , \wishbone_bd_ram_mem0_reg[25][2]/P0001  , \wishbone_bd_ram_mem0_reg[25][3]/P0001  , \wishbone_bd_ram_mem0_reg[25][4]/P0001  , \wishbone_bd_ram_mem0_reg[25][5]/P0001  , \wishbone_bd_ram_mem0_reg[25][6]/P0001  , \wishbone_bd_ram_mem0_reg[25][7]/P0001  , \wishbone_bd_ram_mem0_reg[26][0]/P0001  , \wishbone_bd_ram_mem0_reg[26][1]/P0001  , \wishbone_bd_ram_mem0_reg[26][2]/P0001  , \wishbone_bd_ram_mem0_reg[26][3]/P0001  , \wishbone_bd_ram_mem0_reg[26][4]/P0001  , \wishbone_bd_ram_mem0_reg[26][5]/P0001  , \wishbone_bd_ram_mem0_reg[26][6]/P0001  , \wishbone_bd_ram_mem0_reg[26][7]/P0001  , \wishbone_bd_ram_mem0_reg[27][0]/P0001  , \wishbone_bd_ram_mem0_reg[27][1]/P0001  , \wishbone_bd_ram_mem0_reg[27][2]/P0001  , \wishbone_bd_ram_mem0_reg[27][3]/P0001  , \wishbone_bd_ram_mem0_reg[27][4]/P0001  , \wishbone_bd_ram_mem0_reg[27][5]/P0001  , \wishbone_bd_ram_mem0_reg[27][6]/P0001  , \wishbone_bd_ram_mem0_reg[27][7]/P0001  , \wishbone_bd_ram_mem0_reg[28][0]/P0001  , \wishbone_bd_ram_mem0_reg[28][1]/P0001  , \wishbone_bd_ram_mem0_reg[28][2]/P0001  , \wishbone_bd_ram_mem0_reg[28][3]/P0001  , \wishbone_bd_ram_mem0_reg[28][4]/P0001  , \wishbone_bd_ram_mem0_reg[28][5]/P0001  , \wishbone_bd_ram_mem0_reg[28][6]/P0001  , \wishbone_bd_ram_mem0_reg[28][7]/P0001  , \wishbone_bd_ram_mem0_reg[29][0]/P0001  , \wishbone_bd_ram_mem0_reg[29][1]/P0001  , \wishbone_bd_ram_mem0_reg[29][2]/P0001  , \wishbone_bd_ram_mem0_reg[29][3]/P0001  , \wishbone_bd_ram_mem0_reg[29][4]/P0001  , \wishbone_bd_ram_mem0_reg[29][5]/P0001  , \wishbone_bd_ram_mem0_reg[29][6]/P0001  , \wishbone_bd_ram_mem0_reg[29][7]/P0001  , \wishbone_bd_ram_mem0_reg[2][0]/P0001  , \wishbone_bd_ram_mem0_reg[2][1]/P0001  , \wishbone_bd_ram_mem0_reg[2][2]/P0001  , \wishbone_bd_ram_mem0_reg[2][3]/P0001  , \wishbone_bd_ram_mem0_reg[2][4]/P0001  , \wishbone_bd_ram_mem0_reg[2][5]/P0001  , \wishbone_bd_ram_mem0_reg[2][6]/P0001  , \wishbone_bd_ram_mem0_reg[2][7]/P0001  , \wishbone_bd_ram_mem0_reg[30][0]/P0001  , \wishbone_bd_ram_mem0_reg[30][1]/P0001  , \wishbone_bd_ram_mem0_reg[30][2]/P0001  , \wishbone_bd_ram_mem0_reg[30][3]/P0001  , \wishbone_bd_ram_mem0_reg[30][4]/P0001  , \wishbone_bd_ram_mem0_reg[30][5]/P0001  , \wishbone_bd_ram_mem0_reg[30][6]/P0001  , \wishbone_bd_ram_mem0_reg[30][7]/P0001  , \wishbone_bd_ram_mem0_reg[31][0]/P0001  , \wishbone_bd_ram_mem0_reg[31][1]/P0001  , \wishbone_bd_ram_mem0_reg[31][2]/P0001  , \wishbone_bd_ram_mem0_reg[31][3]/P0001  , \wishbone_bd_ram_mem0_reg[31][4]/P0001  , \wishbone_bd_ram_mem0_reg[31][5]/P0001  , \wishbone_bd_ram_mem0_reg[31][6]/P0001  , \wishbone_bd_ram_mem0_reg[31][7]/P0001  , \wishbone_bd_ram_mem0_reg[32][0]/P0001  , \wishbone_bd_ram_mem0_reg[32][1]/P0001  , \wishbone_bd_ram_mem0_reg[32][2]/P0001  , \wishbone_bd_ram_mem0_reg[32][3]/P0001  , \wishbone_bd_ram_mem0_reg[32][4]/P0001  , \wishbone_bd_ram_mem0_reg[32][5]/P0001  , \wishbone_bd_ram_mem0_reg[32][6]/P0001  , \wishbone_bd_ram_mem0_reg[32][7]/P0001  , \wishbone_bd_ram_mem0_reg[33][0]/P0001  , \wishbone_bd_ram_mem0_reg[33][1]/P0001  , \wishbone_bd_ram_mem0_reg[33][2]/P0001  , \wishbone_bd_ram_mem0_reg[33][3]/P0001  , \wishbone_bd_ram_mem0_reg[33][4]/P0001  , \wishbone_bd_ram_mem0_reg[33][5]/P0001  , \wishbone_bd_ram_mem0_reg[33][6]/P0001  , \wishbone_bd_ram_mem0_reg[33][7]/P0001  , \wishbone_bd_ram_mem0_reg[34][0]/P0001  , \wishbone_bd_ram_mem0_reg[34][1]/P0001  , \wishbone_bd_ram_mem0_reg[34][2]/P0001  , \wishbone_bd_ram_mem0_reg[34][3]/P0001  , \wishbone_bd_ram_mem0_reg[34][4]/P0001  , \wishbone_bd_ram_mem0_reg[34][5]/P0001  , \wishbone_bd_ram_mem0_reg[34][6]/P0001  , \wishbone_bd_ram_mem0_reg[34][7]/P0001  , \wishbone_bd_ram_mem0_reg[35][0]/P0001  , \wishbone_bd_ram_mem0_reg[35][1]/P0001  , \wishbone_bd_ram_mem0_reg[35][2]/P0001  , \wishbone_bd_ram_mem0_reg[35][3]/P0001  , \wishbone_bd_ram_mem0_reg[35][4]/P0001  , \wishbone_bd_ram_mem0_reg[35][5]/P0001  , \wishbone_bd_ram_mem0_reg[35][6]/P0001  , \wishbone_bd_ram_mem0_reg[35][7]/P0001  , \wishbone_bd_ram_mem0_reg[36][0]/P0001  , \wishbone_bd_ram_mem0_reg[36][1]/P0001  , \wishbone_bd_ram_mem0_reg[36][2]/P0001  , \wishbone_bd_ram_mem0_reg[36][3]/P0001  , \wishbone_bd_ram_mem0_reg[36][4]/P0001  , \wishbone_bd_ram_mem0_reg[36][5]/P0001  , \wishbone_bd_ram_mem0_reg[36][6]/P0001  , \wishbone_bd_ram_mem0_reg[36][7]/P0001  , \wishbone_bd_ram_mem0_reg[37][0]/P0001  , \wishbone_bd_ram_mem0_reg[37][1]/P0001  , \wishbone_bd_ram_mem0_reg[37][2]/P0001  , \wishbone_bd_ram_mem0_reg[37][3]/P0001  , \wishbone_bd_ram_mem0_reg[37][4]/P0001  , \wishbone_bd_ram_mem0_reg[37][5]/P0001  , \wishbone_bd_ram_mem0_reg[37][6]/P0001  , \wishbone_bd_ram_mem0_reg[37][7]/P0001  , \wishbone_bd_ram_mem0_reg[38][0]/P0001  , \wishbone_bd_ram_mem0_reg[38][1]/P0001  , \wishbone_bd_ram_mem0_reg[38][2]/P0001  , \wishbone_bd_ram_mem0_reg[38][3]/P0001  , \wishbone_bd_ram_mem0_reg[38][4]/P0001  , \wishbone_bd_ram_mem0_reg[38][5]/P0001  , \wishbone_bd_ram_mem0_reg[38][6]/P0001  , \wishbone_bd_ram_mem0_reg[38][7]/P0001  , \wishbone_bd_ram_mem0_reg[39][0]/P0001  , \wishbone_bd_ram_mem0_reg[39][1]/P0001  , \wishbone_bd_ram_mem0_reg[39][2]/P0001  , \wishbone_bd_ram_mem0_reg[39][3]/P0001  , \wishbone_bd_ram_mem0_reg[39][4]/P0001  , \wishbone_bd_ram_mem0_reg[39][5]/P0001  , \wishbone_bd_ram_mem0_reg[39][6]/P0001  , \wishbone_bd_ram_mem0_reg[39][7]/P0001  , \wishbone_bd_ram_mem0_reg[3][0]/P0001  , \wishbone_bd_ram_mem0_reg[3][1]/P0001  , \wishbone_bd_ram_mem0_reg[3][2]/P0001  , \wishbone_bd_ram_mem0_reg[3][3]/P0001  , \wishbone_bd_ram_mem0_reg[3][4]/P0001  , \wishbone_bd_ram_mem0_reg[3][5]/P0001  , \wishbone_bd_ram_mem0_reg[3][6]/P0001  , \wishbone_bd_ram_mem0_reg[3][7]/P0001  , \wishbone_bd_ram_mem0_reg[40][0]/P0001  , \wishbone_bd_ram_mem0_reg[40][1]/P0001  , \wishbone_bd_ram_mem0_reg[40][2]/P0001  , \wishbone_bd_ram_mem0_reg[40][3]/P0001  , \wishbone_bd_ram_mem0_reg[40][4]/P0001  , \wishbone_bd_ram_mem0_reg[40][5]/P0001  , \wishbone_bd_ram_mem0_reg[40][6]/P0001  , \wishbone_bd_ram_mem0_reg[40][7]/P0001  , \wishbone_bd_ram_mem0_reg[41][0]/P0001  , \wishbone_bd_ram_mem0_reg[41][1]/P0001  , \wishbone_bd_ram_mem0_reg[41][2]/P0001  , \wishbone_bd_ram_mem0_reg[41][3]/P0001  , \wishbone_bd_ram_mem0_reg[41][4]/P0001  , \wishbone_bd_ram_mem0_reg[41][5]/P0001  , \wishbone_bd_ram_mem0_reg[41][6]/P0001  , \wishbone_bd_ram_mem0_reg[41][7]/P0001  , \wishbone_bd_ram_mem0_reg[42][0]/P0001  , \wishbone_bd_ram_mem0_reg[42][1]/P0001  , \wishbone_bd_ram_mem0_reg[42][2]/P0001  , \wishbone_bd_ram_mem0_reg[42][3]/P0001  , \wishbone_bd_ram_mem0_reg[42][4]/P0001  , \wishbone_bd_ram_mem0_reg[42][5]/P0001  , \wishbone_bd_ram_mem0_reg[42][6]/P0001  , \wishbone_bd_ram_mem0_reg[42][7]/P0001  , \wishbone_bd_ram_mem0_reg[43][0]/P0001  , \wishbone_bd_ram_mem0_reg[43][1]/P0001  , \wishbone_bd_ram_mem0_reg[43][2]/P0001  , \wishbone_bd_ram_mem0_reg[43][3]/P0001  , \wishbone_bd_ram_mem0_reg[43][4]/P0001  , \wishbone_bd_ram_mem0_reg[43][5]/P0001  , \wishbone_bd_ram_mem0_reg[43][6]/P0001  , \wishbone_bd_ram_mem0_reg[43][7]/P0001  , \wishbone_bd_ram_mem0_reg[44][0]/P0001  , \wishbone_bd_ram_mem0_reg[44][1]/P0001  , \wishbone_bd_ram_mem0_reg[44][2]/P0001  , \wishbone_bd_ram_mem0_reg[44][3]/P0001  , \wishbone_bd_ram_mem0_reg[44][4]/P0001  , \wishbone_bd_ram_mem0_reg[44][5]/P0001  , \wishbone_bd_ram_mem0_reg[44][6]/P0001  , \wishbone_bd_ram_mem0_reg[44][7]/P0001  , \wishbone_bd_ram_mem0_reg[45][0]/P0001  , \wishbone_bd_ram_mem0_reg[45][1]/P0001  , \wishbone_bd_ram_mem0_reg[45][2]/P0001  , \wishbone_bd_ram_mem0_reg[45][3]/P0001  , \wishbone_bd_ram_mem0_reg[45][4]/P0001  , \wishbone_bd_ram_mem0_reg[45][5]/P0001  , \wishbone_bd_ram_mem0_reg[45][6]/P0001  , \wishbone_bd_ram_mem0_reg[45][7]/P0001  , \wishbone_bd_ram_mem0_reg[46][0]/P0001  , \wishbone_bd_ram_mem0_reg[46][1]/P0001  , \wishbone_bd_ram_mem0_reg[46][2]/P0001  , \wishbone_bd_ram_mem0_reg[46][3]/P0001  , \wishbone_bd_ram_mem0_reg[46][4]/P0001  , \wishbone_bd_ram_mem0_reg[46][5]/P0001  , \wishbone_bd_ram_mem0_reg[46][6]/P0001  , \wishbone_bd_ram_mem0_reg[46][7]/P0001  , \wishbone_bd_ram_mem0_reg[47][0]/P0001  , \wishbone_bd_ram_mem0_reg[47][1]/P0001  , \wishbone_bd_ram_mem0_reg[47][2]/P0001  , \wishbone_bd_ram_mem0_reg[47][3]/P0001  , \wishbone_bd_ram_mem0_reg[47][4]/P0001  , \wishbone_bd_ram_mem0_reg[47][5]/P0001  , \wishbone_bd_ram_mem0_reg[47][6]/P0001  , \wishbone_bd_ram_mem0_reg[47][7]/P0001  , \wishbone_bd_ram_mem0_reg[48][0]/P0001  , \wishbone_bd_ram_mem0_reg[48][1]/P0001  , \wishbone_bd_ram_mem0_reg[48][2]/P0001  , \wishbone_bd_ram_mem0_reg[48][3]/P0001  , \wishbone_bd_ram_mem0_reg[48][4]/P0001  , \wishbone_bd_ram_mem0_reg[48][5]/P0001  , \wishbone_bd_ram_mem0_reg[48][6]/P0001  , \wishbone_bd_ram_mem0_reg[48][7]/P0001  , \wishbone_bd_ram_mem0_reg[49][0]/P0001  , \wishbone_bd_ram_mem0_reg[49][1]/P0001  , \wishbone_bd_ram_mem0_reg[49][2]/P0001  , \wishbone_bd_ram_mem0_reg[49][3]/P0001  , \wishbone_bd_ram_mem0_reg[49][4]/P0001  , \wishbone_bd_ram_mem0_reg[49][5]/P0001  , \wishbone_bd_ram_mem0_reg[49][6]/P0001  , \wishbone_bd_ram_mem0_reg[49][7]/P0001  , \wishbone_bd_ram_mem0_reg[4][0]/P0001  , \wishbone_bd_ram_mem0_reg[4][1]/P0001  , \wishbone_bd_ram_mem0_reg[4][2]/P0001  , \wishbone_bd_ram_mem0_reg[4][3]/P0001  , \wishbone_bd_ram_mem0_reg[4][4]/P0001  , \wishbone_bd_ram_mem0_reg[4][5]/P0001  , \wishbone_bd_ram_mem0_reg[4][6]/P0001  , \wishbone_bd_ram_mem0_reg[4][7]/P0001  , \wishbone_bd_ram_mem0_reg[50][0]/P0001  , \wishbone_bd_ram_mem0_reg[50][1]/P0001  , \wishbone_bd_ram_mem0_reg[50][2]/P0001  , \wishbone_bd_ram_mem0_reg[50][3]/P0001  , \wishbone_bd_ram_mem0_reg[50][4]/P0001  , \wishbone_bd_ram_mem0_reg[50][5]/P0001  , \wishbone_bd_ram_mem0_reg[50][6]/P0001  , \wishbone_bd_ram_mem0_reg[50][7]/P0001  , \wishbone_bd_ram_mem0_reg[51][0]/P0001  , \wishbone_bd_ram_mem0_reg[51][1]/P0001  , \wishbone_bd_ram_mem0_reg[51][2]/P0001  , \wishbone_bd_ram_mem0_reg[51][3]/P0001  , \wishbone_bd_ram_mem0_reg[51][4]/P0001  , \wishbone_bd_ram_mem0_reg[51][5]/P0001  , \wishbone_bd_ram_mem0_reg[51][6]/P0001  , \wishbone_bd_ram_mem0_reg[51][7]/P0001  , \wishbone_bd_ram_mem0_reg[52][0]/P0001  , \wishbone_bd_ram_mem0_reg[52][1]/P0001  , \wishbone_bd_ram_mem0_reg[52][2]/P0001  , \wishbone_bd_ram_mem0_reg[52][3]/P0001  , \wishbone_bd_ram_mem0_reg[52][4]/P0001  , \wishbone_bd_ram_mem0_reg[52][5]/P0001  , \wishbone_bd_ram_mem0_reg[52][6]/P0001  , \wishbone_bd_ram_mem0_reg[52][7]/P0001  , \wishbone_bd_ram_mem0_reg[53][0]/P0001  , \wishbone_bd_ram_mem0_reg[53][1]/P0001  , \wishbone_bd_ram_mem0_reg[53][2]/P0001  , \wishbone_bd_ram_mem0_reg[53][3]/P0001  , \wishbone_bd_ram_mem0_reg[53][4]/P0001  , \wishbone_bd_ram_mem0_reg[53][5]/P0001  , \wishbone_bd_ram_mem0_reg[53][6]/P0001  , \wishbone_bd_ram_mem0_reg[53][7]/P0001  , \wishbone_bd_ram_mem0_reg[54][0]/P0001  , \wishbone_bd_ram_mem0_reg[54][1]/P0001  , \wishbone_bd_ram_mem0_reg[54][2]/P0001  , \wishbone_bd_ram_mem0_reg[54][3]/P0001  , \wishbone_bd_ram_mem0_reg[54][4]/P0001  , \wishbone_bd_ram_mem0_reg[54][5]/P0001  , \wishbone_bd_ram_mem0_reg[54][6]/P0001  , \wishbone_bd_ram_mem0_reg[54][7]/P0001  , \wishbone_bd_ram_mem0_reg[55][0]/P0001  , \wishbone_bd_ram_mem0_reg[55][1]/P0001  , \wishbone_bd_ram_mem0_reg[55][2]/P0001  , \wishbone_bd_ram_mem0_reg[55][3]/P0001  , \wishbone_bd_ram_mem0_reg[55][4]/P0001  , \wishbone_bd_ram_mem0_reg[55][5]/P0001  , \wishbone_bd_ram_mem0_reg[55][6]/P0001  , \wishbone_bd_ram_mem0_reg[55][7]/P0001  , \wishbone_bd_ram_mem0_reg[56][0]/P0001  , \wishbone_bd_ram_mem0_reg[56][1]/P0001  , \wishbone_bd_ram_mem0_reg[56][2]/P0001  , \wishbone_bd_ram_mem0_reg[56][3]/P0001  , \wishbone_bd_ram_mem0_reg[56][4]/P0001  , \wishbone_bd_ram_mem0_reg[56][5]/P0001  , \wishbone_bd_ram_mem0_reg[56][6]/P0001  , \wishbone_bd_ram_mem0_reg[56][7]/P0001  , \wishbone_bd_ram_mem0_reg[57][0]/P0001  , \wishbone_bd_ram_mem0_reg[57][1]/P0001  , \wishbone_bd_ram_mem0_reg[57][2]/P0001  , \wishbone_bd_ram_mem0_reg[57][3]/P0001  , \wishbone_bd_ram_mem0_reg[57][4]/P0001  , \wishbone_bd_ram_mem0_reg[57][5]/P0001  , \wishbone_bd_ram_mem0_reg[57][6]/P0001  , \wishbone_bd_ram_mem0_reg[57][7]/P0001  , \wishbone_bd_ram_mem0_reg[58][0]/P0001  , \wishbone_bd_ram_mem0_reg[58][1]/P0001  , \wishbone_bd_ram_mem0_reg[58][2]/P0001  , \wishbone_bd_ram_mem0_reg[58][3]/P0001  , \wishbone_bd_ram_mem0_reg[58][4]/P0001  , \wishbone_bd_ram_mem0_reg[58][5]/P0001  , \wishbone_bd_ram_mem0_reg[58][6]/P0001  , \wishbone_bd_ram_mem0_reg[58][7]/P0001  , \wishbone_bd_ram_mem0_reg[59][0]/P0001  , \wishbone_bd_ram_mem0_reg[59][1]/P0001  , \wishbone_bd_ram_mem0_reg[59][2]/P0001  , \wishbone_bd_ram_mem0_reg[59][3]/P0001  , \wishbone_bd_ram_mem0_reg[59][4]/P0001  , \wishbone_bd_ram_mem0_reg[59][5]/P0001  , \wishbone_bd_ram_mem0_reg[59][6]/P0001  , \wishbone_bd_ram_mem0_reg[59][7]/P0001  , \wishbone_bd_ram_mem0_reg[5][0]/P0001  , \wishbone_bd_ram_mem0_reg[5][1]/P0001  , \wishbone_bd_ram_mem0_reg[5][2]/P0001  , \wishbone_bd_ram_mem0_reg[5][3]/P0001  , \wishbone_bd_ram_mem0_reg[5][4]/P0001  , \wishbone_bd_ram_mem0_reg[5][5]/P0001  , \wishbone_bd_ram_mem0_reg[5][6]/P0001  , \wishbone_bd_ram_mem0_reg[5][7]/P0001  , \wishbone_bd_ram_mem0_reg[60][0]/P0001  , \wishbone_bd_ram_mem0_reg[60][1]/P0001  , \wishbone_bd_ram_mem0_reg[60][2]/P0001  , \wishbone_bd_ram_mem0_reg[60][3]/P0001  , \wishbone_bd_ram_mem0_reg[60][4]/P0001  , \wishbone_bd_ram_mem0_reg[60][5]/P0001  , \wishbone_bd_ram_mem0_reg[60][6]/P0001  , \wishbone_bd_ram_mem0_reg[60][7]/P0001  , \wishbone_bd_ram_mem0_reg[61][0]/P0001  , \wishbone_bd_ram_mem0_reg[61][1]/P0001  , \wishbone_bd_ram_mem0_reg[61][2]/P0001  , \wishbone_bd_ram_mem0_reg[61][3]/P0001  , \wishbone_bd_ram_mem0_reg[61][4]/P0001  , \wishbone_bd_ram_mem0_reg[61][5]/P0001  , \wishbone_bd_ram_mem0_reg[61][6]/P0001  , \wishbone_bd_ram_mem0_reg[61][7]/P0001  , \wishbone_bd_ram_mem0_reg[62][0]/P0001  , \wishbone_bd_ram_mem0_reg[62][1]/P0001  , \wishbone_bd_ram_mem0_reg[62][2]/P0001  , \wishbone_bd_ram_mem0_reg[62][3]/P0001  , \wishbone_bd_ram_mem0_reg[62][4]/P0001  , \wishbone_bd_ram_mem0_reg[62][5]/P0001  , \wishbone_bd_ram_mem0_reg[62][6]/P0001  , \wishbone_bd_ram_mem0_reg[62][7]/P0001  , \wishbone_bd_ram_mem0_reg[63][0]/P0001  , \wishbone_bd_ram_mem0_reg[63][1]/P0001  , \wishbone_bd_ram_mem0_reg[63][2]/P0001  , \wishbone_bd_ram_mem0_reg[63][3]/P0001  , \wishbone_bd_ram_mem0_reg[63][4]/P0001  , \wishbone_bd_ram_mem0_reg[63][5]/P0001  , \wishbone_bd_ram_mem0_reg[63][6]/P0001  , \wishbone_bd_ram_mem0_reg[63][7]/P0001  , \wishbone_bd_ram_mem0_reg[64][0]/P0001  , \wishbone_bd_ram_mem0_reg[64][1]/P0001  , \wishbone_bd_ram_mem0_reg[64][2]/P0001  , \wishbone_bd_ram_mem0_reg[64][3]/P0001  , \wishbone_bd_ram_mem0_reg[64][4]/P0001  , \wishbone_bd_ram_mem0_reg[64][5]/P0001  , \wishbone_bd_ram_mem0_reg[64][6]/P0001  , \wishbone_bd_ram_mem0_reg[64][7]/P0001  , \wishbone_bd_ram_mem0_reg[65][0]/P0001  , \wishbone_bd_ram_mem0_reg[65][1]/P0001  , \wishbone_bd_ram_mem0_reg[65][2]/P0001  , \wishbone_bd_ram_mem0_reg[65][3]/P0001  , \wishbone_bd_ram_mem0_reg[65][4]/P0001  , \wishbone_bd_ram_mem0_reg[65][5]/P0001  , \wishbone_bd_ram_mem0_reg[65][6]/P0001  , \wishbone_bd_ram_mem0_reg[65][7]/P0001  , \wishbone_bd_ram_mem0_reg[66][0]/P0001  , \wishbone_bd_ram_mem0_reg[66][1]/P0001  , \wishbone_bd_ram_mem0_reg[66][2]/P0001  , \wishbone_bd_ram_mem0_reg[66][3]/P0001  , \wishbone_bd_ram_mem0_reg[66][4]/P0001  , \wishbone_bd_ram_mem0_reg[66][5]/P0001  , \wishbone_bd_ram_mem0_reg[66][6]/P0001  , \wishbone_bd_ram_mem0_reg[66][7]/P0001  , \wishbone_bd_ram_mem0_reg[67][0]/P0001  , \wishbone_bd_ram_mem0_reg[67][1]/P0001  , \wishbone_bd_ram_mem0_reg[67][2]/P0001  , \wishbone_bd_ram_mem0_reg[67][3]/P0001  , \wishbone_bd_ram_mem0_reg[67][4]/P0001  , \wishbone_bd_ram_mem0_reg[67][5]/P0001  , \wishbone_bd_ram_mem0_reg[67][6]/P0001  , \wishbone_bd_ram_mem0_reg[67][7]/P0001  , \wishbone_bd_ram_mem0_reg[68][0]/P0001  , \wishbone_bd_ram_mem0_reg[68][1]/P0001  , \wishbone_bd_ram_mem0_reg[68][2]/P0001  , \wishbone_bd_ram_mem0_reg[68][3]/P0001  , \wishbone_bd_ram_mem0_reg[68][4]/P0001  , \wishbone_bd_ram_mem0_reg[68][5]/P0001  , \wishbone_bd_ram_mem0_reg[68][6]/P0001  , \wishbone_bd_ram_mem0_reg[68][7]/P0001  , \wishbone_bd_ram_mem0_reg[69][0]/P0001  , \wishbone_bd_ram_mem0_reg[69][1]/P0001  , \wishbone_bd_ram_mem0_reg[69][2]/P0001  , \wishbone_bd_ram_mem0_reg[69][3]/P0001  , \wishbone_bd_ram_mem0_reg[69][4]/P0001  , \wishbone_bd_ram_mem0_reg[69][5]/P0001  , \wishbone_bd_ram_mem0_reg[69][6]/P0001  , \wishbone_bd_ram_mem0_reg[69][7]/P0001  , \wishbone_bd_ram_mem0_reg[6][0]/P0001  , \wishbone_bd_ram_mem0_reg[6][1]/P0001  , \wishbone_bd_ram_mem0_reg[6][2]/P0001  , \wishbone_bd_ram_mem0_reg[6][3]/P0001  , \wishbone_bd_ram_mem0_reg[6][4]/P0001  , \wishbone_bd_ram_mem0_reg[6][5]/P0001  , \wishbone_bd_ram_mem0_reg[6][6]/P0001  , \wishbone_bd_ram_mem0_reg[6][7]/P0001  , \wishbone_bd_ram_mem0_reg[70][0]/P0001  , \wishbone_bd_ram_mem0_reg[70][1]/P0001  , \wishbone_bd_ram_mem0_reg[70][2]/P0001  , \wishbone_bd_ram_mem0_reg[70][3]/P0001  , \wishbone_bd_ram_mem0_reg[70][4]/P0001  , \wishbone_bd_ram_mem0_reg[70][5]/P0001  , \wishbone_bd_ram_mem0_reg[70][6]/P0001  , \wishbone_bd_ram_mem0_reg[70][7]/P0001  , \wishbone_bd_ram_mem0_reg[71][0]/P0001  , \wishbone_bd_ram_mem0_reg[71][1]/P0001  , \wishbone_bd_ram_mem0_reg[71][2]/P0001  , \wishbone_bd_ram_mem0_reg[71][3]/P0001  , \wishbone_bd_ram_mem0_reg[71][4]/P0001  , \wishbone_bd_ram_mem0_reg[71][5]/P0001  , \wishbone_bd_ram_mem0_reg[71][6]/P0001  , \wishbone_bd_ram_mem0_reg[71][7]/P0001  , \wishbone_bd_ram_mem0_reg[72][0]/P0001  , \wishbone_bd_ram_mem0_reg[72][1]/P0001  , \wishbone_bd_ram_mem0_reg[72][2]/P0001  , \wishbone_bd_ram_mem0_reg[72][3]/P0001  , \wishbone_bd_ram_mem0_reg[72][4]/P0001  , \wishbone_bd_ram_mem0_reg[72][5]/P0001  , \wishbone_bd_ram_mem0_reg[72][6]/P0001  , \wishbone_bd_ram_mem0_reg[72][7]/P0001  , \wishbone_bd_ram_mem0_reg[73][0]/P0001  , \wishbone_bd_ram_mem0_reg[73][1]/P0001  , \wishbone_bd_ram_mem0_reg[73][2]/P0001  , \wishbone_bd_ram_mem0_reg[73][3]/P0001  , \wishbone_bd_ram_mem0_reg[73][4]/P0001  , \wishbone_bd_ram_mem0_reg[73][5]/P0001  , \wishbone_bd_ram_mem0_reg[73][6]/P0001  , \wishbone_bd_ram_mem0_reg[73][7]/P0001  , \wishbone_bd_ram_mem0_reg[74][0]/P0001  , \wishbone_bd_ram_mem0_reg[74][1]/P0001  , \wishbone_bd_ram_mem0_reg[74][2]/P0001  , \wishbone_bd_ram_mem0_reg[74][3]/P0001  , \wishbone_bd_ram_mem0_reg[74][4]/P0001  , \wishbone_bd_ram_mem0_reg[74][5]/P0001  , \wishbone_bd_ram_mem0_reg[74][6]/P0001  , \wishbone_bd_ram_mem0_reg[74][7]/P0001  , \wishbone_bd_ram_mem0_reg[75][0]/P0001  , \wishbone_bd_ram_mem0_reg[75][1]/P0001  , \wishbone_bd_ram_mem0_reg[75][2]/P0001  , \wishbone_bd_ram_mem0_reg[75][3]/P0001  , \wishbone_bd_ram_mem0_reg[75][4]/P0001  , \wishbone_bd_ram_mem0_reg[75][5]/P0001  , \wishbone_bd_ram_mem0_reg[75][6]/P0001  , \wishbone_bd_ram_mem0_reg[75][7]/P0001  , \wishbone_bd_ram_mem0_reg[76][0]/P0001  , \wishbone_bd_ram_mem0_reg[76][1]/P0001  , \wishbone_bd_ram_mem0_reg[76][2]/P0001  , \wishbone_bd_ram_mem0_reg[76][3]/P0001  , \wishbone_bd_ram_mem0_reg[76][4]/P0001  , \wishbone_bd_ram_mem0_reg[76][5]/P0001  , \wishbone_bd_ram_mem0_reg[76][6]/P0001  , \wishbone_bd_ram_mem0_reg[76][7]/P0001  , \wishbone_bd_ram_mem0_reg[77][0]/P0001  , \wishbone_bd_ram_mem0_reg[77][1]/P0001  , \wishbone_bd_ram_mem0_reg[77][2]/P0001  , \wishbone_bd_ram_mem0_reg[77][3]/P0001  , \wishbone_bd_ram_mem0_reg[77][4]/P0001  , \wishbone_bd_ram_mem0_reg[77][5]/P0001  , \wishbone_bd_ram_mem0_reg[77][6]/P0001  , \wishbone_bd_ram_mem0_reg[77][7]/P0001  , \wishbone_bd_ram_mem0_reg[78][0]/P0001  , \wishbone_bd_ram_mem0_reg[78][1]/P0001  , \wishbone_bd_ram_mem0_reg[78][2]/P0001  , \wishbone_bd_ram_mem0_reg[78][3]/P0001  , \wishbone_bd_ram_mem0_reg[78][4]/P0001  , \wishbone_bd_ram_mem0_reg[78][5]/P0001  , \wishbone_bd_ram_mem0_reg[78][6]/P0001  , \wishbone_bd_ram_mem0_reg[78][7]/P0001  , \wishbone_bd_ram_mem0_reg[79][0]/P0001  , \wishbone_bd_ram_mem0_reg[79][1]/P0001  , \wishbone_bd_ram_mem0_reg[79][2]/P0001  , \wishbone_bd_ram_mem0_reg[79][3]/P0001  , \wishbone_bd_ram_mem0_reg[79][4]/P0001  , \wishbone_bd_ram_mem0_reg[79][5]/P0001  , \wishbone_bd_ram_mem0_reg[79][6]/P0001  , \wishbone_bd_ram_mem0_reg[79][7]/P0001  , \wishbone_bd_ram_mem0_reg[7][0]/P0001  , \wishbone_bd_ram_mem0_reg[7][1]/P0001  , \wishbone_bd_ram_mem0_reg[7][2]/P0001  , \wishbone_bd_ram_mem0_reg[7][3]/P0001  , \wishbone_bd_ram_mem0_reg[7][4]/P0001  , \wishbone_bd_ram_mem0_reg[7][5]/P0001  , \wishbone_bd_ram_mem0_reg[7][6]/P0001  , \wishbone_bd_ram_mem0_reg[7][7]/P0001  , \wishbone_bd_ram_mem0_reg[80][0]/P0001  , \wishbone_bd_ram_mem0_reg[80][1]/P0001  , \wishbone_bd_ram_mem0_reg[80][2]/P0001  , \wishbone_bd_ram_mem0_reg[80][3]/P0001  , \wishbone_bd_ram_mem0_reg[80][4]/P0001  , \wishbone_bd_ram_mem0_reg[80][5]/P0001  , \wishbone_bd_ram_mem0_reg[80][6]/P0001  , \wishbone_bd_ram_mem0_reg[80][7]/P0001  , \wishbone_bd_ram_mem0_reg[81][0]/P0001  , \wishbone_bd_ram_mem0_reg[81][1]/P0001  , \wishbone_bd_ram_mem0_reg[81][2]/P0001  , \wishbone_bd_ram_mem0_reg[81][3]/P0001  , \wishbone_bd_ram_mem0_reg[81][4]/P0001  , \wishbone_bd_ram_mem0_reg[81][5]/P0001  , \wishbone_bd_ram_mem0_reg[81][6]/P0001  , \wishbone_bd_ram_mem0_reg[81][7]/P0001  , \wishbone_bd_ram_mem0_reg[82][0]/P0001  , \wishbone_bd_ram_mem0_reg[82][1]/P0001  , \wishbone_bd_ram_mem0_reg[82][2]/P0001  , \wishbone_bd_ram_mem0_reg[82][3]/P0001  , \wishbone_bd_ram_mem0_reg[82][4]/P0001  , \wishbone_bd_ram_mem0_reg[82][5]/P0001  , \wishbone_bd_ram_mem0_reg[82][6]/P0001  , \wishbone_bd_ram_mem0_reg[82][7]/P0001  , \wishbone_bd_ram_mem0_reg[83][0]/P0001  , \wishbone_bd_ram_mem0_reg[83][1]/P0001  , \wishbone_bd_ram_mem0_reg[83][2]/P0001  , \wishbone_bd_ram_mem0_reg[83][3]/P0001  , \wishbone_bd_ram_mem0_reg[83][4]/P0001  , \wishbone_bd_ram_mem0_reg[83][5]/P0001  , \wishbone_bd_ram_mem0_reg[83][6]/P0001  , \wishbone_bd_ram_mem0_reg[83][7]/P0001  , \wishbone_bd_ram_mem0_reg[84][0]/P0001  , \wishbone_bd_ram_mem0_reg[84][1]/P0001  , \wishbone_bd_ram_mem0_reg[84][2]/P0001  , \wishbone_bd_ram_mem0_reg[84][3]/P0001  , \wishbone_bd_ram_mem0_reg[84][4]/P0001  , \wishbone_bd_ram_mem0_reg[84][5]/P0001  , \wishbone_bd_ram_mem0_reg[84][6]/P0001  , \wishbone_bd_ram_mem0_reg[84][7]/P0001  , \wishbone_bd_ram_mem0_reg[85][0]/P0001  , \wishbone_bd_ram_mem0_reg[85][1]/P0001  , \wishbone_bd_ram_mem0_reg[85][2]/P0001  , \wishbone_bd_ram_mem0_reg[85][3]/P0001  , \wishbone_bd_ram_mem0_reg[85][4]/P0001  , \wishbone_bd_ram_mem0_reg[85][5]/P0001  , \wishbone_bd_ram_mem0_reg[85][6]/P0001  , \wishbone_bd_ram_mem0_reg[85][7]/P0001  , \wishbone_bd_ram_mem0_reg[86][0]/P0001  , \wishbone_bd_ram_mem0_reg[86][1]/P0001  , \wishbone_bd_ram_mem0_reg[86][2]/P0001  , \wishbone_bd_ram_mem0_reg[86][3]/P0001  , \wishbone_bd_ram_mem0_reg[86][4]/P0001  , \wishbone_bd_ram_mem0_reg[86][5]/P0001  , \wishbone_bd_ram_mem0_reg[86][6]/P0001  , \wishbone_bd_ram_mem0_reg[86][7]/P0001  , \wishbone_bd_ram_mem0_reg[87][0]/P0001  , \wishbone_bd_ram_mem0_reg[87][1]/P0001  , \wishbone_bd_ram_mem0_reg[87][2]/P0001  , \wishbone_bd_ram_mem0_reg[87][3]/P0001  , \wishbone_bd_ram_mem0_reg[87][4]/P0001  , \wishbone_bd_ram_mem0_reg[87][5]/P0001  , \wishbone_bd_ram_mem0_reg[87][6]/P0001  , \wishbone_bd_ram_mem0_reg[87][7]/P0001  , \wishbone_bd_ram_mem0_reg[88][0]/P0001  , \wishbone_bd_ram_mem0_reg[88][1]/P0001  , \wishbone_bd_ram_mem0_reg[88][2]/P0001  , \wishbone_bd_ram_mem0_reg[88][3]/P0001  , \wishbone_bd_ram_mem0_reg[88][4]/P0001  , \wishbone_bd_ram_mem0_reg[88][5]/P0001  , \wishbone_bd_ram_mem0_reg[88][6]/P0001  , \wishbone_bd_ram_mem0_reg[88][7]/P0001  , \wishbone_bd_ram_mem0_reg[89][0]/P0001  , \wishbone_bd_ram_mem0_reg[89][1]/P0001  , \wishbone_bd_ram_mem0_reg[89][2]/P0001  , \wishbone_bd_ram_mem0_reg[89][3]/P0001  , \wishbone_bd_ram_mem0_reg[89][4]/P0001  , \wishbone_bd_ram_mem0_reg[89][5]/P0001  , \wishbone_bd_ram_mem0_reg[89][6]/P0001  , \wishbone_bd_ram_mem0_reg[89][7]/P0001  , \wishbone_bd_ram_mem0_reg[8][0]/P0001  , \wishbone_bd_ram_mem0_reg[8][1]/P0001  , \wishbone_bd_ram_mem0_reg[8][2]/P0001  , \wishbone_bd_ram_mem0_reg[8][3]/P0001  , \wishbone_bd_ram_mem0_reg[8][4]/P0001  , \wishbone_bd_ram_mem0_reg[8][5]/P0001  , \wishbone_bd_ram_mem0_reg[8][6]/P0001  , \wishbone_bd_ram_mem0_reg[8][7]/P0001  , \wishbone_bd_ram_mem0_reg[90][0]/P0001  , \wishbone_bd_ram_mem0_reg[90][1]/P0001  , \wishbone_bd_ram_mem0_reg[90][2]/P0001  , \wishbone_bd_ram_mem0_reg[90][3]/P0001  , \wishbone_bd_ram_mem0_reg[90][4]/P0001  , \wishbone_bd_ram_mem0_reg[90][5]/P0001  , \wishbone_bd_ram_mem0_reg[90][6]/P0001  , \wishbone_bd_ram_mem0_reg[90][7]/P0001  , \wishbone_bd_ram_mem0_reg[91][0]/P0001  , \wishbone_bd_ram_mem0_reg[91][1]/P0001  , \wishbone_bd_ram_mem0_reg[91][2]/P0001  , \wishbone_bd_ram_mem0_reg[91][3]/P0001  , \wishbone_bd_ram_mem0_reg[91][4]/P0001  , \wishbone_bd_ram_mem0_reg[91][5]/P0001  , \wishbone_bd_ram_mem0_reg[91][6]/P0001  , \wishbone_bd_ram_mem0_reg[91][7]/P0001  , \wishbone_bd_ram_mem0_reg[92][0]/P0001  , \wishbone_bd_ram_mem0_reg[92][1]/P0001  , \wishbone_bd_ram_mem0_reg[92][2]/P0001  , \wishbone_bd_ram_mem0_reg[92][3]/P0001  , \wishbone_bd_ram_mem0_reg[92][4]/P0001  , \wishbone_bd_ram_mem0_reg[92][5]/P0001  , \wishbone_bd_ram_mem0_reg[92][6]/P0001  , \wishbone_bd_ram_mem0_reg[92][7]/P0001  , \wishbone_bd_ram_mem0_reg[93][0]/P0001  , \wishbone_bd_ram_mem0_reg[93][1]/P0001  , \wishbone_bd_ram_mem0_reg[93][2]/P0001  , \wishbone_bd_ram_mem0_reg[93][3]/P0001  , \wishbone_bd_ram_mem0_reg[93][4]/P0001  , \wishbone_bd_ram_mem0_reg[93][5]/P0001  , \wishbone_bd_ram_mem0_reg[93][6]/P0001  , \wishbone_bd_ram_mem0_reg[93][7]/P0001  , \wishbone_bd_ram_mem0_reg[94][0]/P0001  , \wishbone_bd_ram_mem0_reg[94][1]/P0001  , \wishbone_bd_ram_mem0_reg[94][2]/P0001  , \wishbone_bd_ram_mem0_reg[94][3]/P0001  , \wishbone_bd_ram_mem0_reg[94][4]/P0001  , \wishbone_bd_ram_mem0_reg[94][5]/P0001  , \wishbone_bd_ram_mem0_reg[94][6]/P0001  , \wishbone_bd_ram_mem0_reg[94][7]/P0001  , \wishbone_bd_ram_mem0_reg[95][0]/P0001  , \wishbone_bd_ram_mem0_reg[95][1]/P0001  , \wishbone_bd_ram_mem0_reg[95][2]/P0001  , \wishbone_bd_ram_mem0_reg[95][3]/P0001  , \wishbone_bd_ram_mem0_reg[95][4]/P0001  , \wishbone_bd_ram_mem0_reg[95][5]/P0001  , \wishbone_bd_ram_mem0_reg[95][6]/P0001  , \wishbone_bd_ram_mem0_reg[95][7]/P0001  , \wishbone_bd_ram_mem0_reg[96][0]/P0001  , \wishbone_bd_ram_mem0_reg[96][1]/P0001  , \wishbone_bd_ram_mem0_reg[96][2]/P0001  , \wishbone_bd_ram_mem0_reg[96][3]/P0001  , \wishbone_bd_ram_mem0_reg[96][4]/P0001  , \wishbone_bd_ram_mem0_reg[96][5]/P0001  , \wishbone_bd_ram_mem0_reg[96][6]/P0001  , \wishbone_bd_ram_mem0_reg[96][7]/P0001  , \wishbone_bd_ram_mem0_reg[97][0]/P0001  , \wishbone_bd_ram_mem0_reg[97][1]/P0001  , \wishbone_bd_ram_mem0_reg[97][2]/P0001  , \wishbone_bd_ram_mem0_reg[97][3]/P0001  , \wishbone_bd_ram_mem0_reg[97][4]/P0001  , \wishbone_bd_ram_mem0_reg[97][5]/P0001  , \wishbone_bd_ram_mem0_reg[97][6]/P0001  , \wishbone_bd_ram_mem0_reg[97][7]/P0001  , \wishbone_bd_ram_mem0_reg[98][0]/P0001  , \wishbone_bd_ram_mem0_reg[98][1]/P0001  , \wishbone_bd_ram_mem0_reg[98][2]/P0001  , \wishbone_bd_ram_mem0_reg[98][3]/P0001  , \wishbone_bd_ram_mem0_reg[98][4]/P0001  , \wishbone_bd_ram_mem0_reg[98][5]/P0001  , \wishbone_bd_ram_mem0_reg[98][6]/P0001  , \wishbone_bd_ram_mem0_reg[98][7]/P0001  , \wishbone_bd_ram_mem0_reg[99][0]/P0001  , \wishbone_bd_ram_mem0_reg[99][1]/P0001  , \wishbone_bd_ram_mem0_reg[99][2]/P0001  , \wishbone_bd_ram_mem0_reg[99][3]/P0001  , \wishbone_bd_ram_mem0_reg[99][4]/P0001  , \wishbone_bd_ram_mem0_reg[99][5]/P0001  , \wishbone_bd_ram_mem0_reg[99][6]/P0001  , \wishbone_bd_ram_mem0_reg[99][7]/P0001  , \wishbone_bd_ram_mem0_reg[9][0]/P0001  , \wishbone_bd_ram_mem0_reg[9][1]/P0001  , \wishbone_bd_ram_mem0_reg[9][2]/P0001  , \wishbone_bd_ram_mem0_reg[9][3]/P0001  , \wishbone_bd_ram_mem0_reg[9][4]/P0001  , \wishbone_bd_ram_mem0_reg[9][5]/P0001  , \wishbone_bd_ram_mem0_reg[9][6]/P0001  , \wishbone_bd_ram_mem0_reg[9][7]/P0001  , \wishbone_bd_ram_mem1_reg[0][10]/P0001  , \wishbone_bd_ram_mem1_reg[0][11]/P0001  , \wishbone_bd_ram_mem1_reg[0][12]/P0001  , \wishbone_bd_ram_mem1_reg[0][13]/P0001  , \wishbone_bd_ram_mem1_reg[0][14]/P0001  , \wishbone_bd_ram_mem1_reg[0][15]/P0001  , \wishbone_bd_ram_mem1_reg[0][8]/P0001  , \wishbone_bd_ram_mem1_reg[0][9]/P0001  , \wishbone_bd_ram_mem1_reg[100][10]/P0001  , \wishbone_bd_ram_mem1_reg[100][11]/P0001  , \wishbone_bd_ram_mem1_reg[100][12]/P0001  , \wishbone_bd_ram_mem1_reg[100][13]/P0001  , \wishbone_bd_ram_mem1_reg[100][14]/P0001  , \wishbone_bd_ram_mem1_reg[100][15]/P0001  , \wishbone_bd_ram_mem1_reg[100][8]/P0001  , \wishbone_bd_ram_mem1_reg[100][9]/P0001  , \wishbone_bd_ram_mem1_reg[101][10]/P0001  , \wishbone_bd_ram_mem1_reg[101][11]/P0001  , \wishbone_bd_ram_mem1_reg[101][12]/P0001  , \wishbone_bd_ram_mem1_reg[101][13]/P0001  , \wishbone_bd_ram_mem1_reg[101][14]/P0001  , \wishbone_bd_ram_mem1_reg[101][15]/P0001  , \wishbone_bd_ram_mem1_reg[101][8]/P0001  , \wishbone_bd_ram_mem1_reg[101][9]/P0001  , \wishbone_bd_ram_mem1_reg[102][10]/P0001  , \wishbone_bd_ram_mem1_reg[102][11]/P0001  , \wishbone_bd_ram_mem1_reg[102][12]/P0001  , \wishbone_bd_ram_mem1_reg[102][13]/P0001  , \wishbone_bd_ram_mem1_reg[102][14]/P0001  , \wishbone_bd_ram_mem1_reg[102][15]/P0001  , \wishbone_bd_ram_mem1_reg[102][8]/P0001  , \wishbone_bd_ram_mem1_reg[102][9]/P0001  , \wishbone_bd_ram_mem1_reg[103][10]/P0001  , \wishbone_bd_ram_mem1_reg[103][11]/P0001  , \wishbone_bd_ram_mem1_reg[103][12]/P0001  , \wishbone_bd_ram_mem1_reg[103][13]/P0001  , \wishbone_bd_ram_mem1_reg[103][14]/P0001  , \wishbone_bd_ram_mem1_reg[103][15]/P0001  , \wishbone_bd_ram_mem1_reg[103][8]/P0001  , \wishbone_bd_ram_mem1_reg[103][9]/P0001  , \wishbone_bd_ram_mem1_reg[104][10]/P0001  , \wishbone_bd_ram_mem1_reg[104][11]/P0001  , \wishbone_bd_ram_mem1_reg[104][12]/P0001  , \wishbone_bd_ram_mem1_reg[104][13]/P0001  , \wishbone_bd_ram_mem1_reg[104][14]/P0001  , \wishbone_bd_ram_mem1_reg[104][15]/P0001  , \wishbone_bd_ram_mem1_reg[104][8]/P0001  , \wishbone_bd_ram_mem1_reg[104][9]/P0001  , \wishbone_bd_ram_mem1_reg[105][10]/P0001  , \wishbone_bd_ram_mem1_reg[105][11]/P0001  , \wishbone_bd_ram_mem1_reg[105][12]/P0001  , \wishbone_bd_ram_mem1_reg[105][13]/P0001  , \wishbone_bd_ram_mem1_reg[105][14]/P0001  , \wishbone_bd_ram_mem1_reg[105][15]/P0001  , \wishbone_bd_ram_mem1_reg[105][8]/P0001  , \wishbone_bd_ram_mem1_reg[105][9]/P0001  , \wishbone_bd_ram_mem1_reg[106][10]/P0001  , \wishbone_bd_ram_mem1_reg[106][11]/P0001  , \wishbone_bd_ram_mem1_reg[106][12]/P0001  , \wishbone_bd_ram_mem1_reg[106][13]/P0001  , \wishbone_bd_ram_mem1_reg[106][14]/P0001  , \wishbone_bd_ram_mem1_reg[106][15]/P0001  , \wishbone_bd_ram_mem1_reg[106][8]/P0001  , \wishbone_bd_ram_mem1_reg[106][9]/P0001  , \wishbone_bd_ram_mem1_reg[107][10]/P0001  , \wishbone_bd_ram_mem1_reg[107][11]/P0001  , \wishbone_bd_ram_mem1_reg[107][12]/P0001  , \wishbone_bd_ram_mem1_reg[107][13]/P0001  , \wishbone_bd_ram_mem1_reg[107][14]/P0001  , \wishbone_bd_ram_mem1_reg[107][15]/P0001  , \wishbone_bd_ram_mem1_reg[107][8]/P0001  , \wishbone_bd_ram_mem1_reg[107][9]/P0001  , \wishbone_bd_ram_mem1_reg[108][10]/P0001  , \wishbone_bd_ram_mem1_reg[108][11]/P0001  , \wishbone_bd_ram_mem1_reg[108][12]/P0001  , \wishbone_bd_ram_mem1_reg[108][13]/P0001  , \wishbone_bd_ram_mem1_reg[108][14]/P0001  , \wishbone_bd_ram_mem1_reg[108][15]/P0001  , \wishbone_bd_ram_mem1_reg[108][8]/P0001  , \wishbone_bd_ram_mem1_reg[108][9]/P0001  , \wishbone_bd_ram_mem1_reg[109][10]/P0001  , \wishbone_bd_ram_mem1_reg[109][11]/P0001  , \wishbone_bd_ram_mem1_reg[109][12]/P0001  , \wishbone_bd_ram_mem1_reg[109][13]/P0001  , \wishbone_bd_ram_mem1_reg[109][14]/P0001  , \wishbone_bd_ram_mem1_reg[109][15]/P0001  , \wishbone_bd_ram_mem1_reg[109][8]/P0001  , \wishbone_bd_ram_mem1_reg[109][9]/P0001  , \wishbone_bd_ram_mem1_reg[10][10]/P0001  , \wishbone_bd_ram_mem1_reg[10][11]/P0001  , \wishbone_bd_ram_mem1_reg[10][12]/P0001  , \wishbone_bd_ram_mem1_reg[10][13]/P0001  , \wishbone_bd_ram_mem1_reg[10][14]/P0001  , \wishbone_bd_ram_mem1_reg[10][15]/P0001  , \wishbone_bd_ram_mem1_reg[10][8]/P0001  , \wishbone_bd_ram_mem1_reg[10][9]/P0001  , \wishbone_bd_ram_mem1_reg[110][10]/P0001  , \wishbone_bd_ram_mem1_reg[110][11]/P0001  , \wishbone_bd_ram_mem1_reg[110][12]/P0001  , \wishbone_bd_ram_mem1_reg[110][13]/P0001  , \wishbone_bd_ram_mem1_reg[110][14]/P0001  , \wishbone_bd_ram_mem1_reg[110][15]/P0001  , \wishbone_bd_ram_mem1_reg[110][8]/P0001  , \wishbone_bd_ram_mem1_reg[110][9]/P0001  , \wishbone_bd_ram_mem1_reg[111][10]/P0001  , \wishbone_bd_ram_mem1_reg[111][11]/P0001  , \wishbone_bd_ram_mem1_reg[111][12]/P0001  , \wishbone_bd_ram_mem1_reg[111][13]/P0001  , \wishbone_bd_ram_mem1_reg[111][14]/P0001  , \wishbone_bd_ram_mem1_reg[111][15]/P0001  , \wishbone_bd_ram_mem1_reg[111][8]/P0001  , \wishbone_bd_ram_mem1_reg[111][9]/P0001  , \wishbone_bd_ram_mem1_reg[112][10]/P0001  , \wishbone_bd_ram_mem1_reg[112][11]/P0001  , \wishbone_bd_ram_mem1_reg[112][12]/P0001  , \wishbone_bd_ram_mem1_reg[112][13]/P0001  , \wishbone_bd_ram_mem1_reg[112][14]/P0001  , \wishbone_bd_ram_mem1_reg[112][15]/P0001  , \wishbone_bd_ram_mem1_reg[112][8]/P0001  , \wishbone_bd_ram_mem1_reg[112][9]/P0001  , \wishbone_bd_ram_mem1_reg[113][10]/P0001  , \wishbone_bd_ram_mem1_reg[113][11]/P0001  , \wishbone_bd_ram_mem1_reg[113][12]/P0001  , \wishbone_bd_ram_mem1_reg[113][13]/P0001  , \wishbone_bd_ram_mem1_reg[113][14]/P0001  , \wishbone_bd_ram_mem1_reg[113][15]/P0001  , \wishbone_bd_ram_mem1_reg[113][8]/P0001  , \wishbone_bd_ram_mem1_reg[113][9]/P0001  , \wishbone_bd_ram_mem1_reg[114][10]/P0001  , \wishbone_bd_ram_mem1_reg[114][11]/P0001  , \wishbone_bd_ram_mem1_reg[114][12]/P0001  , \wishbone_bd_ram_mem1_reg[114][13]/P0001  , \wishbone_bd_ram_mem1_reg[114][14]/P0001  , \wishbone_bd_ram_mem1_reg[114][15]/P0001  , \wishbone_bd_ram_mem1_reg[114][8]/P0001  , \wishbone_bd_ram_mem1_reg[114][9]/P0001  , \wishbone_bd_ram_mem1_reg[115][10]/P0001  , \wishbone_bd_ram_mem1_reg[115][11]/P0001  , \wishbone_bd_ram_mem1_reg[115][12]/P0001  , \wishbone_bd_ram_mem1_reg[115][13]/P0001  , \wishbone_bd_ram_mem1_reg[115][14]/P0001  , \wishbone_bd_ram_mem1_reg[115][15]/P0001  , \wishbone_bd_ram_mem1_reg[115][8]/P0001  , \wishbone_bd_ram_mem1_reg[115][9]/P0001  , \wishbone_bd_ram_mem1_reg[116][10]/P0001  , \wishbone_bd_ram_mem1_reg[116][11]/P0001  , \wishbone_bd_ram_mem1_reg[116][12]/P0001  , \wishbone_bd_ram_mem1_reg[116][13]/P0001  , \wishbone_bd_ram_mem1_reg[116][14]/P0001  , \wishbone_bd_ram_mem1_reg[116][15]/P0001  , \wishbone_bd_ram_mem1_reg[116][8]/P0001  , \wishbone_bd_ram_mem1_reg[116][9]/P0001  , \wishbone_bd_ram_mem1_reg[117][10]/P0001  , \wishbone_bd_ram_mem1_reg[117][11]/P0001  , \wishbone_bd_ram_mem1_reg[117][12]/P0001  , \wishbone_bd_ram_mem1_reg[117][13]/P0001  , \wishbone_bd_ram_mem1_reg[117][14]/P0001  , \wishbone_bd_ram_mem1_reg[117][15]/P0001  , \wishbone_bd_ram_mem1_reg[117][8]/P0001  , \wishbone_bd_ram_mem1_reg[117][9]/P0001  , \wishbone_bd_ram_mem1_reg[118][10]/P0001  , \wishbone_bd_ram_mem1_reg[118][11]/P0001  , \wishbone_bd_ram_mem1_reg[118][12]/P0001  , \wishbone_bd_ram_mem1_reg[118][13]/P0001  , \wishbone_bd_ram_mem1_reg[118][14]/P0001  , \wishbone_bd_ram_mem1_reg[118][15]/P0001  , \wishbone_bd_ram_mem1_reg[118][8]/P0001  , \wishbone_bd_ram_mem1_reg[118][9]/P0001  , \wishbone_bd_ram_mem1_reg[119][10]/P0001  , \wishbone_bd_ram_mem1_reg[119][11]/P0001  , \wishbone_bd_ram_mem1_reg[119][12]/P0001  , \wishbone_bd_ram_mem1_reg[119][13]/P0001  , \wishbone_bd_ram_mem1_reg[119][14]/P0001  , \wishbone_bd_ram_mem1_reg[119][15]/P0001  , \wishbone_bd_ram_mem1_reg[119][8]/P0001  , \wishbone_bd_ram_mem1_reg[119][9]/P0001  , \wishbone_bd_ram_mem1_reg[11][10]/P0001  , \wishbone_bd_ram_mem1_reg[11][11]/P0001  , \wishbone_bd_ram_mem1_reg[11][12]/P0001  , \wishbone_bd_ram_mem1_reg[11][13]/P0001  , \wishbone_bd_ram_mem1_reg[11][14]/P0001  , \wishbone_bd_ram_mem1_reg[11][15]/P0001  , \wishbone_bd_ram_mem1_reg[11][8]/P0001  , \wishbone_bd_ram_mem1_reg[11][9]/P0001  , \wishbone_bd_ram_mem1_reg[120][10]/P0001  , \wishbone_bd_ram_mem1_reg[120][11]/P0001  , \wishbone_bd_ram_mem1_reg[120][12]/P0001  , \wishbone_bd_ram_mem1_reg[120][13]/P0001  , \wishbone_bd_ram_mem1_reg[120][14]/P0001  , \wishbone_bd_ram_mem1_reg[120][15]/P0001  , \wishbone_bd_ram_mem1_reg[120][8]/P0001  , \wishbone_bd_ram_mem1_reg[120][9]/P0001  , \wishbone_bd_ram_mem1_reg[121][10]/P0001  , \wishbone_bd_ram_mem1_reg[121][11]/P0001  , \wishbone_bd_ram_mem1_reg[121][12]/P0001  , \wishbone_bd_ram_mem1_reg[121][13]/P0001  , \wishbone_bd_ram_mem1_reg[121][14]/P0001  , \wishbone_bd_ram_mem1_reg[121][15]/P0001  , \wishbone_bd_ram_mem1_reg[121][8]/P0001  , \wishbone_bd_ram_mem1_reg[121][9]/P0001  , \wishbone_bd_ram_mem1_reg[122][10]/P0001  , \wishbone_bd_ram_mem1_reg[122][11]/P0001  , \wishbone_bd_ram_mem1_reg[122][12]/P0001  , \wishbone_bd_ram_mem1_reg[122][13]/P0001  , \wishbone_bd_ram_mem1_reg[122][14]/P0001  , \wishbone_bd_ram_mem1_reg[122][15]/P0001  , \wishbone_bd_ram_mem1_reg[122][8]/P0001  , \wishbone_bd_ram_mem1_reg[122][9]/P0001  , \wishbone_bd_ram_mem1_reg[123][10]/P0001  , \wishbone_bd_ram_mem1_reg[123][11]/P0001  , \wishbone_bd_ram_mem1_reg[123][12]/P0001  , \wishbone_bd_ram_mem1_reg[123][13]/P0001  , \wishbone_bd_ram_mem1_reg[123][14]/P0001  , \wishbone_bd_ram_mem1_reg[123][15]/P0001  , \wishbone_bd_ram_mem1_reg[123][8]/P0001  , \wishbone_bd_ram_mem1_reg[123][9]/P0001  , \wishbone_bd_ram_mem1_reg[124][10]/P0001  , \wishbone_bd_ram_mem1_reg[124][11]/P0001  , \wishbone_bd_ram_mem1_reg[124][12]/P0001  , \wishbone_bd_ram_mem1_reg[124][13]/P0001  , \wishbone_bd_ram_mem1_reg[124][14]/P0001  , \wishbone_bd_ram_mem1_reg[124][15]/P0001  , \wishbone_bd_ram_mem1_reg[124][8]/P0001  , \wishbone_bd_ram_mem1_reg[124][9]/P0001  , \wishbone_bd_ram_mem1_reg[125][10]/P0001  , \wishbone_bd_ram_mem1_reg[125][11]/P0001  , \wishbone_bd_ram_mem1_reg[125][12]/P0001  , \wishbone_bd_ram_mem1_reg[125][13]/P0001  , \wishbone_bd_ram_mem1_reg[125][14]/P0001  , \wishbone_bd_ram_mem1_reg[125][15]/P0001  , \wishbone_bd_ram_mem1_reg[125][8]/P0001  , \wishbone_bd_ram_mem1_reg[125][9]/P0001  , \wishbone_bd_ram_mem1_reg[126][10]/P0001  , \wishbone_bd_ram_mem1_reg[126][11]/P0001  , \wishbone_bd_ram_mem1_reg[126][12]/P0001  , \wishbone_bd_ram_mem1_reg[126][13]/P0001  , \wishbone_bd_ram_mem1_reg[126][14]/P0001  , \wishbone_bd_ram_mem1_reg[126][15]/P0001  , \wishbone_bd_ram_mem1_reg[126][8]/P0001  , \wishbone_bd_ram_mem1_reg[126][9]/P0001  , \wishbone_bd_ram_mem1_reg[127][10]/P0001  , \wishbone_bd_ram_mem1_reg[127][11]/P0001  , \wishbone_bd_ram_mem1_reg[127][12]/P0001  , \wishbone_bd_ram_mem1_reg[127][13]/P0001  , \wishbone_bd_ram_mem1_reg[127][14]/P0001  , \wishbone_bd_ram_mem1_reg[127][15]/P0001  , \wishbone_bd_ram_mem1_reg[127][8]/P0001  , \wishbone_bd_ram_mem1_reg[127][9]/P0001  , \wishbone_bd_ram_mem1_reg[128][10]/P0001  , \wishbone_bd_ram_mem1_reg[128][11]/P0001  , \wishbone_bd_ram_mem1_reg[128][12]/P0001  , \wishbone_bd_ram_mem1_reg[128][13]/P0001  , \wishbone_bd_ram_mem1_reg[128][14]/P0001  , \wishbone_bd_ram_mem1_reg[128][15]/P0001  , \wishbone_bd_ram_mem1_reg[128][8]/P0001  , \wishbone_bd_ram_mem1_reg[128][9]/P0001  , \wishbone_bd_ram_mem1_reg[129][10]/P0001  , \wishbone_bd_ram_mem1_reg[129][11]/P0001  , \wishbone_bd_ram_mem1_reg[129][12]/P0001  , \wishbone_bd_ram_mem1_reg[129][13]/P0001  , \wishbone_bd_ram_mem1_reg[129][14]/P0001  , \wishbone_bd_ram_mem1_reg[129][15]/P0001  , \wishbone_bd_ram_mem1_reg[129][8]/P0001  , \wishbone_bd_ram_mem1_reg[129][9]/P0001  , \wishbone_bd_ram_mem1_reg[12][10]/P0001  , \wishbone_bd_ram_mem1_reg[12][11]/P0001  , \wishbone_bd_ram_mem1_reg[12][12]/P0001  , \wishbone_bd_ram_mem1_reg[12][13]/P0001  , \wishbone_bd_ram_mem1_reg[12][14]/P0001  , \wishbone_bd_ram_mem1_reg[12][15]/P0001  , \wishbone_bd_ram_mem1_reg[12][8]/P0001  , \wishbone_bd_ram_mem1_reg[12][9]/P0001  , \wishbone_bd_ram_mem1_reg[130][10]/P0001  , \wishbone_bd_ram_mem1_reg[130][11]/P0001  , \wishbone_bd_ram_mem1_reg[130][12]/P0001  , \wishbone_bd_ram_mem1_reg[130][13]/P0001  , \wishbone_bd_ram_mem1_reg[130][14]/P0001  , \wishbone_bd_ram_mem1_reg[130][15]/P0001  , \wishbone_bd_ram_mem1_reg[130][8]/P0001  , \wishbone_bd_ram_mem1_reg[130][9]/P0001  , \wishbone_bd_ram_mem1_reg[131][10]/P0001  , \wishbone_bd_ram_mem1_reg[131][11]/P0001  , \wishbone_bd_ram_mem1_reg[131][12]/P0001  , \wishbone_bd_ram_mem1_reg[131][13]/P0001  , \wishbone_bd_ram_mem1_reg[131][14]/P0001  , \wishbone_bd_ram_mem1_reg[131][15]/P0001  , \wishbone_bd_ram_mem1_reg[131][8]/P0001  , \wishbone_bd_ram_mem1_reg[131][9]/P0001  , \wishbone_bd_ram_mem1_reg[132][10]/P0001  , \wishbone_bd_ram_mem1_reg[132][11]/P0001  , \wishbone_bd_ram_mem1_reg[132][12]/P0001  , \wishbone_bd_ram_mem1_reg[132][13]/P0001  , \wishbone_bd_ram_mem1_reg[132][14]/P0001  , \wishbone_bd_ram_mem1_reg[132][15]/P0001  , \wishbone_bd_ram_mem1_reg[132][8]/P0001  , \wishbone_bd_ram_mem1_reg[132][9]/P0001  , \wishbone_bd_ram_mem1_reg[133][10]/P0001  , \wishbone_bd_ram_mem1_reg[133][11]/P0001  , \wishbone_bd_ram_mem1_reg[133][12]/P0001  , \wishbone_bd_ram_mem1_reg[133][13]/P0001  , \wishbone_bd_ram_mem1_reg[133][14]/P0001  , \wishbone_bd_ram_mem1_reg[133][15]/P0001  , \wishbone_bd_ram_mem1_reg[133][8]/P0001  , \wishbone_bd_ram_mem1_reg[133][9]/P0001  , \wishbone_bd_ram_mem1_reg[134][10]/P0001  , \wishbone_bd_ram_mem1_reg[134][11]/P0001  , \wishbone_bd_ram_mem1_reg[134][12]/P0001  , \wishbone_bd_ram_mem1_reg[134][13]/P0001  , \wishbone_bd_ram_mem1_reg[134][14]/P0001  , \wishbone_bd_ram_mem1_reg[134][15]/P0001  , \wishbone_bd_ram_mem1_reg[134][8]/P0001  , \wishbone_bd_ram_mem1_reg[134][9]/P0001  , \wishbone_bd_ram_mem1_reg[135][10]/P0001  , \wishbone_bd_ram_mem1_reg[135][11]/P0001  , \wishbone_bd_ram_mem1_reg[135][12]/P0001  , \wishbone_bd_ram_mem1_reg[135][13]/P0001  , \wishbone_bd_ram_mem1_reg[135][14]/P0001  , \wishbone_bd_ram_mem1_reg[135][15]/P0001  , \wishbone_bd_ram_mem1_reg[135][8]/P0001  , \wishbone_bd_ram_mem1_reg[135][9]/P0001  , \wishbone_bd_ram_mem1_reg[136][10]/P0001  , \wishbone_bd_ram_mem1_reg[136][11]/P0001  , \wishbone_bd_ram_mem1_reg[136][12]/P0001  , \wishbone_bd_ram_mem1_reg[136][13]/P0001  , \wishbone_bd_ram_mem1_reg[136][14]/P0001  , \wishbone_bd_ram_mem1_reg[136][15]/P0001  , \wishbone_bd_ram_mem1_reg[136][8]/P0001  , \wishbone_bd_ram_mem1_reg[136][9]/P0001  , \wishbone_bd_ram_mem1_reg[137][10]/P0001  , \wishbone_bd_ram_mem1_reg[137][11]/P0001  , \wishbone_bd_ram_mem1_reg[137][12]/P0001  , \wishbone_bd_ram_mem1_reg[137][13]/P0001  , \wishbone_bd_ram_mem1_reg[137][14]/P0001  , \wishbone_bd_ram_mem1_reg[137][15]/P0001  , \wishbone_bd_ram_mem1_reg[137][8]/P0001  , \wishbone_bd_ram_mem1_reg[137][9]/P0001  , \wishbone_bd_ram_mem1_reg[138][10]/P0001  , \wishbone_bd_ram_mem1_reg[138][11]/P0001  , \wishbone_bd_ram_mem1_reg[138][12]/P0001  , \wishbone_bd_ram_mem1_reg[138][13]/P0001  , \wishbone_bd_ram_mem1_reg[138][14]/P0001  , \wishbone_bd_ram_mem1_reg[138][15]/P0001  , \wishbone_bd_ram_mem1_reg[138][8]/P0001  , \wishbone_bd_ram_mem1_reg[138][9]/P0001  , \wishbone_bd_ram_mem1_reg[139][10]/P0001  , \wishbone_bd_ram_mem1_reg[139][11]/P0001  , \wishbone_bd_ram_mem1_reg[139][12]/P0001  , \wishbone_bd_ram_mem1_reg[139][13]/P0001  , \wishbone_bd_ram_mem1_reg[139][14]/P0001  , \wishbone_bd_ram_mem1_reg[139][15]/P0001  , \wishbone_bd_ram_mem1_reg[139][8]/P0001  , \wishbone_bd_ram_mem1_reg[139][9]/P0001  , \wishbone_bd_ram_mem1_reg[13][10]/P0001  , \wishbone_bd_ram_mem1_reg[13][11]/P0001  , \wishbone_bd_ram_mem1_reg[13][12]/P0001  , \wishbone_bd_ram_mem1_reg[13][13]/P0001  , \wishbone_bd_ram_mem1_reg[13][14]/P0001  , \wishbone_bd_ram_mem1_reg[13][15]/P0001  , \wishbone_bd_ram_mem1_reg[13][8]/P0001  , \wishbone_bd_ram_mem1_reg[13][9]/P0001  , \wishbone_bd_ram_mem1_reg[140][10]/P0001  , \wishbone_bd_ram_mem1_reg[140][11]/P0001  , \wishbone_bd_ram_mem1_reg[140][12]/P0001  , \wishbone_bd_ram_mem1_reg[140][13]/P0001  , \wishbone_bd_ram_mem1_reg[140][14]/P0001  , \wishbone_bd_ram_mem1_reg[140][15]/P0001  , \wishbone_bd_ram_mem1_reg[140][8]/P0001  , \wishbone_bd_ram_mem1_reg[140][9]/P0001  , \wishbone_bd_ram_mem1_reg[141][10]/P0001  , \wishbone_bd_ram_mem1_reg[141][11]/P0001  , \wishbone_bd_ram_mem1_reg[141][12]/P0001  , \wishbone_bd_ram_mem1_reg[141][13]/P0001  , \wishbone_bd_ram_mem1_reg[141][14]/P0001  , \wishbone_bd_ram_mem1_reg[141][15]/P0001  , \wishbone_bd_ram_mem1_reg[141][8]/P0001  , \wishbone_bd_ram_mem1_reg[141][9]/P0001  , \wishbone_bd_ram_mem1_reg[142][10]/P0001  , \wishbone_bd_ram_mem1_reg[142][11]/P0001  , \wishbone_bd_ram_mem1_reg[142][12]/P0001  , \wishbone_bd_ram_mem1_reg[142][13]/P0001  , \wishbone_bd_ram_mem1_reg[142][14]/P0001  , \wishbone_bd_ram_mem1_reg[142][15]/P0001  , \wishbone_bd_ram_mem1_reg[142][8]/P0001  , \wishbone_bd_ram_mem1_reg[142][9]/P0001  , \wishbone_bd_ram_mem1_reg[143][10]/P0001  , \wishbone_bd_ram_mem1_reg[143][11]/P0001  , \wishbone_bd_ram_mem1_reg[143][12]/P0001  , \wishbone_bd_ram_mem1_reg[143][13]/P0001  , \wishbone_bd_ram_mem1_reg[143][14]/P0001  , \wishbone_bd_ram_mem1_reg[143][15]/P0001  , \wishbone_bd_ram_mem1_reg[143][8]/P0001  , \wishbone_bd_ram_mem1_reg[143][9]/P0001  , \wishbone_bd_ram_mem1_reg[144][10]/P0001  , \wishbone_bd_ram_mem1_reg[144][11]/P0001  , \wishbone_bd_ram_mem1_reg[144][12]/P0001  , \wishbone_bd_ram_mem1_reg[144][13]/P0001  , \wishbone_bd_ram_mem1_reg[144][14]/P0001  , \wishbone_bd_ram_mem1_reg[144][15]/P0001  , \wishbone_bd_ram_mem1_reg[144][8]/P0001  , \wishbone_bd_ram_mem1_reg[144][9]/P0001  , \wishbone_bd_ram_mem1_reg[145][10]/P0001  , \wishbone_bd_ram_mem1_reg[145][11]/P0001  , \wishbone_bd_ram_mem1_reg[145][12]/P0001  , \wishbone_bd_ram_mem1_reg[145][13]/P0001  , \wishbone_bd_ram_mem1_reg[145][14]/P0001  , \wishbone_bd_ram_mem1_reg[145][15]/P0001  , \wishbone_bd_ram_mem1_reg[145][8]/P0001  , \wishbone_bd_ram_mem1_reg[145][9]/P0001  , \wishbone_bd_ram_mem1_reg[146][10]/P0001  , \wishbone_bd_ram_mem1_reg[146][11]/P0001  , \wishbone_bd_ram_mem1_reg[146][12]/P0001  , \wishbone_bd_ram_mem1_reg[146][13]/P0001  , \wishbone_bd_ram_mem1_reg[146][14]/P0001  , \wishbone_bd_ram_mem1_reg[146][15]/P0001  , \wishbone_bd_ram_mem1_reg[146][8]/P0001  , \wishbone_bd_ram_mem1_reg[146][9]/P0001  , \wishbone_bd_ram_mem1_reg[147][10]/P0001  , \wishbone_bd_ram_mem1_reg[147][11]/P0001  , \wishbone_bd_ram_mem1_reg[147][12]/P0001  , \wishbone_bd_ram_mem1_reg[147][13]/P0001  , \wishbone_bd_ram_mem1_reg[147][14]/P0001  , \wishbone_bd_ram_mem1_reg[147][15]/P0001  , \wishbone_bd_ram_mem1_reg[147][8]/P0001  , \wishbone_bd_ram_mem1_reg[147][9]/P0001  , \wishbone_bd_ram_mem1_reg[148][10]/P0001  , \wishbone_bd_ram_mem1_reg[148][11]/P0001  , \wishbone_bd_ram_mem1_reg[148][12]/P0001  , \wishbone_bd_ram_mem1_reg[148][13]/P0001  , \wishbone_bd_ram_mem1_reg[148][14]/P0001  , \wishbone_bd_ram_mem1_reg[148][15]/P0001  , \wishbone_bd_ram_mem1_reg[148][8]/P0001  , \wishbone_bd_ram_mem1_reg[148][9]/P0001  , \wishbone_bd_ram_mem1_reg[149][10]/P0001  , \wishbone_bd_ram_mem1_reg[149][11]/P0001  , \wishbone_bd_ram_mem1_reg[149][12]/P0001  , \wishbone_bd_ram_mem1_reg[149][13]/P0001  , \wishbone_bd_ram_mem1_reg[149][14]/P0001  , \wishbone_bd_ram_mem1_reg[149][15]/P0001  , \wishbone_bd_ram_mem1_reg[149][8]/P0001  , \wishbone_bd_ram_mem1_reg[149][9]/P0001  , \wishbone_bd_ram_mem1_reg[14][10]/P0001  , \wishbone_bd_ram_mem1_reg[14][11]/P0001  , \wishbone_bd_ram_mem1_reg[14][12]/P0001  , \wishbone_bd_ram_mem1_reg[14][13]/P0001  , \wishbone_bd_ram_mem1_reg[14][14]/P0001  , \wishbone_bd_ram_mem1_reg[14][15]/P0001  , \wishbone_bd_ram_mem1_reg[14][8]/P0001  , \wishbone_bd_ram_mem1_reg[14][9]/P0001  , \wishbone_bd_ram_mem1_reg[150][10]/P0001  , \wishbone_bd_ram_mem1_reg[150][11]/P0001  , \wishbone_bd_ram_mem1_reg[150][12]/P0001  , \wishbone_bd_ram_mem1_reg[150][13]/P0001  , \wishbone_bd_ram_mem1_reg[150][14]/P0001  , \wishbone_bd_ram_mem1_reg[150][15]/P0001  , \wishbone_bd_ram_mem1_reg[150][8]/P0001  , \wishbone_bd_ram_mem1_reg[150][9]/P0001  , \wishbone_bd_ram_mem1_reg[151][10]/P0001  , \wishbone_bd_ram_mem1_reg[151][11]/P0001  , \wishbone_bd_ram_mem1_reg[151][12]/P0001  , \wishbone_bd_ram_mem1_reg[151][13]/P0001  , \wishbone_bd_ram_mem1_reg[151][14]/P0001  , \wishbone_bd_ram_mem1_reg[151][15]/P0001  , \wishbone_bd_ram_mem1_reg[151][8]/P0001  , \wishbone_bd_ram_mem1_reg[151][9]/P0001  , \wishbone_bd_ram_mem1_reg[152][10]/P0001  , \wishbone_bd_ram_mem1_reg[152][11]/P0001  , \wishbone_bd_ram_mem1_reg[152][12]/P0001  , \wishbone_bd_ram_mem1_reg[152][13]/P0001  , \wishbone_bd_ram_mem1_reg[152][14]/P0001  , \wishbone_bd_ram_mem1_reg[152][15]/P0001  , \wishbone_bd_ram_mem1_reg[152][8]/P0001  , \wishbone_bd_ram_mem1_reg[152][9]/P0001  , \wishbone_bd_ram_mem1_reg[153][10]/P0001  , \wishbone_bd_ram_mem1_reg[153][11]/P0001  , \wishbone_bd_ram_mem1_reg[153][12]/P0001  , \wishbone_bd_ram_mem1_reg[153][13]/P0001  , \wishbone_bd_ram_mem1_reg[153][14]/P0001  , \wishbone_bd_ram_mem1_reg[153][15]/P0001  , \wishbone_bd_ram_mem1_reg[153][8]/P0001  , \wishbone_bd_ram_mem1_reg[153][9]/P0001  , \wishbone_bd_ram_mem1_reg[154][10]/P0001  , \wishbone_bd_ram_mem1_reg[154][11]/P0001  , \wishbone_bd_ram_mem1_reg[154][12]/P0001  , \wishbone_bd_ram_mem1_reg[154][13]/P0001  , \wishbone_bd_ram_mem1_reg[154][14]/P0001  , \wishbone_bd_ram_mem1_reg[154][15]/P0001  , \wishbone_bd_ram_mem1_reg[154][8]/P0001  , \wishbone_bd_ram_mem1_reg[154][9]/P0001  , \wishbone_bd_ram_mem1_reg[155][10]/P0001  , \wishbone_bd_ram_mem1_reg[155][11]/P0001  , \wishbone_bd_ram_mem1_reg[155][12]/P0001  , \wishbone_bd_ram_mem1_reg[155][13]/P0001  , \wishbone_bd_ram_mem1_reg[155][14]/P0001  , \wishbone_bd_ram_mem1_reg[155][15]/P0001  , \wishbone_bd_ram_mem1_reg[155][8]/P0001  , \wishbone_bd_ram_mem1_reg[155][9]/P0001  , \wishbone_bd_ram_mem1_reg[156][10]/P0001  , \wishbone_bd_ram_mem1_reg[156][11]/P0001  , \wishbone_bd_ram_mem1_reg[156][12]/P0001  , \wishbone_bd_ram_mem1_reg[156][13]/P0001  , \wishbone_bd_ram_mem1_reg[156][14]/P0001  , \wishbone_bd_ram_mem1_reg[156][15]/P0001  , \wishbone_bd_ram_mem1_reg[156][8]/P0001  , \wishbone_bd_ram_mem1_reg[156][9]/P0001  , \wishbone_bd_ram_mem1_reg[157][10]/P0001  , \wishbone_bd_ram_mem1_reg[157][11]/P0001  , \wishbone_bd_ram_mem1_reg[157][12]/P0001  , \wishbone_bd_ram_mem1_reg[157][13]/P0001  , \wishbone_bd_ram_mem1_reg[157][14]/P0001  , \wishbone_bd_ram_mem1_reg[157][15]/P0001  , \wishbone_bd_ram_mem1_reg[157][8]/P0001  , \wishbone_bd_ram_mem1_reg[157][9]/P0001  , \wishbone_bd_ram_mem1_reg[158][10]/P0001  , \wishbone_bd_ram_mem1_reg[158][11]/P0001  , \wishbone_bd_ram_mem1_reg[158][12]/P0001  , \wishbone_bd_ram_mem1_reg[158][13]/P0001  , \wishbone_bd_ram_mem1_reg[158][14]/P0001  , \wishbone_bd_ram_mem1_reg[158][15]/P0001  , \wishbone_bd_ram_mem1_reg[158][8]/P0001  , \wishbone_bd_ram_mem1_reg[158][9]/P0001  , \wishbone_bd_ram_mem1_reg[159][10]/P0001  , \wishbone_bd_ram_mem1_reg[159][11]/P0001  , \wishbone_bd_ram_mem1_reg[159][12]/P0001  , \wishbone_bd_ram_mem1_reg[159][13]/P0001  , \wishbone_bd_ram_mem1_reg[159][14]/P0001  , \wishbone_bd_ram_mem1_reg[159][15]/P0001  , \wishbone_bd_ram_mem1_reg[159][8]/P0001  , \wishbone_bd_ram_mem1_reg[159][9]/P0001  , \wishbone_bd_ram_mem1_reg[15][10]/P0001  , \wishbone_bd_ram_mem1_reg[15][11]/P0001  , \wishbone_bd_ram_mem1_reg[15][12]/P0001  , \wishbone_bd_ram_mem1_reg[15][13]/P0001  , \wishbone_bd_ram_mem1_reg[15][14]/P0001  , \wishbone_bd_ram_mem1_reg[15][15]/P0001  , \wishbone_bd_ram_mem1_reg[15][8]/P0001  , \wishbone_bd_ram_mem1_reg[15][9]/P0001  , \wishbone_bd_ram_mem1_reg[160][10]/P0001  , \wishbone_bd_ram_mem1_reg[160][11]/P0001  , \wishbone_bd_ram_mem1_reg[160][12]/P0001  , \wishbone_bd_ram_mem1_reg[160][13]/P0001  , \wishbone_bd_ram_mem1_reg[160][14]/P0001  , \wishbone_bd_ram_mem1_reg[160][15]/P0001  , \wishbone_bd_ram_mem1_reg[160][8]/P0001  , \wishbone_bd_ram_mem1_reg[160][9]/P0001  , \wishbone_bd_ram_mem1_reg[161][10]/P0001  , \wishbone_bd_ram_mem1_reg[161][11]/P0001  , \wishbone_bd_ram_mem1_reg[161][12]/P0001  , \wishbone_bd_ram_mem1_reg[161][13]/P0001  , \wishbone_bd_ram_mem1_reg[161][14]/P0001  , \wishbone_bd_ram_mem1_reg[161][15]/P0001  , \wishbone_bd_ram_mem1_reg[161][8]/P0001  , \wishbone_bd_ram_mem1_reg[161][9]/P0001  , \wishbone_bd_ram_mem1_reg[162][10]/P0001  , \wishbone_bd_ram_mem1_reg[162][11]/P0001  , \wishbone_bd_ram_mem1_reg[162][12]/P0001  , \wishbone_bd_ram_mem1_reg[162][13]/P0001  , \wishbone_bd_ram_mem1_reg[162][14]/P0001  , \wishbone_bd_ram_mem1_reg[162][15]/P0001  , \wishbone_bd_ram_mem1_reg[162][8]/P0001  , \wishbone_bd_ram_mem1_reg[162][9]/P0001  , \wishbone_bd_ram_mem1_reg[163][10]/P0001  , \wishbone_bd_ram_mem1_reg[163][11]/P0001  , \wishbone_bd_ram_mem1_reg[163][12]/P0001  , \wishbone_bd_ram_mem1_reg[163][13]/P0001  , \wishbone_bd_ram_mem1_reg[163][14]/P0001  , \wishbone_bd_ram_mem1_reg[163][15]/P0001  , \wishbone_bd_ram_mem1_reg[163][8]/P0001  , \wishbone_bd_ram_mem1_reg[163][9]/P0001  , \wishbone_bd_ram_mem1_reg[164][10]/P0001  , \wishbone_bd_ram_mem1_reg[164][11]/P0001  , \wishbone_bd_ram_mem1_reg[164][12]/P0001  , \wishbone_bd_ram_mem1_reg[164][13]/P0001  , \wishbone_bd_ram_mem1_reg[164][14]/P0001  , \wishbone_bd_ram_mem1_reg[164][15]/P0001  , \wishbone_bd_ram_mem1_reg[164][8]/P0001  , \wishbone_bd_ram_mem1_reg[164][9]/P0001  , \wishbone_bd_ram_mem1_reg[165][10]/P0001  , \wishbone_bd_ram_mem1_reg[165][11]/P0001  , \wishbone_bd_ram_mem1_reg[165][12]/P0001  , \wishbone_bd_ram_mem1_reg[165][13]/P0001  , \wishbone_bd_ram_mem1_reg[165][14]/P0001  , \wishbone_bd_ram_mem1_reg[165][15]/P0001  , \wishbone_bd_ram_mem1_reg[165][8]/P0001  , \wishbone_bd_ram_mem1_reg[165][9]/P0001  , \wishbone_bd_ram_mem1_reg[166][10]/P0001  , \wishbone_bd_ram_mem1_reg[166][11]/P0001  , \wishbone_bd_ram_mem1_reg[166][12]/P0001  , \wishbone_bd_ram_mem1_reg[166][13]/P0001  , \wishbone_bd_ram_mem1_reg[166][14]/P0001  , \wishbone_bd_ram_mem1_reg[166][15]/P0001  , \wishbone_bd_ram_mem1_reg[166][8]/P0001  , \wishbone_bd_ram_mem1_reg[166][9]/P0001  , \wishbone_bd_ram_mem1_reg[167][10]/P0001  , \wishbone_bd_ram_mem1_reg[167][11]/P0001  , \wishbone_bd_ram_mem1_reg[167][12]/P0001  , \wishbone_bd_ram_mem1_reg[167][13]/P0001  , \wishbone_bd_ram_mem1_reg[167][14]/P0001  , \wishbone_bd_ram_mem1_reg[167][15]/P0001  , \wishbone_bd_ram_mem1_reg[167][8]/P0001  , \wishbone_bd_ram_mem1_reg[167][9]/P0001  , \wishbone_bd_ram_mem1_reg[168][10]/P0001  , \wishbone_bd_ram_mem1_reg[168][11]/P0001  , \wishbone_bd_ram_mem1_reg[168][12]/P0001  , \wishbone_bd_ram_mem1_reg[168][13]/P0001  , \wishbone_bd_ram_mem1_reg[168][14]/P0001  , \wishbone_bd_ram_mem1_reg[168][15]/P0001  , \wishbone_bd_ram_mem1_reg[168][8]/P0001  , \wishbone_bd_ram_mem1_reg[168][9]/P0001  , \wishbone_bd_ram_mem1_reg[169][10]/P0001  , \wishbone_bd_ram_mem1_reg[169][11]/P0001  , \wishbone_bd_ram_mem1_reg[169][12]/P0001  , \wishbone_bd_ram_mem1_reg[169][13]/P0001  , \wishbone_bd_ram_mem1_reg[169][14]/P0001  , \wishbone_bd_ram_mem1_reg[169][15]/P0001  , \wishbone_bd_ram_mem1_reg[169][8]/P0001  , \wishbone_bd_ram_mem1_reg[169][9]/P0001  , \wishbone_bd_ram_mem1_reg[16][10]/P0001  , \wishbone_bd_ram_mem1_reg[16][11]/P0001  , \wishbone_bd_ram_mem1_reg[16][12]/P0001  , \wishbone_bd_ram_mem1_reg[16][13]/P0001  , \wishbone_bd_ram_mem1_reg[16][14]/P0001  , \wishbone_bd_ram_mem1_reg[16][15]/P0001  , \wishbone_bd_ram_mem1_reg[16][8]/P0001  , \wishbone_bd_ram_mem1_reg[16][9]/P0001  , \wishbone_bd_ram_mem1_reg[170][10]/P0001  , \wishbone_bd_ram_mem1_reg[170][11]/P0001  , \wishbone_bd_ram_mem1_reg[170][12]/P0001  , \wishbone_bd_ram_mem1_reg[170][13]/P0001  , \wishbone_bd_ram_mem1_reg[170][14]/P0001  , \wishbone_bd_ram_mem1_reg[170][15]/P0001  , \wishbone_bd_ram_mem1_reg[170][8]/P0001  , \wishbone_bd_ram_mem1_reg[170][9]/P0001  , \wishbone_bd_ram_mem1_reg[171][10]/P0001  , \wishbone_bd_ram_mem1_reg[171][11]/P0001  , \wishbone_bd_ram_mem1_reg[171][12]/P0001  , \wishbone_bd_ram_mem1_reg[171][13]/P0001  , \wishbone_bd_ram_mem1_reg[171][14]/P0001  , \wishbone_bd_ram_mem1_reg[171][15]/P0001  , \wishbone_bd_ram_mem1_reg[171][8]/P0001  , \wishbone_bd_ram_mem1_reg[171][9]/P0001  , \wishbone_bd_ram_mem1_reg[172][10]/P0001  , \wishbone_bd_ram_mem1_reg[172][11]/P0001  , \wishbone_bd_ram_mem1_reg[172][12]/P0001  , \wishbone_bd_ram_mem1_reg[172][13]/P0001  , \wishbone_bd_ram_mem1_reg[172][14]/P0001  , \wishbone_bd_ram_mem1_reg[172][15]/P0001  , \wishbone_bd_ram_mem1_reg[172][8]/P0001  , \wishbone_bd_ram_mem1_reg[172][9]/P0001  , \wishbone_bd_ram_mem1_reg[173][10]/P0001  , \wishbone_bd_ram_mem1_reg[173][11]/P0001  , \wishbone_bd_ram_mem1_reg[173][12]/P0001  , \wishbone_bd_ram_mem1_reg[173][13]/P0001  , \wishbone_bd_ram_mem1_reg[173][14]/P0001  , \wishbone_bd_ram_mem1_reg[173][15]/P0001  , \wishbone_bd_ram_mem1_reg[173][8]/P0001  , \wishbone_bd_ram_mem1_reg[173][9]/P0001  , \wishbone_bd_ram_mem1_reg[174][10]/P0001  , \wishbone_bd_ram_mem1_reg[174][11]/P0001  , \wishbone_bd_ram_mem1_reg[174][12]/P0001  , \wishbone_bd_ram_mem1_reg[174][13]/P0001  , \wishbone_bd_ram_mem1_reg[174][14]/P0001  , \wishbone_bd_ram_mem1_reg[174][15]/P0001  , \wishbone_bd_ram_mem1_reg[174][8]/P0001  , \wishbone_bd_ram_mem1_reg[174][9]/P0001  , \wishbone_bd_ram_mem1_reg[175][10]/P0001  , \wishbone_bd_ram_mem1_reg[175][11]/P0001  , \wishbone_bd_ram_mem1_reg[175][12]/P0001  , \wishbone_bd_ram_mem1_reg[175][13]/P0001  , \wishbone_bd_ram_mem1_reg[175][14]/P0001  , \wishbone_bd_ram_mem1_reg[175][15]/P0001  , \wishbone_bd_ram_mem1_reg[175][8]/P0001  , \wishbone_bd_ram_mem1_reg[175][9]/P0001  , \wishbone_bd_ram_mem1_reg[176][10]/P0001  , \wishbone_bd_ram_mem1_reg[176][11]/P0001  , \wishbone_bd_ram_mem1_reg[176][12]/P0001  , \wishbone_bd_ram_mem1_reg[176][13]/P0001  , \wishbone_bd_ram_mem1_reg[176][14]/P0001  , \wishbone_bd_ram_mem1_reg[176][15]/P0001  , \wishbone_bd_ram_mem1_reg[176][8]/P0001  , \wishbone_bd_ram_mem1_reg[176][9]/P0001  , \wishbone_bd_ram_mem1_reg[177][10]/P0001  , \wishbone_bd_ram_mem1_reg[177][11]/P0001  , \wishbone_bd_ram_mem1_reg[177][12]/P0001  , \wishbone_bd_ram_mem1_reg[177][13]/P0001  , \wishbone_bd_ram_mem1_reg[177][14]/P0001  , \wishbone_bd_ram_mem1_reg[177][15]/P0001  , \wishbone_bd_ram_mem1_reg[177][8]/P0001  , \wishbone_bd_ram_mem1_reg[177][9]/P0001  , \wishbone_bd_ram_mem1_reg[178][10]/P0001  , \wishbone_bd_ram_mem1_reg[178][11]/P0001  , \wishbone_bd_ram_mem1_reg[178][12]/P0001  , \wishbone_bd_ram_mem1_reg[178][13]/P0001  , \wishbone_bd_ram_mem1_reg[178][14]/P0001  , \wishbone_bd_ram_mem1_reg[178][15]/P0001  , \wishbone_bd_ram_mem1_reg[178][8]/P0001  , \wishbone_bd_ram_mem1_reg[178][9]/P0001  , \wishbone_bd_ram_mem1_reg[179][10]/P0001  , \wishbone_bd_ram_mem1_reg[179][11]/P0001  , \wishbone_bd_ram_mem1_reg[179][12]/P0001  , \wishbone_bd_ram_mem1_reg[179][13]/P0001  , \wishbone_bd_ram_mem1_reg[179][14]/P0001  , \wishbone_bd_ram_mem1_reg[179][15]/P0001  , \wishbone_bd_ram_mem1_reg[179][8]/P0001  , \wishbone_bd_ram_mem1_reg[179][9]/P0001  , \wishbone_bd_ram_mem1_reg[17][10]/P0001  , \wishbone_bd_ram_mem1_reg[17][11]/P0001  , \wishbone_bd_ram_mem1_reg[17][12]/P0001  , \wishbone_bd_ram_mem1_reg[17][13]/P0001  , \wishbone_bd_ram_mem1_reg[17][14]/P0001  , \wishbone_bd_ram_mem1_reg[17][15]/P0001  , \wishbone_bd_ram_mem1_reg[17][8]/P0001  , \wishbone_bd_ram_mem1_reg[17][9]/P0001  , \wishbone_bd_ram_mem1_reg[180][10]/P0001  , \wishbone_bd_ram_mem1_reg[180][11]/P0001  , \wishbone_bd_ram_mem1_reg[180][12]/P0001  , \wishbone_bd_ram_mem1_reg[180][13]/P0001  , \wishbone_bd_ram_mem1_reg[180][14]/P0001  , \wishbone_bd_ram_mem1_reg[180][15]/P0001  , \wishbone_bd_ram_mem1_reg[180][8]/P0001  , \wishbone_bd_ram_mem1_reg[180][9]/P0001  , \wishbone_bd_ram_mem1_reg[181][10]/P0001  , \wishbone_bd_ram_mem1_reg[181][11]/P0001  , \wishbone_bd_ram_mem1_reg[181][12]/P0001  , \wishbone_bd_ram_mem1_reg[181][13]/P0001  , \wishbone_bd_ram_mem1_reg[181][14]/P0001  , \wishbone_bd_ram_mem1_reg[181][15]/P0001  , \wishbone_bd_ram_mem1_reg[181][8]/P0001  , \wishbone_bd_ram_mem1_reg[181][9]/P0001  , \wishbone_bd_ram_mem1_reg[182][10]/P0001  , \wishbone_bd_ram_mem1_reg[182][11]/P0001  , \wishbone_bd_ram_mem1_reg[182][12]/P0001  , \wishbone_bd_ram_mem1_reg[182][13]/P0001  , \wishbone_bd_ram_mem1_reg[182][14]/P0001  , \wishbone_bd_ram_mem1_reg[182][15]/P0001  , \wishbone_bd_ram_mem1_reg[182][8]/P0001  , \wishbone_bd_ram_mem1_reg[182][9]/P0001  , \wishbone_bd_ram_mem1_reg[183][10]/P0001  , \wishbone_bd_ram_mem1_reg[183][11]/P0001  , \wishbone_bd_ram_mem1_reg[183][12]/P0001  , \wishbone_bd_ram_mem1_reg[183][13]/P0001  , \wishbone_bd_ram_mem1_reg[183][14]/P0001  , \wishbone_bd_ram_mem1_reg[183][15]/P0001  , \wishbone_bd_ram_mem1_reg[183][8]/P0001  , \wishbone_bd_ram_mem1_reg[183][9]/P0001  , \wishbone_bd_ram_mem1_reg[184][10]/P0001  , \wishbone_bd_ram_mem1_reg[184][11]/P0001  , \wishbone_bd_ram_mem1_reg[184][12]/P0001  , \wishbone_bd_ram_mem1_reg[184][13]/P0001  , \wishbone_bd_ram_mem1_reg[184][14]/P0001  , \wishbone_bd_ram_mem1_reg[184][15]/P0001  , \wishbone_bd_ram_mem1_reg[184][8]/P0001  , \wishbone_bd_ram_mem1_reg[184][9]/P0001  , \wishbone_bd_ram_mem1_reg[185][10]/P0001  , \wishbone_bd_ram_mem1_reg[185][11]/P0001  , \wishbone_bd_ram_mem1_reg[185][12]/P0001  , \wishbone_bd_ram_mem1_reg[185][13]/P0001  , \wishbone_bd_ram_mem1_reg[185][14]/P0001  , \wishbone_bd_ram_mem1_reg[185][15]/P0001  , \wishbone_bd_ram_mem1_reg[185][8]/P0001  , \wishbone_bd_ram_mem1_reg[185][9]/P0001  , \wishbone_bd_ram_mem1_reg[186][10]/P0001  , \wishbone_bd_ram_mem1_reg[186][11]/P0001  , \wishbone_bd_ram_mem1_reg[186][12]/P0001  , \wishbone_bd_ram_mem1_reg[186][13]/P0001  , \wishbone_bd_ram_mem1_reg[186][14]/P0001  , \wishbone_bd_ram_mem1_reg[186][15]/P0001  , \wishbone_bd_ram_mem1_reg[186][8]/P0001  , \wishbone_bd_ram_mem1_reg[186][9]/P0001  , \wishbone_bd_ram_mem1_reg[187][10]/P0001  , \wishbone_bd_ram_mem1_reg[187][11]/P0001  , \wishbone_bd_ram_mem1_reg[187][12]/P0001  , \wishbone_bd_ram_mem1_reg[187][13]/P0001  , \wishbone_bd_ram_mem1_reg[187][14]/P0001  , \wishbone_bd_ram_mem1_reg[187][15]/P0001  , \wishbone_bd_ram_mem1_reg[187][8]/P0001  , \wishbone_bd_ram_mem1_reg[187][9]/P0001  , \wishbone_bd_ram_mem1_reg[188][10]/P0001  , \wishbone_bd_ram_mem1_reg[188][11]/P0001  , \wishbone_bd_ram_mem1_reg[188][12]/P0001  , \wishbone_bd_ram_mem1_reg[188][13]/P0001  , \wishbone_bd_ram_mem1_reg[188][14]/P0001  , \wishbone_bd_ram_mem1_reg[188][15]/P0001  , \wishbone_bd_ram_mem1_reg[188][8]/P0001  , \wishbone_bd_ram_mem1_reg[188][9]/P0001  , \wishbone_bd_ram_mem1_reg[189][10]/P0001  , \wishbone_bd_ram_mem1_reg[189][11]/P0001  , \wishbone_bd_ram_mem1_reg[189][12]/P0001  , \wishbone_bd_ram_mem1_reg[189][13]/P0001  , \wishbone_bd_ram_mem1_reg[189][14]/P0001  , \wishbone_bd_ram_mem1_reg[189][15]/P0001  , \wishbone_bd_ram_mem1_reg[189][8]/P0001  , \wishbone_bd_ram_mem1_reg[189][9]/P0001  , \wishbone_bd_ram_mem1_reg[18][10]/P0001  , \wishbone_bd_ram_mem1_reg[18][11]/P0001  , \wishbone_bd_ram_mem1_reg[18][12]/P0001  , \wishbone_bd_ram_mem1_reg[18][13]/P0001  , \wishbone_bd_ram_mem1_reg[18][14]/P0001  , \wishbone_bd_ram_mem1_reg[18][15]/P0001  , \wishbone_bd_ram_mem1_reg[18][8]/P0001  , \wishbone_bd_ram_mem1_reg[18][9]/P0001  , \wishbone_bd_ram_mem1_reg[190][10]/P0001  , \wishbone_bd_ram_mem1_reg[190][11]/P0001  , \wishbone_bd_ram_mem1_reg[190][12]/P0001  , \wishbone_bd_ram_mem1_reg[190][13]/P0001  , \wishbone_bd_ram_mem1_reg[190][14]/P0001  , \wishbone_bd_ram_mem1_reg[190][15]/P0001  , \wishbone_bd_ram_mem1_reg[190][8]/P0001  , \wishbone_bd_ram_mem1_reg[190][9]/P0001  , \wishbone_bd_ram_mem1_reg[191][10]/P0001  , \wishbone_bd_ram_mem1_reg[191][11]/P0001  , \wishbone_bd_ram_mem1_reg[191][12]/P0001  , \wishbone_bd_ram_mem1_reg[191][13]/P0001  , \wishbone_bd_ram_mem1_reg[191][14]/P0001  , \wishbone_bd_ram_mem1_reg[191][15]/P0001  , \wishbone_bd_ram_mem1_reg[191][8]/P0001  , \wishbone_bd_ram_mem1_reg[191][9]/P0001  , \wishbone_bd_ram_mem1_reg[192][10]/P0001  , \wishbone_bd_ram_mem1_reg[192][11]/P0001  , \wishbone_bd_ram_mem1_reg[192][12]/P0001  , \wishbone_bd_ram_mem1_reg[192][13]/P0001  , \wishbone_bd_ram_mem1_reg[192][14]/P0001  , \wishbone_bd_ram_mem1_reg[192][15]/P0001  , \wishbone_bd_ram_mem1_reg[192][8]/P0001  , \wishbone_bd_ram_mem1_reg[192][9]/P0001  , \wishbone_bd_ram_mem1_reg[193][10]/P0001  , \wishbone_bd_ram_mem1_reg[193][11]/P0001  , \wishbone_bd_ram_mem1_reg[193][12]/P0001  , \wishbone_bd_ram_mem1_reg[193][13]/P0001  , \wishbone_bd_ram_mem1_reg[193][14]/P0001  , \wishbone_bd_ram_mem1_reg[193][15]/P0001  , \wishbone_bd_ram_mem1_reg[193][8]/P0001  , \wishbone_bd_ram_mem1_reg[193][9]/P0001  , \wishbone_bd_ram_mem1_reg[194][10]/P0001  , \wishbone_bd_ram_mem1_reg[194][11]/P0001  , \wishbone_bd_ram_mem1_reg[194][12]/P0001  , \wishbone_bd_ram_mem1_reg[194][13]/P0001  , \wishbone_bd_ram_mem1_reg[194][14]/P0001  , \wishbone_bd_ram_mem1_reg[194][15]/P0001  , \wishbone_bd_ram_mem1_reg[194][8]/P0001  , \wishbone_bd_ram_mem1_reg[194][9]/P0001  , \wishbone_bd_ram_mem1_reg[195][10]/P0001  , \wishbone_bd_ram_mem1_reg[195][11]/P0001  , \wishbone_bd_ram_mem1_reg[195][12]/P0001  , \wishbone_bd_ram_mem1_reg[195][13]/P0001  , \wishbone_bd_ram_mem1_reg[195][14]/P0001  , \wishbone_bd_ram_mem1_reg[195][15]/P0001  , \wishbone_bd_ram_mem1_reg[195][8]/P0001  , \wishbone_bd_ram_mem1_reg[195][9]/P0001  , \wishbone_bd_ram_mem1_reg[196][10]/P0001  , \wishbone_bd_ram_mem1_reg[196][11]/P0001  , \wishbone_bd_ram_mem1_reg[196][12]/P0001  , \wishbone_bd_ram_mem1_reg[196][13]/P0001  , \wishbone_bd_ram_mem1_reg[196][14]/P0001  , \wishbone_bd_ram_mem1_reg[196][15]/P0001  , \wishbone_bd_ram_mem1_reg[196][8]/P0001  , \wishbone_bd_ram_mem1_reg[196][9]/P0001  , \wishbone_bd_ram_mem1_reg[197][10]/P0001  , \wishbone_bd_ram_mem1_reg[197][11]/P0001  , \wishbone_bd_ram_mem1_reg[197][12]/P0001  , \wishbone_bd_ram_mem1_reg[197][13]/P0001  , \wishbone_bd_ram_mem1_reg[197][14]/P0001  , \wishbone_bd_ram_mem1_reg[197][15]/P0001  , \wishbone_bd_ram_mem1_reg[197][8]/P0001  , \wishbone_bd_ram_mem1_reg[197][9]/P0001  , \wishbone_bd_ram_mem1_reg[198][10]/P0001  , \wishbone_bd_ram_mem1_reg[198][11]/P0001  , \wishbone_bd_ram_mem1_reg[198][12]/P0001  , \wishbone_bd_ram_mem1_reg[198][13]/P0001  , \wishbone_bd_ram_mem1_reg[198][14]/P0001  , \wishbone_bd_ram_mem1_reg[198][15]/P0001  , \wishbone_bd_ram_mem1_reg[198][8]/P0001  , \wishbone_bd_ram_mem1_reg[198][9]/P0001  , \wishbone_bd_ram_mem1_reg[199][10]/P0001  , \wishbone_bd_ram_mem1_reg[199][11]/P0001  , \wishbone_bd_ram_mem1_reg[199][12]/P0001  , \wishbone_bd_ram_mem1_reg[199][13]/P0001  , \wishbone_bd_ram_mem1_reg[199][14]/P0001  , \wishbone_bd_ram_mem1_reg[199][15]/P0001  , \wishbone_bd_ram_mem1_reg[199][8]/P0001  , \wishbone_bd_ram_mem1_reg[199][9]/P0001  , \wishbone_bd_ram_mem1_reg[19][10]/P0001  , \wishbone_bd_ram_mem1_reg[19][11]/P0001  , \wishbone_bd_ram_mem1_reg[19][12]/P0001  , \wishbone_bd_ram_mem1_reg[19][13]/P0001  , \wishbone_bd_ram_mem1_reg[19][14]/P0001  , \wishbone_bd_ram_mem1_reg[19][15]/P0001  , \wishbone_bd_ram_mem1_reg[19][8]/P0001  , \wishbone_bd_ram_mem1_reg[19][9]/P0001  , \wishbone_bd_ram_mem1_reg[1][10]/P0001  , \wishbone_bd_ram_mem1_reg[1][11]/P0001  , \wishbone_bd_ram_mem1_reg[1][12]/P0001  , \wishbone_bd_ram_mem1_reg[1][13]/P0001  , \wishbone_bd_ram_mem1_reg[1][14]/P0001  , \wishbone_bd_ram_mem1_reg[1][15]/P0001  , \wishbone_bd_ram_mem1_reg[1][8]/P0001  , \wishbone_bd_ram_mem1_reg[1][9]/P0001  , \wishbone_bd_ram_mem1_reg[200][10]/P0001  , \wishbone_bd_ram_mem1_reg[200][11]/P0001  , \wishbone_bd_ram_mem1_reg[200][12]/P0001  , \wishbone_bd_ram_mem1_reg[200][13]/P0001  , \wishbone_bd_ram_mem1_reg[200][14]/P0001  , \wishbone_bd_ram_mem1_reg[200][15]/P0001  , \wishbone_bd_ram_mem1_reg[200][8]/P0001  , \wishbone_bd_ram_mem1_reg[200][9]/P0001  , \wishbone_bd_ram_mem1_reg[201][10]/P0001  , \wishbone_bd_ram_mem1_reg[201][11]/P0001  , \wishbone_bd_ram_mem1_reg[201][12]/P0001  , \wishbone_bd_ram_mem1_reg[201][13]/P0001  , \wishbone_bd_ram_mem1_reg[201][14]/P0001  , \wishbone_bd_ram_mem1_reg[201][15]/P0001  , \wishbone_bd_ram_mem1_reg[201][8]/P0001  , \wishbone_bd_ram_mem1_reg[201][9]/P0001  , \wishbone_bd_ram_mem1_reg[202][10]/P0001  , \wishbone_bd_ram_mem1_reg[202][11]/P0001  , \wishbone_bd_ram_mem1_reg[202][12]/P0001  , \wishbone_bd_ram_mem1_reg[202][13]/P0001  , \wishbone_bd_ram_mem1_reg[202][14]/P0001  , \wishbone_bd_ram_mem1_reg[202][15]/P0001  , \wishbone_bd_ram_mem1_reg[202][8]/P0001  , \wishbone_bd_ram_mem1_reg[202][9]/P0001  , \wishbone_bd_ram_mem1_reg[203][10]/P0001  , \wishbone_bd_ram_mem1_reg[203][11]/P0001  , \wishbone_bd_ram_mem1_reg[203][12]/P0001  , \wishbone_bd_ram_mem1_reg[203][13]/P0001  , \wishbone_bd_ram_mem1_reg[203][14]/P0001  , \wishbone_bd_ram_mem1_reg[203][15]/P0001  , \wishbone_bd_ram_mem1_reg[203][8]/P0001  , \wishbone_bd_ram_mem1_reg[203][9]/P0001  , \wishbone_bd_ram_mem1_reg[204][10]/P0001  , \wishbone_bd_ram_mem1_reg[204][11]/P0001  , \wishbone_bd_ram_mem1_reg[204][12]/P0001  , \wishbone_bd_ram_mem1_reg[204][13]/P0001  , \wishbone_bd_ram_mem1_reg[204][14]/P0001  , \wishbone_bd_ram_mem1_reg[204][15]/P0001  , \wishbone_bd_ram_mem1_reg[204][8]/P0001  , \wishbone_bd_ram_mem1_reg[204][9]/P0001  , \wishbone_bd_ram_mem1_reg[205][10]/P0001  , \wishbone_bd_ram_mem1_reg[205][11]/P0001  , \wishbone_bd_ram_mem1_reg[205][12]/P0001  , \wishbone_bd_ram_mem1_reg[205][13]/P0001  , \wishbone_bd_ram_mem1_reg[205][14]/P0001  , \wishbone_bd_ram_mem1_reg[205][15]/P0001  , \wishbone_bd_ram_mem1_reg[205][8]/P0001  , \wishbone_bd_ram_mem1_reg[205][9]/P0001  , \wishbone_bd_ram_mem1_reg[206][10]/P0001  , \wishbone_bd_ram_mem1_reg[206][11]/P0001  , \wishbone_bd_ram_mem1_reg[206][12]/P0001  , \wishbone_bd_ram_mem1_reg[206][13]/P0001  , \wishbone_bd_ram_mem1_reg[206][14]/P0001  , \wishbone_bd_ram_mem1_reg[206][15]/P0001  , \wishbone_bd_ram_mem1_reg[206][8]/P0001  , \wishbone_bd_ram_mem1_reg[206][9]/P0001  , \wishbone_bd_ram_mem1_reg[207][10]/P0001  , \wishbone_bd_ram_mem1_reg[207][11]/P0001  , \wishbone_bd_ram_mem1_reg[207][12]/P0001  , \wishbone_bd_ram_mem1_reg[207][13]/P0001  , \wishbone_bd_ram_mem1_reg[207][14]/P0001  , \wishbone_bd_ram_mem1_reg[207][15]/P0001  , \wishbone_bd_ram_mem1_reg[207][8]/P0001  , \wishbone_bd_ram_mem1_reg[207][9]/P0001  , \wishbone_bd_ram_mem1_reg[208][10]/P0001  , \wishbone_bd_ram_mem1_reg[208][11]/P0001  , \wishbone_bd_ram_mem1_reg[208][12]/P0001  , \wishbone_bd_ram_mem1_reg[208][13]/P0001  , \wishbone_bd_ram_mem1_reg[208][14]/P0001  , \wishbone_bd_ram_mem1_reg[208][15]/P0001  , \wishbone_bd_ram_mem1_reg[208][8]/P0001  , \wishbone_bd_ram_mem1_reg[208][9]/P0001  , \wishbone_bd_ram_mem1_reg[209][10]/P0001  , \wishbone_bd_ram_mem1_reg[209][11]/P0001  , \wishbone_bd_ram_mem1_reg[209][12]/P0001  , \wishbone_bd_ram_mem1_reg[209][13]/P0001  , \wishbone_bd_ram_mem1_reg[209][14]/P0001  , \wishbone_bd_ram_mem1_reg[209][15]/P0001  , \wishbone_bd_ram_mem1_reg[209][8]/P0001  , \wishbone_bd_ram_mem1_reg[209][9]/P0001  , \wishbone_bd_ram_mem1_reg[20][10]/P0001  , \wishbone_bd_ram_mem1_reg[20][11]/P0001  , \wishbone_bd_ram_mem1_reg[20][12]/P0001  , \wishbone_bd_ram_mem1_reg[20][13]/P0001  , \wishbone_bd_ram_mem1_reg[20][14]/P0001  , \wishbone_bd_ram_mem1_reg[20][15]/P0001  , \wishbone_bd_ram_mem1_reg[20][8]/P0001  , \wishbone_bd_ram_mem1_reg[20][9]/P0001  , \wishbone_bd_ram_mem1_reg[210][10]/P0001  , \wishbone_bd_ram_mem1_reg[210][11]/P0001  , \wishbone_bd_ram_mem1_reg[210][12]/P0001  , \wishbone_bd_ram_mem1_reg[210][13]/P0001  , \wishbone_bd_ram_mem1_reg[210][14]/P0001  , \wishbone_bd_ram_mem1_reg[210][15]/P0001  , \wishbone_bd_ram_mem1_reg[210][8]/P0001  , \wishbone_bd_ram_mem1_reg[210][9]/P0001  , \wishbone_bd_ram_mem1_reg[211][10]/P0001  , \wishbone_bd_ram_mem1_reg[211][11]/P0001  , \wishbone_bd_ram_mem1_reg[211][12]/P0001  , \wishbone_bd_ram_mem1_reg[211][13]/P0001  , \wishbone_bd_ram_mem1_reg[211][14]/P0001  , \wishbone_bd_ram_mem1_reg[211][15]/P0001  , \wishbone_bd_ram_mem1_reg[211][8]/P0001  , \wishbone_bd_ram_mem1_reg[211][9]/P0001  , \wishbone_bd_ram_mem1_reg[212][10]/P0001  , \wishbone_bd_ram_mem1_reg[212][11]/P0001  , \wishbone_bd_ram_mem1_reg[212][12]/P0001  , \wishbone_bd_ram_mem1_reg[212][13]/P0001  , \wishbone_bd_ram_mem1_reg[212][14]/P0001  , \wishbone_bd_ram_mem1_reg[212][15]/P0001  , \wishbone_bd_ram_mem1_reg[212][8]/P0001  , \wishbone_bd_ram_mem1_reg[212][9]/P0001  , \wishbone_bd_ram_mem1_reg[213][10]/P0001  , \wishbone_bd_ram_mem1_reg[213][11]/P0001  , \wishbone_bd_ram_mem1_reg[213][12]/P0001  , \wishbone_bd_ram_mem1_reg[213][13]/P0001  , \wishbone_bd_ram_mem1_reg[213][14]/P0001  , \wishbone_bd_ram_mem1_reg[213][15]/P0001  , \wishbone_bd_ram_mem1_reg[213][8]/P0001  , \wishbone_bd_ram_mem1_reg[213][9]/P0001  , \wishbone_bd_ram_mem1_reg[214][10]/P0001  , \wishbone_bd_ram_mem1_reg[214][11]/P0001  , \wishbone_bd_ram_mem1_reg[214][12]/P0001  , \wishbone_bd_ram_mem1_reg[214][13]/P0001  , \wishbone_bd_ram_mem1_reg[214][14]/P0001  , \wishbone_bd_ram_mem1_reg[214][15]/P0001  , \wishbone_bd_ram_mem1_reg[214][8]/P0001  , \wishbone_bd_ram_mem1_reg[214][9]/P0001  , \wishbone_bd_ram_mem1_reg[215][10]/P0001  , \wishbone_bd_ram_mem1_reg[215][11]/P0001  , \wishbone_bd_ram_mem1_reg[215][12]/P0001  , \wishbone_bd_ram_mem1_reg[215][13]/P0001  , \wishbone_bd_ram_mem1_reg[215][14]/P0001  , \wishbone_bd_ram_mem1_reg[215][15]/P0001  , \wishbone_bd_ram_mem1_reg[215][8]/P0001  , \wishbone_bd_ram_mem1_reg[215][9]/P0001  , \wishbone_bd_ram_mem1_reg[216][10]/P0001  , \wishbone_bd_ram_mem1_reg[216][11]/P0001  , \wishbone_bd_ram_mem1_reg[216][12]/P0001  , \wishbone_bd_ram_mem1_reg[216][13]/P0001  , \wishbone_bd_ram_mem1_reg[216][14]/P0001  , \wishbone_bd_ram_mem1_reg[216][15]/P0001  , \wishbone_bd_ram_mem1_reg[216][8]/P0001  , \wishbone_bd_ram_mem1_reg[216][9]/P0001  , \wishbone_bd_ram_mem1_reg[217][10]/P0001  , \wishbone_bd_ram_mem1_reg[217][11]/P0001  , \wishbone_bd_ram_mem1_reg[217][12]/P0001  , \wishbone_bd_ram_mem1_reg[217][13]/P0001  , \wishbone_bd_ram_mem1_reg[217][14]/P0001  , \wishbone_bd_ram_mem1_reg[217][15]/P0001  , \wishbone_bd_ram_mem1_reg[217][8]/P0001  , \wishbone_bd_ram_mem1_reg[217][9]/P0001  , \wishbone_bd_ram_mem1_reg[218][10]/P0001  , \wishbone_bd_ram_mem1_reg[218][11]/P0001  , \wishbone_bd_ram_mem1_reg[218][12]/P0001  , \wishbone_bd_ram_mem1_reg[218][13]/P0001  , \wishbone_bd_ram_mem1_reg[218][14]/P0001  , \wishbone_bd_ram_mem1_reg[218][15]/P0001  , \wishbone_bd_ram_mem1_reg[218][8]/P0001  , \wishbone_bd_ram_mem1_reg[218][9]/P0001  , \wishbone_bd_ram_mem1_reg[219][10]/P0001  , \wishbone_bd_ram_mem1_reg[219][11]/P0001  , \wishbone_bd_ram_mem1_reg[219][12]/P0001  , \wishbone_bd_ram_mem1_reg[219][13]/P0001  , \wishbone_bd_ram_mem1_reg[219][14]/P0001  , \wishbone_bd_ram_mem1_reg[219][15]/P0001  , \wishbone_bd_ram_mem1_reg[219][8]/P0001  , \wishbone_bd_ram_mem1_reg[219][9]/P0001  , \wishbone_bd_ram_mem1_reg[21][10]/P0001  , \wishbone_bd_ram_mem1_reg[21][11]/P0001  , \wishbone_bd_ram_mem1_reg[21][12]/P0001  , \wishbone_bd_ram_mem1_reg[21][13]/P0001  , \wishbone_bd_ram_mem1_reg[21][14]/P0001  , \wishbone_bd_ram_mem1_reg[21][15]/P0001  , \wishbone_bd_ram_mem1_reg[21][8]/P0001  , \wishbone_bd_ram_mem1_reg[21][9]/P0001  , \wishbone_bd_ram_mem1_reg[220][10]/P0001  , \wishbone_bd_ram_mem1_reg[220][11]/P0001  , \wishbone_bd_ram_mem1_reg[220][12]/P0001  , \wishbone_bd_ram_mem1_reg[220][13]/P0001  , \wishbone_bd_ram_mem1_reg[220][14]/P0001  , \wishbone_bd_ram_mem1_reg[220][15]/P0001  , \wishbone_bd_ram_mem1_reg[220][8]/P0001  , \wishbone_bd_ram_mem1_reg[220][9]/P0001  , \wishbone_bd_ram_mem1_reg[221][10]/P0001  , \wishbone_bd_ram_mem1_reg[221][11]/P0001  , \wishbone_bd_ram_mem1_reg[221][12]/P0001  , \wishbone_bd_ram_mem1_reg[221][13]/P0001  , \wishbone_bd_ram_mem1_reg[221][14]/P0001  , \wishbone_bd_ram_mem1_reg[221][15]/P0001  , \wishbone_bd_ram_mem1_reg[221][8]/P0001  , \wishbone_bd_ram_mem1_reg[221][9]/P0001  , \wishbone_bd_ram_mem1_reg[222][10]/P0001  , \wishbone_bd_ram_mem1_reg[222][11]/P0001  , \wishbone_bd_ram_mem1_reg[222][12]/P0001  , \wishbone_bd_ram_mem1_reg[222][13]/P0001  , \wishbone_bd_ram_mem1_reg[222][14]/P0001  , \wishbone_bd_ram_mem1_reg[222][15]/P0001  , \wishbone_bd_ram_mem1_reg[222][8]/P0001  , \wishbone_bd_ram_mem1_reg[222][9]/P0001  , \wishbone_bd_ram_mem1_reg[223][10]/P0001  , \wishbone_bd_ram_mem1_reg[223][11]/P0001  , \wishbone_bd_ram_mem1_reg[223][12]/P0001  , \wishbone_bd_ram_mem1_reg[223][13]/P0001  , \wishbone_bd_ram_mem1_reg[223][14]/P0001  , \wishbone_bd_ram_mem1_reg[223][15]/P0001  , \wishbone_bd_ram_mem1_reg[223][8]/P0001  , \wishbone_bd_ram_mem1_reg[223][9]/P0001  , \wishbone_bd_ram_mem1_reg[224][10]/P0001  , \wishbone_bd_ram_mem1_reg[224][11]/P0001  , \wishbone_bd_ram_mem1_reg[224][12]/P0001  , \wishbone_bd_ram_mem1_reg[224][13]/P0001  , \wishbone_bd_ram_mem1_reg[224][14]/P0001  , \wishbone_bd_ram_mem1_reg[224][15]/P0001  , \wishbone_bd_ram_mem1_reg[224][8]/P0001  , \wishbone_bd_ram_mem1_reg[224][9]/P0001  , \wishbone_bd_ram_mem1_reg[225][10]/P0001  , \wishbone_bd_ram_mem1_reg[225][11]/P0001  , \wishbone_bd_ram_mem1_reg[225][12]/P0001  , \wishbone_bd_ram_mem1_reg[225][13]/P0001  , \wishbone_bd_ram_mem1_reg[225][14]/P0001  , \wishbone_bd_ram_mem1_reg[225][15]/P0001  , \wishbone_bd_ram_mem1_reg[225][8]/P0001  , \wishbone_bd_ram_mem1_reg[225][9]/P0001  , \wishbone_bd_ram_mem1_reg[226][10]/P0001  , \wishbone_bd_ram_mem1_reg[226][11]/P0001  , \wishbone_bd_ram_mem1_reg[226][12]/P0001  , \wishbone_bd_ram_mem1_reg[226][13]/P0001  , \wishbone_bd_ram_mem1_reg[226][14]/P0001  , \wishbone_bd_ram_mem1_reg[226][15]/P0001  , \wishbone_bd_ram_mem1_reg[226][8]/P0001  , \wishbone_bd_ram_mem1_reg[226][9]/P0001  , \wishbone_bd_ram_mem1_reg[227][10]/P0001  , \wishbone_bd_ram_mem1_reg[227][11]/P0001  , \wishbone_bd_ram_mem1_reg[227][12]/P0001  , \wishbone_bd_ram_mem1_reg[227][13]/P0001  , \wishbone_bd_ram_mem1_reg[227][14]/P0001  , \wishbone_bd_ram_mem1_reg[227][15]/P0001  , \wishbone_bd_ram_mem1_reg[227][8]/P0001  , \wishbone_bd_ram_mem1_reg[227][9]/P0001  , \wishbone_bd_ram_mem1_reg[228][10]/P0001  , \wishbone_bd_ram_mem1_reg[228][11]/P0001  , \wishbone_bd_ram_mem1_reg[228][12]/P0001  , \wishbone_bd_ram_mem1_reg[228][13]/P0001  , \wishbone_bd_ram_mem1_reg[228][14]/P0001  , \wishbone_bd_ram_mem1_reg[228][15]/P0001  , \wishbone_bd_ram_mem1_reg[228][8]/P0001  , \wishbone_bd_ram_mem1_reg[228][9]/P0001  , \wishbone_bd_ram_mem1_reg[229][10]/P0001  , \wishbone_bd_ram_mem1_reg[229][11]/P0001  , \wishbone_bd_ram_mem1_reg[229][12]/P0001  , \wishbone_bd_ram_mem1_reg[229][13]/P0001  , \wishbone_bd_ram_mem1_reg[229][14]/P0001  , \wishbone_bd_ram_mem1_reg[229][15]/P0001  , \wishbone_bd_ram_mem1_reg[229][8]/P0001  , \wishbone_bd_ram_mem1_reg[229][9]/P0001  , \wishbone_bd_ram_mem1_reg[22][10]/P0001  , \wishbone_bd_ram_mem1_reg[22][11]/P0001  , \wishbone_bd_ram_mem1_reg[22][12]/P0001  , \wishbone_bd_ram_mem1_reg[22][13]/P0001  , \wishbone_bd_ram_mem1_reg[22][14]/P0001  , \wishbone_bd_ram_mem1_reg[22][15]/P0001  , \wishbone_bd_ram_mem1_reg[22][8]/P0001  , \wishbone_bd_ram_mem1_reg[22][9]/P0001  , \wishbone_bd_ram_mem1_reg[230][10]/P0001  , \wishbone_bd_ram_mem1_reg[230][11]/P0001  , \wishbone_bd_ram_mem1_reg[230][12]/P0001  , \wishbone_bd_ram_mem1_reg[230][13]/P0001  , \wishbone_bd_ram_mem1_reg[230][14]/P0001  , \wishbone_bd_ram_mem1_reg[230][15]/P0001  , \wishbone_bd_ram_mem1_reg[230][8]/P0001  , \wishbone_bd_ram_mem1_reg[230][9]/P0001  , \wishbone_bd_ram_mem1_reg[231][10]/P0001  , \wishbone_bd_ram_mem1_reg[231][11]/P0001  , \wishbone_bd_ram_mem1_reg[231][12]/P0001  , \wishbone_bd_ram_mem1_reg[231][13]/P0001  , \wishbone_bd_ram_mem1_reg[231][14]/P0001  , \wishbone_bd_ram_mem1_reg[231][15]/P0001  , \wishbone_bd_ram_mem1_reg[231][8]/P0001  , \wishbone_bd_ram_mem1_reg[231][9]/P0001  , \wishbone_bd_ram_mem1_reg[232][10]/P0001  , \wishbone_bd_ram_mem1_reg[232][11]/P0001  , \wishbone_bd_ram_mem1_reg[232][12]/P0001  , \wishbone_bd_ram_mem1_reg[232][13]/P0001  , \wishbone_bd_ram_mem1_reg[232][14]/P0001  , \wishbone_bd_ram_mem1_reg[232][15]/P0001  , \wishbone_bd_ram_mem1_reg[232][8]/P0001  , \wishbone_bd_ram_mem1_reg[232][9]/P0001  , \wishbone_bd_ram_mem1_reg[233][10]/P0001  , \wishbone_bd_ram_mem1_reg[233][11]/P0001  , \wishbone_bd_ram_mem1_reg[233][12]/P0001  , \wishbone_bd_ram_mem1_reg[233][13]/P0001  , \wishbone_bd_ram_mem1_reg[233][14]/P0001  , \wishbone_bd_ram_mem1_reg[233][15]/P0001  , \wishbone_bd_ram_mem1_reg[233][8]/P0001  , \wishbone_bd_ram_mem1_reg[233][9]/P0001  , \wishbone_bd_ram_mem1_reg[234][10]/P0001  , \wishbone_bd_ram_mem1_reg[234][11]/P0001  , \wishbone_bd_ram_mem1_reg[234][12]/P0001  , \wishbone_bd_ram_mem1_reg[234][13]/P0001  , \wishbone_bd_ram_mem1_reg[234][14]/P0001  , \wishbone_bd_ram_mem1_reg[234][15]/P0001  , \wishbone_bd_ram_mem1_reg[234][8]/P0001  , \wishbone_bd_ram_mem1_reg[234][9]/P0001  , \wishbone_bd_ram_mem1_reg[235][10]/P0001  , \wishbone_bd_ram_mem1_reg[235][11]/P0001  , \wishbone_bd_ram_mem1_reg[235][12]/P0001  , \wishbone_bd_ram_mem1_reg[235][13]/P0001  , \wishbone_bd_ram_mem1_reg[235][14]/P0001  , \wishbone_bd_ram_mem1_reg[235][15]/P0001  , \wishbone_bd_ram_mem1_reg[235][8]/P0001  , \wishbone_bd_ram_mem1_reg[235][9]/P0001  , \wishbone_bd_ram_mem1_reg[236][10]/P0001  , \wishbone_bd_ram_mem1_reg[236][11]/P0001  , \wishbone_bd_ram_mem1_reg[236][12]/P0001  , \wishbone_bd_ram_mem1_reg[236][13]/P0001  , \wishbone_bd_ram_mem1_reg[236][14]/P0001  , \wishbone_bd_ram_mem1_reg[236][15]/P0001  , \wishbone_bd_ram_mem1_reg[236][8]/P0001  , \wishbone_bd_ram_mem1_reg[236][9]/P0001  , \wishbone_bd_ram_mem1_reg[237][10]/P0001  , \wishbone_bd_ram_mem1_reg[237][11]/P0001  , \wishbone_bd_ram_mem1_reg[237][12]/P0001  , \wishbone_bd_ram_mem1_reg[237][13]/P0001  , \wishbone_bd_ram_mem1_reg[237][14]/P0001  , \wishbone_bd_ram_mem1_reg[237][15]/P0001  , \wishbone_bd_ram_mem1_reg[237][8]/P0001  , \wishbone_bd_ram_mem1_reg[237][9]/P0001  , \wishbone_bd_ram_mem1_reg[238][10]/P0001  , \wishbone_bd_ram_mem1_reg[238][11]/P0001  , \wishbone_bd_ram_mem1_reg[238][12]/P0001  , \wishbone_bd_ram_mem1_reg[238][13]/P0001  , \wishbone_bd_ram_mem1_reg[238][14]/P0001  , \wishbone_bd_ram_mem1_reg[238][15]/P0001  , \wishbone_bd_ram_mem1_reg[238][8]/P0001  , \wishbone_bd_ram_mem1_reg[238][9]/P0001  , \wishbone_bd_ram_mem1_reg[239][10]/P0001  , \wishbone_bd_ram_mem1_reg[239][11]/P0001  , \wishbone_bd_ram_mem1_reg[239][12]/P0001  , \wishbone_bd_ram_mem1_reg[239][13]/P0001  , \wishbone_bd_ram_mem1_reg[239][14]/P0001  , \wishbone_bd_ram_mem1_reg[239][15]/P0001  , \wishbone_bd_ram_mem1_reg[239][8]/P0001  , \wishbone_bd_ram_mem1_reg[239][9]/P0001  , \wishbone_bd_ram_mem1_reg[23][10]/P0001  , \wishbone_bd_ram_mem1_reg[23][11]/P0001  , \wishbone_bd_ram_mem1_reg[23][12]/P0001  , \wishbone_bd_ram_mem1_reg[23][13]/P0001  , \wishbone_bd_ram_mem1_reg[23][14]/P0001  , \wishbone_bd_ram_mem1_reg[23][15]/P0001  , \wishbone_bd_ram_mem1_reg[23][8]/P0001  , \wishbone_bd_ram_mem1_reg[23][9]/P0001  , \wishbone_bd_ram_mem1_reg[240][10]/P0001  , \wishbone_bd_ram_mem1_reg[240][11]/P0001  , \wishbone_bd_ram_mem1_reg[240][12]/P0001  , \wishbone_bd_ram_mem1_reg[240][13]/P0001  , \wishbone_bd_ram_mem1_reg[240][14]/P0001  , \wishbone_bd_ram_mem1_reg[240][15]/P0001  , \wishbone_bd_ram_mem1_reg[240][8]/P0001  , \wishbone_bd_ram_mem1_reg[240][9]/P0001  , \wishbone_bd_ram_mem1_reg[241][10]/P0001  , \wishbone_bd_ram_mem1_reg[241][11]/P0001  , \wishbone_bd_ram_mem1_reg[241][12]/P0001  , \wishbone_bd_ram_mem1_reg[241][13]/P0001  , \wishbone_bd_ram_mem1_reg[241][14]/P0001  , \wishbone_bd_ram_mem1_reg[241][15]/P0001  , \wishbone_bd_ram_mem1_reg[241][8]/P0001  , \wishbone_bd_ram_mem1_reg[241][9]/P0001  , \wishbone_bd_ram_mem1_reg[242][10]/P0001  , \wishbone_bd_ram_mem1_reg[242][11]/P0001  , \wishbone_bd_ram_mem1_reg[242][12]/P0001  , \wishbone_bd_ram_mem1_reg[242][13]/P0001  , \wishbone_bd_ram_mem1_reg[242][14]/P0001  , \wishbone_bd_ram_mem1_reg[242][15]/P0001  , \wishbone_bd_ram_mem1_reg[242][8]/P0001  , \wishbone_bd_ram_mem1_reg[242][9]/P0001  , \wishbone_bd_ram_mem1_reg[243][10]/P0001  , \wishbone_bd_ram_mem1_reg[243][11]/P0001  , \wishbone_bd_ram_mem1_reg[243][12]/P0001  , \wishbone_bd_ram_mem1_reg[243][13]/P0001  , \wishbone_bd_ram_mem1_reg[243][14]/P0001  , \wishbone_bd_ram_mem1_reg[243][15]/P0001  , \wishbone_bd_ram_mem1_reg[243][8]/P0001  , \wishbone_bd_ram_mem1_reg[243][9]/P0001  , \wishbone_bd_ram_mem1_reg[244][10]/P0001  , \wishbone_bd_ram_mem1_reg[244][11]/P0001  , \wishbone_bd_ram_mem1_reg[244][12]/P0001  , \wishbone_bd_ram_mem1_reg[244][13]/P0001  , \wishbone_bd_ram_mem1_reg[244][14]/P0001  , \wishbone_bd_ram_mem1_reg[244][15]/P0001  , \wishbone_bd_ram_mem1_reg[244][8]/P0001  , \wishbone_bd_ram_mem1_reg[244][9]/P0001  , \wishbone_bd_ram_mem1_reg[245][10]/P0001  , \wishbone_bd_ram_mem1_reg[245][11]/P0001  , \wishbone_bd_ram_mem1_reg[245][12]/P0001  , \wishbone_bd_ram_mem1_reg[245][13]/P0001  , \wishbone_bd_ram_mem1_reg[245][14]/P0001  , \wishbone_bd_ram_mem1_reg[245][15]/P0001  , \wishbone_bd_ram_mem1_reg[245][8]/P0001  , \wishbone_bd_ram_mem1_reg[245][9]/P0001  , \wishbone_bd_ram_mem1_reg[246][10]/P0001  , \wishbone_bd_ram_mem1_reg[246][11]/P0001  , \wishbone_bd_ram_mem1_reg[246][12]/P0001  , \wishbone_bd_ram_mem1_reg[246][13]/P0001  , \wishbone_bd_ram_mem1_reg[246][14]/P0001  , \wishbone_bd_ram_mem1_reg[246][15]/P0001  , \wishbone_bd_ram_mem1_reg[246][8]/P0001  , \wishbone_bd_ram_mem1_reg[246][9]/P0001  , \wishbone_bd_ram_mem1_reg[247][10]/P0001  , \wishbone_bd_ram_mem1_reg[247][11]/P0001  , \wishbone_bd_ram_mem1_reg[247][12]/P0001  , \wishbone_bd_ram_mem1_reg[247][13]/P0001  , \wishbone_bd_ram_mem1_reg[247][14]/P0001  , \wishbone_bd_ram_mem1_reg[247][15]/P0001  , \wishbone_bd_ram_mem1_reg[247][8]/P0001  , \wishbone_bd_ram_mem1_reg[247][9]/P0001  , \wishbone_bd_ram_mem1_reg[248][10]/P0001  , \wishbone_bd_ram_mem1_reg[248][11]/P0001  , \wishbone_bd_ram_mem1_reg[248][12]/P0001  , \wishbone_bd_ram_mem1_reg[248][13]/P0001  , \wishbone_bd_ram_mem1_reg[248][14]/P0001  , \wishbone_bd_ram_mem1_reg[248][15]/P0001  , \wishbone_bd_ram_mem1_reg[248][8]/P0001  , \wishbone_bd_ram_mem1_reg[248][9]/P0001  , \wishbone_bd_ram_mem1_reg[249][10]/P0001  , \wishbone_bd_ram_mem1_reg[249][11]/P0001  , \wishbone_bd_ram_mem1_reg[249][12]/P0001  , \wishbone_bd_ram_mem1_reg[249][13]/P0001  , \wishbone_bd_ram_mem1_reg[249][14]/P0001  , \wishbone_bd_ram_mem1_reg[249][15]/P0001  , \wishbone_bd_ram_mem1_reg[249][8]/P0001  , \wishbone_bd_ram_mem1_reg[249][9]/P0001  , \wishbone_bd_ram_mem1_reg[24][10]/P0001  , \wishbone_bd_ram_mem1_reg[24][11]/P0001  , \wishbone_bd_ram_mem1_reg[24][12]/P0001  , \wishbone_bd_ram_mem1_reg[24][13]/P0001  , \wishbone_bd_ram_mem1_reg[24][14]/P0001  , \wishbone_bd_ram_mem1_reg[24][15]/P0001  , \wishbone_bd_ram_mem1_reg[24][8]/P0001  , \wishbone_bd_ram_mem1_reg[24][9]/P0001  , \wishbone_bd_ram_mem1_reg[250][10]/P0001  , \wishbone_bd_ram_mem1_reg[250][11]/P0001  , \wishbone_bd_ram_mem1_reg[250][12]/P0001  , \wishbone_bd_ram_mem1_reg[250][13]/P0001  , \wishbone_bd_ram_mem1_reg[250][14]/P0001  , \wishbone_bd_ram_mem1_reg[250][15]/P0001  , \wishbone_bd_ram_mem1_reg[250][8]/P0001  , \wishbone_bd_ram_mem1_reg[250][9]/P0001  , \wishbone_bd_ram_mem1_reg[251][10]/P0001  , \wishbone_bd_ram_mem1_reg[251][11]/P0001  , \wishbone_bd_ram_mem1_reg[251][12]/P0001  , \wishbone_bd_ram_mem1_reg[251][13]/P0001  , \wishbone_bd_ram_mem1_reg[251][14]/P0001  , \wishbone_bd_ram_mem1_reg[251][15]/P0001  , \wishbone_bd_ram_mem1_reg[251][8]/P0001  , \wishbone_bd_ram_mem1_reg[251][9]/P0001  , \wishbone_bd_ram_mem1_reg[252][10]/P0001  , \wishbone_bd_ram_mem1_reg[252][11]/P0001  , \wishbone_bd_ram_mem1_reg[252][12]/P0001  , \wishbone_bd_ram_mem1_reg[252][13]/P0001  , \wishbone_bd_ram_mem1_reg[252][14]/P0001  , \wishbone_bd_ram_mem1_reg[252][15]/P0001  , \wishbone_bd_ram_mem1_reg[252][8]/P0001  , \wishbone_bd_ram_mem1_reg[252][9]/P0001  , \wishbone_bd_ram_mem1_reg[253][10]/P0001  , \wishbone_bd_ram_mem1_reg[253][11]/P0001  , \wishbone_bd_ram_mem1_reg[253][12]/P0001  , \wishbone_bd_ram_mem1_reg[253][13]/P0001  , \wishbone_bd_ram_mem1_reg[253][14]/P0001  , \wishbone_bd_ram_mem1_reg[253][15]/P0001  , \wishbone_bd_ram_mem1_reg[253][8]/P0001  , \wishbone_bd_ram_mem1_reg[253][9]/P0001  , \wishbone_bd_ram_mem1_reg[254][10]/P0001  , \wishbone_bd_ram_mem1_reg[254][11]/P0001  , \wishbone_bd_ram_mem1_reg[254][12]/P0001  , \wishbone_bd_ram_mem1_reg[254][13]/P0001  , \wishbone_bd_ram_mem1_reg[254][14]/P0001  , \wishbone_bd_ram_mem1_reg[254][15]/P0001  , \wishbone_bd_ram_mem1_reg[254][8]/P0001  , \wishbone_bd_ram_mem1_reg[254][9]/P0001  , \wishbone_bd_ram_mem1_reg[255][10]/P0001  , \wishbone_bd_ram_mem1_reg[255][11]/P0001  , \wishbone_bd_ram_mem1_reg[255][12]/P0001  , \wishbone_bd_ram_mem1_reg[255][13]/P0001  , \wishbone_bd_ram_mem1_reg[255][14]/P0001  , \wishbone_bd_ram_mem1_reg[255][15]/P0001  , \wishbone_bd_ram_mem1_reg[255][8]/P0001  , \wishbone_bd_ram_mem1_reg[255][9]/P0001  , \wishbone_bd_ram_mem1_reg[25][10]/P0001  , \wishbone_bd_ram_mem1_reg[25][11]/P0001  , \wishbone_bd_ram_mem1_reg[25][12]/P0001  , \wishbone_bd_ram_mem1_reg[25][13]/P0001  , \wishbone_bd_ram_mem1_reg[25][14]/P0001  , \wishbone_bd_ram_mem1_reg[25][15]/P0001  , \wishbone_bd_ram_mem1_reg[25][8]/P0001  , \wishbone_bd_ram_mem1_reg[25][9]/P0001  , \wishbone_bd_ram_mem1_reg[26][10]/P0001  , \wishbone_bd_ram_mem1_reg[26][11]/P0001  , \wishbone_bd_ram_mem1_reg[26][12]/P0001  , \wishbone_bd_ram_mem1_reg[26][13]/P0001  , \wishbone_bd_ram_mem1_reg[26][14]/P0001  , \wishbone_bd_ram_mem1_reg[26][15]/P0001  , \wishbone_bd_ram_mem1_reg[26][8]/P0001  , \wishbone_bd_ram_mem1_reg[26][9]/P0001  , \wishbone_bd_ram_mem1_reg[27][10]/P0001  , \wishbone_bd_ram_mem1_reg[27][11]/P0001  , \wishbone_bd_ram_mem1_reg[27][12]/P0001  , \wishbone_bd_ram_mem1_reg[27][13]/P0001  , \wishbone_bd_ram_mem1_reg[27][14]/P0001  , \wishbone_bd_ram_mem1_reg[27][15]/P0001  , \wishbone_bd_ram_mem1_reg[27][8]/P0001  , \wishbone_bd_ram_mem1_reg[27][9]/P0001  , \wishbone_bd_ram_mem1_reg[28][10]/P0001  , \wishbone_bd_ram_mem1_reg[28][11]/P0001  , \wishbone_bd_ram_mem1_reg[28][12]/P0001  , \wishbone_bd_ram_mem1_reg[28][13]/P0001  , \wishbone_bd_ram_mem1_reg[28][14]/P0001  , \wishbone_bd_ram_mem1_reg[28][15]/P0001  , \wishbone_bd_ram_mem1_reg[28][8]/P0001  , \wishbone_bd_ram_mem1_reg[28][9]/P0001  , \wishbone_bd_ram_mem1_reg[29][10]/P0001  , \wishbone_bd_ram_mem1_reg[29][11]/P0001  , \wishbone_bd_ram_mem1_reg[29][12]/P0001  , \wishbone_bd_ram_mem1_reg[29][13]/P0001  , \wishbone_bd_ram_mem1_reg[29][14]/P0001  , \wishbone_bd_ram_mem1_reg[29][15]/P0001  , \wishbone_bd_ram_mem1_reg[29][8]/P0001  , \wishbone_bd_ram_mem1_reg[29][9]/P0001  , \wishbone_bd_ram_mem1_reg[2][10]/P0001  , \wishbone_bd_ram_mem1_reg[2][11]/P0001  , \wishbone_bd_ram_mem1_reg[2][12]/P0001  , \wishbone_bd_ram_mem1_reg[2][13]/P0001  , \wishbone_bd_ram_mem1_reg[2][14]/P0001  , \wishbone_bd_ram_mem1_reg[2][15]/P0001  , \wishbone_bd_ram_mem1_reg[2][8]/P0001  , \wishbone_bd_ram_mem1_reg[2][9]/P0001  , \wishbone_bd_ram_mem1_reg[30][10]/P0001  , \wishbone_bd_ram_mem1_reg[30][11]/P0001  , \wishbone_bd_ram_mem1_reg[30][12]/P0001  , \wishbone_bd_ram_mem1_reg[30][13]/P0001  , \wishbone_bd_ram_mem1_reg[30][14]/P0001  , \wishbone_bd_ram_mem1_reg[30][15]/P0001  , \wishbone_bd_ram_mem1_reg[30][8]/P0001  , \wishbone_bd_ram_mem1_reg[30][9]/P0001  , \wishbone_bd_ram_mem1_reg[31][10]/P0001  , \wishbone_bd_ram_mem1_reg[31][11]/P0001  , \wishbone_bd_ram_mem1_reg[31][12]/P0001  , \wishbone_bd_ram_mem1_reg[31][13]/P0001  , \wishbone_bd_ram_mem1_reg[31][14]/P0001  , \wishbone_bd_ram_mem1_reg[31][15]/P0001  , \wishbone_bd_ram_mem1_reg[31][8]/P0001  , \wishbone_bd_ram_mem1_reg[31][9]/P0001  , \wishbone_bd_ram_mem1_reg[32][10]/P0001  , \wishbone_bd_ram_mem1_reg[32][11]/P0001  , \wishbone_bd_ram_mem1_reg[32][12]/P0001  , \wishbone_bd_ram_mem1_reg[32][13]/P0001  , \wishbone_bd_ram_mem1_reg[32][14]/P0001  , \wishbone_bd_ram_mem1_reg[32][15]/P0001  , \wishbone_bd_ram_mem1_reg[32][8]/P0001  , \wishbone_bd_ram_mem1_reg[32][9]/P0001  , \wishbone_bd_ram_mem1_reg[33][10]/P0001  , \wishbone_bd_ram_mem1_reg[33][11]/P0001  , \wishbone_bd_ram_mem1_reg[33][12]/P0001  , \wishbone_bd_ram_mem1_reg[33][13]/P0001  , \wishbone_bd_ram_mem1_reg[33][14]/P0001  , \wishbone_bd_ram_mem1_reg[33][15]/P0001  , \wishbone_bd_ram_mem1_reg[33][8]/P0001  , \wishbone_bd_ram_mem1_reg[33][9]/P0001  , \wishbone_bd_ram_mem1_reg[34][10]/P0001  , \wishbone_bd_ram_mem1_reg[34][11]/P0001  , \wishbone_bd_ram_mem1_reg[34][12]/P0001  , \wishbone_bd_ram_mem1_reg[34][13]/P0001  , \wishbone_bd_ram_mem1_reg[34][14]/P0001  , \wishbone_bd_ram_mem1_reg[34][15]/P0001  , \wishbone_bd_ram_mem1_reg[34][8]/P0001  , \wishbone_bd_ram_mem1_reg[34][9]/P0001  , \wishbone_bd_ram_mem1_reg[35][10]/P0001  , \wishbone_bd_ram_mem1_reg[35][11]/P0001  , \wishbone_bd_ram_mem1_reg[35][12]/P0001  , \wishbone_bd_ram_mem1_reg[35][13]/P0001  , \wishbone_bd_ram_mem1_reg[35][14]/P0001  , \wishbone_bd_ram_mem1_reg[35][15]/P0001  , \wishbone_bd_ram_mem1_reg[35][8]/P0001  , \wishbone_bd_ram_mem1_reg[35][9]/P0001  , \wishbone_bd_ram_mem1_reg[36][10]/P0001  , \wishbone_bd_ram_mem1_reg[36][11]/P0001  , \wishbone_bd_ram_mem1_reg[36][12]/P0001  , \wishbone_bd_ram_mem1_reg[36][13]/P0001  , \wishbone_bd_ram_mem1_reg[36][14]/P0001  , \wishbone_bd_ram_mem1_reg[36][15]/P0001  , \wishbone_bd_ram_mem1_reg[36][8]/P0001  , \wishbone_bd_ram_mem1_reg[36][9]/P0001  , \wishbone_bd_ram_mem1_reg[37][10]/P0001  , \wishbone_bd_ram_mem1_reg[37][11]/P0001  , \wishbone_bd_ram_mem1_reg[37][12]/P0001  , \wishbone_bd_ram_mem1_reg[37][13]/P0001  , \wishbone_bd_ram_mem1_reg[37][14]/P0001  , \wishbone_bd_ram_mem1_reg[37][15]/P0001  , \wishbone_bd_ram_mem1_reg[37][8]/P0001  , \wishbone_bd_ram_mem1_reg[37][9]/P0001  , \wishbone_bd_ram_mem1_reg[38][10]/P0001  , \wishbone_bd_ram_mem1_reg[38][11]/P0001  , \wishbone_bd_ram_mem1_reg[38][12]/P0001  , \wishbone_bd_ram_mem1_reg[38][13]/P0001  , \wishbone_bd_ram_mem1_reg[38][14]/P0001  , \wishbone_bd_ram_mem1_reg[38][15]/P0001  , \wishbone_bd_ram_mem1_reg[38][8]/P0001  , \wishbone_bd_ram_mem1_reg[38][9]/P0001  , \wishbone_bd_ram_mem1_reg[39][10]/P0001  , \wishbone_bd_ram_mem1_reg[39][11]/P0001  , \wishbone_bd_ram_mem1_reg[39][12]/P0001  , \wishbone_bd_ram_mem1_reg[39][13]/P0001  , \wishbone_bd_ram_mem1_reg[39][14]/P0001  , \wishbone_bd_ram_mem1_reg[39][15]/P0001  , \wishbone_bd_ram_mem1_reg[39][8]/P0001  , \wishbone_bd_ram_mem1_reg[39][9]/P0001  , \wishbone_bd_ram_mem1_reg[3][10]/P0001  , \wishbone_bd_ram_mem1_reg[3][11]/P0001  , \wishbone_bd_ram_mem1_reg[3][12]/P0001  , \wishbone_bd_ram_mem1_reg[3][13]/P0001  , \wishbone_bd_ram_mem1_reg[3][14]/P0001  , \wishbone_bd_ram_mem1_reg[3][15]/P0001  , \wishbone_bd_ram_mem1_reg[3][8]/P0001  , \wishbone_bd_ram_mem1_reg[3][9]/P0001  , \wishbone_bd_ram_mem1_reg[40][10]/P0001  , \wishbone_bd_ram_mem1_reg[40][11]/P0001  , \wishbone_bd_ram_mem1_reg[40][12]/P0001  , \wishbone_bd_ram_mem1_reg[40][13]/P0001  , \wishbone_bd_ram_mem1_reg[40][14]/P0001  , \wishbone_bd_ram_mem1_reg[40][15]/P0001  , \wishbone_bd_ram_mem1_reg[40][8]/P0001  , \wishbone_bd_ram_mem1_reg[40][9]/P0001  , \wishbone_bd_ram_mem1_reg[41][10]/P0001  , \wishbone_bd_ram_mem1_reg[41][11]/P0001  , \wishbone_bd_ram_mem1_reg[41][12]/P0001  , \wishbone_bd_ram_mem1_reg[41][13]/P0001  , \wishbone_bd_ram_mem1_reg[41][14]/P0001  , \wishbone_bd_ram_mem1_reg[41][15]/P0001  , \wishbone_bd_ram_mem1_reg[41][8]/P0001  , \wishbone_bd_ram_mem1_reg[41][9]/P0001  , \wishbone_bd_ram_mem1_reg[42][10]/P0001  , \wishbone_bd_ram_mem1_reg[42][11]/P0001  , \wishbone_bd_ram_mem1_reg[42][12]/P0001  , \wishbone_bd_ram_mem1_reg[42][13]/P0001  , \wishbone_bd_ram_mem1_reg[42][14]/P0001  , \wishbone_bd_ram_mem1_reg[42][15]/P0001  , \wishbone_bd_ram_mem1_reg[42][8]/P0001  , \wishbone_bd_ram_mem1_reg[42][9]/P0001  , \wishbone_bd_ram_mem1_reg[43][10]/P0001  , \wishbone_bd_ram_mem1_reg[43][11]/P0001  , \wishbone_bd_ram_mem1_reg[43][12]/P0001  , \wishbone_bd_ram_mem1_reg[43][13]/P0001  , \wishbone_bd_ram_mem1_reg[43][14]/P0001  , \wishbone_bd_ram_mem1_reg[43][15]/P0001  , \wishbone_bd_ram_mem1_reg[43][8]/P0001  , \wishbone_bd_ram_mem1_reg[43][9]/P0001  , \wishbone_bd_ram_mem1_reg[44][10]/P0001  , \wishbone_bd_ram_mem1_reg[44][11]/P0001  , \wishbone_bd_ram_mem1_reg[44][12]/P0001  , \wishbone_bd_ram_mem1_reg[44][13]/P0001  , \wishbone_bd_ram_mem1_reg[44][14]/P0001  , \wishbone_bd_ram_mem1_reg[44][15]/P0001  , \wishbone_bd_ram_mem1_reg[44][8]/P0001  , \wishbone_bd_ram_mem1_reg[44][9]/P0001  , \wishbone_bd_ram_mem1_reg[45][10]/P0001  , \wishbone_bd_ram_mem1_reg[45][11]/P0001  , \wishbone_bd_ram_mem1_reg[45][12]/P0001  , \wishbone_bd_ram_mem1_reg[45][13]/P0001  , \wishbone_bd_ram_mem1_reg[45][14]/P0001  , \wishbone_bd_ram_mem1_reg[45][15]/P0001  , \wishbone_bd_ram_mem1_reg[45][8]/P0001  , \wishbone_bd_ram_mem1_reg[45][9]/P0001  , \wishbone_bd_ram_mem1_reg[46][10]/P0001  , \wishbone_bd_ram_mem1_reg[46][11]/P0001  , \wishbone_bd_ram_mem1_reg[46][12]/P0001  , \wishbone_bd_ram_mem1_reg[46][13]/P0001  , \wishbone_bd_ram_mem1_reg[46][14]/P0001  , \wishbone_bd_ram_mem1_reg[46][15]/P0001  , \wishbone_bd_ram_mem1_reg[46][8]/P0001  , \wishbone_bd_ram_mem1_reg[46][9]/P0001  , \wishbone_bd_ram_mem1_reg[47][10]/P0001  , \wishbone_bd_ram_mem1_reg[47][11]/P0001  , \wishbone_bd_ram_mem1_reg[47][12]/P0001  , \wishbone_bd_ram_mem1_reg[47][13]/P0001  , \wishbone_bd_ram_mem1_reg[47][14]/P0001  , \wishbone_bd_ram_mem1_reg[47][15]/P0001  , \wishbone_bd_ram_mem1_reg[47][8]/P0001  , \wishbone_bd_ram_mem1_reg[47][9]/P0001  , \wishbone_bd_ram_mem1_reg[48][10]/P0001  , \wishbone_bd_ram_mem1_reg[48][11]/P0001  , \wishbone_bd_ram_mem1_reg[48][12]/P0001  , \wishbone_bd_ram_mem1_reg[48][13]/P0001  , \wishbone_bd_ram_mem1_reg[48][14]/P0001  , \wishbone_bd_ram_mem1_reg[48][15]/P0001  , \wishbone_bd_ram_mem1_reg[48][8]/P0001  , \wishbone_bd_ram_mem1_reg[48][9]/P0001  , \wishbone_bd_ram_mem1_reg[49][10]/P0001  , \wishbone_bd_ram_mem1_reg[49][11]/P0001  , \wishbone_bd_ram_mem1_reg[49][12]/P0001  , \wishbone_bd_ram_mem1_reg[49][13]/P0001  , \wishbone_bd_ram_mem1_reg[49][14]/P0001  , \wishbone_bd_ram_mem1_reg[49][15]/P0001  , \wishbone_bd_ram_mem1_reg[49][8]/P0001  , \wishbone_bd_ram_mem1_reg[49][9]/P0001  , \wishbone_bd_ram_mem1_reg[4][10]/P0001  , \wishbone_bd_ram_mem1_reg[4][11]/P0001  , \wishbone_bd_ram_mem1_reg[4][12]/P0001  , \wishbone_bd_ram_mem1_reg[4][13]/P0001  , \wishbone_bd_ram_mem1_reg[4][14]/P0001  , \wishbone_bd_ram_mem1_reg[4][15]/P0001  , \wishbone_bd_ram_mem1_reg[4][8]/P0001  , \wishbone_bd_ram_mem1_reg[4][9]/P0001  , \wishbone_bd_ram_mem1_reg[50][10]/P0001  , \wishbone_bd_ram_mem1_reg[50][11]/P0001  , \wishbone_bd_ram_mem1_reg[50][12]/P0001  , \wishbone_bd_ram_mem1_reg[50][13]/P0001  , \wishbone_bd_ram_mem1_reg[50][14]/P0001  , \wishbone_bd_ram_mem1_reg[50][15]/P0001  , \wishbone_bd_ram_mem1_reg[50][8]/P0001  , \wishbone_bd_ram_mem1_reg[50][9]/P0001  , \wishbone_bd_ram_mem1_reg[51][10]/P0001  , \wishbone_bd_ram_mem1_reg[51][11]/P0001  , \wishbone_bd_ram_mem1_reg[51][12]/P0001  , \wishbone_bd_ram_mem1_reg[51][13]/P0001  , \wishbone_bd_ram_mem1_reg[51][14]/P0001  , \wishbone_bd_ram_mem1_reg[51][15]/P0001  , \wishbone_bd_ram_mem1_reg[51][8]/P0001  , \wishbone_bd_ram_mem1_reg[51][9]/P0001  , \wishbone_bd_ram_mem1_reg[52][10]/P0001  , \wishbone_bd_ram_mem1_reg[52][11]/P0001  , \wishbone_bd_ram_mem1_reg[52][12]/P0001  , \wishbone_bd_ram_mem1_reg[52][13]/P0001  , \wishbone_bd_ram_mem1_reg[52][14]/P0001  , \wishbone_bd_ram_mem1_reg[52][15]/P0001  , \wishbone_bd_ram_mem1_reg[52][8]/P0001  , \wishbone_bd_ram_mem1_reg[52][9]/P0001  , \wishbone_bd_ram_mem1_reg[53][10]/P0001  , \wishbone_bd_ram_mem1_reg[53][11]/P0001  , \wishbone_bd_ram_mem1_reg[53][12]/P0001  , \wishbone_bd_ram_mem1_reg[53][13]/P0001  , \wishbone_bd_ram_mem1_reg[53][14]/P0001  , \wishbone_bd_ram_mem1_reg[53][15]/P0001  , \wishbone_bd_ram_mem1_reg[53][8]/P0001  , \wishbone_bd_ram_mem1_reg[53][9]/P0001  , \wishbone_bd_ram_mem1_reg[54][10]/P0001  , \wishbone_bd_ram_mem1_reg[54][11]/P0001  , \wishbone_bd_ram_mem1_reg[54][12]/P0001  , \wishbone_bd_ram_mem1_reg[54][13]/P0001  , \wishbone_bd_ram_mem1_reg[54][14]/P0001  , \wishbone_bd_ram_mem1_reg[54][15]/P0001  , \wishbone_bd_ram_mem1_reg[54][8]/P0001  , \wishbone_bd_ram_mem1_reg[54][9]/P0001  , \wishbone_bd_ram_mem1_reg[55][10]/P0001  , \wishbone_bd_ram_mem1_reg[55][11]/P0001  , \wishbone_bd_ram_mem1_reg[55][12]/P0001  , \wishbone_bd_ram_mem1_reg[55][13]/P0001  , \wishbone_bd_ram_mem1_reg[55][14]/P0001  , \wishbone_bd_ram_mem1_reg[55][15]/P0001  , \wishbone_bd_ram_mem1_reg[55][8]/P0001  , \wishbone_bd_ram_mem1_reg[55][9]/P0001  , \wishbone_bd_ram_mem1_reg[56][10]/P0001  , \wishbone_bd_ram_mem1_reg[56][11]/P0001  , \wishbone_bd_ram_mem1_reg[56][12]/P0001  , \wishbone_bd_ram_mem1_reg[56][13]/P0001  , \wishbone_bd_ram_mem1_reg[56][14]/P0001  , \wishbone_bd_ram_mem1_reg[56][15]/P0001  , \wishbone_bd_ram_mem1_reg[56][8]/P0001  , \wishbone_bd_ram_mem1_reg[56][9]/P0001  , \wishbone_bd_ram_mem1_reg[57][10]/P0001  , \wishbone_bd_ram_mem1_reg[57][11]/P0001  , \wishbone_bd_ram_mem1_reg[57][12]/P0001  , \wishbone_bd_ram_mem1_reg[57][13]/P0001  , \wishbone_bd_ram_mem1_reg[57][14]/P0001  , \wishbone_bd_ram_mem1_reg[57][15]/P0001  , \wishbone_bd_ram_mem1_reg[57][8]/P0001  , \wishbone_bd_ram_mem1_reg[57][9]/P0001  , \wishbone_bd_ram_mem1_reg[58][10]/P0001  , \wishbone_bd_ram_mem1_reg[58][11]/P0001  , \wishbone_bd_ram_mem1_reg[58][12]/P0001  , \wishbone_bd_ram_mem1_reg[58][13]/P0001  , \wishbone_bd_ram_mem1_reg[58][14]/P0001  , \wishbone_bd_ram_mem1_reg[58][15]/P0001  , \wishbone_bd_ram_mem1_reg[58][8]/P0001  , \wishbone_bd_ram_mem1_reg[58][9]/P0001  , \wishbone_bd_ram_mem1_reg[59][10]/P0001  , \wishbone_bd_ram_mem1_reg[59][11]/P0001  , \wishbone_bd_ram_mem1_reg[59][12]/P0001  , \wishbone_bd_ram_mem1_reg[59][13]/P0001  , \wishbone_bd_ram_mem1_reg[59][14]/P0001  , \wishbone_bd_ram_mem1_reg[59][15]/P0001  , \wishbone_bd_ram_mem1_reg[59][8]/P0001  , \wishbone_bd_ram_mem1_reg[59][9]/P0001  , \wishbone_bd_ram_mem1_reg[5][10]/P0001  , \wishbone_bd_ram_mem1_reg[5][11]/P0001  , \wishbone_bd_ram_mem1_reg[5][12]/P0001  , \wishbone_bd_ram_mem1_reg[5][13]/P0001  , \wishbone_bd_ram_mem1_reg[5][14]/P0001  , \wishbone_bd_ram_mem1_reg[5][15]/P0001  , \wishbone_bd_ram_mem1_reg[5][8]/P0001  , \wishbone_bd_ram_mem1_reg[5][9]/P0001  , \wishbone_bd_ram_mem1_reg[60][10]/P0001  , \wishbone_bd_ram_mem1_reg[60][11]/P0001  , \wishbone_bd_ram_mem1_reg[60][12]/P0001  , \wishbone_bd_ram_mem1_reg[60][13]/P0001  , \wishbone_bd_ram_mem1_reg[60][14]/P0001  , \wishbone_bd_ram_mem1_reg[60][15]/P0001  , \wishbone_bd_ram_mem1_reg[60][8]/P0001  , \wishbone_bd_ram_mem1_reg[60][9]/P0001  , \wishbone_bd_ram_mem1_reg[61][10]/P0001  , \wishbone_bd_ram_mem1_reg[61][11]/P0001  , \wishbone_bd_ram_mem1_reg[61][12]/P0001  , \wishbone_bd_ram_mem1_reg[61][13]/P0001  , \wishbone_bd_ram_mem1_reg[61][14]/P0001  , \wishbone_bd_ram_mem1_reg[61][15]/P0001  , \wishbone_bd_ram_mem1_reg[61][8]/P0001  , \wishbone_bd_ram_mem1_reg[61][9]/P0001  , \wishbone_bd_ram_mem1_reg[62][10]/P0001  , \wishbone_bd_ram_mem1_reg[62][11]/P0001  , \wishbone_bd_ram_mem1_reg[62][12]/P0001  , \wishbone_bd_ram_mem1_reg[62][13]/P0001  , \wishbone_bd_ram_mem1_reg[62][14]/P0001  , \wishbone_bd_ram_mem1_reg[62][15]/P0001  , \wishbone_bd_ram_mem1_reg[62][8]/P0001  , \wishbone_bd_ram_mem1_reg[62][9]/P0001  , \wishbone_bd_ram_mem1_reg[63][10]/P0001  , \wishbone_bd_ram_mem1_reg[63][11]/P0001  , \wishbone_bd_ram_mem1_reg[63][12]/P0001  , \wishbone_bd_ram_mem1_reg[63][13]/P0001  , \wishbone_bd_ram_mem1_reg[63][14]/P0001  , \wishbone_bd_ram_mem1_reg[63][15]/P0001  , \wishbone_bd_ram_mem1_reg[63][8]/P0001  , \wishbone_bd_ram_mem1_reg[63][9]/P0001  , \wishbone_bd_ram_mem1_reg[64][10]/P0001  , \wishbone_bd_ram_mem1_reg[64][11]/P0001  , \wishbone_bd_ram_mem1_reg[64][12]/P0001  , \wishbone_bd_ram_mem1_reg[64][13]/P0001  , \wishbone_bd_ram_mem1_reg[64][14]/P0001  , \wishbone_bd_ram_mem1_reg[64][15]/P0001  , \wishbone_bd_ram_mem1_reg[64][8]/P0001  , \wishbone_bd_ram_mem1_reg[64][9]/P0001  , \wishbone_bd_ram_mem1_reg[65][10]/P0001  , \wishbone_bd_ram_mem1_reg[65][11]/P0001  , \wishbone_bd_ram_mem1_reg[65][12]/P0001  , \wishbone_bd_ram_mem1_reg[65][13]/P0001  , \wishbone_bd_ram_mem1_reg[65][14]/P0001  , \wishbone_bd_ram_mem1_reg[65][15]/P0001  , \wishbone_bd_ram_mem1_reg[65][8]/P0001  , \wishbone_bd_ram_mem1_reg[65][9]/P0001  , \wishbone_bd_ram_mem1_reg[66][10]/P0001  , \wishbone_bd_ram_mem1_reg[66][11]/P0001  , \wishbone_bd_ram_mem1_reg[66][12]/P0001  , \wishbone_bd_ram_mem1_reg[66][13]/P0001  , \wishbone_bd_ram_mem1_reg[66][14]/P0001  , \wishbone_bd_ram_mem1_reg[66][15]/P0001  , \wishbone_bd_ram_mem1_reg[66][8]/P0001  , \wishbone_bd_ram_mem1_reg[66][9]/P0001  , \wishbone_bd_ram_mem1_reg[67][10]/P0001  , \wishbone_bd_ram_mem1_reg[67][11]/P0001  , \wishbone_bd_ram_mem1_reg[67][12]/P0001  , \wishbone_bd_ram_mem1_reg[67][13]/P0001  , \wishbone_bd_ram_mem1_reg[67][14]/P0001  , \wishbone_bd_ram_mem1_reg[67][15]/P0001  , \wishbone_bd_ram_mem1_reg[67][8]/P0001  , \wishbone_bd_ram_mem1_reg[67][9]/P0001  , \wishbone_bd_ram_mem1_reg[68][10]/P0001  , \wishbone_bd_ram_mem1_reg[68][11]/P0001  , \wishbone_bd_ram_mem1_reg[68][12]/P0001  , \wishbone_bd_ram_mem1_reg[68][13]/P0001  , \wishbone_bd_ram_mem1_reg[68][14]/P0001  , \wishbone_bd_ram_mem1_reg[68][15]/P0001  , \wishbone_bd_ram_mem1_reg[68][8]/P0001  , \wishbone_bd_ram_mem1_reg[68][9]/P0001  , \wishbone_bd_ram_mem1_reg[69][10]/P0001  , \wishbone_bd_ram_mem1_reg[69][11]/P0001  , \wishbone_bd_ram_mem1_reg[69][12]/P0001  , \wishbone_bd_ram_mem1_reg[69][13]/P0001  , \wishbone_bd_ram_mem1_reg[69][14]/P0001  , \wishbone_bd_ram_mem1_reg[69][15]/P0001  , \wishbone_bd_ram_mem1_reg[69][8]/P0001  , \wishbone_bd_ram_mem1_reg[69][9]/P0001  , \wishbone_bd_ram_mem1_reg[6][10]/P0001  , \wishbone_bd_ram_mem1_reg[6][11]/P0001  , \wishbone_bd_ram_mem1_reg[6][12]/P0001  , \wishbone_bd_ram_mem1_reg[6][13]/P0001  , \wishbone_bd_ram_mem1_reg[6][14]/P0001  , \wishbone_bd_ram_mem1_reg[6][15]/P0001  , \wishbone_bd_ram_mem1_reg[6][8]/P0001  , \wishbone_bd_ram_mem1_reg[6][9]/P0001  , \wishbone_bd_ram_mem1_reg[70][10]/P0001  , \wishbone_bd_ram_mem1_reg[70][11]/P0001  , \wishbone_bd_ram_mem1_reg[70][12]/P0001  , \wishbone_bd_ram_mem1_reg[70][13]/P0001  , \wishbone_bd_ram_mem1_reg[70][14]/P0001  , \wishbone_bd_ram_mem1_reg[70][15]/P0001  , \wishbone_bd_ram_mem1_reg[70][8]/P0001  , \wishbone_bd_ram_mem1_reg[70][9]/P0001  , \wishbone_bd_ram_mem1_reg[71][10]/P0001  , \wishbone_bd_ram_mem1_reg[71][11]/P0001  , \wishbone_bd_ram_mem1_reg[71][12]/P0001  , \wishbone_bd_ram_mem1_reg[71][13]/P0001  , \wishbone_bd_ram_mem1_reg[71][14]/P0001  , \wishbone_bd_ram_mem1_reg[71][15]/P0001  , \wishbone_bd_ram_mem1_reg[71][8]/P0001  , \wishbone_bd_ram_mem1_reg[71][9]/P0001  , \wishbone_bd_ram_mem1_reg[72][10]/P0001  , \wishbone_bd_ram_mem1_reg[72][11]/P0001  , \wishbone_bd_ram_mem1_reg[72][12]/P0001  , \wishbone_bd_ram_mem1_reg[72][13]/P0001  , \wishbone_bd_ram_mem1_reg[72][14]/P0001  , \wishbone_bd_ram_mem1_reg[72][15]/P0001  , \wishbone_bd_ram_mem1_reg[72][8]/P0001  , \wishbone_bd_ram_mem1_reg[72][9]/P0001  , \wishbone_bd_ram_mem1_reg[73][10]/P0001  , \wishbone_bd_ram_mem1_reg[73][11]/P0001  , \wishbone_bd_ram_mem1_reg[73][12]/P0001  , \wishbone_bd_ram_mem1_reg[73][13]/P0001  , \wishbone_bd_ram_mem1_reg[73][14]/P0001  , \wishbone_bd_ram_mem1_reg[73][15]/P0001  , \wishbone_bd_ram_mem1_reg[73][8]/P0001  , \wishbone_bd_ram_mem1_reg[73][9]/P0001  , \wishbone_bd_ram_mem1_reg[74][10]/P0001  , \wishbone_bd_ram_mem1_reg[74][11]/P0001  , \wishbone_bd_ram_mem1_reg[74][12]/P0001  , \wishbone_bd_ram_mem1_reg[74][13]/P0001  , \wishbone_bd_ram_mem1_reg[74][14]/P0001  , \wishbone_bd_ram_mem1_reg[74][15]/P0001  , \wishbone_bd_ram_mem1_reg[74][8]/P0001  , \wishbone_bd_ram_mem1_reg[74][9]/P0001  , \wishbone_bd_ram_mem1_reg[75][10]/P0001  , \wishbone_bd_ram_mem1_reg[75][11]/P0001  , \wishbone_bd_ram_mem1_reg[75][12]/P0001  , \wishbone_bd_ram_mem1_reg[75][13]/P0001  , \wishbone_bd_ram_mem1_reg[75][14]/P0001  , \wishbone_bd_ram_mem1_reg[75][15]/P0001  , \wishbone_bd_ram_mem1_reg[75][8]/P0001  , \wishbone_bd_ram_mem1_reg[75][9]/P0001  , \wishbone_bd_ram_mem1_reg[76][10]/P0001  , \wishbone_bd_ram_mem1_reg[76][11]/P0001  , \wishbone_bd_ram_mem1_reg[76][12]/P0001  , \wishbone_bd_ram_mem1_reg[76][13]/P0001  , \wishbone_bd_ram_mem1_reg[76][14]/P0001  , \wishbone_bd_ram_mem1_reg[76][15]/P0001  , \wishbone_bd_ram_mem1_reg[76][8]/P0001  , \wishbone_bd_ram_mem1_reg[76][9]/P0001  , \wishbone_bd_ram_mem1_reg[77][10]/P0001  , \wishbone_bd_ram_mem1_reg[77][11]/P0001  , \wishbone_bd_ram_mem1_reg[77][12]/P0001  , \wishbone_bd_ram_mem1_reg[77][13]/P0001  , \wishbone_bd_ram_mem1_reg[77][14]/P0001  , \wishbone_bd_ram_mem1_reg[77][15]/P0001  , \wishbone_bd_ram_mem1_reg[77][8]/P0001  , \wishbone_bd_ram_mem1_reg[77][9]/P0001  , \wishbone_bd_ram_mem1_reg[78][10]/P0001  , \wishbone_bd_ram_mem1_reg[78][11]/P0001  , \wishbone_bd_ram_mem1_reg[78][12]/P0001  , \wishbone_bd_ram_mem1_reg[78][13]/P0001  , \wishbone_bd_ram_mem1_reg[78][14]/P0001  , \wishbone_bd_ram_mem1_reg[78][15]/P0001  , \wishbone_bd_ram_mem1_reg[78][8]/P0001  , \wishbone_bd_ram_mem1_reg[78][9]/P0001  , \wishbone_bd_ram_mem1_reg[79][10]/P0001  , \wishbone_bd_ram_mem1_reg[79][11]/P0001  , \wishbone_bd_ram_mem1_reg[79][12]/P0001  , \wishbone_bd_ram_mem1_reg[79][13]/P0001  , \wishbone_bd_ram_mem1_reg[79][14]/P0001  , \wishbone_bd_ram_mem1_reg[79][15]/P0001  , \wishbone_bd_ram_mem1_reg[79][8]/P0001  , \wishbone_bd_ram_mem1_reg[79][9]/P0001  , \wishbone_bd_ram_mem1_reg[7][10]/P0001  , \wishbone_bd_ram_mem1_reg[7][11]/P0001  , \wishbone_bd_ram_mem1_reg[7][12]/P0001  , \wishbone_bd_ram_mem1_reg[7][13]/P0001  , \wishbone_bd_ram_mem1_reg[7][14]/P0001  , \wishbone_bd_ram_mem1_reg[7][15]/P0001  , \wishbone_bd_ram_mem1_reg[7][8]/P0001  , \wishbone_bd_ram_mem1_reg[7][9]/P0001  , \wishbone_bd_ram_mem1_reg[80][10]/P0001  , \wishbone_bd_ram_mem1_reg[80][11]/P0001  , \wishbone_bd_ram_mem1_reg[80][12]/P0001  , \wishbone_bd_ram_mem1_reg[80][13]/P0001  , \wishbone_bd_ram_mem1_reg[80][14]/P0001  , \wishbone_bd_ram_mem1_reg[80][15]/P0001  , \wishbone_bd_ram_mem1_reg[80][8]/P0001  , \wishbone_bd_ram_mem1_reg[80][9]/P0001  , \wishbone_bd_ram_mem1_reg[81][10]/P0001  , \wishbone_bd_ram_mem1_reg[81][11]/P0001  , \wishbone_bd_ram_mem1_reg[81][12]/P0001  , \wishbone_bd_ram_mem1_reg[81][13]/P0001  , \wishbone_bd_ram_mem1_reg[81][14]/P0001  , \wishbone_bd_ram_mem1_reg[81][15]/P0001  , \wishbone_bd_ram_mem1_reg[81][8]/P0001  , \wishbone_bd_ram_mem1_reg[81][9]/P0001  , \wishbone_bd_ram_mem1_reg[82][10]/P0001  , \wishbone_bd_ram_mem1_reg[82][11]/P0001  , \wishbone_bd_ram_mem1_reg[82][12]/P0001  , \wishbone_bd_ram_mem1_reg[82][13]/P0001  , \wishbone_bd_ram_mem1_reg[82][14]/P0001  , \wishbone_bd_ram_mem1_reg[82][15]/P0001  , \wishbone_bd_ram_mem1_reg[82][8]/P0001  , \wishbone_bd_ram_mem1_reg[82][9]/P0001  , \wishbone_bd_ram_mem1_reg[83][10]/P0001  , \wishbone_bd_ram_mem1_reg[83][11]/P0001  , \wishbone_bd_ram_mem1_reg[83][12]/P0001  , \wishbone_bd_ram_mem1_reg[83][13]/P0001  , \wishbone_bd_ram_mem1_reg[83][14]/P0001  , \wishbone_bd_ram_mem1_reg[83][15]/P0001  , \wishbone_bd_ram_mem1_reg[83][8]/P0001  , \wishbone_bd_ram_mem1_reg[83][9]/P0001  , \wishbone_bd_ram_mem1_reg[84][10]/P0001  , \wishbone_bd_ram_mem1_reg[84][11]/P0001  , \wishbone_bd_ram_mem1_reg[84][12]/P0001  , \wishbone_bd_ram_mem1_reg[84][13]/P0001  , \wishbone_bd_ram_mem1_reg[84][14]/P0001  , \wishbone_bd_ram_mem1_reg[84][15]/P0001  , \wishbone_bd_ram_mem1_reg[84][8]/P0001  , \wishbone_bd_ram_mem1_reg[84][9]/P0001  , \wishbone_bd_ram_mem1_reg[85][10]/P0001  , \wishbone_bd_ram_mem1_reg[85][11]/P0001  , \wishbone_bd_ram_mem1_reg[85][12]/P0001  , \wishbone_bd_ram_mem1_reg[85][13]/P0001  , \wishbone_bd_ram_mem1_reg[85][14]/P0001  , \wishbone_bd_ram_mem1_reg[85][15]/P0001  , \wishbone_bd_ram_mem1_reg[85][8]/P0001  , \wishbone_bd_ram_mem1_reg[85][9]/P0001  , \wishbone_bd_ram_mem1_reg[86][10]/P0001  , \wishbone_bd_ram_mem1_reg[86][11]/P0001  , \wishbone_bd_ram_mem1_reg[86][12]/P0001  , \wishbone_bd_ram_mem1_reg[86][13]/P0001  , \wishbone_bd_ram_mem1_reg[86][14]/P0001  , \wishbone_bd_ram_mem1_reg[86][15]/P0001  , \wishbone_bd_ram_mem1_reg[86][8]/P0001  , \wishbone_bd_ram_mem1_reg[86][9]/P0001  , \wishbone_bd_ram_mem1_reg[87][10]/P0001  , \wishbone_bd_ram_mem1_reg[87][11]/P0001  , \wishbone_bd_ram_mem1_reg[87][12]/P0001  , \wishbone_bd_ram_mem1_reg[87][13]/P0001  , \wishbone_bd_ram_mem1_reg[87][14]/P0001  , \wishbone_bd_ram_mem1_reg[87][15]/P0001  , \wishbone_bd_ram_mem1_reg[87][8]/P0001  , \wishbone_bd_ram_mem1_reg[87][9]/P0001  , \wishbone_bd_ram_mem1_reg[88][10]/P0001  , \wishbone_bd_ram_mem1_reg[88][11]/P0001  , \wishbone_bd_ram_mem1_reg[88][12]/P0001  , \wishbone_bd_ram_mem1_reg[88][13]/P0001  , \wishbone_bd_ram_mem1_reg[88][14]/P0001  , \wishbone_bd_ram_mem1_reg[88][15]/P0001  , \wishbone_bd_ram_mem1_reg[88][8]/P0001  , \wishbone_bd_ram_mem1_reg[88][9]/P0001  , \wishbone_bd_ram_mem1_reg[89][10]/P0001  , \wishbone_bd_ram_mem1_reg[89][11]/P0001  , \wishbone_bd_ram_mem1_reg[89][12]/P0001  , \wishbone_bd_ram_mem1_reg[89][13]/P0001  , \wishbone_bd_ram_mem1_reg[89][14]/P0001  , \wishbone_bd_ram_mem1_reg[89][15]/P0001  , \wishbone_bd_ram_mem1_reg[89][8]/P0001  , \wishbone_bd_ram_mem1_reg[89][9]/P0001  , \wishbone_bd_ram_mem1_reg[8][10]/P0001  , \wishbone_bd_ram_mem1_reg[8][11]/P0001  , \wishbone_bd_ram_mem1_reg[8][12]/P0001  , \wishbone_bd_ram_mem1_reg[8][13]/P0001  , \wishbone_bd_ram_mem1_reg[8][14]/P0001  , \wishbone_bd_ram_mem1_reg[8][15]/P0001  , \wishbone_bd_ram_mem1_reg[8][8]/P0001  , \wishbone_bd_ram_mem1_reg[8][9]/P0001  , \wishbone_bd_ram_mem1_reg[90][10]/P0001  , \wishbone_bd_ram_mem1_reg[90][11]/P0001  , \wishbone_bd_ram_mem1_reg[90][12]/P0001  , \wishbone_bd_ram_mem1_reg[90][13]/P0001  , \wishbone_bd_ram_mem1_reg[90][14]/P0001  , \wishbone_bd_ram_mem1_reg[90][15]/P0001  , \wishbone_bd_ram_mem1_reg[90][8]/P0001  , \wishbone_bd_ram_mem1_reg[90][9]/P0001  , \wishbone_bd_ram_mem1_reg[91][10]/P0001  , \wishbone_bd_ram_mem1_reg[91][11]/P0001  , \wishbone_bd_ram_mem1_reg[91][12]/P0001  , \wishbone_bd_ram_mem1_reg[91][13]/P0001  , \wishbone_bd_ram_mem1_reg[91][14]/P0001  , \wishbone_bd_ram_mem1_reg[91][15]/P0001  , \wishbone_bd_ram_mem1_reg[91][8]/P0001  , \wishbone_bd_ram_mem1_reg[91][9]/P0001  , \wishbone_bd_ram_mem1_reg[92][10]/P0001  , \wishbone_bd_ram_mem1_reg[92][11]/P0001  , \wishbone_bd_ram_mem1_reg[92][12]/P0001  , \wishbone_bd_ram_mem1_reg[92][13]/P0001  , \wishbone_bd_ram_mem1_reg[92][14]/P0001  , \wishbone_bd_ram_mem1_reg[92][15]/P0001  , \wishbone_bd_ram_mem1_reg[92][8]/P0001  , \wishbone_bd_ram_mem1_reg[92][9]/P0001  , \wishbone_bd_ram_mem1_reg[93][10]/P0001  , \wishbone_bd_ram_mem1_reg[93][11]/P0001  , \wishbone_bd_ram_mem1_reg[93][12]/P0001  , \wishbone_bd_ram_mem1_reg[93][13]/P0001  , \wishbone_bd_ram_mem1_reg[93][14]/P0001  , \wishbone_bd_ram_mem1_reg[93][15]/P0001  , \wishbone_bd_ram_mem1_reg[93][8]/P0001  , \wishbone_bd_ram_mem1_reg[93][9]/P0001  , \wishbone_bd_ram_mem1_reg[94][10]/P0001  , \wishbone_bd_ram_mem1_reg[94][11]/P0001  , \wishbone_bd_ram_mem1_reg[94][12]/P0001  , \wishbone_bd_ram_mem1_reg[94][13]/P0001  , \wishbone_bd_ram_mem1_reg[94][14]/P0001  , \wishbone_bd_ram_mem1_reg[94][15]/P0001  , \wishbone_bd_ram_mem1_reg[94][8]/P0001  , \wishbone_bd_ram_mem1_reg[94][9]/P0001  , \wishbone_bd_ram_mem1_reg[95][10]/P0001  , \wishbone_bd_ram_mem1_reg[95][11]/P0001  , \wishbone_bd_ram_mem1_reg[95][12]/P0001  , \wishbone_bd_ram_mem1_reg[95][13]/P0001  , \wishbone_bd_ram_mem1_reg[95][14]/P0001  , \wishbone_bd_ram_mem1_reg[95][15]/P0001  , \wishbone_bd_ram_mem1_reg[95][8]/P0001  , \wishbone_bd_ram_mem1_reg[95][9]/P0001  , \wishbone_bd_ram_mem1_reg[96][10]/P0001  , \wishbone_bd_ram_mem1_reg[96][11]/P0001  , \wishbone_bd_ram_mem1_reg[96][12]/P0001  , \wishbone_bd_ram_mem1_reg[96][13]/P0001  , \wishbone_bd_ram_mem1_reg[96][14]/P0001  , \wishbone_bd_ram_mem1_reg[96][15]/P0001  , \wishbone_bd_ram_mem1_reg[96][8]/P0001  , \wishbone_bd_ram_mem1_reg[96][9]/P0001  , \wishbone_bd_ram_mem1_reg[97][10]/P0001  , \wishbone_bd_ram_mem1_reg[97][11]/P0001  , \wishbone_bd_ram_mem1_reg[97][12]/P0001  , \wishbone_bd_ram_mem1_reg[97][13]/P0001  , \wishbone_bd_ram_mem1_reg[97][14]/P0001  , \wishbone_bd_ram_mem1_reg[97][15]/P0001  , \wishbone_bd_ram_mem1_reg[97][8]/P0001  , \wishbone_bd_ram_mem1_reg[97][9]/P0001  , \wishbone_bd_ram_mem1_reg[98][10]/P0001  , \wishbone_bd_ram_mem1_reg[98][11]/P0001  , \wishbone_bd_ram_mem1_reg[98][12]/P0001  , \wishbone_bd_ram_mem1_reg[98][13]/P0001  , \wishbone_bd_ram_mem1_reg[98][14]/P0001  , \wishbone_bd_ram_mem1_reg[98][15]/P0001  , \wishbone_bd_ram_mem1_reg[98][8]/P0001  , \wishbone_bd_ram_mem1_reg[98][9]/P0001  , \wishbone_bd_ram_mem1_reg[99][10]/P0001  , \wishbone_bd_ram_mem1_reg[99][11]/P0001  , \wishbone_bd_ram_mem1_reg[99][12]/P0001  , \wishbone_bd_ram_mem1_reg[99][13]/P0001  , \wishbone_bd_ram_mem1_reg[99][14]/P0001  , \wishbone_bd_ram_mem1_reg[99][15]/P0001  , \wishbone_bd_ram_mem1_reg[99][8]/P0001  , \wishbone_bd_ram_mem1_reg[99][9]/P0001  , \wishbone_bd_ram_mem1_reg[9][10]/P0001  , \wishbone_bd_ram_mem1_reg[9][11]/P0001  , \wishbone_bd_ram_mem1_reg[9][12]/P0001  , \wishbone_bd_ram_mem1_reg[9][13]/P0001  , \wishbone_bd_ram_mem1_reg[9][14]/P0001  , \wishbone_bd_ram_mem1_reg[9][15]/P0001  , \wishbone_bd_ram_mem1_reg[9][8]/P0001  , \wishbone_bd_ram_mem1_reg[9][9]/P0001  , \wishbone_bd_ram_mem2_reg[0][16]/P0001  , \wishbone_bd_ram_mem2_reg[0][17]/P0001  , \wishbone_bd_ram_mem2_reg[0][18]/P0001  , \wishbone_bd_ram_mem2_reg[0][19]/P0001  , \wishbone_bd_ram_mem2_reg[0][20]/P0001  , \wishbone_bd_ram_mem2_reg[0][21]/P0001  , \wishbone_bd_ram_mem2_reg[0][22]/P0001  , \wishbone_bd_ram_mem2_reg[0][23]/P0001  , \wishbone_bd_ram_mem2_reg[100][16]/P0001  , \wishbone_bd_ram_mem2_reg[100][17]/P0001  , \wishbone_bd_ram_mem2_reg[100][18]/P0001  , \wishbone_bd_ram_mem2_reg[100][19]/P0001  , \wishbone_bd_ram_mem2_reg[100][20]/P0001  , \wishbone_bd_ram_mem2_reg[100][21]/P0001  , \wishbone_bd_ram_mem2_reg[100][22]/P0001  , \wishbone_bd_ram_mem2_reg[100][23]/P0001  , \wishbone_bd_ram_mem2_reg[101][16]/P0001  , \wishbone_bd_ram_mem2_reg[101][17]/P0001  , \wishbone_bd_ram_mem2_reg[101][18]/P0001  , \wishbone_bd_ram_mem2_reg[101][19]/P0001  , \wishbone_bd_ram_mem2_reg[101][20]/P0001  , \wishbone_bd_ram_mem2_reg[101][21]/P0001  , \wishbone_bd_ram_mem2_reg[101][22]/P0001  , \wishbone_bd_ram_mem2_reg[101][23]/P0001  , \wishbone_bd_ram_mem2_reg[102][16]/P0001  , \wishbone_bd_ram_mem2_reg[102][17]/P0001  , \wishbone_bd_ram_mem2_reg[102][18]/P0001  , \wishbone_bd_ram_mem2_reg[102][19]/P0001  , \wishbone_bd_ram_mem2_reg[102][20]/P0001  , \wishbone_bd_ram_mem2_reg[102][21]/P0001  , \wishbone_bd_ram_mem2_reg[102][22]/P0001  , \wishbone_bd_ram_mem2_reg[102][23]/P0001  , \wishbone_bd_ram_mem2_reg[103][16]/P0001  , \wishbone_bd_ram_mem2_reg[103][17]/P0001  , \wishbone_bd_ram_mem2_reg[103][18]/P0001  , \wishbone_bd_ram_mem2_reg[103][19]/P0001  , \wishbone_bd_ram_mem2_reg[103][20]/P0001  , \wishbone_bd_ram_mem2_reg[103][21]/P0001  , \wishbone_bd_ram_mem2_reg[103][22]/P0001  , \wishbone_bd_ram_mem2_reg[103][23]/P0001  , \wishbone_bd_ram_mem2_reg[104][16]/P0001  , \wishbone_bd_ram_mem2_reg[104][17]/P0001  , \wishbone_bd_ram_mem2_reg[104][18]/P0001  , \wishbone_bd_ram_mem2_reg[104][19]/P0001  , \wishbone_bd_ram_mem2_reg[104][20]/P0001  , \wishbone_bd_ram_mem2_reg[104][21]/P0001  , \wishbone_bd_ram_mem2_reg[104][22]/P0001  , \wishbone_bd_ram_mem2_reg[104][23]/P0001  , \wishbone_bd_ram_mem2_reg[105][16]/P0001  , \wishbone_bd_ram_mem2_reg[105][17]/P0001  , \wishbone_bd_ram_mem2_reg[105][18]/P0001  , \wishbone_bd_ram_mem2_reg[105][19]/P0001  , \wishbone_bd_ram_mem2_reg[105][20]/P0001  , \wishbone_bd_ram_mem2_reg[105][21]/P0001  , \wishbone_bd_ram_mem2_reg[105][22]/P0001  , \wishbone_bd_ram_mem2_reg[105][23]/P0001  , \wishbone_bd_ram_mem2_reg[106][16]/P0001  , \wishbone_bd_ram_mem2_reg[106][17]/P0001  , \wishbone_bd_ram_mem2_reg[106][18]/P0001  , \wishbone_bd_ram_mem2_reg[106][19]/P0001  , \wishbone_bd_ram_mem2_reg[106][20]/P0001  , \wishbone_bd_ram_mem2_reg[106][21]/P0001  , \wishbone_bd_ram_mem2_reg[106][22]/P0001  , \wishbone_bd_ram_mem2_reg[106][23]/P0001  , \wishbone_bd_ram_mem2_reg[107][16]/P0001  , \wishbone_bd_ram_mem2_reg[107][17]/P0001  , \wishbone_bd_ram_mem2_reg[107][18]/P0001  , \wishbone_bd_ram_mem2_reg[107][19]/P0001  , \wishbone_bd_ram_mem2_reg[107][20]/P0001  , \wishbone_bd_ram_mem2_reg[107][21]/P0001  , \wishbone_bd_ram_mem2_reg[107][22]/P0001  , \wishbone_bd_ram_mem2_reg[107][23]/P0001  , \wishbone_bd_ram_mem2_reg[108][16]/P0001  , \wishbone_bd_ram_mem2_reg[108][17]/P0001  , \wishbone_bd_ram_mem2_reg[108][18]/P0001  , \wishbone_bd_ram_mem2_reg[108][19]/P0001  , \wishbone_bd_ram_mem2_reg[108][20]/P0001  , \wishbone_bd_ram_mem2_reg[108][21]/P0001  , \wishbone_bd_ram_mem2_reg[108][22]/P0001  , \wishbone_bd_ram_mem2_reg[108][23]/P0001  , \wishbone_bd_ram_mem2_reg[109][16]/P0001  , \wishbone_bd_ram_mem2_reg[109][17]/P0001  , \wishbone_bd_ram_mem2_reg[109][18]/P0001  , \wishbone_bd_ram_mem2_reg[109][19]/P0001  , \wishbone_bd_ram_mem2_reg[109][20]/P0001  , \wishbone_bd_ram_mem2_reg[109][21]/P0001  , \wishbone_bd_ram_mem2_reg[109][22]/P0001  , \wishbone_bd_ram_mem2_reg[109][23]/P0001  , \wishbone_bd_ram_mem2_reg[10][16]/P0001  , \wishbone_bd_ram_mem2_reg[10][17]/P0001  , \wishbone_bd_ram_mem2_reg[10][18]/P0001  , \wishbone_bd_ram_mem2_reg[10][19]/P0001  , \wishbone_bd_ram_mem2_reg[10][20]/P0001  , \wishbone_bd_ram_mem2_reg[10][21]/P0001  , \wishbone_bd_ram_mem2_reg[10][22]/P0001  , \wishbone_bd_ram_mem2_reg[10][23]/P0001  , \wishbone_bd_ram_mem2_reg[110][16]/P0001  , \wishbone_bd_ram_mem2_reg[110][17]/P0001  , \wishbone_bd_ram_mem2_reg[110][18]/P0001  , \wishbone_bd_ram_mem2_reg[110][19]/P0001  , \wishbone_bd_ram_mem2_reg[110][20]/P0001  , \wishbone_bd_ram_mem2_reg[110][21]/P0001  , \wishbone_bd_ram_mem2_reg[110][22]/P0001  , \wishbone_bd_ram_mem2_reg[110][23]/P0001  , \wishbone_bd_ram_mem2_reg[111][16]/P0001  , \wishbone_bd_ram_mem2_reg[111][17]/P0001  , \wishbone_bd_ram_mem2_reg[111][18]/P0001  , \wishbone_bd_ram_mem2_reg[111][19]/P0001  , \wishbone_bd_ram_mem2_reg[111][20]/P0001  , \wishbone_bd_ram_mem2_reg[111][21]/P0001  , \wishbone_bd_ram_mem2_reg[111][22]/P0001  , \wishbone_bd_ram_mem2_reg[111][23]/P0001  , \wishbone_bd_ram_mem2_reg[112][16]/P0001  , \wishbone_bd_ram_mem2_reg[112][17]/P0001  , \wishbone_bd_ram_mem2_reg[112][18]/P0001  , \wishbone_bd_ram_mem2_reg[112][19]/P0001  , \wishbone_bd_ram_mem2_reg[112][20]/P0001  , \wishbone_bd_ram_mem2_reg[112][21]/P0001  , \wishbone_bd_ram_mem2_reg[112][22]/P0001  , \wishbone_bd_ram_mem2_reg[112][23]/P0001  , \wishbone_bd_ram_mem2_reg[113][16]/P0001  , \wishbone_bd_ram_mem2_reg[113][17]/P0001  , \wishbone_bd_ram_mem2_reg[113][18]/P0001  , \wishbone_bd_ram_mem2_reg[113][19]/P0001  , \wishbone_bd_ram_mem2_reg[113][20]/P0001  , \wishbone_bd_ram_mem2_reg[113][21]/P0001  , \wishbone_bd_ram_mem2_reg[113][22]/P0001  , \wishbone_bd_ram_mem2_reg[113][23]/P0001  , \wishbone_bd_ram_mem2_reg[114][16]/P0001  , \wishbone_bd_ram_mem2_reg[114][17]/P0001  , \wishbone_bd_ram_mem2_reg[114][18]/P0001  , \wishbone_bd_ram_mem2_reg[114][19]/P0001  , \wishbone_bd_ram_mem2_reg[114][20]/P0001  , \wishbone_bd_ram_mem2_reg[114][21]/P0001  , \wishbone_bd_ram_mem2_reg[114][22]/P0001  , \wishbone_bd_ram_mem2_reg[114][23]/P0001  , \wishbone_bd_ram_mem2_reg[115][16]/P0001  , \wishbone_bd_ram_mem2_reg[115][17]/P0001  , \wishbone_bd_ram_mem2_reg[115][18]/P0001  , \wishbone_bd_ram_mem2_reg[115][19]/P0001  , \wishbone_bd_ram_mem2_reg[115][20]/P0001  , \wishbone_bd_ram_mem2_reg[115][21]/P0001  , \wishbone_bd_ram_mem2_reg[115][22]/P0001  , \wishbone_bd_ram_mem2_reg[115][23]/P0001  , \wishbone_bd_ram_mem2_reg[116][16]/P0001  , \wishbone_bd_ram_mem2_reg[116][17]/P0001  , \wishbone_bd_ram_mem2_reg[116][18]/P0001  , \wishbone_bd_ram_mem2_reg[116][19]/P0001  , \wishbone_bd_ram_mem2_reg[116][20]/P0001  , \wishbone_bd_ram_mem2_reg[116][21]/P0001  , \wishbone_bd_ram_mem2_reg[116][22]/P0001  , \wishbone_bd_ram_mem2_reg[116][23]/P0001  , \wishbone_bd_ram_mem2_reg[117][16]/P0001  , \wishbone_bd_ram_mem2_reg[117][17]/P0001  , \wishbone_bd_ram_mem2_reg[117][18]/P0001  , \wishbone_bd_ram_mem2_reg[117][19]/P0001  , \wishbone_bd_ram_mem2_reg[117][20]/P0001  , \wishbone_bd_ram_mem2_reg[117][21]/P0001  , \wishbone_bd_ram_mem2_reg[117][22]/P0001  , \wishbone_bd_ram_mem2_reg[117][23]/P0001  , \wishbone_bd_ram_mem2_reg[118][16]/P0001  , \wishbone_bd_ram_mem2_reg[118][17]/P0001  , \wishbone_bd_ram_mem2_reg[118][18]/P0001  , \wishbone_bd_ram_mem2_reg[118][19]/P0001  , \wishbone_bd_ram_mem2_reg[118][20]/P0001  , \wishbone_bd_ram_mem2_reg[118][21]/P0001  , \wishbone_bd_ram_mem2_reg[118][22]/P0001  , \wishbone_bd_ram_mem2_reg[118][23]/P0001  , \wishbone_bd_ram_mem2_reg[119][16]/P0001  , \wishbone_bd_ram_mem2_reg[119][17]/P0001  , \wishbone_bd_ram_mem2_reg[119][18]/P0001  , \wishbone_bd_ram_mem2_reg[119][19]/P0001  , \wishbone_bd_ram_mem2_reg[119][20]/P0001  , \wishbone_bd_ram_mem2_reg[119][21]/P0001  , \wishbone_bd_ram_mem2_reg[119][22]/P0001  , \wishbone_bd_ram_mem2_reg[119][23]/P0001  , \wishbone_bd_ram_mem2_reg[11][16]/P0001  , \wishbone_bd_ram_mem2_reg[11][17]/P0001  , \wishbone_bd_ram_mem2_reg[11][18]/P0001  , \wishbone_bd_ram_mem2_reg[11][19]/P0001  , \wishbone_bd_ram_mem2_reg[11][20]/P0001  , \wishbone_bd_ram_mem2_reg[11][21]/P0001  , \wishbone_bd_ram_mem2_reg[11][22]/P0001  , \wishbone_bd_ram_mem2_reg[11][23]/P0001  , \wishbone_bd_ram_mem2_reg[120][16]/P0001  , \wishbone_bd_ram_mem2_reg[120][17]/P0001  , \wishbone_bd_ram_mem2_reg[120][18]/P0001  , \wishbone_bd_ram_mem2_reg[120][19]/P0001  , \wishbone_bd_ram_mem2_reg[120][20]/P0001  , \wishbone_bd_ram_mem2_reg[120][21]/P0001  , \wishbone_bd_ram_mem2_reg[120][22]/P0001  , \wishbone_bd_ram_mem2_reg[120][23]/P0001  , \wishbone_bd_ram_mem2_reg[121][16]/P0001  , \wishbone_bd_ram_mem2_reg[121][17]/P0001  , \wishbone_bd_ram_mem2_reg[121][18]/P0001  , \wishbone_bd_ram_mem2_reg[121][19]/P0001  , \wishbone_bd_ram_mem2_reg[121][20]/P0001  , \wishbone_bd_ram_mem2_reg[121][21]/P0001  , \wishbone_bd_ram_mem2_reg[121][22]/P0001  , \wishbone_bd_ram_mem2_reg[121][23]/P0001  , \wishbone_bd_ram_mem2_reg[122][16]/P0001  , \wishbone_bd_ram_mem2_reg[122][17]/P0001  , \wishbone_bd_ram_mem2_reg[122][18]/P0001  , \wishbone_bd_ram_mem2_reg[122][19]/P0001  , \wishbone_bd_ram_mem2_reg[122][20]/P0001  , \wishbone_bd_ram_mem2_reg[122][21]/P0001  , \wishbone_bd_ram_mem2_reg[122][22]/P0001  , \wishbone_bd_ram_mem2_reg[122][23]/P0001  , \wishbone_bd_ram_mem2_reg[123][16]/P0001  , \wishbone_bd_ram_mem2_reg[123][17]/P0001  , \wishbone_bd_ram_mem2_reg[123][18]/P0001  , \wishbone_bd_ram_mem2_reg[123][19]/P0001  , \wishbone_bd_ram_mem2_reg[123][20]/P0001  , \wishbone_bd_ram_mem2_reg[123][21]/P0001  , \wishbone_bd_ram_mem2_reg[123][22]/P0001  , \wishbone_bd_ram_mem2_reg[123][23]/P0001  , \wishbone_bd_ram_mem2_reg[124][16]/P0001  , \wishbone_bd_ram_mem2_reg[124][17]/P0001  , \wishbone_bd_ram_mem2_reg[124][18]/P0001  , \wishbone_bd_ram_mem2_reg[124][19]/P0001  , \wishbone_bd_ram_mem2_reg[124][20]/P0001  , \wishbone_bd_ram_mem2_reg[124][21]/P0001  , \wishbone_bd_ram_mem2_reg[124][22]/P0001  , \wishbone_bd_ram_mem2_reg[124][23]/P0001  , \wishbone_bd_ram_mem2_reg[125][16]/P0001  , \wishbone_bd_ram_mem2_reg[125][17]/P0001  , \wishbone_bd_ram_mem2_reg[125][18]/P0001  , \wishbone_bd_ram_mem2_reg[125][19]/P0001  , \wishbone_bd_ram_mem2_reg[125][20]/P0001  , \wishbone_bd_ram_mem2_reg[125][21]/P0001  , \wishbone_bd_ram_mem2_reg[125][22]/P0001  , \wishbone_bd_ram_mem2_reg[125][23]/P0001  , \wishbone_bd_ram_mem2_reg[126][16]/P0001  , \wishbone_bd_ram_mem2_reg[126][17]/P0001  , \wishbone_bd_ram_mem2_reg[126][18]/P0001  , \wishbone_bd_ram_mem2_reg[126][19]/P0001  , \wishbone_bd_ram_mem2_reg[126][20]/P0001  , \wishbone_bd_ram_mem2_reg[126][21]/P0001  , \wishbone_bd_ram_mem2_reg[126][22]/P0001  , \wishbone_bd_ram_mem2_reg[126][23]/P0001  , \wishbone_bd_ram_mem2_reg[127][16]/P0001  , \wishbone_bd_ram_mem2_reg[127][17]/P0001  , \wishbone_bd_ram_mem2_reg[127][18]/P0001  , \wishbone_bd_ram_mem2_reg[127][19]/P0001  , \wishbone_bd_ram_mem2_reg[127][20]/P0001  , \wishbone_bd_ram_mem2_reg[127][21]/P0001  , \wishbone_bd_ram_mem2_reg[127][22]/P0001  , \wishbone_bd_ram_mem2_reg[127][23]/P0001  , \wishbone_bd_ram_mem2_reg[128][16]/P0001  , \wishbone_bd_ram_mem2_reg[128][17]/P0001  , \wishbone_bd_ram_mem2_reg[128][18]/P0001  , \wishbone_bd_ram_mem2_reg[128][19]/P0001  , \wishbone_bd_ram_mem2_reg[128][20]/P0001  , \wishbone_bd_ram_mem2_reg[128][21]/P0001  , \wishbone_bd_ram_mem2_reg[128][22]/P0001  , \wishbone_bd_ram_mem2_reg[128][23]/P0001  , \wishbone_bd_ram_mem2_reg[129][16]/P0001  , \wishbone_bd_ram_mem2_reg[129][17]/P0001  , \wishbone_bd_ram_mem2_reg[129][18]/P0001  , \wishbone_bd_ram_mem2_reg[129][19]/P0001  , \wishbone_bd_ram_mem2_reg[129][20]/P0001  , \wishbone_bd_ram_mem2_reg[129][21]/P0001  , \wishbone_bd_ram_mem2_reg[129][22]/P0001  , \wishbone_bd_ram_mem2_reg[129][23]/P0001  , \wishbone_bd_ram_mem2_reg[12][16]/P0001  , \wishbone_bd_ram_mem2_reg[12][17]/P0001  , \wishbone_bd_ram_mem2_reg[12][18]/P0001  , \wishbone_bd_ram_mem2_reg[12][19]/P0001  , \wishbone_bd_ram_mem2_reg[12][20]/P0001  , \wishbone_bd_ram_mem2_reg[12][21]/P0001  , \wishbone_bd_ram_mem2_reg[12][22]/P0001  , \wishbone_bd_ram_mem2_reg[12][23]/P0001  , \wishbone_bd_ram_mem2_reg[130][16]/P0001  , \wishbone_bd_ram_mem2_reg[130][17]/P0001  , \wishbone_bd_ram_mem2_reg[130][18]/P0001  , \wishbone_bd_ram_mem2_reg[130][19]/P0001  , \wishbone_bd_ram_mem2_reg[130][20]/P0001  , \wishbone_bd_ram_mem2_reg[130][21]/P0001  , \wishbone_bd_ram_mem2_reg[130][22]/P0001  , \wishbone_bd_ram_mem2_reg[130][23]/P0001  , \wishbone_bd_ram_mem2_reg[131][16]/P0001  , \wishbone_bd_ram_mem2_reg[131][17]/P0001  , \wishbone_bd_ram_mem2_reg[131][18]/P0001  , \wishbone_bd_ram_mem2_reg[131][19]/P0001  , \wishbone_bd_ram_mem2_reg[131][20]/P0001  , \wishbone_bd_ram_mem2_reg[131][21]/P0001  , \wishbone_bd_ram_mem2_reg[131][22]/P0001  , \wishbone_bd_ram_mem2_reg[131][23]/P0001  , \wishbone_bd_ram_mem2_reg[132][16]/P0001  , \wishbone_bd_ram_mem2_reg[132][17]/P0001  , \wishbone_bd_ram_mem2_reg[132][18]/P0001  , \wishbone_bd_ram_mem2_reg[132][19]/P0001  , \wishbone_bd_ram_mem2_reg[132][20]/P0001  , \wishbone_bd_ram_mem2_reg[132][21]/P0001  , \wishbone_bd_ram_mem2_reg[132][22]/P0001  , \wishbone_bd_ram_mem2_reg[132][23]/P0001  , \wishbone_bd_ram_mem2_reg[133][16]/P0001  , \wishbone_bd_ram_mem2_reg[133][17]/P0001  , \wishbone_bd_ram_mem2_reg[133][18]/P0001  , \wishbone_bd_ram_mem2_reg[133][19]/P0001  , \wishbone_bd_ram_mem2_reg[133][20]/P0001  , \wishbone_bd_ram_mem2_reg[133][21]/P0001  , \wishbone_bd_ram_mem2_reg[133][22]/P0001  , \wishbone_bd_ram_mem2_reg[133][23]/P0001  , \wishbone_bd_ram_mem2_reg[134][16]/P0001  , \wishbone_bd_ram_mem2_reg[134][17]/P0001  , \wishbone_bd_ram_mem2_reg[134][18]/P0001  , \wishbone_bd_ram_mem2_reg[134][19]/P0001  , \wishbone_bd_ram_mem2_reg[134][20]/P0001  , \wishbone_bd_ram_mem2_reg[134][21]/P0001  , \wishbone_bd_ram_mem2_reg[134][22]/P0001  , \wishbone_bd_ram_mem2_reg[134][23]/P0001  , \wishbone_bd_ram_mem2_reg[135][16]/P0001  , \wishbone_bd_ram_mem2_reg[135][17]/P0001  , \wishbone_bd_ram_mem2_reg[135][18]/P0001  , \wishbone_bd_ram_mem2_reg[135][19]/P0001  , \wishbone_bd_ram_mem2_reg[135][20]/P0001  , \wishbone_bd_ram_mem2_reg[135][21]/P0001  , \wishbone_bd_ram_mem2_reg[135][22]/P0001  , \wishbone_bd_ram_mem2_reg[135][23]/P0001  , \wishbone_bd_ram_mem2_reg[136][16]/P0001  , \wishbone_bd_ram_mem2_reg[136][17]/P0001  , \wishbone_bd_ram_mem2_reg[136][18]/P0001  , \wishbone_bd_ram_mem2_reg[136][19]/P0001  , \wishbone_bd_ram_mem2_reg[136][20]/P0001  , \wishbone_bd_ram_mem2_reg[136][21]/P0001  , \wishbone_bd_ram_mem2_reg[136][22]/P0001  , \wishbone_bd_ram_mem2_reg[136][23]/P0001  , \wishbone_bd_ram_mem2_reg[137][16]/P0001  , \wishbone_bd_ram_mem2_reg[137][17]/P0001  , \wishbone_bd_ram_mem2_reg[137][18]/P0001  , \wishbone_bd_ram_mem2_reg[137][19]/P0001  , \wishbone_bd_ram_mem2_reg[137][20]/P0001  , \wishbone_bd_ram_mem2_reg[137][21]/P0001  , \wishbone_bd_ram_mem2_reg[137][22]/P0001  , \wishbone_bd_ram_mem2_reg[137][23]/P0001  , \wishbone_bd_ram_mem2_reg[138][16]/P0001  , \wishbone_bd_ram_mem2_reg[138][17]/P0001  , \wishbone_bd_ram_mem2_reg[138][18]/P0001  , \wishbone_bd_ram_mem2_reg[138][19]/P0001  , \wishbone_bd_ram_mem2_reg[138][20]/P0001  , \wishbone_bd_ram_mem2_reg[138][21]/P0001  , \wishbone_bd_ram_mem2_reg[138][22]/P0001  , \wishbone_bd_ram_mem2_reg[138][23]/P0001  , \wishbone_bd_ram_mem2_reg[139][16]/P0001  , \wishbone_bd_ram_mem2_reg[139][17]/P0001  , \wishbone_bd_ram_mem2_reg[139][18]/P0001  , \wishbone_bd_ram_mem2_reg[139][19]/P0001  , \wishbone_bd_ram_mem2_reg[139][20]/P0001  , \wishbone_bd_ram_mem2_reg[139][21]/P0001  , \wishbone_bd_ram_mem2_reg[139][22]/P0001  , \wishbone_bd_ram_mem2_reg[139][23]/P0001  , \wishbone_bd_ram_mem2_reg[13][16]/P0001  , \wishbone_bd_ram_mem2_reg[13][17]/P0001  , \wishbone_bd_ram_mem2_reg[13][18]/P0001  , \wishbone_bd_ram_mem2_reg[13][19]/P0001  , \wishbone_bd_ram_mem2_reg[13][20]/P0001  , \wishbone_bd_ram_mem2_reg[13][21]/P0001  , \wishbone_bd_ram_mem2_reg[13][22]/P0001  , \wishbone_bd_ram_mem2_reg[13][23]/P0001  , \wishbone_bd_ram_mem2_reg[140][16]/P0001  , \wishbone_bd_ram_mem2_reg[140][17]/P0001  , \wishbone_bd_ram_mem2_reg[140][18]/P0001  , \wishbone_bd_ram_mem2_reg[140][19]/P0001  , \wishbone_bd_ram_mem2_reg[140][20]/P0001  , \wishbone_bd_ram_mem2_reg[140][21]/P0001  , \wishbone_bd_ram_mem2_reg[140][22]/P0001  , \wishbone_bd_ram_mem2_reg[140][23]/P0001  , \wishbone_bd_ram_mem2_reg[141][16]/P0001  , \wishbone_bd_ram_mem2_reg[141][17]/P0001  , \wishbone_bd_ram_mem2_reg[141][18]/P0001  , \wishbone_bd_ram_mem2_reg[141][19]/P0001  , \wishbone_bd_ram_mem2_reg[141][20]/P0001  , \wishbone_bd_ram_mem2_reg[141][21]/P0001  , \wishbone_bd_ram_mem2_reg[141][22]/P0001  , \wishbone_bd_ram_mem2_reg[141][23]/P0001  , \wishbone_bd_ram_mem2_reg[142][16]/P0001  , \wishbone_bd_ram_mem2_reg[142][17]/P0001  , \wishbone_bd_ram_mem2_reg[142][18]/P0001  , \wishbone_bd_ram_mem2_reg[142][19]/P0001  , \wishbone_bd_ram_mem2_reg[142][20]/P0001  , \wishbone_bd_ram_mem2_reg[142][21]/P0001  , \wishbone_bd_ram_mem2_reg[142][22]/P0001  , \wishbone_bd_ram_mem2_reg[142][23]/P0001  , \wishbone_bd_ram_mem2_reg[143][16]/P0001  , \wishbone_bd_ram_mem2_reg[143][17]/P0001  , \wishbone_bd_ram_mem2_reg[143][18]/P0001  , \wishbone_bd_ram_mem2_reg[143][19]/P0001  , \wishbone_bd_ram_mem2_reg[143][20]/P0001  , \wishbone_bd_ram_mem2_reg[143][21]/P0001  , \wishbone_bd_ram_mem2_reg[143][22]/P0001  , \wishbone_bd_ram_mem2_reg[143][23]/P0001  , \wishbone_bd_ram_mem2_reg[144][16]/P0001  , \wishbone_bd_ram_mem2_reg[144][17]/P0001  , \wishbone_bd_ram_mem2_reg[144][18]/P0001  , \wishbone_bd_ram_mem2_reg[144][19]/P0001  , \wishbone_bd_ram_mem2_reg[144][20]/P0001  , \wishbone_bd_ram_mem2_reg[144][21]/P0001  , \wishbone_bd_ram_mem2_reg[144][22]/P0001  , \wishbone_bd_ram_mem2_reg[144][23]/P0001  , \wishbone_bd_ram_mem2_reg[145][16]/P0001  , \wishbone_bd_ram_mem2_reg[145][17]/P0001  , \wishbone_bd_ram_mem2_reg[145][18]/P0001  , \wishbone_bd_ram_mem2_reg[145][19]/P0001  , \wishbone_bd_ram_mem2_reg[145][20]/P0001  , \wishbone_bd_ram_mem2_reg[145][21]/P0001  , \wishbone_bd_ram_mem2_reg[145][22]/P0001  , \wishbone_bd_ram_mem2_reg[145][23]/P0001  , \wishbone_bd_ram_mem2_reg[146][16]/P0001  , \wishbone_bd_ram_mem2_reg[146][17]/P0001  , \wishbone_bd_ram_mem2_reg[146][18]/P0001  , \wishbone_bd_ram_mem2_reg[146][19]/P0001  , \wishbone_bd_ram_mem2_reg[146][20]/P0001  , \wishbone_bd_ram_mem2_reg[146][21]/P0001  , \wishbone_bd_ram_mem2_reg[146][22]/P0001  , \wishbone_bd_ram_mem2_reg[146][23]/P0001  , \wishbone_bd_ram_mem2_reg[147][16]/P0001  , \wishbone_bd_ram_mem2_reg[147][17]/P0001  , \wishbone_bd_ram_mem2_reg[147][18]/P0001  , \wishbone_bd_ram_mem2_reg[147][19]/P0001  , \wishbone_bd_ram_mem2_reg[147][20]/P0001  , \wishbone_bd_ram_mem2_reg[147][21]/P0001  , \wishbone_bd_ram_mem2_reg[147][22]/P0001  , \wishbone_bd_ram_mem2_reg[147][23]/P0001  , \wishbone_bd_ram_mem2_reg[148][16]/P0001  , \wishbone_bd_ram_mem2_reg[148][17]/P0001  , \wishbone_bd_ram_mem2_reg[148][18]/P0001  , \wishbone_bd_ram_mem2_reg[148][19]/P0001  , \wishbone_bd_ram_mem2_reg[148][20]/P0001  , \wishbone_bd_ram_mem2_reg[148][21]/P0001  , \wishbone_bd_ram_mem2_reg[148][22]/P0001  , \wishbone_bd_ram_mem2_reg[148][23]/P0001  , \wishbone_bd_ram_mem2_reg[149][16]/P0001  , \wishbone_bd_ram_mem2_reg[149][17]/P0001  , \wishbone_bd_ram_mem2_reg[149][18]/P0001  , \wishbone_bd_ram_mem2_reg[149][19]/P0001  , \wishbone_bd_ram_mem2_reg[149][20]/P0001  , \wishbone_bd_ram_mem2_reg[149][21]/P0001  , \wishbone_bd_ram_mem2_reg[149][22]/P0001  , \wishbone_bd_ram_mem2_reg[149][23]/P0001  , \wishbone_bd_ram_mem2_reg[14][16]/P0001  , \wishbone_bd_ram_mem2_reg[14][17]/P0001  , \wishbone_bd_ram_mem2_reg[14][18]/P0001  , \wishbone_bd_ram_mem2_reg[14][19]/P0001  , \wishbone_bd_ram_mem2_reg[14][20]/P0001  , \wishbone_bd_ram_mem2_reg[14][21]/P0001  , \wishbone_bd_ram_mem2_reg[14][22]/P0001  , \wishbone_bd_ram_mem2_reg[14][23]/P0001  , \wishbone_bd_ram_mem2_reg[150][16]/P0001  , \wishbone_bd_ram_mem2_reg[150][17]/P0001  , \wishbone_bd_ram_mem2_reg[150][18]/P0001  , \wishbone_bd_ram_mem2_reg[150][19]/P0001  , \wishbone_bd_ram_mem2_reg[150][20]/P0001  , \wishbone_bd_ram_mem2_reg[150][21]/P0001  , \wishbone_bd_ram_mem2_reg[150][22]/P0001  , \wishbone_bd_ram_mem2_reg[150][23]/P0001  , \wishbone_bd_ram_mem2_reg[151][16]/P0001  , \wishbone_bd_ram_mem2_reg[151][17]/P0001  , \wishbone_bd_ram_mem2_reg[151][18]/P0001  , \wishbone_bd_ram_mem2_reg[151][19]/P0001  , \wishbone_bd_ram_mem2_reg[151][20]/P0001  , \wishbone_bd_ram_mem2_reg[151][21]/P0001  , \wishbone_bd_ram_mem2_reg[151][22]/P0001  , \wishbone_bd_ram_mem2_reg[151][23]/P0001  , \wishbone_bd_ram_mem2_reg[152][16]/P0001  , \wishbone_bd_ram_mem2_reg[152][17]/P0001  , \wishbone_bd_ram_mem2_reg[152][18]/P0001  , \wishbone_bd_ram_mem2_reg[152][19]/P0001  , \wishbone_bd_ram_mem2_reg[152][20]/P0001  , \wishbone_bd_ram_mem2_reg[152][21]/P0001  , \wishbone_bd_ram_mem2_reg[152][22]/P0001  , \wishbone_bd_ram_mem2_reg[152][23]/P0001  , \wishbone_bd_ram_mem2_reg[153][16]/P0001  , \wishbone_bd_ram_mem2_reg[153][17]/P0001  , \wishbone_bd_ram_mem2_reg[153][18]/P0001  , \wishbone_bd_ram_mem2_reg[153][19]/P0001  , \wishbone_bd_ram_mem2_reg[153][20]/P0001  , \wishbone_bd_ram_mem2_reg[153][21]/P0001  , \wishbone_bd_ram_mem2_reg[153][22]/P0001  , \wishbone_bd_ram_mem2_reg[153][23]/P0001  , \wishbone_bd_ram_mem2_reg[154][16]/P0001  , \wishbone_bd_ram_mem2_reg[154][17]/P0001  , \wishbone_bd_ram_mem2_reg[154][18]/P0001  , \wishbone_bd_ram_mem2_reg[154][19]/P0001  , \wishbone_bd_ram_mem2_reg[154][20]/P0001  , \wishbone_bd_ram_mem2_reg[154][21]/P0001  , \wishbone_bd_ram_mem2_reg[154][22]/P0001  , \wishbone_bd_ram_mem2_reg[154][23]/P0001  , \wishbone_bd_ram_mem2_reg[155][16]/P0001  , \wishbone_bd_ram_mem2_reg[155][17]/P0001  , \wishbone_bd_ram_mem2_reg[155][18]/P0001  , \wishbone_bd_ram_mem2_reg[155][19]/P0001  , \wishbone_bd_ram_mem2_reg[155][20]/P0001  , \wishbone_bd_ram_mem2_reg[155][21]/P0001  , \wishbone_bd_ram_mem2_reg[155][22]/P0001  , \wishbone_bd_ram_mem2_reg[155][23]/P0001  , \wishbone_bd_ram_mem2_reg[156][16]/P0001  , \wishbone_bd_ram_mem2_reg[156][17]/P0001  , \wishbone_bd_ram_mem2_reg[156][18]/P0001  , \wishbone_bd_ram_mem2_reg[156][19]/P0001  , \wishbone_bd_ram_mem2_reg[156][20]/P0001  , \wishbone_bd_ram_mem2_reg[156][21]/P0001  , \wishbone_bd_ram_mem2_reg[156][22]/P0001  , \wishbone_bd_ram_mem2_reg[156][23]/P0001  , \wishbone_bd_ram_mem2_reg[157][16]/P0001  , \wishbone_bd_ram_mem2_reg[157][17]/P0001  , \wishbone_bd_ram_mem2_reg[157][18]/P0001  , \wishbone_bd_ram_mem2_reg[157][19]/P0001  , \wishbone_bd_ram_mem2_reg[157][20]/P0001  , \wishbone_bd_ram_mem2_reg[157][21]/P0001  , \wishbone_bd_ram_mem2_reg[157][22]/P0001  , \wishbone_bd_ram_mem2_reg[157][23]/P0001  , \wishbone_bd_ram_mem2_reg[158][16]/P0001  , \wishbone_bd_ram_mem2_reg[158][17]/P0001  , \wishbone_bd_ram_mem2_reg[158][18]/P0001  , \wishbone_bd_ram_mem2_reg[158][19]/P0001  , \wishbone_bd_ram_mem2_reg[158][20]/P0001  , \wishbone_bd_ram_mem2_reg[158][21]/P0001  , \wishbone_bd_ram_mem2_reg[158][22]/P0001  , \wishbone_bd_ram_mem2_reg[158][23]/P0001  , \wishbone_bd_ram_mem2_reg[159][16]/P0001  , \wishbone_bd_ram_mem2_reg[159][17]/P0001  , \wishbone_bd_ram_mem2_reg[159][18]/P0001  , \wishbone_bd_ram_mem2_reg[159][19]/P0001  , \wishbone_bd_ram_mem2_reg[159][20]/P0001  , \wishbone_bd_ram_mem2_reg[159][21]/P0001  , \wishbone_bd_ram_mem2_reg[159][22]/P0001  , \wishbone_bd_ram_mem2_reg[159][23]/P0001  , \wishbone_bd_ram_mem2_reg[15][16]/P0001  , \wishbone_bd_ram_mem2_reg[15][17]/P0001  , \wishbone_bd_ram_mem2_reg[15][18]/P0001  , \wishbone_bd_ram_mem2_reg[15][19]/P0001  , \wishbone_bd_ram_mem2_reg[15][20]/P0001  , \wishbone_bd_ram_mem2_reg[15][21]/P0001  , \wishbone_bd_ram_mem2_reg[15][22]/P0001  , \wishbone_bd_ram_mem2_reg[15][23]/P0001  , \wishbone_bd_ram_mem2_reg[160][16]/P0001  , \wishbone_bd_ram_mem2_reg[160][17]/P0001  , \wishbone_bd_ram_mem2_reg[160][18]/P0001  , \wishbone_bd_ram_mem2_reg[160][19]/P0001  , \wishbone_bd_ram_mem2_reg[160][20]/P0001  , \wishbone_bd_ram_mem2_reg[160][21]/P0001  , \wishbone_bd_ram_mem2_reg[160][22]/P0001  , \wishbone_bd_ram_mem2_reg[160][23]/P0001  , \wishbone_bd_ram_mem2_reg[161][16]/P0001  , \wishbone_bd_ram_mem2_reg[161][17]/P0001  , \wishbone_bd_ram_mem2_reg[161][18]/P0001  , \wishbone_bd_ram_mem2_reg[161][19]/P0001  , \wishbone_bd_ram_mem2_reg[161][20]/P0001  , \wishbone_bd_ram_mem2_reg[161][21]/P0001  , \wishbone_bd_ram_mem2_reg[161][22]/P0001  , \wishbone_bd_ram_mem2_reg[161][23]/P0001  , \wishbone_bd_ram_mem2_reg[162][16]/P0001  , \wishbone_bd_ram_mem2_reg[162][17]/P0001  , \wishbone_bd_ram_mem2_reg[162][18]/P0001  , \wishbone_bd_ram_mem2_reg[162][19]/P0001  , \wishbone_bd_ram_mem2_reg[162][20]/P0001  , \wishbone_bd_ram_mem2_reg[162][21]/P0001  , \wishbone_bd_ram_mem2_reg[162][22]/P0001  , \wishbone_bd_ram_mem2_reg[162][23]/P0001  , \wishbone_bd_ram_mem2_reg[163][16]/P0001  , \wishbone_bd_ram_mem2_reg[163][17]/P0001  , \wishbone_bd_ram_mem2_reg[163][18]/P0001  , \wishbone_bd_ram_mem2_reg[163][19]/P0001  , \wishbone_bd_ram_mem2_reg[163][20]/P0001  , \wishbone_bd_ram_mem2_reg[163][21]/P0001  , \wishbone_bd_ram_mem2_reg[163][22]/P0001  , \wishbone_bd_ram_mem2_reg[163][23]/P0001  , \wishbone_bd_ram_mem2_reg[164][16]/P0001  , \wishbone_bd_ram_mem2_reg[164][17]/P0001  , \wishbone_bd_ram_mem2_reg[164][18]/P0001  , \wishbone_bd_ram_mem2_reg[164][19]/P0001  , \wishbone_bd_ram_mem2_reg[164][20]/P0001  , \wishbone_bd_ram_mem2_reg[164][21]/P0001  , \wishbone_bd_ram_mem2_reg[164][22]/P0001  , \wishbone_bd_ram_mem2_reg[164][23]/P0001  , \wishbone_bd_ram_mem2_reg[165][16]/P0001  , \wishbone_bd_ram_mem2_reg[165][17]/P0001  , \wishbone_bd_ram_mem2_reg[165][18]/P0001  , \wishbone_bd_ram_mem2_reg[165][19]/P0001  , \wishbone_bd_ram_mem2_reg[165][20]/P0001  , \wishbone_bd_ram_mem2_reg[165][21]/P0001  , \wishbone_bd_ram_mem2_reg[165][22]/P0001  , \wishbone_bd_ram_mem2_reg[165][23]/P0001  , \wishbone_bd_ram_mem2_reg[166][16]/P0001  , \wishbone_bd_ram_mem2_reg[166][17]/P0001  , \wishbone_bd_ram_mem2_reg[166][18]/P0001  , \wishbone_bd_ram_mem2_reg[166][19]/P0001  , \wishbone_bd_ram_mem2_reg[166][20]/P0001  , \wishbone_bd_ram_mem2_reg[166][21]/P0001  , \wishbone_bd_ram_mem2_reg[166][22]/P0001  , \wishbone_bd_ram_mem2_reg[166][23]/P0001  , \wishbone_bd_ram_mem2_reg[167][16]/P0001  , \wishbone_bd_ram_mem2_reg[167][17]/P0001  , \wishbone_bd_ram_mem2_reg[167][18]/P0001  , \wishbone_bd_ram_mem2_reg[167][19]/P0001  , \wishbone_bd_ram_mem2_reg[167][20]/P0001  , \wishbone_bd_ram_mem2_reg[167][21]/P0001  , \wishbone_bd_ram_mem2_reg[167][22]/P0001  , \wishbone_bd_ram_mem2_reg[167][23]/P0001  , \wishbone_bd_ram_mem2_reg[168][16]/P0001  , \wishbone_bd_ram_mem2_reg[168][17]/P0001  , \wishbone_bd_ram_mem2_reg[168][18]/P0001  , \wishbone_bd_ram_mem2_reg[168][19]/P0001  , \wishbone_bd_ram_mem2_reg[168][20]/P0001  , \wishbone_bd_ram_mem2_reg[168][21]/P0001  , \wishbone_bd_ram_mem2_reg[168][22]/P0001  , \wishbone_bd_ram_mem2_reg[168][23]/P0001  , \wishbone_bd_ram_mem2_reg[169][16]/P0001  , \wishbone_bd_ram_mem2_reg[169][17]/P0001  , \wishbone_bd_ram_mem2_reg[169][18]/P0001  , \wishbone_bd_ram_mem2_reg[169][19]/P0001  , \wishbone_bd_ram_mem2_reg[169][20]/P0001  , \wishbone_bd_ram_mem2_reg[169][21]/P0001  , \wishbone_bd_ram_mem2_reg[169][22]/P0001  , \wishbone_bd_ram_mem2_reg[169][23]/P0001  , \wishbone_bd_ram_mem2_reg[16][16]/P0001  , \wishbone_bd_ram_mem2_reg[16][17]/P0001  , \wishbone_bd_ram_mem2_reg[16][18]/P0001  , \wishbone_bd_ram_mem2_reg[16][19]/P0001  , \wishbone_bd_ram_mem2_reg[16][20]/P0001  , \wishbone_bd_ram_mem2_reg[16][21]/P0001  , \wishbone_bd_ram_mem2_reg[16][22]/P0001  , \wishbone_bd_ram_mem2_reg[16][23]/P0001  , \wishbone_bd_ram_mem2_reg[170][16]/P0001  , \wishbone_bd_ram_mem2_reg[170][17]/P0001  , \wishbone_bd_ram_mem2_reg[170][18]/P0001  , \wishbone_bd_ram_mem2_reg[170][19]/P0001  , \wishbone_bd_ram_mem2_reg[170][20]/P0001  , \wishbone_bd_ram_mem2_reg[170][21]/P0001  , \wishbone_bd_ram_mem2_reg[170][22]/P0001  , \wishbone_bd_ram_mem2_reg[170][23]/P0001  , \wishbone_bd_ram_mem2_reg[171][16]/P0001  , \wishbone_bd_ram_mem2_reg[171][17]/P0001  , \wishbone_bd_ram_mem2_reg[171][18]/P0001  , \wishbone_bd_ram_mem2_reg[171][19]/P0001  , \wishbone_bd_ram_mem2_reg[171][20]/P0001  , \wishbone_bd_ram_mem2_reg[171][21]/P0001  , \wishbone_bd_ram_mem2_reg[171][22]/P0001  , \wishbone_bd_ram_mem2_reg[171][23]/P0001  , \wishbone_bd_ram_mem2_reg[172][16]/P0001  , \wishbone_bd_ram_mem2_reg[172][17]/P0001  , \wishbone_bd_ram_mem2_reg[172][18]/P0001  , \wishbone_bd_ram_mem2_reg[172][19]/P0001  , \wishbone_bd_ram_mem2_reg[172][20]/P0001  , \wishbone_bd_ram_mem2_reg[172][21]/P0001  , \wishbone_bd_ram_mem2_reg[172][22]/P0001  , \wishbone_bd_ram_mem2_reg[172][23]/P0001  , \wishbone_bd_ram_mem2_reg[173][16]/P0001  , \wishbone_bd_ram_mem2_reg[173][17]/P0001  , \wishbone_bd_ram_mem2_reg[173][18]/P0001  , \wishbone_bd_ram_mem2_reg[173][19]/P0001  , \wishbone_bd_ram_mem2_reg[173][20]/P0001  , \wishbone_bd_ram_mem2_reg[173][21]/P0001  , \wishbone_bd_ram_mem2_reg[173][22]/P0001  , \wishbone_bd_ram_mem2_reg[173][23]/P0001  , \wishbone_bd_ram_mem2_reg[174][16]/P0001  , \wishbone_bd_ram_mem2_reg[174][17]/P0001  , \wishbone_bd_ram_mem2_reg[174][18]/P0001  , \wishbone_bd_ram_mem2_reg[174][19]/P0001  , \wishbone_bd_ram_mem2_reg[174][20]/P0001  , \wishbone_bd_ram_mem2_reg[174][21]/P0001  , \wishbone_bd_ram_mem2_reg[174][22]/P0001  , \wishbone_bd_ram_mem2_reg[174][23]/P0001  , \wishbone_bd_ram_mem2_reg[175][16]/P0001  , \wishbone_bd_ram_mem2_reg[175][17]/P0001  , \wishbone_bd_ram_mem2_reg[175][18]/P0001  , \wishbone_bd_ram_mem2_reg[175][19]/P0001  , \wishbone_bd_ram_mem2_reg[175][20]/P0001  , \wishbone_bd_ram_mem2_reg[175][21]/P0001  , \wishbone_bd_ram_mem2_reg[175][22]/P0001  , \wishbone_bd_ram_mem2_reg[175][23]/P0001  , \wishbone_bd_ram_mem2_reg[176][16]/P0001  , \wishbone_bd_ram_mem2_reg[176][17]/P0001  , \wishbone_bd_ram_mem2_reg[176][18]/P0001  , \wishbone_bd_ram_mem2_reg[176][19]/P0001  , \wishbone_bd_ram_mem2_reg[176][20]/P0001  , \wishbone_bd_ram_mem2_reg[176][21]/P0001  , \wishbone_bd_ram_mem2_reg[176][22]/P0001  , \wishbone_bd_ram_mem2_reg[176][23]/P0001  , \wishbone_bd_ram_mem2_reg[177][16]/P0001  , \wishbone_bd_ram_mem2_reg[177][17]/P0001  , \wishbone_bd_ram_mem2_reg[177][18]/P0001  , \wishbone_bd_ram_mem2_reg[177][19]/P0001  , \wishbone_bd_ram_mem2_reg[177][20]/P0001  , \wishbone_bd_ram_mem2_reg[177][21]/P0001  , \wishbone_bd_ram_mem2_reg[177][22]/P0001  , \wishbone_bd_ram_mem2_reg[177][23]/P0001  , \wishbone_bd_ram_mem2_reg[178][16]/P0001  , \wishbone_bd_ram_mem2_reg[178][17]/P0001  , \wishbone_bd_ram_mem2_reg[178][18]/P0001  , \wishbone_bd_ram_mem2_reg[178][19]/P0001  , \wishbone_bd_ram_mem2_reg[178][20]/P0001  , \wishbone_bd_ram_mem2_reg[178][21]/P0001  , \wishbone_bd_ram_mem2_reg[178][22]/P0001  , \wishbone_bd_ram_mem2_reg[178][23]/P0001  , \wishbone_bd_ram_mem2_reg[179][16]/P0001  , \wishbone_bd_ram_mem2_reg[179][17]/P0001  , \wishbone_bd_ram_mem2_reg[179][18]/P0001  , \wishbone_bd_ram_mem2_reg[179][19]/P0001  , \wishbone_bd_ram_mem2_reg[179][20]/P0001  , \wishbone_bd_ram_mem2_reg[179][21]/P0001  , \wishbone_bd_ram_mem2_reg[179][22]/P0001  , \wishbone_bd_ram_mem2_reg[179][23]/P0001  , \wishbone_bd_ram_mem2_reg[17][16]/P0001  , \wishbone_bd_ram_mem2_reg[17][17]/P0001  , \wishbone_bd_ram_mem2_reg[17][18]/P0001  , \wishbone_bd_ram_mem2_reg[17][19]/P0001  , \wishbone_bd_ram_mem2_reg[17][20]/P0001  , \wishbone_bd_ram_mem2_reg[17][21]/P0001  , \wishbone_bd_ram_mem2_reg[17][22]/P0001  , \wishbone_bd_ram_mem2_reg[17][23]/P0001  , \wishbone_bd_ram_mem2_reg[180][16]/P0001  , \wishbone_bd_ram_mem2_reg[180][17]/P0001  , \wishbone_bd_ram_mem2_reg[180][18]/P0001  , \wishbone_bd_ram_mem2_reg[180][19]/P0001  , \wishbone_bd_ram_mem2_reg[180][20]/P0001  , \wishbone_bd_ram_mem2_reg[180][21]/P0001  , \wishbone_bd_ram_mem2_reg[180][22]/P0001  , \wishbone_bd_ram_mem2_reg[180][23]/P0001  , \wishbone_bd_ram_mem2_reg[181][16]/P0001  , \wishbone_bd_ram_mem2_reg[181][17]/P0001  , \wishbone_bd_ram_mem2_reg[181][18]/P0001  , \wishbone_bd_ram_mem2_reg[181][19]/P0001  , \wishbone_bd_ram_mem2_reg[181][20]/P0001  , \wishbone_bd_ram_mem2_reg[181][21]/P0001  , \wishbone_bd_ram_mem2_reg[181][22]/P0001  , \wishbone_bd_ram_mem2_reg[181][23]/P0001  , \wishbone_bd_ram_mem2_reg[182][16]/P0001  , \wishbone_bd_ram_mem2_reg[182][17]/P0001  , \wishbone_bd_ram_mem2_reg[182][18]/P0001  , \wishbone_bd_ram_mem2_reg[182][19]/P0001  , \wishbone_bd_ram_mem2_reg[182][20]/P0001  , \wishbone_bd_ram_mem2_reg[182][21]/P0001  , \wishbone_bd_ram_mem2_reg[182][22]/P0001  , \wishbone_bd_ram_mem2_reg[182][23]/P0001  , \wishbone_bd_ram_mem2_reg[183][16]/P0001  , \wishbone_bd_ram_mem2_reg[183][17]/P0001  , \wishbone_bd_ram_mem2_reg[183][18]/P0001  , \wishbone_bd_ram_mem2_reg[183][19]/P0001  , \wishbone_bd_ram_mem2_reg[183][20]/P0001  , \wishbone_bd_ram_mem2_reg[183][21]/P0001  , \wishbone_bd_ram_mem2_reg[183][22]/P0001  , \wishbone_bd_ram_mem2_reg[183][23]/P0001  , \wishbone_bd_ram_mem2_reg[184][16]/P0001  , \wishbone_bd_ram_mem2_reg[184][17]/P0001  , \wishbone_bd_ram_mem2_reg[184][18]/P0001  , \wishbone_bd_ram_mem2_reg[184][19]/P0001  , \wishbone_bd_ram_mem2_reg[184][20]/P0001  , \wishbone_bd_ram_mem2_reg[184][21]/P0001  , \wishbone_bd_ram_mem2_reg[184][22]/P0001  , \wishbone_bd_ram_mem2_reg[184][23]/P0001  , \wishbone_bd_ram_mem2_reg[185][16]/P0001  , \wishbone_bd_ram_mem2_reg[185][17]/P0001  , \wishbone_bd_ram_mem2_reg[185][18]/P0001  , \wishbone_bd_ram_mem2_reg[185][19]/P0001  , \wishbone_bd_ram_mem2_reg[185][20]/P0001  , \wishbone_bd_ram_mem2_reg[185][21]/P0001  , \wishbone_bd_ram_mem2_reg[185][22]/P0001  , \wishbone_bd_ram_mem2_reg[185][23]/P0001  , \wishbone_bd_ram_mem2_reg[186][16]/P0001  , \wishbone_bd_ram_mem2_reg[186][17]/P0001  , \wishbone_bd_ram_mem2_reg[186][18]/P0001  , \wishbone_bd_ram_mem2_reg[186][19]/P0001  , \wishbone_bd_ram_mem2_reg[186][20]/P0001  , \wishbone_bd_ram_mem2_reg[186][21]/P0001  , \wishbone_bd_ram_mem2_reg[186][22]/P0001  , \wishbone_bd_ram_mem2_reg[186][23]/P0001  , \wishbone_bd_ram_mem2_reg[187][16]/P0001  , \wishbone_bd_ram_mem2_reg[187][17]/P0001  , \wishbone_bd_ram_mem2_reg[187][18]/P0001  , \wishbone_bd_ram_mem2_reg[187][19]/P0001  , \wishbone_bd_ram_mem2_reg[187][20]/P0001  , \wishbone_bd_ram_mem2_reg[187][21]/P0001  , \wishbone_bd_ram_mem2_reg[187][22]/P0001  , \wishbone_bd_ram_mem2_reg[187][23]/P0001  , \wishbone_bd_ram_mem2_reg[188][16]/P0001  , \wishbone_bd_ram_mem2_reg[188][17]/P0001  , \wishbone_bd_ram_mem2_reg[188][18]/P0001  , \wishbone_bd_ram_mem2_reg[188][19]/P0001  , \wishbone_bd_ram_mem2_reg[188][20]/P0001  , \wishbone_bd_ram_mem2_reg[188][21]/P0001  , \wishbone_bd_ram_mem2_reg[188][22]/P0001  , \wishbone_bd_ram_mem2_reg[188][23]/P0001  , \wishbone_bd_ram_mem2_reg[189][16]/P0001  , \wishbone_bd_ram_mem2_reg[189][17]/P0001  , \wishbone_bd_ram_mem2_reg[189][18]/P0001  , \wishbone_bd_ram_mem2_reg[189][19]/P0001  , \wishbone_bd_ram_mem2_reg[189][20]/P0001  , \wishbone_bd_ram_mem2_reg[189][21]/P0001  , \wishbone_bd_ram_mem2_reg[189][22]/P0001  , \wishbone_bd_ram_mem2_reg[189][23]/P0001  , \wishbone_bd_ram_mem2_reg[18][16]/P0001  , \wishbone_bd_ram_mem2_reg[18][17]/P0001  , \wishbone_bd_ram_mem2_reg[18][18]/P0001  , \wishbone_bd_ram_mem2_reg[18][19]/P0001  , \wishbone_bd_ram_mem2_reg[18][20]/P0001  , \wishbone_bd_ram_mem2_reg[18][21]/P0001  , \wishbone_bd_ram_mem2_reg[18][22]/P0001  , \wishbone_bd_ram_mem2_reg[18][23]/P0001  , \wishbone_bd_ram_mem2_reg[190][16]/P0001  , \wishbone_bd_ram_mem2_reg[190][17]/P0001  , \wishbone_bd_ram_mem2_reg[190][18]/P0001  , \wishbone_bd_ram_mem2_reg[190][19]/P0001  , \wishbone_bd_ram_mem2_reg[190][20]/P0001  , \wishbone_bd_ram_mem2_reg[190][21]/P0001  , \wishbone_bd_ram_mem2_reg[190][22]/P0001  , \wishbone_bd_ram_mem2_reg[190][23]/P0001  , \wishbone_bd_ram_mem2_reg[191][16]/P0001  , \wishbone_bd_ram_mem2_reg[191][17]/P0001  , \wishbone_bd_ram_mem2_reg[191][18]/P0001  , \wishbone_bd_ram_mem2_reg[191][19]/P0001  , \wishbone_bd_ram_mem2_reg[191][20]/P0001  , \wishbone_bd_ram_mem2_reg[191][21]/P0001  , \wishbone_bd_ram_mem2_reg[191][22]/P0001  , \wishbone_bd_ram_mem2_reg[191][23]/P0001  , \wishbone_bd_ram_mem2_reg[192][16]/P0001  , \wishbone_bd_ram_mem2_reg[192][17]/P0001  , \wishbone_bd_ram_mem2_reg[192][18]/P0001  , \wishbone_bd_ram_mem2_reg[192][19]/P0001  , \wishbone_bd_ram_mem2_reg[192][20]/P0001  , \wishbone_bd_ram_mem2_reg[192][21]/P0001  , \wishbone_bd_ram_mem2_reg[192][22]/P0001  , \wishbone_bd_ram_mem2_reg[192][23]/P0001  , \wishbone_bd_ram_mem2_reg[193][16]/P0001  , \wishbone_bd_ram_mem2_reg[193][17]/P0001  , \wishbone_bd_ram_mem2_reg[193][18]/P0001  , \wishbone_bd_ram_mem2_reg[193][19]/P0001  , \wishbone_bd_ram_mem2_reg[193][20]/P0001  , \wishbone_bd_ram_mem2_reg[193][21]/P0001  , \wishbone_bd_ram_mem2_reg[193][22]/P0001  , \wishbone_bd_ram_mem2_reg[193][23]/P0001  , \wishbone_bd_ram_mem2_reg[194][16]/P0001  , \wishbone_bd_ram_mem2_reg[194][17]/P0001  , \wishbone_bd_ram_mem2_reg[194][18]/P0001  , \wishbone_bd_ram_mem2_reg[194][19]/P0001  , \wishbone_bd_ram_mem2_reg[194][20]/P0001  , \wishbone_bd_ram_mem2_reg[194][21]/P0001  , \wishbone_bd_ram_mem2_reg[194][22]/P0001  , \wishbone_bd_ram_mem2_reg[194][23]/P0001  , \wishbone_bd_ram_mem2_reg[195][16]/P0001  , \wishbone_bd_ram_mem2_reg[195][17]/P0001  , \wishbone_bd_ram_mem2_reg[195][18]/P0001  , \wishbone_bd_ram_mem2_reg[195][19]/P0001  , \wishbone_bd_ram_mem2_reg[195][20]/P0001  , \wishbone_bd_ram_mem2_reg[195][21]/P0001  , \wishbone_bd_ram_mem2_reg[195][22]/P0001  , \wishbone_bd_ram_mem2_reg[195][23]/P0001  , \wishbone_bd_ram_mem2_reg[196][16]/P0001  , \wishbone_bd_ram_mem2_reg[196][17]/P0001  , \wishbone_bd_ram_mem2_reg[196][18]/P0001  , \wishbone_bd_ram_mem2_reg[196][19]/P0001  , \wishbone_bd_ram_mem2_reg[196][20]/P0001  , \wishbone_bd_ram_mem2_reg[196][21]/P0001  , \wishbone_bd_ram_mem2_reg[196][22]/P0001  , \wishbone_bd_ram_mem2_reg[196][23]/P0001  , \wishbone_bd_ram_mem2_reg[197][16]/P0001  , \wishbone_bd_ram_mem2_reg[197][17]/P0001  , \wishbone_bd_ram_mem2_reg[197][18]/P0001  , \wishbone_bd_ram_mem2_reg[197][19]/P0001  , \wishbone_bd_ram_mem2_reg[197][20]/P0001  , \wishbone_bd_ram_mem2_reg[197][21]/P0001  , \wishbone_bd_ram_mem2_reg[197][22]/P0001  , \wishbone_bd_ram_mem2_reg[197][23]/P0001  , \wishbone_bd_ram_mem2_reg[198][16]/P0001  , \wishbone_bd_ram_mem2_reg[198][17]/P0001  , \wishbone_bd_ram_mem2_reg[198][18]/P0001  , \wishbone_bd_ram_mem2_reg[198][19]/P0001  , \wishbone_bd_ram_mem2_reg[198][20]/P0001  , \wishbone_bd_ram_mem2_reg[198][21]/P0001  , \wishbone_bd_ram_mem2_reg[198][22]/P0001  , \wishbone_bd_ram_mem2_reg[198][23]/P0001  , \wishbone_bd_ram_mem2_reg[199][16]/P0001  , \wishbone_bd_ram_mem2_reg[199][17]/P0001  , \wishbone_bd_ram_mem2_reg[199][18]/P0001  , \wishbone_bd_ram_mem2_reg[199][19]/P0001  , \wishbone_bd_ram_mem2_reg[199][20]/P0001  , \wishbone_bd_ram_mem2_reg[199][21]/P0001  , \wishbone_bd_ram_mem2_reg[199][22]/P0001  , \wishbone_bd_ram_mem2_reg[199][23]/P0001  , \wishbone_bd_ram_mem2_reg[19][16]/P0001  , \wishbone_bd_ram_mem2_reg[19][17]/P0001  , \wishbone_bd_ram_mem2_reg[19][18]/P0001  , \wishbone_bd_ram_mem2_reg[19][19]/P0001  , \wishbone_bd_ram_mem2_reg[19][20]/P0001  , \wishbone_bd_ram_mem2_reg[19][21]/P0001  , \wishbone_bd_ram_mem2_reg[19][22]/P0001  , \wishbone_bd_ram_mem2_reg[19][23]/P0001  , \wishbone_bd_ram_mem2_reg[1][16]/P0001  , \wishbone_bd_ram_mem2_reg[1][17]/P0001  , \wishbone_bd_ram_mem2_reg[1][18]/P0001  , \wishbone_bd_ram_mem2_reg[1][19]/P0001  , \wishbone_bd_ram_mem2_reg[1][20]/P0001  , \wishbone_bd_ram_mem2_reg[1][21]/P0001  , \wishbone_bd_ram_mem2_reg[1][22]/P0001  , \wishbone_bd_ram_mem2_reg[1][23]/P0001  , \wishbone_bd_ram_mem2_reg[200][16]/P0001  , \wishbone_bd_ram_mem2_reg[200][17]/P0001  , \wishbone_bd_ram_mem2_reg[200][18]/P0001  , \wishbone_bd_ram_mem2_reg[200][19]/P0001  , \wishbone_bd_ram_mem2_reg[200][20]/P0001  , \wishbone_bd_ram_mem2_reg[200][21]/P0001  , \wishbone_bd_ram_mem2_reg[200][22]/P0001  , \wishbone_bd_ram_mem2_reg[200][23]/P0001  , \wishbone_bd_ram_mem2_reg[201][16]/P0001  , \wishbone_bd_ram_mem2_reg[201][17]/P0001  , \wishbone_bd_ram_mem2_reg[201][18]/P0001  , \wishbone_bd_ram_mem2_reg[201][19]/P0001  , \wishbone_bd_ram_mem2_reg[201][20]/P0001  , \wishbone_bd_ram_mem2_reg[201][21]/P0001  , \wishbone_bd_ram_mem2_reg[201][22]/P0001  , \wishbone_bd_ram_mem2_reg[201][23]/P0001  , \wishbone_bd_ram_mem2_reg[202][16]/P0001  , \wishbone_bd_ram_mem2_reg[202][17]/P0001  , \wishbone_bd_ram_mem2_reg[202][18]/P0001  , \wishbone_bd_ram_mem2_reg[202][19]/P0001  , \wishbone_bd_ram_mem2_reg[202][20]/P0001  , \wishbone_bd_ram_mem2_reg[202][21]/P0001  , \wishbone_bd_ram_mem2_reg[202][22]/P0001  , \wishbone_bd_ram_mem2_reg[202][23]/P0001  , \wishbone_bd_ram_mem2_reg[203][16]/P0001  , \wishbone_bd_ram_mem2_reg[203][17]/P0001  , \wishbone_bd_ram_mem2_reg[203][18]/P0001  , \wishbone_bd_ram_mem2_reg[203][19]/P0001  , \wishbone_bd_ram_mem2_reg[203][20]/P0001  , \wishbone_bd_ram_mem2_reg[203][21]/P0001  , \wishbone_bd_ram_mem2_reg[203][22]/P0001  , \wishbone_bd_ram_mem2_reg[203][23]/P0001  , \wishbone_bd_ram_mem2_reg[204][16]/P0001  , \wishbone_bd_ram_mem2_reg[204][17]/P0001  , \wishbone_bd_ram_mem2_reg[204][18]/P0001  , \wishbone_bd_ram_mem2_reg[204][19]/P0001  , \wishbone_bd_ram_mem2_reg[204][20]/P0001  , \wishbone_bd_ram_mem2_reg[204][21]/P0001  , \wishbone_bd_ram_mem2_reg[204][22]/P0001  , \wishbone_bd_ram_mem2_reg[204][23]/P0001  , \wishbone_bd_ram_mem2_reg[205][16]/P0001  , \wishbone_bd_ram_mem2_reg[205][17]/P0001  , \wishbone_bd_ram_mem2_reg[205][18]/P0001  , \wishbone_bd_ram_mem2_reg[205][19]/P0001  , \wishbone_bd_ram_mem2_reg[205][20]/P0001  , \wishbone_bd_ram_mem2_reg[205][21]/P0001  , \wishbone_bd_ram_mem2_reg[205][22]/P0001  , \wishbone_bd_ram_mem2_reg[205][23]/P0001  , \wishbone_bd_ram_mem2_reg[206][16]/P0001  , \wishbone_bd_ram_mem2_reg[206][17]/P0001  , \wishbone_bd_ram_mem2_reg[206][18]/P0001  , \wishbone_bd_ram_mem2_reg[206][19]/P0001  , \wishbone_bd_ram_mem2_reg[206][20]/P0001  , \wishbone_bd_ram_mem2_reg[206][21]/P0001  , \wishbone_bd_ram_mem2_reg[206][22]/P0001  , \wishbone_bd_ram_mem2_reg[206][23]/P0001  , \wishbone_bd_ram_mem2_reg[207][16]/P0001  , \wishbone_bd_ram_mem2_reg[207][17]/P0001  , \wishbone_bd_ram_mem2_reg[207][18]/P0001  , \wishbone_bd_ram_mem2_reg[207][19]/P0001  , \wishbone_bd_ram_mem2_reg[207][20]/P0001  , \wishbone_bd_ram_mem2_reg[207][21]/P0001  , \wishbone_bd_ram_mem2_reg[207][22]/P0001  , \wishbone_bd_ram_mem2_reg[207][23]/P0001  , \wishbone_bd_ram_mem2_reg[208][16]/P0001  , \wishbone_bd_ram_mem2_reg[208][17]/P0001  , \wishbone_bd_ram_mem2_reg[208][18]/P0001  , \wishbone_bd_ram_mem2_reg[208][19]/P0001  , \wishbone_bd_ram_mem2_reg[208][20]/P0001  , \wishbone_bd_ram_mem2_reg[208][21]/P0001  , \wishbone_bd_ram_mem2_reg[208][22]/P0001  , \wishbone_bd_ram_mem2_reg[208][23]/P0001  , \wishbone_bd_ram_mem2_reg[209][16]/P0001  , \wishbone_bd_ram_mem2_reg[209][17]/P0001  , \wishbone_bd_ram_mem2_reg[209][18]/P0001  , \wishbone_bd_ram_mem2_reg[209][19]/P0001  , \wishbone_bd_ram_mem2_reg[209][20]/P0001  , \wishbone_bd_ram_mem2_reg[209][21]/P0001  , \wishbone_bd_ram_mem2_reg[209][22]/P0001  , \wishbone_bd_ram_mem2_reg[209][23]/P0001  , \wishbone_bd_ram_mem2_reg[20][16]/P0001  , \wishbone_bd_ram_mem2_reg[20][17]/P0001  , \wishbone_bd_ram_mem2_reg[20][18]/P0001  , \wishbone_bd_ram_mem2_reg[20][19]/P0001  , \wishbone_bd_ram_mem2_reg[20][20]/P0001  , \wishbone_bd_ram_mem2_reg[20][21]/P0001  , \wishbone_bd_ram_mem2_reg[20][22]/P0001  , \wishbone_bd_ram_mem2_reg[20][23]/P0001  , \wishbone_bd_ram_mem2_reg[210][16]/P0001  , \wishbone_bd_ram_mem2_reg[210][17]/P0001  , \wishbone_bd_ram_mem2_reg[210][18]/P0001  , \wishbone_bd_ram_mem2_reg[210][19]/P0001  , \wishbone_bd_ram_mem2_reg[210][20]/P0001  , \wishbone_bd_ram_mem2_reg[210][21]/P0001  , \wishbone_bd_ram_mem2_reg[210][22]/P0001  , \wishbone_bd_ram_mem2_reg[210][23]/P0001  , \wishbone_bd_ram_mem2_reg[211][16]/P0001  , \wishbone_bd_ram_mem2_reg[211][17]/P0001  , \wishbone_bd_ram_mem2_reg[211][18]/P0001  , \wishbone_bd_ram_mem2_reg[211][19]/P0001  , \wishbone_bd_ram_mem2_reg[211][20]/P0001  , \wishbone_bd_ram_mem2_reg[211][21]/P0001  , \wishbone_bd_ram_mem2_reg[211][22]/P0001  , \wishbone_bd_ram_mem2_reg[211][23]/P0001  , \wishbone_bd_ram_mem2_reg[212][16]/P0001  , \wishbone_bd_ram_mem2_reg[212][17]/P0001  , \wishbone_bd_ram_mem2_reg[212][18]/P0001  , \wishbone_bd_ram_mem2_reg[212][19]/P0001  , \wishbone_bd_ram_mem2_reg[212][20]/P0001  , \wishbone_bd_ram_mem2_reg[212][21]/P0001  , \wishbone_bd_ram_mem2_reg[212][22]/P0001  , \wishbone_bd_ram_mem2_reg[212][23]/P0001  , \wishbone_bd_ram_mem2_reg[213][16]/P0001  , \wishbone_bd_ram_mem2_reg[213][17]/P0001  , \wishbone_bd_ram_mem2_reg[213][18]/P0001  , \wishbone_bd_ram_mem2_reg[213][19]/P0001  , \wishbone_bd_ram_mem2_reg[213][20]/P0001  , \wishbone_bd_ram_mem2_reg[213][21]/P0001  , \wishbone_bd_ram_mem2_reg[213][22]/P0001  , \wishbone_bd_ram_mem2_reg[213][23]/P0001  , \wishbone_bd_ram_mem2_reg[214][16]/P0001  , \wishbone_bd_ram_mem2_reg[214][17]/P0001  , \wishbone_bd_ram_mem2_reg[214][18]/P0001  , \wishbone_bd_ram_mem2_reg[214][19]/P0001  , \wishbone_bd_ram_mem2_reg[214][20]/P0001  , \wishbone_bd_ram_mem2_reg[214][21]/P0001  , \wishbone_bd_ram_mem2_reg[214][22]/P0001  , \wishbone_bd_ram_mem2_reg[214][23]/P0001  , \wishbone_bd_ram_mem2_reg[215][16]/P0001  , \wishbone_bd_ram_mem2_reg[215][17]/P0001  , \wishbone_bd_ram_mem2_reg[215][18]/P0001  , \wishbone_bd_ram_mem2_reg[215][19]/P0001  , \wishbone_bd_ram_mem2_reg[215][20]/P0001  , \wishbone_bd_ram_mem2_reg[215][21]/P0001  , \wishbone_bd_ram_mem2_reg[215][22]/P0001  , \wishbone_bd_ram_mem2_reg[215][23]/P0001  , \wishbone_bd_ram_mem2_reg[216][16]/P0001  , \wishbone_bd_ram_mem2_reg[216][17]/P0001  , \wishbone_bd_ram_mem2_reg[216][18]/P0001  , \wishbone_bd_ram_mem2_reg[216][19]/P0001  , \wishbone_bd_ram_mem2_reg[216][20]/P0001  , \wishbone_bd_ram_mem2_reg[216][21]/P0001  , \wishbone_bd_ram_mem2_reg[216][22]/P0001  , \wishbone_bd_ram_mem2_reg[216][23]/P0001  , \wishbone_bd_ram_mem2_reg[217][16]/P0001  , \wishbone_bd_ram_mem2_reg[217][17]/P0001  , \wishbone_bd_ram_mem2_reg[217][18]/P0001  , \wishbone_bd_ram_mem2_reg[217][19]/P0001  , \wishbone_bd_ram_mem2_reg[217][20]/P0001  , \wishbone_bd_ram_mem2_reg[217][21]/P0001  , \wishbone_bd_ram_mem2_reg[217][22]/P0001  , \wishbone_bd_ram_mem2_reg[217][23]/P0001  , \wishbone_bd_ram_mem2_reg[218][16]/P0001  , \wishbone_bd_ram_mem2_reg[218][17]/P0001  , \wishbone_bd_ram_mem2_reg[218][18]/P0001  , \wishbone_bd_ram_mem2_reg[218][19]/P0001  , \wishbone_bd_ram_mem2_reg[218][20]/P0001  , \wishbone_bd_ram_mem2_reg[218][21]/P0001  , \wishbone_bd_ram_mem2_reg[218][22]/P0001  , \wishbone_bd_ram_mem2_reg[218][23]/P0001  , \wishbone_bd_ram_mem2_reg[219][16]/P0001  , \wishbone_bd_ram_mem2_reg[219][17]/P0001  , \wishbone_bd_ram_mem2_reg[219][18]/P0001  , \wishbone_bd_ram_mem2_reg[219][19]/P0001  , \wishbone_bd_ram_mem2_reg[219][20]/P0001  , \wishbone_bd_ram_mem2_reg[219][21]/P0001  , \wishbone_bd_ram_mem2_reg[219][22]/P0001  , \wishbone_bd_ram_mem2_reg[219][23]/P0001  , \wishbone_bd_ram_mem2_reg[21][16]/P0001  , \wishbone_bd_ram_mem2_reg[21][17]/P0001  , \wishbone_bd_ram_mem2_reg[21][18]/P0001  , \wishbone_bd_ram_mem2_reg[21][19]/P0001  , \wishbone_bd_ram_mem2_reg[21][20]/P0001  , \wishbone_bd_ram_mem2_reg[21][21]/P0001  , \wishbone_bd_ram_mem2_reg[21][22]/P0001  , \wishbone_bd_ram_mem2_reg[21][23]/P0001  , \wishbone_bd_ram_mem2_reg[220][16]/P0001  , \wishbone_bd_ram_mem2_reg[220][17]/P0001  , \wishbone_bd_ram_mem2_reg[220][18]/P0001  , \wishbone_bd_ram_mem2_reg[220][19]/P0001  , \wishbone_bd_ram_mem2_reg[220][20]/P0001  , \wishbone_bd_ram_mem2_reg[220][21]/P0001  , \wishbone_bd_ram_mem2_reg[220][22]/P0001  , \wishbone_bd_ram_mem2_reg[220][23]/P0001  , \wishbone_bd_ram_mem2_reg[221][16]/P0001  , \wishbone_bd_ram_mem2_reg[221][17]/P0001  , \wishbone_bd_ram_mem2_reg[221][18]/P0001  , \wishbone_bd_ram_mem2_reg[221][19]/P0001  , \wishbone_bd_ram_mem2_reg[221][20]/P0001  , \wishbone_bd_ram_mem2_reg[221][21]/P0001  , \wishbone_bd_ram_mem2_reg[221][22]/P0001  , \wishbone_bd_ram_mem2_reg[221][23]/P0001  , \wishbone_bd_ram_mem2_reg[222][16]/P0001  , \wishbone_bd_ram_mem2_reg[222][17]/P0001  , \wishbone_bd_ram_mem2_reg[222][18]/P0001  , \wishbone_bd_ram_mem2_reg[222][19]/P0001  , \wishbone_bd_ram_mem2_reg[222][20]/P0001  , \wishbone_bd_ram_mem2_reg[222][21]/P0001  , \wishbone_bd_ram_mem2_reg[222][22]/P0001  , \wishbone_bd_ram_mem2_reg[222][23]/P0001  , \wishbone_bd_ram_mem2_reg[223][16]/P0001  , \wishbone_bd_ram_mem2_reg[223][17]/P0001  , \wishbone_bd_ram_mem2_reg[223][18]/P0001  , \wishbone_bd_ram_mem2_reg[223][19]/P0001  , \wishbone_bd_ram_mem2_reg[223][20]/P0001  , \wishbone_bd_ram_mem2_reg[223][21]/P0001  , \wishbone_bd_ram_mem2_reg[223][22]/P0001  , \wishbone_bd_ram_mem2_reg[223][23]/P0001  , \wishbone_bd_ram_mem2_reg[224][16]/P0001  , \wishbone_bd_ram_mem2_reg[224][17]/P0001  , \wishbone_bd_ram_mem2_reg[224][18]/P0001  , \wishbone_bd_ram_mem2_reg[224][19]/P0001  , \wishbone_bd_ram_mem2_reg[224][20]/P0001  , \wishbone_bd_ram_mem2_reg[224][21]/P0001  , \wishbone_bd_ram_mem2_reg[224][22]/P0001  , \wishbone_bd_ram_mem2_reg[224][23]/P0001  , \wishbone_bd_ram_mem2_reg[225][16]/P0001  , \wishbone_bd_ram_mem2_reg[225][17]/P0001  , \wishbone_bd_ram_mem2_reg[225][18]/P0001  , \wishbone_bd_ram_mem2_reg[225][19]/P0001  , \wishbone_bd_ram_mem2_reg[225][20]/P0001  , \wishbone_bd_ram_mem2_reg[225][21]/P0001  , \wishbone_bd_ram_mem2_reg[225][22]/P0001  , \wishbone_bd_ram_mem2_reg[225][23]/P0001  , \wishbone_bd_ram_mem2_reg[226][16]/P0001  , \wishbone_bd_ram_mem2_reg[226][17]/P0001  , \wishbone_bd_ram_mem2_reg[226][18]/P0001  , \wishbone_bd_ram_mem2_reg[226][19]/P0001  , \wishbone_bd_ram_mem2_reg[226][20]/P0001  , \wishbone_bd_ram_mem2_reg[226][21]/P0001  , \wishbone_bd_ram_mem2_reg[226][22]/P0001  , \wishbone_bd_ram_mem2_reg[226][23]/P0001  , \wishbone_bd_ram_mem2_reg[227][16]/P0001  , \wishbone_bd_ram_mem2_reg[227][17]/P0001  , \wishbone_bd_ram_mem2_reg[227][18]/P0001  , \wishbone_bd_ram_mem2_reg[227][19]/P0001  , \wishbone_bd_ram_mem2_reg[227][20]/P0001  , \wishbone_bd_ram_mem2_reg[227][21]/P0001  , \wishbone_bd_ram_mem2_reg[227][22]/P0001  , \wishbone_bd_ram_mem2_reg[227][23]/P0001  , \wishbone_bd_ram_mem2_reg[228][16]/P0001  , \wishbone_bd_ram_mem2_reg[228][17]/P0001  , \wishbone_bd_ram_mem2_reg[228][18]/P0001  , \wishbone_bd_ram_mem2_reg[228][19]/P0001  , \wishbone_bd_ram_mem2_reg[228][20]/P0001  , \wishbone_bd_ram_mem2_reg[228][21]/P0001  , \wishbone_bd_ram_mem2_reg[228][22]/P0001  , \wishbone_bd_ram_mem2_reg[228][23]/P0001  , \wishbone_bd_ram_mem2_reg[229][16]/P0001  , \wishbone_bd_ram_mem2_reg[229][17]/P0001  , \wishbone_bd_ram_mem2_reg[229][18]/P0001  , \wishbone_bd_ram_mem2_reg[229][19]/P0001  , \wishbone_bd_ram_mem2_reg[229][20]/P0001  , \wishbone_bd_ram_mem2_reg[229][21]/P0001  , \wishbone_bd_ram_mem2_reg[229][22]/P0001  , \wishbone_bd_ram_mem2_reg[229][23]/P0001  , \wishbone_bd_ram_mem2_reg[22][16]/P0001  , \wishbone_bd_ram_mem2_reg[22][17]/P0001  , \wishbone_bd_ram_mem2_reg[22][18]/P0001  , \wishbone_bd_ram_mem2_reg[22][19]/P0001  , \wishbone_bd_ram_mem2_reg[22][20]/P0001  , \wishbone_bd_ram_mem2_reg[22][21]/P0001  , \wishbone_bd_ram_mem2_reg[22][22]/P0001  , \wishbone_bd_ram_mem2_reg[22][23]/P0001  , \wishbone_bd_ram_mem2_reg[230][16]/P0001  , \wishbone_bd_ram_mem2_reg[230][17]/P0001  , \wishbone_bd_ram_mem2_reg[230][18]/P0001  , \wishbone_bd_ram_mem2_reg[230][19]/P0001  , \wishbone_bd_ram_mem2_reg[230][20]/P0001  , \wishbone_bd_ram_mem2_reg[230][21]/P0001  , \wishbone_bd_ram_mem2_reg[230][22]/P0001  , \wishbone_bd_ram_mem2_reg[230][23]/P0001  , \wishbone_bd_ram_mem2_reg[231][16]/P0001  , \wishbone_bd_ram_mem2_reg[231][17]/P0001  , \wishbone_bd_ram_mem2_reg[231][18]/P0001  , \wishbone_bd_ram_mem2_reg[231][19]/P0001  , \wishbone_bd_ram_mem2_reg[231][20]/P0001  , \wishbone_bd_ram_mem2_reg[231][21]/P0001  , \wishbone_bd_ram_mem2_reg[231][22]/P0001  , \wishbone_bd_ram_mem2_reg[231][23]/P0001  , \wishbone_bd_ram_mem2_reg[232][16]/P0001  , \wishbone_bd_ram_mem2_reg[232][17]/P0001  , \wishbone_bd_ram_mem2_reg[232][18]/P0001  , \wishbone_bd_ram_mem2_reg[232][19]/P0001  , \wishbone_bd_ram_mem2_reg[232][20]/P0001  , \wishbone_bd_ram_mem2_reg[232][21]/P0001  , \wishbone_bd_ram_mem2_reg[232][22]/P0001  , \wishbone_bd_ram_mem2_reg[232][23]/P0001  , \wishbone_bd_ram_mem2_reg[233][16]/P0001  , \wishbone_bd_ram_mem2_reg[233][17]/P0001  , \wishbone_bd_ram_mem2_reg[233][18]/P0001  , \wishbone_bd_ram_mem2_reg[233][19]/P0001  , \wishbone_bd_ram_mem2_reg[233][20]/P0001  , \wishbone_bd_ram_mem2_reg[233][21]/P0001  , \wishbone_bd_ram_mem2_reg[233][22]/P0001  , \wishbone_bd_ram_mem2_reg[233][23]/P0001  , \wishbone_bd_ram_mem2_reg[234][16]/P0001  , \wishbone_bd_ram_mem2_reg[234][17]/P0001  , \wishbone_bd_ram_mem2_reg[234][18]/P0001  , \wishbone_bd_ram_mem2_reg[234][19]/P0001  , \wishbone_bd_ram_mem2_reg[234][20]/P0001  , \wishbone_bd_ram_mem2_reg[234][21]/P0001  , \wishbone_bd_ram_mem2_reg[234][22]/P0001  , \wishbone_bd_ram_mem2_reg[234][23]/P0001  , \wishbone_bd_ram_mem2_reg[235][16]/P0001  , \wishbone_bd_ram_mem2_reg[235][17]/P0001  , \wishbone_bd_ram_mem2_reg[235][18]/P0001  , \wishbone_bd_ram_mem2_reg[235][19]/P0001  , \wishbone_bd_ram_mem2_reg[235][20]/P0001  , \wishbone_bd_ram_mem2_reg[235][21]/P0001  , \wishbone_bd_ram_mem2_reg[235][22]/P0001  , \wishbone_bd_ram_mem2_reg[235][23]/P0001  , \wishbone_bd_ram_mem2_reg[236][16]/P0001  , \wishbone_bd_ram_mem2_reg[236][17]/P0001  , \wishbone_bd_ram_mem2_reg[236][18]/P0001  , \wishbone_bd_ram_mem2_reg[236][19]/P0001  , \wishbone_bd_ram_mem2_reg[236][20]/P0001  , \wishbone_bd_ram_mem2_reg[236][21]/P0001  , \wishbone_bd_ram_mem2_reg[236][22]/P0001  , \wishbone_bd_ram_mem2_reg[236][23]/P0001  , \wishbone_bd_ram_mem2_reg[237][16]/P0001  , \wishbone_bd_ram_mem2_reg[237][17]/P0001  , \wishbone_bd_ram_mem2_reg[237][18]/P0001  , \wishbone_bd_ram_mem2_reg[237][19]/P0001  , \wishbone_bd_ram_mem2_reg[237][20]/P0001  , \wishbone_bd_ram_mem2_reg[237][21]/P0001  , \wishbone_bd_ram_mem2_reg[237][22]/P0001  , \wishbone_bd_ram_mem2_reg[237][23]/P0001  , \wishbone_bd_ram_mem2_reg[238][16]/P0001  , \wishbone_bd_ram_mem2_reg[238][17]/P0001  , \wishbone_bd_ram_mem2_reg[238][18]/P0001  , \wishbone_bd_ram_mem2_reg[238][19]/P0001  , \wishbone_bd_ram_mem2_reg[238][20]/P0001  , \wishbone_bd_ram_mem2_reg[238][21]/P0001  , \wishbone_bd_ram_mem2_reg[238][22]/P0001  , \wishbone_bd_ram_mem2_reg[238][23]/P0001  , \wishbone_bd_ram_mem2_reg[239][16]/P0001  , \wishbone_bd_ram_mem2_reg[239][17]/P0001  , \wishbone_bd_ram_mem2_reg[239][18]/P0001  , \wishbone_bd_ram_mem2_reg[239][19]/P0001  , \wishbone_bd_ram_mem2_reg[239][20]/P0001  , \wishbone_bd_ram_mem2_reg[239][21]/P0001  , \wishbone_bd_ram_mem2_reg[239][22]/P0001  , \wishbone_bd_ram_mem2_reg[239][23]/P0001  , \wishbone_bd_ram_mem2_reg[23][16]/P0001  , \wishbone_bd_ram_mem2_reg[23][17]/P0001  , \wishbone_bd_ram_mem2_reg[23][18]/P0001  , \wishbone_bd_ram_mem2_reg[23][19]/P0001  , \wishbone_bd_ram_mem2_reg[23][20]/P0001  , \wishbone_bd_ram_mem2_reg[23][21]/P0001  , \wishbone_bd_ram_mem2_reg[23][22]/P0001  , \wishbone_bd_ram_mem2_reg[23][23]/P0001  , \wishbone_bd_ram_mem2_reg[240][16]/P0001  , \wishbone_bd_ram_mem2_reg[240][17]/P0001  , \wishbone_bd_ram_mem2_reg[240][18]/P0001  , \wishbone_bd_ram_mem2_reg[240][19]/P0001  , \wishbone_bd_ram_mem2_reg[240][20]/P0001  , \wishbone_bd_ram_mem2_reg[240][21]/P0001  , \wishbone_bd_ram_mem2_reg[240][22]/P0001  , \wishbone_bd_ram_mem2_reg[240][23]/P0001  , \wishbone_bd_ram_mem2_reg[241][16]/P0001  , \wishbone_bd_ram_mem2_reg[241][17]/P0001  , \wishbone_bd_ram_mem2_reg[241][18]/P0001  , \wishbone_bd_ram_mem2_reg[241][19]/P0001  , \wishbone_bd_ram_mem2_reg[241][20]/P0001  , \wishbone_bd_ram_mem2_reg[241][21]/P0001  , \wishbone_bd_ram_mem2_reg[241][22]/P0001  , \wishbone_bd_ram_mem2_reg[241][23]/P0001  , \wishbone_bd_ram_mem2_reg[242][16]/P0001  , \wishbone_bd_ram_mem2_reg[242][17]/P0001  , \wishbone_bd_ram_mem2_reg[242][18]/P0001  , \wishbone_bd_ram_mem2_reg[242][19]/P0001  , \wishbone_bd_ram_mem2_reg[242][20]/P0001  , \wishbone_bd_ram_mem2_reg[242][21]/P0001  , \wishbone_bd_ram_mem2_reg[242][22]/P0001  , \wishbone_bd_ram_mem2_reg[242][23]/P0001  , \wishbone_bd_ram_mem2_reg[243][16]/P0001  , \wishbone_bd_ram_mem2_reg[243][17]/P0001  , \wishbone_bd_ram_mem2_reg[243][18]/P0001  , \wishbone_bd_ram_mem2_reg[243][19]/P0001  , \wishbone_bd_ram_mem2_reg[243][20]/P0001  , \wishbone_bd_ram_mem2_reg[243][21]/P0001  , \wishbone_bd_ram_mem2_reg[243][22]/P0001  , \wishbone_bd_ram_mem2_reg[243][23]/P0001  , \wishbone_bd_ram_mem2_reg[244][16]/P0001  , \wishbone_bd_ram_mem2_reg[244][17]/P0001  , \wishbone_bd_ram_mem2_reg[244][18]/P0001  , \wishbone_bd_ram_mem2_reg[244][19]/P0001  , \wishbone_bd_ram_mem2_reg[244][20]/P0001  , \wishbone_bd_ram_mem2_reg[244][21]/P0001  , \wishbone_bd_ram_mem2_reg[244][22]/P0001  , \wishbone_bd_ram_mem2_reg[244][23]/P0001  , \wishbone_bd_ram_mem2_reg[245][16]/P0001  , \wishbone_bd_ram_mem2_reg[245][17]/P0001  , \wishbone_bd_ram_mem2_reg[245][18]/P0001  , \wishbone_bd_ram_mem2_reg[245][19]/P0001  , \wishbone_bd_ram_mem2_reg[245][20]/P0001  , \wishbone_bd_ram_mem2_reg[245][21]/P0001  , \wishbone_bd_ram_mem2_reg[245][22]/P0001  , \wishbone_bd_ram_mem2_reg[245][23]/P0001  , \wishbone_bd_ram_mem2_reg[246][16]/P0001  , \wishbone_bd_ram_mem2_reg[246][17]/P0001  , \wishbone_bd_ram_mem2_reg[246][18]/P0001  , \wishbone_bd_ram_mem2_reg[246][19]/P0001  , \wishbone_bd_ram_mem2_reg[246][20]/P0001  , \wishbone_bd_ram_mem2_reg[246][21]/P0001  , \wishbone_bd_ram_mem2_reg[246][22]/P0001  , \wishbone_bd_ram_mem2_reg[246][23]/P0001  , \wishbone_bd_ram_mem2_reg[247][16]/P0001  , \wishbone_bd_ram_mem2_reg[247][17]/P0001  , \wishbone_bd_ram_mem2_reg[247][18]/P0001  , \wishbone_bd_ram_mem2_reg[247][19]/P0001  , \wishbone_bd_ram_mem2_reg[247][20]/P0001  , \wishbone_bd_ram_mem2_reg[247][21]/P0001  , \wishbone_bd_ram_mem2_reg[247][22]/P0001  , \wishbone_bd_ram_mem2_reg[247][23]/P0001  , \wishbone_bd_ram_mem2_reg[248][16]/P0001  , \wishbone_bd_ram_mem2_reg[248][17]/P0001  , \wishbone_bd_ram_mem2_reg[248][18]/P0001  , \wishbone_bd_ram_mem2_reg[248][19]/P0001  , \wishbone_bd_ram_mem2_reg[248][20]/P0001  , \wishbone_bd_ram_mem2_reg[248][21]/P0001  , \wishbone_bd_ram_mem2_reg[248][22]/P0001  , \wishbone_bd_ram_mem2_reg[248][23]/P0001  , \wishbone_bd_ram_mem2_reg[249][16]/P0001  , \wishbone_bd_ram_mem2_reg[249][17]/P0001  , \wishbone_bd_ram_mem2_reg[249][18]/P0001  , \wishbone_bd_ram_mem2_reg[249][19]/P0001  , \wishbone_bd_ram_mem2_reg[249][20]/P0001  , \wishbone_bd_ram_mem2_reg[249][21]/P0001  , \wishbone_bd_ram_mem2_reg[249][22]/P0001  , \wishbone_bd_ram_mem2_reg[249][23]/P0001  , \wishbone_bd_ram_mem2_reg[24][16]/P0001  , \wishbone_bd_ram_mem2_reg[24][17]/P0001  , \wishbone_bd_ram_mem2_reg[24][18]/P0001  , \wishbone_bd_ram_mem2_reg[24][19]/P0001  , \wishbone_bd_ram_mem2_reg[24][20]/P0001  , \wishbone_bd_ram_mem2_reg[24][21]/P0001  , \wishbone_bd_ram_mem2_reg[24][22]/P0001  , \wishbone_bd_ram_mem2_reg[24][23]/P0001  , \wishbone_bd_ram_mem2_reg[250][16]/P0001  , \wishbone_bd_ram_mem2_reg[250][17]/P0001  , \wishbone_bd_ram_mem2_reg[250][18]/P0001  , \wishbone_bd_ram_mem2_reg[250][19]/P0001  , \wishbone_bd_ram_mem2_reg[250][20]/P0001  , \wishbone_bd_ram_mem2_reg[250][21]/P0001  , \wishbone_bd_ram_mem2_reg[250][22]/P0001  , \wishbone_bd_ram_mem2_reg[250][23]/P0001  , \wishbone_bd_ram_mem2_reg[251][16]/P0001  , \wishbone_bd_ram_mem2_reg[251][17]/P0001  , \wishbone_bd_ram_mem2_reg[251][18]/P0001  , \wishbone_bd_ram_mem2_reg[251][19]/P0001  , \wishbone_bd_ram_mem2_reg[251][20]/P0001  , \wishbone_bd_ram_mem2_reg[251][21]/P0001  , \wishbone_bd_ram_mem2_reg[251][22]/P0001  , \wishbone_bd_ram_mem2_reg[251][23]/P0001  , \wishbone_bd_ram_mem2_reg[252][16]/P0001  , \wishbone_bd_ram_mem2_reg[252][17]/P0001  , \wishbone_bd_ram_mem2_reg[252][18]/P0001  , \wishbone_bd_ram_mem2_reg[252][19]/P0001  , \wishbone_bd_ram_mem2_reg[252][20]/P0001  , \wishbone_bd_ram_mem2_reg[252][21]/P0001  , \wishbone_bd_ram_mem2_reg[252][22]/P0001  , \wishbone_bd_ram_mem2_reg[252][23]/P0001  , \wishbone_bd_ram_mem2_reg[253][16]/P0001  , \wishbone_bd_ram_mem2_reg[253][17]/P0001  , \wishbone_bd_ram_mem2_reg[253][18]/P0001  , \wishbone_bd_ram_mem2_reg[253][19]/P0001  , \wishbone_bd_ram_mem2_reg[253][20]/P0001  , \wishbone_bd_ram_mem2_reg[253][21]/P0001  , \wishbone_bd_ram_mem2_reg[253][22]/P0001  , \wishbone_bd_ram_mem2_reg[253][23]/P0001  , \wishbone_bd_ram_mem2_reg[254][16]/P0001  , \wishbone_bd_ram_mem2_reg[254][17]/P0001  , \wishbone_bd_ram_mem2_reg[254][18]/P0001  , \wishbone_bd_ram_mem2_reg[254][19]/P0001  , \wishbone_bd_ram_mem2_reg[254][20]/P0001  , \wishbone_bd_ram_mem2_reg[254][21]/P0001  , \wishbone_bd_ram_mem2_reg[254][22]/P0001  , \wishbone_bd_ram_mem2_reg[254][23]/P0001  , \wishbone_bd_ram_mem2_reg[255][16]/P0001  , \wishbone_bd_ram_mem2_reg[255][17]/P0001  , \wishbone_bd_ram_mem2_reg[255][18]/P0001  , \wishbone_bd_ram_mem2_reg[255][19]/P0001  , \wishbone_bd_ram_mem2_reg[255][20]/P0001  , \wishbone_bd_ram_mem2_reg[255][21]/P0001  , \wishbone_bd_ram_mem2_reg[255][22]/P0001  , \wishbone_bd_ram_mem2_reg[255][23]/P0001  , \wishbone_bd_ram_mem2_reg[25][16]/P0001  , \wishbone_bd_ram_mem2_reg[25][17]/P0001  , \wishbone_bd_ram_mem2_reg[25][18]/P0001  , \wishbone_bd_ram_mem2_reg[25][19]/P0001  , \wishbone_bd_ram_mem2_reg[25][20]/P0001  , \wishbone_bd_ram_mem2_reg[25][21]/P0001  , \wishbone_bd_ram_mem2_reg[25][22]/P0001  , \wishbone_bd_ram_mem2_reg[25][23]/P0001  , \wishbone_bd_ram_mem2_reg[26][16]/P0001  , \wishbone_bd_ram_mem2_reg[26][17]/P0001  , \wishbone_bd_ram_mem2_reg[26][18]/P0001  , \wishbone_bd_ram_mem2_reg[26][19]/P0001  , \wishbone_bd_ram_mem2_reg[26][20]/P0001  , \wishbone_bd_ram_mem2_reg[26][21]/P0001  , \wishbone_bd_ram_mem2_reg[26][22]/P0001  , \wishbone_bd_ram_mem2_reg[26][23]/P0001  , \wishbone_bd_ram_mem2_reg[27][16]/P0001  , \wishbone_bd_ram_mem2_reg[27][17]/P0001  , \wishbone_bd_ram_mem2_reg[27][18]/P0001  , \wishbone_bd_ram_mem2_reg[27][19]/P0001  , \wishbone_bd_ram_mem2_reg[27][20]/P0001  , \wishbone_bd_ram_mem2_reg[27][21]/P0001  , \wishbone_bd_ram_mem2_reg[27][22]/P0001  , \wishbone_bd_ram_mem2_reg[27][23]/P0001  , \wishbone_bd_ram_mem2_reg[28][16]/P0001  , \wishbone_bd_ram_mem2_reg[28][17]/P0001  , \wishbone_bd_ram_mem2_reg[28][18]/P0001  , \wishbone_bd_ram_mem2_reg[28][19]/P0001  , \wishbone_bd_ram_mem2_reg[28][20]/P0001  , \wishbone_bd_ram_mem2_reg[28][21]/P0001  , \wishbone_bd_ram_mem2_reg[28][22]/P0001  , \wishbone_bd_ram_mem2_reg[28][23]/P0001  , \wishbone_bd_ram_mem2_reg[29][16]/P0001  , \wishbone_bd_ram_mem2_reg[29][17]/P0001  , \wishbone_bd_ram_mem2_reg[29][18]/P0001  , \wishbone_bd_ram_mem2_reg[29][19]/P0001  , \wishbone_bd_ram_mem2_reg[29][20]/P0001  , \wishbone_bd_ram_mem2_reg[29][21]/P0001  , \wishbone_bd_ram_mem2_reg[29][22]/P0001  , \wishbone_bd_ram_mem2_reg[29][23]/P0001  , \wishbone_bd_ram_mem2_reg[2][16]/P0001  , \wishbone_bd_ram_mem2_reg[2][17]/P0001  , \wishbone_bd_ram_mem2_reg[2][18]/P0001  , \wishbone_bd_ram_mem2_reg[2][19]/P0001  , \wishbone_bd_ram_mem2_reg[2][20]/P0001  , \wishbone_bd_ram_mem2_reg[2][21]/P0001  , \wishbone_bd_ram_mem2_reg[2][22]/P0001  , \wishbone_bd_ram_mem2_reg[2][23]/P0001  , \wishbone_bd_ram_mem2_reg[30][16]/P0001  , \wishbone_bd_ram_mem2_reg[30][17]/P0001  , \wishbone_bd_ram_mem2_reg[30][18]/P0001  , \wishbone_bd_ram_mem2_reg[30][19]/P0001  , \wishbone_bd_ram_mem2_reg[30][20]/P0001  , \wishbone_bd_ram_mem2_reg[30][21]/P0001  , \wishbone_bd_ram_mem2_reg[30][22]/P0001  , \wishbone_bd_ram_mem2_reg[30][23]/P0001  , \wishbone_bd_ram_mem2_reg[31][16]/P0001  , \wishbone_bd_ram_mem2_reg[31][17]/P0001  , \wishbone_bd_ram_mem2_reg[31][18]/P0001  , \wishbone_bd_ram_mem2_reg[31][19]/P0001  , \wishbone_bd_ram_mem2_reg[31][20]/P0001  , \wishbone_bd_ram_mem2_reg[31][21]/P0001  , \wishbone_bd_ram_mem2_reg[31][22]/P0001  , \wishbone_bd_ram_mem2_reg[31][23]/P0001  , \wishbone_bd_ram_mem2_reg[32][16]/P0001  , \wishbone_bd_ram_mem2_reg[32][17]/P0001  , \wishbone_bd_ram_mem2_reg[32][18]/P0001  , \wishbone_bd_ram_mem2_reg[32][19]/P0001  , \wishbone_bd_ram_mem2_reg[32][20]/P0001  , \wishbone_bd_ram_mem2_reg[32][21]/P0001  , \wishbone_bd_ram_mem2_reg[32][22]/P0001  , \wishbone_bd_ram_mem2_reg[32][23]/P0001  , \wishbone_bd_ram_mem2_reg[33][16]/P0001  , \wishbone_bd_ram_mem2_reg[33][17]/P0001  , \wishbone_bd_ram_mem2_reg[33][18]/P0001  , \wishbone_bd_ram_mem2_reg[33][19]/P0001  , \wishbone_bd_ram_mem2_reg[33][20]/P0001  , \wishbone_bd_ram_mem2_reg[33][21]/P0001  , \wishbone_bd_ram_mem2_reg[33][22]/P0001  , \wishbone_bd_ram_mem2_reg[33][23]/P0001  , \wishbone_bd_ram_mem2_reg[34][16]/P0001  , \wishbone_bd_ram_mem2_reg[34][17]/P0001  , \wishbone_bd_ram_mem2_reg[34][18]/P0001  , \wishbone_bd_ram_mem2_reg[34][19]/P0001  , \wishbone_bd_ram_mem2_reg[34][20]/P0001  , \wishbone_bd_ram_mem2_reg[34][21]/P0001  , \wishbone_bd_ram_mem2_reg[34][22]/P0001  , \wishbone_bd_ram_mem2_reg[34][23]/P0001  , \wishbone_bd_ram_mem2_reg[35][16]/P0001  , \wishbone_bd_ram_mem2_reg[35][17]/P0001  , \wishbone_bd_ram_mem2_reg[35][18]/P0001  , \wishbone_bd_ram_mem2_reg[35][19]/P0001  , \wishbone_bd_ram_mem2_reg[35][20]/P0001  , \wishbone_bd_ram_mem2_reg[35][21]/P0001  , \wishbone_bd_ram_mem2_reg[35][22]/P0001  , \wishbone_bd_ram_mem2_reg[35][23]/P0001  , \wishbone_bd_ram_mem2_reg[36][16]/P0001  , \wishbone_bd_ram_mem2_reg[36][17]/P0001  , \wishbone_bd_ram_mem2_reg[36][18]/P0001  , \wishbone_bd_ram_mem2_reg[36][19]/P0001  , \wishbone_bd_ram_mem2_reg[36][20]/P0001  , \wishbone_bd_ram_mem2_reg[36][21]/P0001  , \wishbone_bd_ram_mem2_reg[36][22]/P0001  , \wishbone_bd_ram_mem2_reg[36][23]/P0001  , \wishbone_bd_ram_mem2_reg[37][16]/P0001  , \wishbone_bd_ram_mem2_reg[37][17]/P0001  , \wishbone_bd_ram_mem2_reg[37][18]/P0001  , \wishbone_bd_ram_mem2_reg[37][19]/P0001  , \wishbone_bd_ram_mem2_reg[37][20]/P0001  , \wishbone_bd_ram_mem2_reg[37][21]/P0001  , \wishbone_bd_ram_mem2_reg[37][22]/P0001  , \wishbone_bd_ram_mem2_reg[37][23]/P0001  , \wishbone_bd_ram_mem2_reg[38][16]/P0001  , \wishbone_bd_ram_mem2_reg[38][17]/P0001  , \wishbone_bd_ram_mem2_reg[38][18]/P0001  , \wishbone_bd_ram_mem2_reg[38][19]/P0001  , \wishbone_bd_ram_mem2_reg[38][20]/P0001  , \wishbone_bd_ram_mem2_reg[38][21]/P0001  , \wishbone_bd_ram_mem2_reg[38][22]/P0001  , \wishbone_bd_ram_mem2_reg[38][23]/P0001  , \wishbone_bd_ram_mem2_reg[39][16]/P0001  , \wishbone_bd_ram_mem2_reg[39][17]/P0001  , \wishbone_bd_ram_mem2_reg[39][18]/P0001  , \wishbone_bd_ram_mem2_reg[39][19]/P0001  , \wishbone_bd_ram_mem2_reg[39][20]/P0001  , \wishbone_bd_ram_mem2_reg[39][21]/P0001  , \wishbone_bd_ram_mem2_reg[39][22]/P0001  , \wishbone_bd_ram_mem2_reg[39][23]/P0001  , \wishbone_bd_ram_mem2_reg[3][16]/P0001  , \wishbone_bd_ram_mem2_reg[3][17]/P0001  , \wishbone_bd_ram_mem2_reg[3][18]/P0001  , \wishbone_bd_ram_mem2_reg[3][19]/P0001  , \wishbone_bd_ram_mem2_reg[3][20]/P0001  , \wishbone_bd_ram_mem2_reg[3][21]/P0001  , \wishbone_bd_ram_mem2_reg[3][22]/P0001  , \wishbone_bd_ram_mem2_reg[3][23]/P0001  , \wishbone_bd_ram_mem2_reg[40][16]/P0001  , \wishbone_bd_ram_mem2_reg[40][17]/P0001  , \wishbone_bd_ram_mem2_reg[40][18]/P0001  , \wishbone_bd_ram_mem2_reg[40][19]/P0001  , \wishbone_bd_ram_mem2_reg[40][20]/P0001  , \wishbone_bd_ram_mem2_reg[40][21]/P0001  , \wishbone_bd_ram_mem2_reg[40][22]/P0001  , \wishbone_bd_ram_mem2_reg[40][23]/P0001  , \wishbone_bd_ram_mem2_reg[41][16]/P0001  , \wishbone_bd_ram_mem2_reg[41][17]/P0001  , \wishbone_bd_ram_mem2_reg[41][18]/P0001  , \wishbone_bd_ram_mem2_reg[41][19]/P0001  , \wishbone_bd_ram_mem2_reg[41][20]/P0001  , \wishbone_bd_ram_mem2_reg[41][21]/P0001  , \wishbone_bd_ram_mem2_reg[41][22]/P0001  , \wishbone_bd_ram_mem2_reg[41][23]/P0001  , \wishbone_bd_ram_mem2_reg[42][16]/P0001  , \wishbone_bd_ram_mem2_reg[42][17]/P0001  , \wishbone_bd_ram_mem2_reg[42][18]/P0001  , \wishbone_bd_ram_mem2_reg[42][19]/P0001  , \wishbone_bd_ram_mem2_reg[42][20]/P0001  , \wishbone_bd_ram_mem2_reg[42][21]/P0001  , \wishbone_bd_ram_mem2_reg[42][22]/P0001  , \wishbone_bd_ram_mem2_reg[42][23]/P0001  , \wishbone_bd_ram_mem2_reg[43][16]/P0001  , \wishbone_bd_ram_mem2_reg[43][17]/P0001  , \wishbone_bd_ram_mem2_reg[43][18]/P0001  , \wishbone_bd_ram_mem2_reg[43][19]/P0001  , \wishbone_bd_ram_mem2_reg[43][20]/P0001  , \wishbone_bd_ram_mem2_reg[43][21]/P0001  , \wishbone_bd_ram_mem2_reg[43][22]/P0001  , \wishbone_bd_ram_mem2_reg[43][23]/P0001  , \wishbone_bd_ram_mem2_reg[44][16]/P0001  , \wishbone_bd_ram_mem2_reg[44][17]/P0001  , \wishbone_bd_ram_mem2_reg[44][18]/P0001  , \wishbone_bd_ram_mem2_reg[44][19]/P0001  , \wishbone_bd_ram_mem2_reg[44][20]/P0001  , \wishbone_bd_ram_mem2_reg[44][21]/P0001  , \wishbone_bd_ram_mem2_reg[44][22]/P0001  , \wishbone_bd_ram_mem2_reg[44][23]/P0001  , \wishbone_bd_ram_mem2_reg[45][16]/P0001  , \wishbone_bd_ram_mem2_reg[45][17]/P0001  , \wishbone_bd_ram_mem2_reg[45][18]/P0001  , \wishbone_bd_ram_mem2_reg[45][19]/P0001  , \wishbone_bd_ram_mem2_reg[45][20]/P0001  , \wishbone_bd_ram_mem2_reg[45][21]/P0001  , \wishbone_bd_ram_mem2_reg[45][22]/P0001  , \wishbone_bd_ram_mem2_reg[45][23]/P0001  , \wishbone_bd_ram_mem2_reg[46][16]/P0001  , \wishbone_bd_ram_mem2_reg[46][17]/P0001  , \wishbone_bd_ram_mem2_reg[46][18]/P0001  , \wishbone_bd_ram_mem2_reg[46][19]/P0001  , \wishbone_bd_ram_mem2_reg[46][20]/P0001  , \wishbone_bd_ram_mem2_reg[46][21]/P0001  , \wishbone_bd_ram_mem2_reg[46][22]/P0001  , \wishbone_bd_ram_mem2_reg[46][23]/P0001  , \wishbone_bd_ram_mem2_reg[47][16]/P0001  , \wishbone_bd_ram_mem2_reg[47][17]/P0001  , \wishbone_bd_ram_mem2_reg[47][18]/P0001  , \wishbone_bd_ram_mem2_reg[47][19]/P0001  , \wishbone_bd_ram_mem2_reg[47][20]/P0001  , \wishbone_bd_ram_mem2_reg[47][21]/P0001  , \wishbone_bd_ram_mem2_reg[47][22]/P0001  , \wishbone_bd_ram_mem2_reg[47][23]/P0001  , \wishbone_bd_ram_mem2_reg[48][16]/P0001  , \wishbone_bd_ram_mem2_reg[48][17]/P0001  , \wishbone_bd_ram_mem2_reg[48][18]/P0001  , \wishbone_bd_ram_mem2_reg[48][19]/P0001  , \wishbone_bd_ram_mem2_reg[48][20]/P0001  , \wishbone_bd_ram_mem2_reg[48][21]/P0001  , \wishbone_bd_ram_mem2_reg[48][22]/P0001  , \wishbone_bd_ram_mem2_reg[48][23]/P0001  , \wishbone_bd_ram_mem2_reg[49][16]/P0001  , \wishbone_bd_ram_mem2_reg[49][17]/P0001  , \wishbone_bd_ram_mem2_reg[49][18]/P0001  , \wishbone_bd_ram_mem2_reg[49][19]/P0001  , \wishbone_bd_ram_mem2_reg[49][20]/P0001  , \wishbone_bd_ram_mem2_reg[49][21]/P0001  , \wishbone_bd_ram_mem2_reg[49][22]/P0001  , \wishbone_bd_ram_mem2_reg[49][23]/P0001  , \wishbone_bd_ram_mem2_reg[4][16]/P0001  , \wishbone_bd_ram_mem2_reg[4][17]/P0001  , \wishbone_bd_ram_mem2_reg[4][18]/P0001  , \wishbone_bd_ram_mem2_reg[4][19]/P0001  , \wishbone_bd_ram_mem2_reg[4][20]/P0001  , \wishbone_bd_ram_mem2_reg[4][21]/P0001  , \wishbone_bd_ram_mem2_reg[4][22]/P0001  , \wishbone_bd_ram_mem2_reg[4][23]/P0001  , \wishbone_bd_ram_mem2_reg[50][16]/P0001  , \wishbone_bd_ram_mem2_reg[50][17]/P0001  , \wishbone_bd_ram_mem2_reg[50][18]/P0001  , \wishbone_bd_ram_mem2_reg[50][19]/P0001  , \wishbone_bd_ram_mem2_reg[50][20]/P0001  , \wishbone_bd_ram_mem2_reg[50][21]/P0001  , \wishbone_bd_ram_mem2_reg[50][22]/P0001  , \wishbone_bd_ram_mem2_reg[50][23]/P0001  , \wishbone_bd_ram_mem2_reg[51][16]/P0001  , \wishbone_bd_ram_mem2_reg[51][17]/P0001  , \wishbone_bd_ram_mem2_reg[51][18]/P0001  , \wishbone_bd_ram_mem2_reg[51][19]/P0001  , \wishbone_bd_ram_mem2_reg[51][20]/P0001  , \wishbone_bd_ram_mem2_reg[51][21]/P0001  , \wishbone_bd_ram_mem2_reg[51][22]/P0001  , \wishbone_bd_ram_mem2_reg[51][23]/P0001  , \wishbone_bd_ram_mem2_reg[52][16]/P0001  , \wishbone_bd_ram_mem2_reg[52][17]/P0001  , \wishbone_bd_ram_mem2_reg[52][18]/P0001  , \wishbone_bd_ram_mem2_reg[52][19]/P0001  , \wishbone_bd_ram_mem2_reg[52][20]/P0001  , \wishbone_bd_ram_mem2_reg[52][21]/P0001  , \wishbone_bd_ram_mem2_reg[52][22]/P0001  , \wishbone_bd_ram_mem2_reg[52][23]/P0001  , \wishbone_bd_ram_mem2_reg[53][16]/P0001  , \wishbone_bd_ram_mem2_reg[53][17]/P0001  , \wishbone_bd_ram_mem2_reg[53][18]/P0001  , \wishbone_bd_ram_mem2_reg[53][19]/P0001  , \wishbone_bd_ram_mem2_reg[53][20]/P0001  , \wishbone_bd_ram_mem2_reg[53][21]/P0001  , \wishbone_bd_ram_mem2_reg[53][22]/P0001  , \wishbone_bd_ram_mem2_reg[53][23]/P0001  , \wishbone_bd_ram_mem2_reg[54][16]/P0001  , \wishbone_bd_ram_mem2_reg[54][17]/P0001  , \wishbone_bd_ram_mem2_reg[54][18]/P0001  , \wishbone_bd_ram_mem2_reg[54][19]/P0001  , \wishbone_bd_ram_mem2_reg[54][20]/P0001  , \wishbone_bd_ram_mem2_reg[54][21]/P0001  , \wishbone_bd_ram_mem2_reg[54][22]/P0001  , \wishbone_bd_ram_mem2_reg[54][23]/P0001  , \wishbone_bd_ram_mem2_reg[55][16]/P0001  , \wishbone_bd_ram_mem2_reg[55][17]/P0001  , \wishbone_bd_ram_mem2_reg[55][18]/P0001  , \wishbone_bd_ram_mem2_reg[55][19]/P0001  , \wishbone_bd_ram_mem2_reg[55][20]/P0001  , \wishbone_bd_ram_mem2_reg[55][21]/P0001  , \wishbone_bd_ram_mem2_reg[55][22]/P0001  , \wishbone_bd_ram_mem2_reg[55][23]/P0001  , \wishbone_bd_ram_mem2_reg[56][16]/P0001  , \wishbone_bd_ram_mem2_reg[56][17]/P0001  , \wishbone_bd_ram_mem2_reg[56][18]/P0001  , \wishbone_bd_ram_mem2_reg[56][19]/P0001  , \wishbone_bd_ram_mem2_reg[56][20]/P0001  , \wishbone_bd_ram_mem2_reg[56][21]/P0001  , \wishbone_bd_ram_mem2_reg[56][22]/P0001  , \wishbone_bd_ram_mem2_reg[56][23]/P0001  , \wishbone_bd_ram_mem2_reg[57][16]/P0001  , \wishbone_bd_ram_mem2_reg[57][17]/P0001  , \wishbone_bd_ram_mem2_reg[57][18]/P0001  , \wishbone_bd_ram_mem2_reg[57][19]/P0001  , \wishbone_bd_ram_mem2_reg[57][20]/P0001  , \wishbone_bd_ram_mem2_reg[57][21]/P0001  , \wishbone_bd_ram_mem2_reg[57][22]/P0001  , \wishbone_bd_ram_mem2_reg[57][23]/P0001  , \wishbone_bd_ram_mem2_reg[58][16]/P0001  , \wishbone_bd_ram_mem2_reg[58][17]/P0001  , \wishbone_bd_ram_mem2_reg[58][18]/P0001  , \wishbone_bd_ram_mem2_reg[58][19]/P0001  , \wishbone_bd_ram_mem2_reg[58][20]/P0001  , \wishbone_bd_ram_mem2_reg[58][21]/P0001  , \wishbone_bd_ram_mem2_reg[58][22]/P0001  , \wishbone_bd_ram_mem2_reg[58][23]/P0001  , \wishbone_bd_ram_mem2_reg[59][16]/P0001  , \wishbone_bd_ram_mem2_reg[59][17]/P0001  , \wishbone_bd_ram_mem2_reg[59][18]/P0001  , \wishbone_bd_ram_mem2_reg[59][19]/P0001  , \wishbone_bd_ram_mem2_reg[59][20]/P0001  , \wishbone_bd_ram_mem2_reg[59][21]/P0001  , \wishbone_bd_ram_mem2_reg[59][22]/P0001  , \wishbone_bd_ram_mem2_reg[59][23]/P0001  , \wishbone_bd_ram_mem2_reg[5][16]/P0001  , \wishbone_bd_ram_mem2_reg[5][17]/P0001  , \wishbone_bd_ram_mem2_reg[5][18]/P0001  , \wishbone_bd_ram_mem2_reg[5][19]/P0001  , \wishbone_bd_ram_mem2_reg[5][20]/P0001  , \wishbone_bd_ram_mem2_reg[5][21]/P0001  , \wishbone_bd_ram_mem2_reg[5][22]/P0001  , \wishbone_bd_ram_mem2_reg[5][23]/P0001  , \wishbone_bd_ram_mem2_reg[60][16]/P0001  , \wishbone_bd_ram_mem2_reg[60][17]/P0001  , \wishbone_bd_ram_mem2_reg[60][18]/P0001  , \wishbone_bd_ram_mem2_reg[60][19]/P0001  , \wishbone_bd_ram_mem2_reg[60][20]/P0001  , \wishbone_bd_ram_mem2_reg[60][21]/P0001  , \wishbone_bd_ram_mem2_reg[60][22]/P0001  , \wishbone_bd_ram_mem2_reg[60][23]/P0001  , \wishbone_bd_ram_mem2_reg[61][16]/P0001  , \wishbone_bd_ram_mem2_reg[61][17]/P0001  , \wishbone_bd_ram_mem2_reg[61][18]/P0001  , \wishbone_bd_ram_mem2_reg[61][19]/P0001  , \wishbone_bd_ram_mem2_reg[61][20]/P0001  , \wishbone_bd_ram_mem2_reg[61][21]/P0001  , \wishbone_bd_ram_mem2_reg[61][22]/P0001  , \wishbone_bd_ram_mem2_reg[61][23]/P0001  , \wishbone_bd_ram_mem2_reg[62][16]/P0001  , \wishbone_bd_ram_mem2_reg[62][17]/P0001  , \wishbone_bd_ram_mem2_reg[62][18]/P0001  , \wishbone_bd_ram_mem2_reg[62][19]/P0001  , \wishbone_bd_ram_mem2_reg[62][20]/P0001  , \wishbone_bd_ram_mem2_reg[62][21]/P0001  , \wishbone_bd_ram_mem2_reg[62][22]/P0001  , \wishbone_bd_ram_mem2_reg[62][23]/P0001  , \wishbone_bd_ram_mem2_reg[63][16]/P0001  , \wishbone_bd_ram_mem2_reg[63][17]/P0001  , \wishbone_bd_ram_mem2_reg[63][18]/P0001  , \wishbone_bd_ram_mem2_reg[63][19]/P0001  , \wishbone_bd_ram_mem2_reg[63][20]/P0001  , \wishbone_bd_ram_mem2_reg[63][21]/P0001  , \wishbone_bd_ram_mem2_reg[63][22]/P0001  , \wishbone_bd_ram_mem2_reg[63][23]/P0001  , \wishbone_bd_ram_mem2_reg[64][16]/P0001  , \wishbone_bd_ram_mem2_reg[64][17]/P0001  , \wishbone_bd_ram_mem2_reg[64][18]/P0001  , \wishbone_bd_ram_mem2_reg[64][19]/P0001  , \wishbone_bd_ram_mem2_reg[64][20]/P0001  , \wishbone_bd_ram_mem2_reg[64][21]/P0001  , \wishbone_bd_ram_mem2_reg[64][22]/P0001  , \wishbone_bd_ram_mem2_reg[64][23]/P0001  , \wishbone_bd_ram_mem2_reg[65][16]/P0001  , \wishbone_bd_ram_mem2_reg[65][17]/P0001  , \wishbone_bd_ram_mem2_reg[65][18]/P0001  , \wishbone_bd_ram_mem2_reg[65][19]/P0001  , \wishbone_bd_ram_mem2_reg[65][20]/P0001  , \wishbone_bd_ram_mem2_reg[65][21]/P0001  , \wishbone_bd_ram_mem2_reg[65][22]/P0001  , \wishbone_bd_ram_mem2_reg[65][23]/P0001  , \wishbone_bd_ram_mem2_reg[66][16]/P0001  , \wishbone_bd_ram_mem2_reg[66][17]/P0001  , \wishbone_bd_ram_mem2_reg[66][18]/P0001  , \wishbone_bd_ram_mem2_reg[66][19]/P0001  , \wishbone_bd_ram_mem2_reg[66][20]/P0001  , \wishbone_bd_ram_mem2_reg[66][21]/P0001  , \wishbone_bd_ram_mem2_reg[66][22]/P0001  , \wishbone_bd_ram_mem2_reg[66][23]/P0001  , \wishbone_bd_ram_mem2_reg[67][16]/P0001  , \wishbone_bd_ram_mem2_reg[67][17]/P0001  , \wishbone_bd_ram_mem2_reg[67][18]/P0001  , \wishbone_bd_ram_mem2_reg[67][19]/P0001  , \wishbone_bd_ram_mem2_reg[67][20]/P0001  , \wishbone_bd_ram_mem2_reg[67][21]/P0001  , \wishbone_bd_ram_mem2_reg[67][22]/P0001  , \wishbone_bd_ram_mem2_reg[67][23]/P0001  , \wishbone_bd_ram_mem2_reg[68][16]/P0001  , \wishbone_bd_ram_mem2_reg[68][17]/P0001  , \wishbone_bd_ram_mem2_reg[68][18]/P0001  , \wishbone_bd_ram_mem2_reg[68][19]/P0001  , \wishbone_bd_ram_mem2_reg[68][20]/P0001  , \wishbone_bd_ram_mem2_reg[68][21]/P0001  , \wishbone_bd_ram_mem2_reg[68][22]/P0001  , \wishbone_bd_ram_mem2_reg[68][23]/P0001  , \wishbone_bd_ram_mem2_reg[69][16]/P0001  , \wishbone_bd_ram_mem2_reg[69][17]/P0001  , \wishbone_bd_ram_mem2_reg[69][18]/P0001  , \wishbone_bd_ram_mem2_reg[69][19]/P0001  , \wishbone_bd_ram_mem2_reg[69][20]/P0001  , \wishbone_bd_ram_mem2_reg[69][21]/P0001  , \wishbone_bd_ram_mem2_reg[69][22]/P0001  , \wishbone_bd_ram_mem2_reg[69][23]/P0001  , \wishbone_bd_ram_mem2_reg[6][16]/P0001  , \wishbone_bd_ram_mem2_reg[6][17]/P0001  , \wishbone_bd_ram_mem2_reg[6][18]/P0001  , \wishbone_bd_ram_mem2_reg[6][19]/P0001  , \wishbone_bd_ram_mem2_reg[6][20]/P0001  , \wishbone_bd_ram_mem2_reg[6][21]/P0001  , \wishbone_bd_ram_mem2_reg[6][22]/P0001  , \wishbone_bd_ram_mem2_reg[6][23]/P0001  , \wishbone_bd_ram_mem2_reg[70][16]/P0001  , \wishbone_bd_ram_mem2_reg[70][17]/P0001  , \wishbone_bd_ram_mem2_reg[70][18]/P0001  , \wishbone_bd_ram_mem2_reg[70][19]/P0001  , \wishbone_bd_ram_mem2_reg[70][20]/P0001  , \wishbone_bd_ram_mem2_reg[70][21]/P0001  , \wishbone_bd_ram_mem2_reg[70][22]/P0001  , \wishbone_bd_ram_mem2_reg[70][23]/P0001  , \wishbone_bd_ram_mem2_reg[71][16]/P0001  , \wishbone_bd_ram_mem2_reg[71][17]/P0001  , \wishbone_bd_ram_mem2_reg[71][18]/P0001  , \wishbone_bd_ram_mem2_reg[71][19]/P0001  , \wishbone_bd_ram_mem2_reg[71][20]/P0001  , \wishbone_bd_ram_mem2_reg[71][21]/P0001  , \wishbone_bd_ram_mem2_reg[71][22]/P0001  , \wishbone_bd_ram_mem2_reg[71][23]/P0001  , \wishbone_bd_ram_mem2_reg[72][16]/P0001  , \wishbone_bd_ram_mem2_reg[72][17]/P0001  , \wishbone_bd_ram_mem2_reg[72][18]/P0001  , \wishbone_bd_ram_mem2_reg[72][19]/P0001  , \wishbone_bd_ram_mem2_reg[72][20]/P0001  , \wishbone_bd_ram_mem2_reg[72][21]/P0001  , \wishbone_bd_ram_mem2_reg[72][22]/P0001  , \wishbone_bd_ram_mem2_reg[72][23]/P0001  , \wishbone_bd_ram_mem2_reg[73][16]/P0001  , \wishbone_bd_ram_mem2_reg[73][17]/P0001  , \wishbone_bd_ram_mem2_reg[73][18]/P0001  , \wishbone_bd_ram_mem2_reg[73][19]/P0001  , \wishbone_bd_ram_mem2_reg[73][20]/P0001  , \wishbone_bd_ram_mem2_reg[73][21]/P0001  , \wishbone_bd_ram_mem2_reg[73][22]/P0001  , \wishbone_bd_ram_mem2_reg[73][23]/P0001  , \wishbone_bd_ram_mem2_reg[74][16]/P0001  , \wishbone_bd_ram_mem2_reg[74][17]/P0001  , \wishbone_bd_ram_mem2_reg[74][18]/P0001  , \wishbone_bd_ram_mem2_reg[74][19]/P0001  , \wishbone_bd_ram_mem2_reg[74][20]/P0001  , \wishbone_bd_ram_mem2_reg[74][21]/P0001  , \wishbone_bd_ram_mem2_reg[74][22]/P0001  , \wishbone_bd_ram_mem2_reg[74][23]/P0001  , \wishbone_bd_ram_mem2_reg[75][16]/P0001  , \wishbone_bd_ram_mem2_reg[75][17]/P0001  , \wishbone_bd_ram_mem2_reg[75][18]/P0001  , \wishbone_bd_ram_mem2_reg[75][19]/P0001  , \wishbone_bd_ram_mem2_reg[75][20]/P0001  , \wishbone_bd_ram_mem2_reg[75][21]/P0001  , \wishbone_bd_ram_mem2_reg[75][22]/P0001  , \wishbone_bd_ram_mem2_reg[75][23]/P0001  , \wishbone_bd_ram_mem2_reg[76][16]/P0001  , \wishbone_bd_ram_mem2_reg[76][17]/P0001  , \wishbone_bd_ram_mem2_reg[76][18]/P0001  , \wishbone_bd_ram_mem2_reg[76][19]/P0001  , \wishbone_bd_ram_mem2_reg[76][20]/P0001  , \wishbone_bd_ram_mem2_reg[76][21]/P0001  , \wishbone_bd_ram_mem2_reg[76][22]/P0001  , \wishbone_bd_ram_mem2_reg[76][23]/P0001  , \wishbone_bd_ram_mem2_reg[77][16]/P0001  , \wishbone_bd_ram_mem2_reg[77][17]/P0001  , \wishbone_bd_ram_mem2_reg[77][18]/P0001  , \wishbone_bd_ram_mem2_reg[77][19]/P0001  , \wishbone_bd_ram_mem2_reg[77][20]/P0001  , \wishbone_bd_ram_mem2_reg[77][21]/P0001  , \wishbone_bd_ram_mem2_reg[77][22]/P0001  , \wishbone_bd_ram_mem2_reg[77][23]/P0001  , \wishbone_bd_ram_mem2_reg[78][16]/P0001  , \wishbone_bd_ram_mem2_reg[78][17]/P0001  , \wishbone_bd_ram_mem2_reg[78][18]/P0001  , \wishbone_bd_ram_mem2_reg[78][19]/P0001  , \wishbone_bd_ram_mem2_reg[78][20]/P0001  , \wishbone_bd_ram_mem2_reg[78][21]/P0001  , \wishbone_bd_ram_mem2_reg[78][22]/P0001  , \wishbone_bd_ram_mem2_reg[78][23]/P0001  , \wishbone_bd_ram_mem2_reg[79][16]/P0001  , \wishbone_bd_ram_mem2_reg[79][17]/P0001  , \wishbone_bd_ram_mem2_reg[79][18]/P0001  , \wishbone_bd_ram_mem2_reg[79][19]/P0001  , \wishbone_bd_ram_mem2_reg[79][20]/P0001  , \wishbone_bd_ram_mem2_reg[79][21]/P0001  , \wishbone_bd_ram_mem2_reg[79][22]/P0001  , \wishbone_bd_ram_mem2_reg[79][23]/P0001  , \wishbone_bd_ram_mem2_reg[7][16]/P0001  , \wishbone_bd_ram_mem2_reg[7][17]/P0001  , \wishbone_bd_ram_mem2_reg[7][18]/P0001  , \wishbone_bd_ram_mem2_reg[7][19]/P0001  , \wishbone_bd_ram_mem2_reg[7][20]/P0001  , \wishbone_bd_ram_mem2_reg[7][21]/P0001  , \wishbone_bd_ram_mem2_reg[7][22]/P0001  , \wishbone_bd_ram_mem2_reg[7][23]/P0001  , \wishbone_bd_ram_mem2_reg[80][16]/P0001  , \wishbone_bd_ram_mem2_reg[80][17]/P0001  , \wishbone_bd_ram_mem2_reg[80][18]/P0001  , \wishbone_bd_ram_mem2_reg[80][19]/P0001  , \wishbone_bd_ram_mem2_reg[80][20]/P0001  , \wishbone_bd_ram_mem2_reg[80][21]/P0001  , \wishbone_bd_ram_mem2_reg[80][22]/P0001  , \wishbone_bd_ram_mem2_reg[80][23]/P0001  , \wishbone_bd_ram_mem2_reg[81][16]/P0001  , \wishbone_bd_ram_mem2_reg[81][17]/P0001  , \wishbone_bd_ram_mem2_reg[81][18]/P0001  , \wishbone_bd_ram_mem2_reg[81][19]/P0001  , \wishbone_bd_ram_mem2_reg[81][20]/P0001  , \wishbone_bd_ram_mem2_reg[81][21]/P0001  , \wishbone_bd_ram_mem2_reg[81][22]/P0001  , \wishbone_bd_ram_mem2_reg[81][23]/P0001  , \wishbone_bd_ram_mem2_reg[82][16]/P0001  , \wishbone_bd_ram_mem2_reg[82][17]/P0001  , \wishbone_bd_ram_mem2_reg[82][18]/P0001  , \wishbone_bd_ram_mem2_reg[82][19]/P0001  , \wishbone_bd_ram_mem2_reg[82][20]/P0001  , \wishbone_bd_ram_mem2_reg[82][21]/P0001  , \wishbone_bd_ram_mem2_reg[82][22]/P0001  , \wishbone_bd_ram_mem2_reg[82][23]/P0001  , \wishbone_bd_ram_mem2_reg[83][16]/P0001  , \wishbone_bd_ram_mem2_reg[83][17]/P0001  , \wishbone_bd_ram_mem2_reg[83][18]/P0001  , \wishbone_bd_ram_mem2_reg[83][19]/P0001  , \wishbone_bd_ram_mem2_reg[83][20]/P0001  , \wishbone_bd_ram_mem2_reg[83][21]/P0001  , \wishbone_bd_ram_mem2_reg[83][22]/P0001  , \wishbone_bd_ram_mem2_reg[83][23]/P0001  , \wishbone_bd_ram_mem2_reg[84][16]/P0001  , \wishbone_bd_ram_mem2_reg[84][17]/P0001  , \wishbone_bd_ram_mem2_reg[84][18]/P0001  , \wishbone_bd_ram_mem2_reg[84][19]/P0001  , \wishbone_bd_ram_mem2_reg[84][20]/P0001  , \wishbone_bd_ram_mem2_reg[84][21]/P0001  , \wishbone_bd_ram_mem2_reg[84][22]/P0001  , \wishbone_bd_ram_mem2_reg[84][23]/P0001  , \wishbone_bd_ram_mem2_reg[85][16]/P0001  , \wishbone_bd_ram_mem2_reg[85][17]/P0001  , \wishbone_bd_ram_mem2_reg[85][18]/P0001  , \wishbone_bd_ram_mem2_reg[85][19]/P0001  , \wishbone_bd_ram_mem2_reg[85][20]/P0001  , \wishbone_bd_ram_mem2_reg[85][21]/P0001  , \wishbone_bd_ram_mem2_reg[85][22]/P0001  , \wishbone_bd_ram_mem2_reg[85][23]/P0001  , \wishbone_bd_ram_mem2_reg[86][16]/P0001  , \wishbone_bd_ram_mem2_reg[86][17]/P0001  , \wishbone_bd_ram_mem2_reg[86][18]/P0001  , \wishbone_bd_ram_mem2_reg[86][19]/P0001  , \wishbone_bd_ram_mem2_reg[86][20]/P0001  , \wishbone_bd_ram_mem2_reg[86][21]/P0001  , \wishbone_bd_ram_mem2_reg[86][22]/P0001  , \wishbone_bd_ram_mem2_reg[86][23]/P0001  , \wishbone_bd_ram_mem2_reg[87][16]/P0001  , \wishbone_bd_ram_mem2_reg[87][17]/P0001  , \wishbone_bd_ram_mem2_reg[87][18]/P0001  , \wishbone_bd_ram_mem2_reg[87][19]/P0001  , \wishbone_bd_ram_mem2_reg[87][20]/P0001  , \wishbone_bd_ram_mem2_reg[87][21]/P0001  , \wishbone_bd_ram_mem2_reg[87][22]/P0001  , \wishbone_bd_ram_mem2_reg[87][23]/P0001  , \wishbone_bd_ram_mem2_reg[88][16]/P0001  , \wishbone_bd_ram_mem2_reg[88][17]/P0001  , \wishbone_bd_ram_mem2_reg[88][18]/P0001  , \wishbone_bd_ram_mem2_reg[88][19]/P0001  , \wishbone_bd_ram_mem2_reg[88][20]/P0001  , \wishbone_bd_ram_mem2_reg[88][21]/P0001  , \wishbone_bd_ram_mem2_reg[88][22]/P0001  , \wishbone_bd_ram_mem2_reg[88][23]/P0001  , \wishbone_bd_ram_mem2_reg[89][16]/P0001  , \wishbone_bd_ram_mem2_reg[89][17]/P0001  , \wishbone_bd_ram_mem2_reg[89][18]/P0001  , \wishbone_bd_ram_mem2_reg[89][19]/P0001  , \wishbone_bd_ram_mem2_reg[89][20]/P0001  , \wishbone_bd_ram_mem2_reg[89][21]/P0001  , \wishbone_bd_ram_mem2_reg[89][22]/P0001  , \wishbone_bd_ram_mem2_reg[89][23]/P0001  , \wishbone_bd_ram_mem2_reg[8][16]/P0001  , \wishbone_bd_ram_mem2_reg[8][17]/P0001  , \wishbone_bd_ram_mem2_reg[8][18]/P0001  , \wishbone_bd_ram_mem2_reg[8][19]/P0001  , \wishbone_bd_ram_mem2_reg[8][20]/P0001  , \wishbone_bd_ram_mem2_reg[8][21]/P0001  , \wishbone_bd_ram_mem2_reg[8][22]/P0001  , \wishbone_bd_ram_mem2_reg[8][23]/P0001  , \wishbone_bd_ram_mem2_reg[90][16]/P0001  , \wishbone_bd_ram_mem2_reg[90][17]/P0001  , \wishbone_bd_ram_mem2_reg[90][18]/P0001  , \wishbone_bd_ram_mem2_reg[90][19]/P0001  , \wishbone_bd_ram_mem2_reg[90][20]/P0001  , \wishbone_bd_ram_mem2_reg[90][21]/P0001  , \wishbone_bd_ram_mem2_reg[90][22]/P0001  , \wishbone_bd_ram_mem2_reg[90][23]/P0001  , \wishbone_bd_ram_mem2_reg[91][16]/P0001  , \wishbone_bd_ram_mem2_reg[91][17]/P0001  , \wishbone_bd_ram_mem2_reg[91][18]/P0001  , \wishbone_bd_ram_mem2_reg[91][19]/P0001  , \wishbone_bd_ram_mem2_reg[91][20]/P0001  , \wishbone_bd_ram_mem2_reg[91][21]/P0001  , \wishbone_bd_ram_mem2_reg[91][22]/P0001  , \wishbone_bd_ram_mem2_reg[91][23]/P0001  , \wishbone_bd_ram_mem2_reg[92][16]/P0001  , \wishbone_bd_ram_mem2_reg[92][17]/P0001  , \wishbone_bd_ram_mem2_reg[92][18]/P0001  , \wishbone_bd_ram_mem2_reg[92][19]/P0001  , \wishbone_bd_ram_mem2_reg[92][20]/P0001  , \wishbone_bd_ram_mem2_reg[92][21]/P0001  , \wishbone_bd_ram_mem2_reg[92][22]/P0001  , \wishbone_bd_ram_mem2_reg[92][23]/P0001  , \wishbone_bd_ram_mem2_reg[93][16]/P0001  , \wishbone_bd_ram_mem2_reg[93][17]/P0001  , \wishbone_bd_ram_mem2_reg[93][18]/P0001  , \wishbone_bd_ram_mem2_reg[93][19]/P0001  , \wishbone_bd_ram_mem2_reg[93][20]/P0001  , \wishbone_bd_ram_mem2_reg[93][21]/P0001  , \wishbone_bd_ram_mem2_reg[93][22]/P0001  , \wishbone_bd_ram_mem2_reg[93][23]/P0001  , \wishbone_bd_ram_mem2_reg[94][16]/P0001  , \wishbone_bd_ram_mem2_reg[94][17]/P0001  , \wishbone_bd_ram_mem2_reg[94][18]/P0001  , \wishbone_bd_ram_mem2_reg[94][19]/P0001  , \wishbone_bd_ram_mem2_reg[94][20]/P0001  , \wishbone_bd_ram_mem2_reg[94][21]/P0001  , \wishbone_bd_ram_mem2_reg[94][22]/P0001  , \wishbone_bd_ram_mem2_reg[94][23]/P0001  , \wishbone_bd_ram_mem2_reg[95][16]/P0001  , \wishbone_bd_ram_mem2_reg[95][17]/P0001  , \wishbone_bd_ram_mem2_reg[95][18]/P0001  , \wishbone_bd_ram_mem2_reg[95][19]/P0001  , \wishbone_bd_ram_mem2_reg[95][20]/P0001  , \wishbone_bd_ram_mem2_reg[95][21]/P0001  , \wishbone_bd_ram_mem2_reg[95][22]/P0001  , \wishbone_bd_ram_mem2_reg[95][23]/P0001  , \wishbone_bd_ram_mem2_reg[96][16]/P0001  , \wishbone_bd_ram_mem2_reg[96][17]/P0001  , \wishbone_bd_ram_mem2_reg[96][18]/P0001  , \wishbone_bd_ram_mem2_reg[96][19]/P0001  , \wishbone_bd_ram_mem2_reg[96][20]/P0001  , \wishbone_bd_ram_mem2_reg[96][21]/P0001  , \wishbone_bd_ram_mem2_reg[96][22]/P0001  , \wishbone_bd_ram_mem2_reg[96][23]/P0001  , \wishbone_bd_ram_mem2_reg[97][16]/P0001  , \wishbone_bd_ram_mem2_reg[97][17]/P0001  , \wishbone_bd_ram_mem2_reg[97][18]/P0001  , \wishbone_bd_ram_mem2_reg[97][19]/P0001  , \wishbone_bd_ram_mem2_reg[97][20]/P0001  , \wishbone_bd_ram_mem2_reg[97][21]/P0001  , \wishbone_bd_ram_mem2_reg[97][22]/P0001  , \wishbone_bd_ram_mem2_reg[97][23]/P0001  , \wishbone_bd_ram_mem2_reg[98][16]/P0001  , \wishbone_bd_ram_mem2_reg[98][17]/P0001  , \wishbone_bd_ram_mem2_reg[98][18]/P0001  , \wishbone_bd_ram_mem2_reg[98][19]/P0001  , \wishbone_bd_ram_mem2_reg[98][20]/P0001  , \wishbone_bd_ram_mem2_reg[98][21]/P0001  , \wishbone_bd_ram_mem2_reg[98][22]/P0001  , \wishbone_bd_ram_mem2_reg[98][23]/P0001  , \wishbone_bd_ram_mem2_reg[99][16]/P0001  , \wishbone_bd_ram_mem2_reg[99][17]/P0001  , \wishbone_bd_ram_mem2_reg[99][18]/P0001  , \wishbone_bd_ram_mem2_reg[99][19]/P0001  , \wishbone_bd_ram_mem2_reg[99][20]/P0001  , \wishbone_bd_ram_mem2_reg[99][21]/P0001  , \wishbone_bd_ram_mem2_reg[99][22]/P0001  , \wishbone_bd_ram_mem2_reg[99][23]/P0001  , \wishbone_bd_ram_mem2_reg[9][16]/P0001  , \wishbone_bd_ram_mem2_reg[9][17]/P0001  , \wishbone_bd_ram_mem2_reg[9][18]/P0001  , \wishbone_bd_ram_mem2_reg[9][19]/P0001  , \wishbone_bd_ram_mem2_reg[9][20]/P0001  , \wishbone_bd_ram_mem2_reg[9][21]/P0001  , \wishbone_bd_ram_mem2_reg[9][22]/P0001  , \wishbone_bd_ram_mem2_reg[9][23]/P0001  , \wishbone_bd_ram_mem3_reg[0][24]/P0001  , \wishbone_bd_ram_mem3_reg[0][25]/P0001  , \wishbone_bd_ram_mem3_reg[0][26]/P0001  , \wishbone_bd_ram_mem3_reg[0][27]/P0001  , \wishbone_bd_ram_mem3_reg[0][28]/P0001  , \wishbone_bd_ram_mem3_reg[0][29]/P0001  , \wishbone_bd_ram_mem3_reg[0][30]/P0001  , \wishbone_bd_ram_mem3_reg[0][31]/P0001  , \wishbone_bd_ram_mem3_reg[100][24]/P0001  , \wishbone_bd_ram_mem3_reg[100][25]/P0001  , \wishbone_bd_ram_mem3_reg[100][26]/P0001  , \wishbone_bd_ram_mem3_reg[100][27]/P0001  , \wishbone_bd_ram_mem3_reg[100][28]/P0001  , \wishbone_bd_ram_mem3_reg[100][29]/P0001  , \wishbone_bd_ram_mem3_reg[100][30]/P0001  , \wishbone_bd_ram_mem3_reg[100][31]/P0001  , \wishbone_bd_ram_mem3_reg[101][24]/P0001  , \wishbone_bd_ram_mem3_reg[101][25]/P0001  , \wishbone_bd_ram_mem3_reg[101][26]/P0001  , \wishbone_bd_ram_mem3_reg[101][27]/P0001  , \wishbone_bd_ram_mem3_reg[101][28]/P0001  , \wishbone_bd_ram_mem3_reg[101][29]/P0001  , \wishbone_bd_ram_mem3_reg[101][30]/P0001  , \wishbone_bd_ram_mem3_reg[101][31]/P0001  , \wishbone_bd_ram_mem3_reg[102][24]/P0001  , \wishbone_bd_ram_mem3_reg[102][25]/P0001  , \wishbone_bd_ram_mem3_reg[102][26]/P0001  , \wishbone_bd_ram_mem3_reg[102][27]/P0001  , \wishbone_bd_ram_mem3_reg[102][28]/P0001  , \wishbone_bd_ram_mem3_reg[102][29]/P0001  , \wishbone_bd_ram_mem3_reg[102][30]/P0001  , \wishbone_bd_ram_mem3_reg[102][31]/P0001  , \wishbone_bd_ram_mem3_reg[103][24]/P0001  , \wishbone_bd_ram_mem3_reg[103][25]/P0001  , \wishbone_bd_ram_mem3_reg[103][26]/P0001  , \wishbone_bd_ram_mem3_reg[103][27]/P0001  , \wishbone_bd_ram_mem3_reg[103][28]/P0001  , \wishbone_bd_ram_mem3_reg[103][29]/P0001  , \wishbone_bd_ram_mem3_reg[103][30]/P0001  , \wishbone_bd_ram_mem3_reg[103][31]/P0001  , \wishbone_bd_ram_mem3_reg[104][24]/P0001  , \wishbone_bd_ram_mem3_reg[104][25]/P0001  , \wishbone_bd_ram_mem3_reg[104][26]/P0001  , \wishbone_bd_ram_mem3_reg[104][27]/P0001  , \wishbone_bd_ram_mem3_reg[104][28]/P0001  , \wishbone_bd_ram_mem3_reg[104][29]/P0001  , \wishbone_bd_ram_mem3_reg[104][30]/P0001  , \wishbone_bd_ram_mem3_reg[104][31]/P0001  , \wishbone_bd_ram_mem3_reg[105][24]/P0001  , \wishbone_bd_ram_mem3_reg[105][25]/P0001  , \wishbone_bd_ram_mem3_reg[105][26]/P0001  , \wishbone_bd_ram_mem3_reg[105][27]/P0001  , \wishbone_bd_ram_mem3_reg[105][28]/P0001  , \wishbone_bd_ram_mem3_reg[105][29]/P0001  , \wishbone_bd_ram_mem3_reg[105][30]/P0001  , \wishbone_bd_ram_mem3_reg[105][31]/P0001  , \wishbone_bd_ram_mem3_reg[106][24]/P0001  , \wishbone_bd_ram_mem3_reg[106][25]/P0001  , \wishbone_bd_ram_mem3_reg[106][26]/P0001  , \wishbone_bd_ram_mem3_reg[106][27]/P0001  , \wishbone_bd_ram_mem3_reg[106][28]/P0001  , \wishbone_bd_ram_mem3_reg[106][29]/P0001  , \wishbone_bd_ram_mem3_reg[106][30]/P0001  , \wishbone_bd_ram_mem3_reg[106][31]/P0001  , \wishbone_bd_ram_mem3_reg[107][24]/P0001  , \wishbone_bd_ram_mem3_reg[107][25]/P0001  , \wishbone_bd_ram_mem3_reg[107][26]/P0001  , \wishbone_bd_ram_mem3_reg[107][27]/P0001  , \wishbone_bd_ram_mem3_reg[107][28]/P0001  , \wishbone_bd_ram_mem3_reg[107][29]/P0001  , \wishbone_bd_ram_mem3_reg[107][30]/P0001  , \wishbone_bd_ram_mem3_reg[107][31]/P0001  , \wishbone_bd_ram_mem3_reg[108][24]/P0001  , \wishbone_bd_ram_mem3_reg[108][25]/P0001  , \wishbone_bd_ram_mem3_reg[108][26]/P0001  , \wishbone_bd_ram_mem3_reg[108][27]/P0001  , \wishbone_bd_ram_mem3_reg[108][28]/P0001  , \wishbone_bd_ram_mem3_reg[108][29]/P0001  , \wishbone_bd_ram_mem3_reg[108][30]/P0001  , \wishbone_bd_ram_mem3_reg[108][31]/P0001  , \wishbone_bd_ram_mem3_reg[109][24]/P0001  , \wishbone_bd_ram_mem3_reg[109][25]/P0001  , \wishbone_bd_ram_mem3_reg[109][26]/P0001  , \wishbone_bd_ram_mem3_reg[109][27]/P0001  , \wishbone_bd_ram_mem3_reg[109][28]/P0001  , \wishbone_bd_ram_mem3_reg[109][29]/P0001  , \wishbone_bd_ram_mem3_reg[109][30]/P0001  , \wishbone_bd_ram_mem3_reg[109][31]/P0001  , \wishbone_bd_ram_mem3_reg[10][24]/P0001  , \wishbone_bd_ram_mem3_reg[10][25]/P0001  , \wishbone_bd_ram_mem3_reg[10][26]/P0001  , \wishbone_bd_ram_mem3_reg[10][27]/P0001  , \wishbone_bd_ram_mem3_reg[10][28]/P0001  , \wishbone_bd_ram_mem3_reg[10][29]/P0001  , \wishbone_bd_ram_mem3_reg[10][30]/P0001  , \wishbone_bd_ram_mem3_reg[10][31]/P0001  , \wishbone_bd_ram_mem3_reg[110][24]/P0001  , \wishbone_bd_ram_mem3_reg[110][25]/P0001  , \wishbone_bd_ram_mem3_reg[110][26]/P0001  , \wishbone_bd_ram_mem3_reg[110][27]/P0001  , \wishbone_bd_ram_mem3_reg[110][28]/P0001  , \wishbone_bd_ram_mem3_reg[110][29]/P0001  , \wishbone_bd_ram_mem3_reg[110][30]/P0001  , \wishbone_bd_ram_mem3_reg[110][31]/P0001  , \wishbone_bd_ram_mem3_reg[111][24]/P0001  , \wishbone_bd_ram_mem3_reg[111][25]/P0001  , \wishbone_bd_ram_mem3_reg[111][26]/P0001  , \wishbone_bd_ram_mem3_reg[111][27]/P0001  , \wishbone_bd_ram_mem3_reg[111][28]/P0001  , \wishbone_bd_ram_mem3_reg[111][29]/P0001  , \wishbone_bd_ram_mem3_reg[111][30]/P0001  , \wishbone_bd_ram_mem3_reg[111][31]/P0001  , \wishbone_bd_ram_mem3_reg[112][24]/P0001  , \wishbone_bd_ram_mem3_reg[112][25]/P0001  , \wishbone_bd_ram_mem3_reg[112][26]/P0001  , \wishbone_bd_ram_mem3_reg[112][27]/P0001  , \wishbone_bd_ram_mem3_reg[112][28]/P0001  , \wishbone_bd_ram_mem3_reg[112][29]/P0001  , \wishbone_bd_ram_mem3_reg[112][30]/P0001  , \wishbone_bd_ram_mem3_reg[112][31]/P0001  , \wishbone_bd_ram_mem3_reg[113][24]/P0001  , \wishbone_bd_ram_mem3_reg[113][25]/P0001  , \wishbone_bd_ram_mem3_reg[113][26]/P0001  , \wishbone_bd_ram_mem3_reg[113][27]/P0001  , \wishbone_bd_ram_mem3_reg[113][28]/P0001  , \wishbone_bd_ram_mem3_reg[113][29]/P0001  , \wishbone_bd_ram_mem3_reg[113][30]/P0001  , \wishbone_bd_ram_mem3_reg[113][31]/P0001  , \wishbone_bd_ram_mem3_reg[114][24]/P0001  , \wishbone_bd_ram_mem3_reg[114][25]/P0001  , \wishbone_bd_ram_mem3_reg[114][26]/P0001  , \wishbone_bd_ram_mem3_reg[114][27]/P0001  , \wishbone_bd_ram_mem3_reg[114][28]/P0001  , \wishbone_bd_ram_mem3_reg[114][29]/P0001  , \wishbone_bd_ram_mem3_reg[114][30]/P0001  , \wishbone_bd_ram_mem3_reg[114][31]/P0001  , \wishbone_bd_ram_mem3_reg[115][24]/P0001  , \wishbone_bd_ram_mem3_reg[115][25]/P0001  , \wishbone_bd_ram_mem3_reg[115][26]/P0001  , \wishbone_bd_ram_mem3_reg[115][27]/P0001  , \wishbone_bd_ram_mem3_reg[115][28]/P0001  , \wishbone_bd_ram_mem3_reg[115][29]/P0001  , \wishbone_bd_ram_mem3_reg[115][30]/P0001  , \wishbone_bd_ram_mem3_reg[115][31]/P0001  , \wishbone_bd_ram_mem3_reg[116][24]/P0001  , \wishbone_bd_ram_mem3_reg[116][25]/P0001  , \wishbone_bd_ram_mem3_reg[116][26]/P0001  , \wishbone_bd_ram_mem3_reg[116][27]/P0001  , \wishbone_bd_ram_mem3_reg[116][28]/P0001  , \wishbone_bd_ram_mem3_reg[116][29]/P0001  , \wishbone_bd_ram_mem3_reg[116][30]/P0001  , \wishbone_bd_ram_mem3_reg[116][31]/P0001  , \wishbone_bd_ram_mem3_reg[117][24]/P0001  , \wishbone_bd_ram_mem3_reg[117][25]/P0001  , \wishbone_bd_ram_mem3_reg[117][26]/P0001  , \wishbone_bd_ram_mem3_reg[117][27]/P0001  , \wishbone_bd_ram_mem3_reg[117][28]/P0001  , \wishbone_bd_ram_mem3_reg[117][29]/P0001  , \wishbone_bd_ram_mem3_reg[117][30]/P0001  , \wishbone_bd_ram_mem3_reg[117][31]/P0001  , \wishbone_bd_ram_mem3_reg[118][24]/P0001  , \wishbone_bd_ram_mem3_reg[118][25]/P0001  , \wishbone_bd_ram_mem3_reg[118][26]/P0001  , \wishbone_bd_ram_mem3_reg[118][27]/P0001  , \wishbone_bd_ram_mem3_reg[118][28]/P0001  , \wishbone_bd_ram_mem3_reg[118][29]/P0001  , \wishbone_bd_ram_mem3_reg[118][30]/P0001  , \wishbone_bd_ram_mem3_reg[118][31]/P0001  , \wishbone_bd_ram_mem3_reg[119][24]/P0001  , \wishbone_bd_ram_mem3_reg[119][25]/P0001  , \wishbone_bd_ram_mem3_reg[119][26]/P0001  , \wishbone_bd_ram_mem3_reg[119][27]/P0001  , \wishbone_bd_ram_mem3_reg[119][28]/P0001  , \wishbone_bd_ram_mem3_reg[119][29]/P0001  , \wishbone_bd_ram_mem3_reg[119][30]/P0001  , \wishbone_bd_ram_mem3_reg[119][31]/P0001  , \wishbone_bd_ram_mem3_reg[11][24]/P0001  , \wishbone_bd_ram_mem3_reg[11][25]/P0001  , \wishbone_bd_ram_mem3_reg[11][26]/P0001  , \wishbone_bd_ram_mem3_reg[11][27]/P0001  , \wishbone_bd_ram_mem3_reg[11][28]/P0001  , \wishbone_bd_ram_mem3_reg[11][29]/P0001  , \wishbone_bd_ram_mem3_reg[11][30]/P0001  , \wishbone_bd_ram_mem3_reg[11][31]/P0001  , \wishbone_bd_ram_mem3_reg[120][24]/P0001  , \wishbone_bd_ram_mem3_reg[120][25]/P0001  , \wishbone_bd_ram_mem3_reg[120][26]/P0001  , \wishbone_bd_ram_mem3_reg[120][27]/P0001  , \wishbone_bd_ram_mem3_reg[120][28]/P0001  , \wishbone_bd_ram_mem3_reg[120][29]/P0001  , \wishbone_bd_ram_mem3_reg[120][30]/P0001  , \wishbone_bd_ram_mem3_reg[120][31]/P0001  , \wishbone_bd_ram_mem3_reg[121][24]/P0001  , \wishbone_bd_ram_mem3_reg[121][25]/P0001  , \wishbone_bd_ram_mem3_reg[121][26]/P0001  , \wishbone_bd_ram_mem3_reg[121][27]/P0001  , \wishbone_bd_ram_mem3_reg[121][28]/P0001  , \wishbone_bd_ram_mem3_reg[121][29]/P0001  , \wishbone_bd_ram_mem3_reg[121][30]/P0001  , \wishbone_bd_ram_mem3_reg[121][31]/P0001  , \wishbone_bd_ram_mem3_reg[122][24]/P0001  , \wishbone_bd_ram_mem3_reg[122][25]/P0001  , \wishbone_bd_ram_mem3_reg[122][26]/P0001  , \wishbone_bd_ram_mem3_reg[122][27]/P0001  , \wishbone_bd_ram_mem3_reg[122][28]/P0001  , \wishbone_bd_ram_mem3_reg[122][29]/P0001  , \wishbone_bd_ram_mem3_reg[122][30]/P0001  , \wishbone_bd_ram_mem3_reg[122][31]/P0001  , \wishbone_bd_ram_mem3_reg[123][24]/P0001  , \wishbone_bd_ram_mem3_reg[123][25]/P0001  , \wishbone_bd_ram_mem3_reg[123][26]/P0001  , \wishbone_bd_ram_mem3_reg[123][27]/P0001  , \wishbone_bd_ram_mem3_reg[123][28]/P0001  , \wishbone_bd_ram_mem3_reg[123][29]/P0001  , \wishbone_bd_ram_mem3_reg[123][30]/P0001  , \wishbone_bd_ram_mem3_reg[123][31]/P0001  , \wishbone_bd_ram_mem3_reg[124][24]/P0001  , \wishbone_bd_ram_mem3_reg[124][25]/P0001  , \wishbone_bd_ram_mem3_reg[124][26]/P0001  , \wishbone_bd_ram_mem3_reg[124][27]/P0001  , \wishbone_bd_ram_mem3_reg[124][28]/P0001  , \wishbone_bd_ram_mem3_reg[124][29]/P0001  , \wishbone_bd_ram_mem3_reg[124][30]/P0001  , \wishbone_bd_ram_mem3_reg[124][31]/P0001  , \wishbone_bd_ram_mem3_reg[125][24]/P0001  , \wishbone_bd_ram_mem3_reg[125][25]/P0001  , \wishbone_bd_ram_mem3_reg[125][26]/P0001  , \wishbone_bd_ram_mem3_reg[125][27]/P0001  , \wishbone_bd_ram_mem3_reg[125][28]/P0001  , \wishbone_bd_ram_mem3_reg[125][29]/P0001  , \wishbone_bd_ram_mem3_reg[125][30]/P0001  , \wishbone_bd_ram_mem3_reg[125][31]/P0001  , \wishbone_bd_ram_mem3_reg[126][24]/P0001  , \wishbone_bd_ram_mem3_reg[126][25]/P0001  , \wishbone_bd_ram_mem3_reg[126][26]/P0001  , \wishbone_bd_ram_mem3_reg[126][27]/P0001  , \wishbone_bd_ram_mem3_reg[126][28]/P0001  , \wishbone_bd_ram_mem3_reg[126][29]/P0001  , \wishbone_bd_ram_mem3_reg[126][30]/P0001  , \wishbone_bd_ram_mem3_reg[126][31]/P0001  , \wishbone_bd_ram_mem3_reg[127][24]/P0001  , \wishbone_bd_ram_mem3_reg[127][25]/P0001  , \wishbone_bd_ram_mem3_reg[127][26]/P0001  , \wishbone_bd_ram_mem3_reg[127][27]/P0001  , \wishbone_bd_ram_mem3_reg[127][28]/P0001  , \wishbone_bd_ram_mem3_reg[127][29]/P0001  , \wishbone_bd_ram_mem3_reg[127][30]/P0001  , \wishbone_bd_ram_mem3_reg[127][31]/P0001  , \wishbone_bd_ram_mem3_reg[128][24]/P0001  , \wishbone_bd_ram_mem3_reg[128][25]/P0001  , \wishbone_bd_ram_mem3_reg[128][26]/P0001  , \wishbone_bd_ram_mem3_reg[128][27]/P0001  , \wishbone_bd_ram_mem3_reg[128][28]/P0001  , \wishbone_bd_ram_mem3_reg[128][29]/P0001  , \wishbone_bd_ram_mem3_reg[128][30]/P0001  , \wishbone_bd_ram_mem3_reg[128][31]/P0001  , \wishbone_bd_ram_mem3_reg[129][24]/P0001  , \wishbone_bd_ram_mem3_reg[129][25]/P0001  , \wishbone_bd_ram_mem3_reg[129][26]/P0001  , \wishbone_bd_ram_mem3_reg[129][27]/P0001  , \wishbone_bd_ram_mem3_reg[129][28]/P0001  , \wishbone_bd_ram_mem3_reg[129][29]/P0001  , \wishbone_bd_ram_mem3_reg[129][30]/P0001  , \wishbone_bd_ram_mem3_reg[129][31]/P0001  , \wishbone_bd_ram_mem3_reg[12][24]/P0001  , \wishbone_bd_ram_mem3_reg[12][25]/P0001  , \wishbone_bd_ram_mem3_reg[12][26]/P0001  , \wishbone_bd_ram_mem3_reg[12][27]/P0001  , \wishbone_bd_ram_mem3_reg[12][28]/P0001  , \wishbone_bd_ram_mem3_reg[12][29]/P0001  , \wishbone_bd_ram_mem3_reg[12][30]/P0001  , \wishbone_bd_ram_mem3_reg[12][31]/P0001  , \wishbone_bd_ram_mem3_reg[130][24]/P0001  , \wishbone_bd_ram_mem3_reg[130][25]/P0001  , \wishbone_bd_ram_mem3_reg[130][26]/P0001  , \wishbone_bd_ram_mem3_reg[130][27]/P0001  , \wishbone_bd_ram_mem3_reg[130][28]/P0001  , \wishbone_bd_ram_mem3_reg[130][29]/P0001  , \wishbone_bd_ram_mem3_reg[130][30]/P0001  , \wishbone_bd_ram_mem3_reg[130][31]/P0001  , \wishbone_bd_ram_mem3_reg[131][24]/P0001  , \wishbone_bd_ram_mem3_reg[131][25]/P0001  , \wishbone_bd_ram_mem3_reg[131][26]/P0001  , \wishbone_bd_ram_mem3_reg[131][27]/P0001  , \wishbone_bd_ram_mem3_reg[131][28]/P0001  , \wishbone_bd_ram_mem3_reg[131][29]/P0001  , \wishbone_bd_ram_mem3_reg[131][30]/P0001  , \wishbone_bd_ram_mem3_reg[131][31]/P0001  , \wishbone_bd_ram_mem3_reg[132][24]/P0001  , \wishbone_bd_ram_mem3_reg[132][25]/P0001  , \wishbone_bd_ram_mem3_reg[132][26]/P0001  , \wishbone_bd_ram_mem3_reg[132][27]/P0001  , \wishbone_bd_ram_mem3_reg[132][28]/P0001  , \wishbone_bd_ram_mem3_reg[132][29]/P0001  , \wishbone_bd_ram_mem3_reg[132][30]/P0001  , \wishbone_bd_ram_mem3_reg[132][31]/P0001  , \wishbone_bd_ram_mem3_reg[133][24]/P0001  , \wishbone_bd_ram_mem3_reg[133][25]/P0001  , \wishbone_bd_ram_mem3_reg[133][26]/P0001  , \wishbone_bd_ram_mem3_reg[133][27]/P0001  , \wishbone_bd_ram_mem3_reg[133][28]/P0001  , \wishbone_bd_ram_mem3_reg[133][29]/P0001  , \wishbone_bd_ram_mem3_reg[133][30]/P0001  , \wishbone_bd_ram_mem3_reg[133][31]/P0001  , \wishbone_bd_ram_mem3_reg[134][24]/P0001  , \wishbone_bd_ram_mem3_reg[134][25]/P0001  , \wishbone_bd_ram_mem3_reg[134][26]/P0001  , \wishbone_bd_ram_mem3_reg[134][27]/P0001  , \wishbone_bd_ram_mem3_reg[134][28]/P0001  , \wishbone_bd_ram_mem3_reg[134][29]/P0001  , \wishbone_bd_ram_mem3_reg[134][30]/P0001  , \wishbone_bd_ram_mem3_reg[134][31]/P0001  , \wishbone_bd_ram_mem3_reg[135][24]/P0001  , \wishbone_bd_ram_mem3_reg[135][25]/P0001  , \wishbone_bd_ram_mem3_reg[135][26]/P0001  , \wishbone_bd_ram_mem3_reg[135][27]/P0001  , \wishbone_bd_ram_mem3_reg[135][28]/P0001  , \wishbone_bd_ram_mem3_reg[135][29]/P0001  , \wishbone_bd_ram_mem3_reg[135][30]/P0001  , \wishbone_bd_ram_mem3_reg[135][31]/P0001  , \wishbone_bd_ram_mem3_reg[136][24]/P0001  , \wishbone_bd_ram_mem3_reg[136][25]/P0001  , \wishbone_bd_ram_mem3_reg[136][26]/P0001  , \wishbone_bd_ram_mem3_reg[136][27]/P0001  , \wishbone_bd_ram_mem3_reg[136][28]/P0001  , \wishbone_bd_ram_mem3_reg[136][29]/P0001  , \wishbone_bd_ram_mem3_reg[136][30]/P0001  , \wishbone_bd_ram_mem3_reg[136][31]/P0001  , \wishbone_bd_ram_mem3_reg[137][24]/P0001  , \wishbone_bd_ram_mem3_reg[137][25]/P0001  , \wishbone_bd_ram_mem3_reg[137][26]/P0001  , \wishbone_bd_ram_mem3_reg[137][27]/P0001  , \wishbone_bd_ram_mem3_reg[137][28]/P0001  , \wishbone_bd_ram_mem3_reg[137][29]/P0001  , \wishbone_bd_ram_mem3_reg[137][30]/P0001  , \wishbone_bd_ram_mem3_reg[137][31]/P0001  , \wishbone_bd_ram_mem3_reg[138][24]/P0001  , \wishbone_bd_ram_mem3_reg[138][25]/P0001  , \wishbone_bd_ram_mem3_reg[138][26]/P0001  , \wishbone_bd_ram_mem3_reg[138][27]/P0001  , \wishbone_bd_ram_mem3_reg[138][28]/P0001  , \wishbone_bd_ram_mem3_reg[138][29]/P0001  , \wishbone_bd_ram_mem3_reg[138][30]/P0001  , \wishbone_bd_ram_mem3_reg[138][31]/P0001  , \wishbone_bd_ram_mem3_reg[139][24]/P0001  , \wishbone_bd_ram_mem3_reg[139][25]/P0001  , \wishbone_bd_ram_mem3_reg[139][26]/P0001  , \wishbone_bd_ram_mem3_reg[139][27]/P0001  , \wishbone_bd_ram_mem3_reg[139][28]/P0001  , \wishbone_bd_ram_mem3_reg[139][29]/P0001  , \wishbone_bd_ram_mem3_reg[139][30]/P0001  , \wishbone_bd_ram_mem3_reg[139][31]/P0001  , \wishbone_bd_ram_mem3_reg[13][24]/P0001  , \wishbone_bd_ram_mem3_reg[13][25]/P0001  , \wishbone_bd_ram_mem3_reg[13][26]/P0001  , \wishbone_bd_ram_mem3_reg[13][27]/P0001  , \wishbone_bd_ram_mem3_reg[13][28]/P0001  , \wishbone_bd_ram_mem3_reg[13][29]/P0001  , \wishbone_bd_ram_mem3_reg[13][30]/P0001  , \wishbone_bd_ram_mem3_reg[13][31]/P0001  , \wishbone_bd_ram_mem3_reg[140][24]/P0001  , \wishbone_bd_ram_mem3_reg[140][25]/P0001  , \wishbone_bd_ram_mem3_reg[140][26]/P0001  , \wishbone_bd_ram_mem3_reg[140][27]/P0001  , \wishbone_bd_ram_mem3_reg[140][28]/P0001  , \wishbone_bd_ram_mem3_reg[140][29]/P0001  , \wishbone_bd_ram_mem3_reg[140][30]/P0001  , \wishbone_bd_ram_mem3_reg[140][31]/P0001  , \wishbone_bd_ram_mem3_reg[141][24]/P0001  , \wishbone_bd_ram_mem3_reg[141][25]/P0001  , \wishbone_bd_ram_mem3_reg[141][26]/P0001  , \wishbone_bd_ram_mem3_reg[141][27]/P0001  , \wishbone_bd_ram_mem3_reg[141][28]/P0001  , \wishbone_bd_ram_mem3_reg[141][29]/P0001  , \wishbone_bd_ram_mem3_reg[141][30]/P0001  , \wishbone_bd_ram_mem3_reg[141][31]/P0001  , \wishbone_bd_ram_mem3_reg[142][24]/P0001  , \wishbone_bd_ram_mem3_reg[142][25]/P0001  , \wishbone_bd_ram_mem3_reg[142][26]/P0001  , \wishbone_bd_ram_mem3_reg[142][27]/P0001  , \wishbone_bd_ram_mem3_reg[142][28]/P0001  , \wishbone_bd_ram_mem3_reg[142][29]/P0001  , \wishbone_bd_ram_mem3_reg[142][30]/P0001  , \wishbone_bd_ram_mem3_reg[142][31]/P0001  , \wishbone_bd_ram_mem3_reg[143][24]/P0001  , \wishbone_bd_ram_mem3_reg[143][25]/P0001  , \wishbone_bd_ram_mem3_reg[143][26]/P0001  , \wishbone_bd_ram_mem3_reg[143][27]/P0001  , \wishbone_bd_ram_mem3_reg[143][28]/P0001  , \wishbone_bd_ram_mem3_reg[143][29]/P0001  , \wishbone_bd_ram_mem3_reg[143][30]/P0001  , \wishbone_bd_ram_mem3_reg[143][31]/P0001  , \wishbone_bd_ram_mem3_reg[144][24]/P0001  , \wishbone_bd_ram_mem3_reg[144][25]/P0001  , \wishbone_bd_ram_mem3_reg[144][26]/P0001  , \wishbone_bd_ram_mem3_reg[144][27]/P0001  , \wishbone_bd_ram_mem3_reg[144][28]/P0001  , \wishbone_bd_ram_mem3_reg[144][29]/P0001  , \wishbone_bd_ram_mem3_reg[144][30]/P0001  , \wishbone_bd_ram_mem3_reg[144][31]/P0001  , \wishbone_bd_ram_mem3_reg[145][24]/P0001  , \wishbone_bd_ram_mem3_reg[145][25]/P0001  , \wishbone_bd_ram_mem3_reg[145][26]/P0001  , \wishbone_bd_ram_mem3_reg[145][27]/P0001  , \wishbone_bd_ram_mem3_reg[145][28]/P0001  , \wishbone_bd_ram_mem3_reg[145][29]/P0001  , \wishbone_bd_ram_mem3_reg[145][30]/P0001  , \wishbone_bd_ram_mem3_reg[145][31]/P0001  , \wishbone_bd_ram_mem3_reg[146][24]/P0001  , \wishbone_bd_ram_mem3_reg[146][25]/P0001  , \wishbone_bd_ram_mem3_reg[146][26]/P0001  , \wishbone_bd_ram_mem3_reg[146][27]/P0001  , \wishbone_bd_ram_mem3_reg[146][28]/P0001  , \wishbone_bd_ram_mem3_reg[146][29]/P0001  , \wishbone_bd_ram_mem3_reg[146][30]/P0001  , \wishbone_bd_ram_mem3_reg[146][31]/P0001  , \wishbone_bd_ram_mem3_reg[147][24]/P0001  , \wishbone_bd_ram_mem3_reg[147][25]/P0001  , \wishbone_bd_ram_mem3_reg[147][26]/P0001  , \wishbone_bd_ram_mem3_reg[147][27]/P0001  , \wishbone_bd_ram_mem3_reg[147][28]/P0001  , \wishbone_bd_ram_mem3_reg[147][29]/P0001  , \wishbone_bd_ram_mem3_reg[147][30]/P0001  , \wishbone_bd_ram_mem3_reg[147][31]/P0001  , \wishbone_bd_ram_mem3_reg[148][24]/P0001  , \wishbone_bd_ram_mem3_reg[148][25]/P0001  , \wishbone_bd_ram_mem3_reg[148][26]/P0001  , \wishbone_bd_ram_mem3_reg[148][27]/P0001  , \wishbone_bd_ram_mem3_reg[148][28]/P0001  , \wishbone_bd_ram_mem3_reg[148][29]/P0001  , \wishbone_bd_ram_mem3_reg[148][30]/P0001  , \wishbone_bd_ram_mem3_reg[148][31]/P0001  , \wishbone_bd_ram_mem3_reg[149][24]/P0001  , \wishbone_bd_ram_mem3_reg[149][25]/P0001  , \wishbone_bd_ram_mem3_reg[149][26]/P0001  , \wishbone_bd_ram_mem3_reg[149][27]/P0001  , \wishbone_bd_ram_mem3_reg[149][28]/P0001  , \wishbone_bd_ram_mem3_reg[149][29]/P0001  , \wishbone_bd_ram_mem3_reg[149][30]/P0001  , \wishbone_bd_ram_mem3_reg[149][31]/P0001  , \wishbone_bd_ram_mem3_reg[14][24]/P0001  , \wishbone_bd_ram_mem3_reg[14][25]/P0001  , \wishbone_bd_ram_mem3_reg[14][26]/P0001  , \wishbone_bd_ram_mem3_reg[14][27]/P0001  , \wishbone_bd_ram_mem3_reg[14][28]/P0001  , \wishbone_bd_ram_mem3_reg[14][29]/P0001  , \wishbone_bd_ram_mem3_reg[14][30]/P0001  , \wishbone_bd_ram_mem3_reg[14][31]/P0001  , \wishbone_bd_ram_mem3_reg[150][24]/P0001  , \wishbone_bd_ram_mem3_reg[150][25]/P0001  , \wishbone_bd_ram_mem3_reg[150][26]/P0001  , \wishbone_bd_ram_mem3_reg[150][27]/P0001  , \wishbone_bd_ram_mem3_reg[150][28]/P0001  , \wishbone_bd_ram_mem3_reg[150][29]/P0001  , \wishbone_bd_ram_mem3_reg[150][30]/P0001  , \wishbone_bd_ram_mem3_reg[150][31]/P0001  , \wishbone_bd_ram_mem3_reg[151][24]/P0001  , \wishbone_bd_ram_mem3_reg[151][25]/P0001  , \wishbone_bd_ram_mem3_reg[151][26]/P0001  , \wishbone_bd_ram_mem3_reg[151][27]/P0001  , \wishbone_bd_ram_mem3_reg[151][28]/P0001  , \wishbone_bd_ram_mem3_reg[151][29]/P0001  , \wishbone_bd_ram_mem3_reg[151][30]/P0001  , \wishbone_bd_ram_mem3_reg[151][31]/P0001  , \wishbone_bd_ram_mem3_reg[152][24]/P0001  , \wishbone_bd_ram_mem3_reg[152][25]/P0001  , \wishbone_bd_ram_mem3_reg[152][26]/P0001  , \wishbone_bd_ram_mem3_reg[152][27]/P0001  , \wishbone_bd_ram_mem3_reg[152][28]/P0001  , \wishbone_bd_ram_mem3_reg[152][29]/P0001  , \wishbone_bd_ram_mem3_reg[152][30]/P0001  , \wishbone_bd_ram_mem3_reg[152][31]/P0001  , \wishbone_bd_ram_mem3_reg[153][24]/P0001  , \wishbone_bd_ram_mem3_reg[153][25]/P0001  , \wishbone_bd_ram_mem3_reg[153][26]/P0001  , \wishbone_bd_ram_mem3_reg[153][27]/P0001  , \wishbone_bd_ram_mem3_reg[153][28]/P0001  , \wishbone_bd_ram_mem3_reg[153][29]/P0001  , \wishbone_bd_ram_mem3_reg[153][30]/P0001  , \wishbone_bd_ram_mem3_reg[153][31]/P0001  , \wishbone_bd_ram_mem3_reg[154][24]/P0001  , \wishbone_bd_ram_mem3_reg[154][25]/P0001  , \wishbone_bd_ram_mem3_reg[154][26]/P0001  , \wishbone_bd_ram_mem3_reg[154][27]/P0001  , \wishbone_bd_ram_mem3_reg[154][28]/P0001  , \wishbone_bd_ram_mem3_reg[154][29]/P0001  , \wishbone_bd_ram_mem3_reg[154][30]/P0001  , \wishbone_bd_ram_mem3_reg[154][31]/P0001  , \wishbone_bd_ram_mem3_reg[155][24]/P0001  , \wishbone_bd_ram_mem3_reg[155][25]/P0001  , \wishbone_bd_ram_mem3_reg[155][26]/P0001  , \wishbone_bd_ram_mem3_reg[155][27]/P0001  , \wishbone_bd_ram_mem3_reg[155][28]/P0001  , \wishbone_bd_ram_mem3_reg[155][29]/P0001  , \wishbone_bd_ram_mem3_reg[155][30]/P0001  , \wishbone_bd_ram_mem3_reg[155][31]/P0001  , \wishbone_bd_ram_mem3_reg[156][24]/P0001  , \wishbone_bd_ram_mem3_reg[156][25]/P0001  , \wishbone_bd_ram_mem3_reg[156][26]/P0001  , \wishbone_bd_ram_mem3_reg[156][27]/P0001  , \wishbone_bd_ram_mem3_reg[156][28]/P0001  , \wishbone_bd_ram_mem3_reg[156][29]/P0001  , \wishbone_bd_ram_mem3_reg[156][30]/P0001  , \wishbone_bd_ram_mem3_reg[156][31]/P0001  , \wishbone_bd_ram_mem3_reg[157][24]/P0001  , \wishbone_bd_ram_mem3_reg[157][25]/P0001  , \wishbone_bd_ram_mem3_reg[157][26]/P0001  , \wishbone_bd_ram_mem3_reg[157][27]/P0001  , \wishbone_bd_ram_mem3_reg[157][28]/P0001  , \wishbone_bd_ram_mem3_reg[157][29]/P0001  , \wishbone_bd_ram_mem3_reg[157][30]/P0001  , \wishbone_bd_ram_mem3_reg[157][31]/P0001  , \wishbone_bd_ram_mem3_reg[158][24]/P0001  , \wishbone_bd_ram_mem3_reg[158][25]/P0001  , \wishbone_bd_ram_mem3_reg[158][26]/P0001  , \wishbone_bd_ram_mem3_reg[158][27]/P0001  , \wishbone_bd_ram_mem3_reg[158][28]/P0001  , \wishbone_bd_ram_mem3_reg[158][29]/P0001  , \wishbone_bd_ram_mem3_reg[158][30]/P0001  , \wishbone_bd_ram_mem3_reg[158][31]/P0001  , \wishbone_bd_ram_mem3_reg[159][24]/P0001  , \wishbone_bd_ram_mem3_reg[159][25]/P0001  , \wishbone_bd_ram_mem3_reg[159][26]/P0001  , \wishbone_bd_ram_mem3_reg[159][27]/P0001  , \wishbone_bd_ram_mem3_reg[159][28]/P0001  , \wishbone_bd_ram_mem3_reg[159][29]/P0001  , \wishbone_bd_ram_mem3_reg[159][30]/P0001  , \wishbone_bd_ram_mem3_reg[159][31]/P0001  , \wishbone_bd_ram_mem3_reg[15][24]/P0001  , \wishbone_bd_ram_mem3_reg[15][25]/P0001  , \wishbone_bd_ram_mem3_reg[15][26]/P0001  , \wishbone_bd_ram_mem3_reg[15][27]/P0001  , \wishbone_bd_ram_mem3_reg[15][28]/P0001  , \wishbone_bd_ram_mem3_reg[15][29]/P0001  , \wishbone_bd_ram_mem3_reg[15][30]/P0001  , \wishbone_bd_ram_mem3_reg[15][31]/P0001  , \wishbone_bd_ram_mem3_reg[160][24]/P0001  , \wishbone_bd_ram_mem3_reg[160][25]/P0001  , \wishbone_bd_ram_mem3_reg[160][26]/P0001  , \wishbone_bd_ram_mem3_reg[160][27]/P0001  , \wishbone_bd_ram_mem3_reg[160][28]/P0001  , \wishbone_bd_ram_mem3_reg[160][29]/P0001  , \wishbone_bd_ram_mem3_reg[160][30]/P0001  , \wishbone_bd_ram_mem3_reg[160][31]/P0001  , \wishbone_bd_ram_mem3_reg[161][24]/P0001  , \wishbone_bd_ram_mem3_reg[161][25]/P0001  , \wishbone_bd_ram_mem3_reg[161][26]/P0001  , \wishbone_bd_ram_mem3_reg[161][27]/P0001  , \wishbone_bd_ram_mem3_reg[161][28]/P0001  , \wishbone_bd_ram_mem3_reg[161][29]/P0001  , \wishbone_bd_ram_mem3_reg[161][30]/P0001  , \wishbone_bd_ram_mem3_reg[161][31]/P0001  , \wishbone_bd_ram_mem3_reg[162][24]/P0001  , \wishbone_bd_ram_mem3_reg[162][25]/P0001  , \wishbone_bd_ram_mem3_reg[162][26]/P0001  , \wishbone_bd_ram_mem3_reg[162][27]/P0001  , \wishbone_bd_ram_mem3_reg[162][28]/P0001  , \wishbone_bd_ram_mem3_reg[162][29]/P0001  , \wishbone_bd_ram_mem3_reg[162][30]/P0001  , \wishbone_bd_ram_mem3_reg[162][31]/P0001  , \wishbone_bd_ram_mem3_reg[163][24]/P0001  , \wishbone_bd_ram_mem3_reg[163][25]/P0001  , \wishbone_bd_ram_mem3_reg[163][26]/P0001  , \wishbone_bd_ram_mem3_reg[163][27]/P0001  , \wishbone_bd_ram_mem3_reg[163][28]/P0001  , \wishbone_bd_ram_mem3_reg[163][29]/P0001  , \wishbone_bd_ram_mem3_reg[163][30]/P0001  , \wishbone_bd_ram_mem3_reg[163][31]/P0001  , \wishbone_bd_ram_mem3_reg[164][24]/P0001  , \wishbone_bd_ram_mem3_reg[164][25]/P0001  , \wishbone_bd_ram_mem3_reg[164][26]/P0001  , \wishbone_bd_ram_mem3_reg[164][27]/P0001  , \wishbone_bd_ram_mem3_reg[164][28]/P0001  , \wishbone_bd_ram_mem3_reg[164][29]/P0001  , \wishbone_bd_ram_mem3_reg[164][30]/P0001  , \wishbone_bd_ram_mem3_reg[164][31]/P0001  , \wishbone_bd_ram_mem3_reg[165][24]/P0001  , \wishbone_bd_ram_mem3_reg[165][25]/P0001  , \wishbone_bd_ram_mem3_reg[165][26]/P0001  , \wishbone_bd_ram_mem3_reg[165][27]/P0001  , \wishbone_bd_ram_mem3_reg[165][28]/P0001  , \wishbone_bd_ram_mem3_reg[165][29]/P0001  , \wishbone_bd_ram_mem3_reg[165][30]/P0001  , \wishbone_bd_ram_mem3_reg[165][31]/P0001  , \wishbone_bd_ram_mem3_reg[166][24]/P0001  , \wishbone_bd_ram_mem3_reg[166][25]/P0001  , \wishbone_bd_ram_mem3_reg[166][26]/P0001  , \wishbone_bd_ram_mem3_reg[166][27]/P0001  , \wishbone_bd_ram_mem3_reg[166][28]/P0001  , \wishbone_bd_ram_mem3_reg[166][29]/P0001  , \wishbone_bd_ram_mem3_reg[166][30]/P0001  , \wishbone_bd_ram_mem3_reg[166][31]/P0001  , \wishbone_bd_ram_mem3_reg[167][24]/P0001  , \wishbone_bd_ram_mem3_reg[167][25]/P0001  , \wishbone_bd_ram_mem3_reg[167][26]/P0001  , \wishbone_bd_ram_mem3_reg[167][27]/P0001  , \wishbone_bd_ram_mem3_reg[167][28]/P0001  , \wishbone_bd_ram_mem3_reg[167][29]/P0001  , \wishbone_bd_ram_mem3_reg[167][30]/P0001  , \wishbone_bd_ram_mem3_reg[167][31]/P0001  , \wishbone_bd_ram_mem3_reg[168][24]/P0001  , \wishbone_bd_ram_mem3_reg[168][25]/P0001  , \wishbone_bd_ram_mem3_reg[168][26]/P0001  , \wishbone_bd_ram_mem3_reg[168][27]/P0001  , \wishbone_bd_ram_mem3_reg[168][28]/P0001  , \wishbone_bd_ram_mem3_reg[168][29]/P0001  , \wishbone_bd_ram_mem3_reg[168][30]/P0001  , \wishbone_bd_ram_mem3_reg[168][31]/P0001  , \wishbone_bd_ram_mem3_reg[169][24]/P0001  , \wishbone_bd_ram_mem3_reg[169][25]/P0001  , \wishbone_bd_ram_mem3_reg[169][26]/P0001  , \wishbone_bd_ram_mem3_reg[169][27]/P0001  , \wishbone_bd_ram_mem3_reg[169][28]/P0001  , \wishbone_bd_ram_mem3_reg[169][29]/P0001  , \wishbone_bd_ram_mem3_reg[169][30]/P0001  , \wishbone_bd_ram_mem3_reg[169][31]/P0001  , \wishbone_bd_ram_mem3_reg[16][24]/P0001  , \wishbone_bd_ram_mem3_reg[16][25]/P0001  , \wishbone_bd_ram_mem3_reg[16][26]/P0001  , \wishbone_bd_ram_mem3_reg[16][27]/P0001  , \wishbone_bd_ram_mem3_reg[16][28]/P0001  , \wishbone_bd_ram_mem3_reg[16][29]/P0001  , \wishbone_bd_ram_mem3_reg[16][30]/P0001  , \wishbone_bd_ram_mem3_reg[16][31]/P0001  , \wishbone_bd_ram_mem3_reg[170][24]/P0001  , \wishbone_bd_ram_mem3_reg[170][25]/P0001  , \wishbone_bd_ram_mem3_reg[170][26]/P0001  , \wishbone_bd_ram_mem3_reg[170][27]/P0001  , \wishbone_bd_ram_mem3_reg[170][28]/P0001  , \wishbone_bd_ram_mem3_reg[170][29]/P0001  , \wishbone_bd_ram_mem3_reg[170][30]/P0001  , \wishbone_bd_ram_mem3_reg[170][31]/P0001  , \wishbone_bd_ram_mem3_reg[171][24]/P0001  , \wishbone_bd_ram_mem3_reg[171][25]/P0001  , \wishbone_bd_ram_mem3_reg[171][26]/P0001  , \wishbone_bd_ram_mem3_reg[171][27]/P0001  , \wishbone_bd_ram_mem3_reg[171][28]/P0001  , \wishbone_bd_ram_mem3_reg[171][29]/P0001  , \wishbone_bd_ram_mem3_reg[171][30]/P0001  , \wishbone_bd_ram_mem3_reg[171][31]/P0001  , \wishbone_bd_ram_mem3_reg[172][24]/P0001  , \wishbone_bd_ram_mem3_reg[172][25]/P0001  , \wishbone_bd_ram_mem3_reg[172][26]/P0001  , \wishbone_bd_ram_mem3_reg[172][27]/P0001  , \wishbone_bd_ram_mem3_reg[172][28]/P0001  , \wishbone_bd_ram_mem3_reg[172][29]/P0001  , \wishbone_bd_ram_mem3_reg[172][30]/P0001  , \wishbone_bd_ram_mem3_reg[172][31]/P0001  , \wishbone_bd_ram_mem3_reg[173][24]/P0001  , \wishbone_bd_ram_mem3_reg[173][25]/P0001  , \wishbone_bd_ram_mem3_reg[173][26]/P0001  , \wishbone_bd_ram_mem3_reg[173][27]/P0001  , \wishbone_bd_ram_mem3_reg[173][28]/P0001  , \wishbone_bd_ram_mem3_reg[173][29]/P0001  , \wishbone_bd_ram_mem3_reg[173][30]/P0001  , \wishbone_bd_ram_mem3_reg[173][31]/P0001  , \wishbone_bd_ram_mem3_reg[174][24]/P0001  , \wishbone_bd_ram_mem3_reg[174][25]/P0001  , \wishbone_bd_ram_mem3_reg[174][26]/P0001  , \wishbone_bd_ram_mem3_reg[174][27]/P0001  , \wishbone_bd_ram_mem3_reg[174][28]/P0001  , \wishbone_bd_ram_mem3_reg[174][29]/P0001  , \wishbone_bd_ram_mem3_reg[174][30]/P0001  , \wishbone_bd_ram_mem3_reg[174][31]/P0001  , \wishbone_bd_ram_mem3_reg[175][24]/P0001  , \wishbone_bd_ram_mem3_reg[175][25]/P0001  , \wishbone_bd_ram_mem3_reg[175][26]/P0001  , \wishbone_bd_ram_mem3_reg[175][27]/P0001  , \wishbone_bd_ram_mem3_reg[175][28]/P0001  , \wishbone_bd_ram_mem3_reg[175][29]/P0001  , \wishbone_bd_ram_mem3_reg[175][30]/P0001  , \wishbone_bd_ram_mem3_reg[175][31]/P0001  , \wishbone_bd_ram_mem3_reg[176][24]/P0001  , \wishbone_bd_ram_mem3_reg[176][25]/P0001  , \wishbone_bd_ram_mem3_reg[176][26]/P0001  , \wishbone_bd_ram_mem3_reg[176][27]/P0001  , \wishbone_bd_ram_mem3_reg[176][28]/P0001  , \wishbone_bd_ram_mem3_reg[176][29]/P0001  , \wishbone_bd_ram_mem3_reg[176][30]/P0001  , \wishbone_bd_ram_mem3_reg[176][31]/P0001  , \wishbone_bd_ram_mem3_reg[177][24]/P0001  , \wishbone_bd_ram_mem3_reg[177][25]/P0001  , \wishbone_bd_ram_mem3_reg[177][26]/P0001  , \wishbone_bd_ram_mem3_reg[177][27]/P0001  , \wishbone_bd_ram_mem3_reg[177][28]/P0001  , \wishbone_bd_ram_mem3_reg[177][29]/P0001  , \wishbone_bd_ram_mem3_reg[177][30]/P0001  , \wishbone_bd_ram_mem3_reg[177][31]/P0001  , \wishbone_bd_ram_mem3_reg[178][24]/P0001  , \wishbone_bd_ram_mem3_reg[178][25]/P0001  , \wishbone_bd_ram_mem3_reg[178][26]/P0001  , \wishbone_bd_ram_mem3_reg[178][27]/P0001  , \wishbone_bd_ram_mem3_reg[178][28]/P0001  , \wishbone_bd_ram_mem3_reg[178][29]/P0001  , \wishbone_bd_ram_mem3_reg[178][30]/P0001  , \wishbone_bd_ram_mem3_reg[178][31]/P0001  , \wishbone_bd_ram_mem3_reg[179][24]/P0001  , \wishbone_bd_ram_mem3_reg[179][25]/P0001  , \wishbone_bd_ram_mem3_reg[179][26]/P0001  , \wishbone_bd_ram_mem3_reg[179][27]/P0001  , \wishbone_bd_ram_mem3_reg[179][28]/P0001  , \wishbone_bd_ram_mem3_reg[179][29]/P0001  , \wishbone_bd_ram_mem3_reg[179][30]/P0001  , \wishbone_bd_ram_mem3_reg[179][31]/P0001  , \wishbone_bd_ram_mem3_reg[17][24]/P0001  , \wishbone_bd_ram_mem3_reg[17][25]/P0001  , \wishbone_bd_ram_mem3_reg[17][26]/P0001  , \wishbone_bd_ram_mem3_reg[17][27]/P0001  , \wishbone_bd_ram_mem3_reg[17][28]/P0001  , \wishbone_bd_ram_mem3_reg[17][29]/P0001  , \wishbone_bd_ram_mem3_reg[17][30]/P0001  , \wishbone_bd_ram_mem3_reg[17][31]/P0001  , \wishbone_bd_ram_mem3_reg[180][24]/P0001  , \wishbone_bd_ram_mem3_reg[180][25]/P0001  , \wishbone_bd_ram_mem3_reg[180][26]/P0001  , \wishbone_bd_ram_mem3_reg[180][27]/P0001  , \wishbone_bd_ram_mem3_reg[180][28]/P0001  , \wishbone_bd_ram_mem3_reg[180][29]/P0001  , \wishbone_bd_ram_mem3_reg[180][30]/P0001  , \wishbone_bd_ram_mem3_reg[180][31]/P0001  , \wishbone_bd_ram_mem3_reg[181][24]/P0001  , \wishbone_bd_ram_mem3_reg[181][25]/P0001  , \wishbone_bd_ram_mem3_reg[181][26]/P0001  , \wishbone_bd_ram_mem3_reg[181][27]/P0001  , \wishbone_bd_ram_mem3_reg[181][28]/P0001  , \wishbone_bd_ram_mem3_reg[181][29]/P0001  , \wishbone_bd_ram_mem3_reg[181][30]/P0001  , \wishbone_bd_ram_mem3_reg[181][31]/P0001  , \wishbone_bd_ram_mem3_reg[182][24]/P0001  , \wishbone_bd_ram_mem3_reg[182][25]/P0001  , \wishbone_bd_ram_mem3_reg[182][26]/P0001  , \wishbone_bd_ram_mem3_reg[182][27]/P0001  , \wishbone_bd_ram_mem3_reg[182][28]/P0001  , \wishbone_bd_ram_mem3_reg[182][29]/P0001  , \wishbone_bd_ram_mem3_reg[182][30]/P0001  , \wishbone_bd_ram_mem3_reg[182][31]/P0001  , \wishbone_bd_ram_mem3_reg[183][24]/P0001  , \wishbone_bd_ram_mem3_reg[183][25]/P0001  , \wishbone_bd_ram_mem3_reg[183][26]/P0001  , \wishbone_bd_ram_mem3_reg[183][27]/P0001  , \wishbone_bd_ram_mem3_reg[183][28]/P0001  , \wishbone_bd_ram_mem3_reg[183][29]/P0001  , \wishbone_bd_ram_mem3_reg[183][30]/P0001  , \wishbone_bd_ram_mem3_reg[183][31]/P0001  , \wishbone_bd_ram_mem3_reg[184][24]/P0001  , \wishbone_bd_ram_mem3_reg[184][25]/P0001  , \wishbone_bd_ram_mem3_reg[184][26]/P0001  , \wishbone_bd_ram_mem3_reg[184][27]/P0001  , \wishbone_bd_ram_mem3_reg[184][28]/P0001  , \wishbone_bd_ram_mem3_reg[184][29]/P0001  , \wishbone_bd_ram_mem3_reg[184][30]/P0001  , \wishbone_bd_ram_mem3_reg[184][31]/P0001  , \wishbone_bd_ram_mem3_reg[185][24]/P0001  , \wishbone_bd_ram_mem3_reg[185][25]/P0001  , \wishbone_bd_ram_mem3_reg[185][26]/P0001  , \wishbone_bd_ram_mem3_reg[185][27]/P0001  , \wishbone_bd_ram_mem3_reg[185][28]/P0001  , \wishbone_bd_ram_mem3_reg[185][29]/P0001  , \wishbone_bd_ram_mem3_reg[185][30]/P0001  , \wishbone_bd_ram_mem3_reg[185][31]/P0001  , \wishbone_bd_ram_mem3_reg[186][24]/P0001  , \wishbone_bd_ram_mem3_reg[186][25]/P0001  , \wishbone_bd_ram_mem3_reg[186][26]/P0001  , \wishbone_bd_ram_mem3_reg[186][27]/P0001  , \wishbone_bd_ram_mem3_reg[186][28]/P0001  , \wishbone_bd_ram_mem3_reg[186][29]/P0001  , \wishbone_bd_ram_mem3_reg[186][30]/P0001  , \wishbone_bd_ram_mem3_reg[186][31]/P0001  , \wishbone_bd_ram_mem3_reg[187][24]/P0001  , \wishbone_bd_ram_mem3_reg[187][25]/P0001  , \wishbone_bd_ram_mem3_reg[187][26]/P0001  , \wishbone_bd_ram_mem3_reg[187][27]/P0001  , \wishbone_bd_ram_mem3_reg[187][28]/P0001  , \wishbone_bd_ram_mem3_reg[187][29]/P0001  , \wishbone_bd_ram_mem3_reg[187][30]/P0001  , \wishbone_bd_ram_mem3_reg[187][31]/P0001  , \wishbone_bd_ram_mem3_reg[188][24]/P0001  , \wishbone_bd_ram_mem3_reg[188][25]/P0001  , \wishbone_bd_ram_mem3_reg[188][26]/P0001  , \wishbone_bd_ram_mem3_reg[188][27]/P0001  , \wishbone_bd_ram_mem3_reg[188][28]/P0001  , \wishbone_bd_ram_mem3_reg[188][29]/P0001  , \wishbone_bd_ram_mem3_reg[188][30]/P0001  , \wishbone_bd_ram_mem3_reg[188][31]/P0001  , \wishbone_bd_ram_mem3_reg[189][24]/P0001  , \wishbone_bd_ram_mem3_reg[189][25]/P0001  , \wishbone_bd_ram_mem3_reg[189][26]/P0001  , \wishbone_bd_ram_mem3_reg[189][27]/P0001  , \wishbone_bd_ram_mem3_reg[189][28]/P0001  , \wishbone_bd_ram_mem3_reg[189][29]/P0001  , \wishbone_bd_ram_mem3_reg[189][30]/P0001  , \wishbone_bd_ram_mem3_reg[189][31]/P0001  , \wishbone_bd_ram_mem3_reg[18][24]/P0001  , \wishbone_bd_ram_mem3_reg[18][25]/P0001  , \wishbone_bd_ram_mem3_reg[18][26]/P0001  , \wishbone_bd_ram_mem3_reg[18][27]/P0001  , \wishbone_bd_ram_mem3_reg[18][28]/P0001  , \wishbone_bd_ram_mem3_reg[18][29]/P0001  , \wishbone_bd_ram_mem3_reg[18][30]/P0001  , \wishbone_bd_ram_mem3_reg[18][31]/P0001  , \wishbone_bd_ram_mem3_reg[190][24]/P0001  , \wishbone_bd_ram_mem3_reg[190][25]/P0001  , \wishbone_bd_ram_mem3_reg[190][26]/P0001  , \wishbone_bd_ram_mem3_reg[190][27]/P0001  , \wishbone_bd_ram_mem3_reg[190][28]/P0001  , \wishbone_bd_ram_mem3_reg[190][29]/P0001  , \wishbone_bd_ram_mem3_reg[190][30]/P0001  , \wishbone_bd_ram_mem3_reg[190][31]/P0001  , \wishbone_bd_ram_mem3_reg[191][24]/P0001  , \wishbone_bd_ram_mem3_reg[191][25]/P0001  , \wishbone_bd_ram_mem3_reg[191][26]/P0001  , \wishbone_bd_ram_mem3_reg[191][27]/P0001  , \wishbone_bd_ram_mem3_reg[191][28]/P0001  , \wishbone_bd_ram_mem3_reg[191][29]/P0001  , \wishbone_bd_ram_mem3_reg[191][30]/P0001  , \wishbone_bd_ram_mem3_reg[191][31]/P0001  , \wishbone_bd_ram_mem3_reg[192][24]/P0001  , \wishbone_bd_ram_mem3_reg[192][25]/P0001  , \wishbone_bd_ram_mem3_reg[192][26]/P0001  , \wishbone_bd_ram_mem3_reg[192][27]/P0001  , \wishbone_bd_ram_mem3_reg[192][28]/P0001  , \wishbone_bd_ram_mem3_reg[192][29]/P0001  , \wishbone_bd_ram_mem3_reg[192][30]/P0001  , \wishbone_bd_ram_mem3_reg[192][31]/P0001  , \wishbone_bd_ram_mem3_reg[193][24]/P0001  , \wishbone_bd_ram_mem3_reg[193][25]/P0001  , \wishbone_bd_ram_mem3_reg[193][26]/P0001  , \wishbone_bd_ram_mem3_reg[193][27]/P0001  , \wishbone_bd_ram_mem3_reg[193][28]/P0001  , \wishbone_bd_ram_mem3_reg[193][29]/P0001  , \wishbone_bd_ram_mem3_reg[193][30]/P0001  , \wishbone_bd_ram_mem3_reg[193][31]/P0001  , \wishbone_bd_ram_mem3_reg[194][24]/P0001  , \wishbone_bd_ram_mem3_reg[194][25]/P0001  , \wishbone_bd_ram_mem3_reg[194][26]/P0001  , \wishbone_bd_ram_mem3_reg[194][27]/P0001  , \wishbone_bd_ram_mem3_reg[194][28]/P0001  , \wishbone_bd_ram_mem3_reg[194][29]/P0001  , \wishbone_bd_ram_mem3_reg[194][30]/P0001  , \wishbone_bd_ram_mem3_reg[194][31]/P0001  , \wishbone_bd_ram_mem3_reg[195][24]/P0001  , \wishbone_bd_ram_mem3_reg[195][25]/P0001  , \wishbone_bd_ram_mem3_reg[195][26]/P0001  , \wishbone_bd_ram_mem3_reg[195][27]/P0001  , \wishbone_bd_ram_mem3_reg[195][28]/P0001  , \wishbone_bd_ram_mem3_reg[195][29]/P0001  , \wishbone_bd_ram_mem3_reg[195][30]/P0001  , \wishbone_bd_ram_mem3_reg[195][31]/P0001  , \wishbone_bd_ram_mem3_reg[196][24]/P0001  , \wishbone_bd_ram_mem3_reg[196][25]/P0001  , \wishbone_bd_ram_mem3_reg[196][26]/P0001  , \wishbone_bd_ram_mem3_reg[196][27]/P0001  , \wishbone_bd_ram_mem3_reg[196][28]/P0001  , \wishbone_bd_ram_mem3_reg[196][29]/P0001  , \wishbone_bd_ram_mem3_reg[196][30]/P0001  , \wishbone_bd_ram_mem3_reg[196][31]/P0001  , \wishbone_bd_ram_mem3_reg[197][24]/P0001  , \wishbone_bd_ram_mem3_reg[197][25]/P0001  , \wishbone_bd_ram_mem3_reg[197][26]/P0001  , \wishbone_bd_ram_mem3_reg[197][27]/P0001  , \wishbone_bd_ram_mem3_reg[197][28]/P0001  , \wishbone_bd_ram_mem3_reg[197][29]/P0001  , \wishbone_bd_ram_mem3_reg[197][30]/P0001  , \wishbone_bd_ram_mem3_reg[197][31]/P0001  , \wishbone_bd_ram_mem3_reg[198][24]/P0001  , \wishbone_bd_ram_mem3_reg[198][25]/P0001  , \wishbone_bd_ram_mem3_reg[198][26]/P0001  , \wishbone_bd_ram_mem3_reg[198][27]/P0001  , \wishbone_bd_ram_mem3_reg[198][28]/P0001  , \wishbone_bd_ram_mem3_reg[198][29]/P0001  , \wishbone_bd_ram_mem3_reg[198][30]/P0001  , \wishbone_bd_ram_mem3_reg[198][31]/P0001  , \wishbone_bd_ram_mem3_reg[199][24]/P0001  , \wishbone_bd_ram_mem3_reg[199][25]/P0001  , \wishbone_bd_ram_mem3_reg[199][26]/P0001  , \wishbone_bd_ram_mem3_reg[199][27]/P0001  , \wishbone_bd_ram_mem3_reg[199][28]/P0001  , \wishbone_bd_ram_mem3_reg[199][29]/P0001  , \wishbone_bd_ram_mem3_reg[199][30]/P0001  , \wishbone_bd_ram_mem3_reg[199][31]/P0001  , \wishbone_bd_ram_mem3_reg[19][24]/P0001  , \wishbone_bd_ram_mem3_reg[19][25]/P0001  , \wishbone_bd_ram_mem3_reg[19][26]/P0001  , \wishbone_bd_ram_mem3_reg[19][27]/P0001  , \wishbone_bd_ram_mem3_reg[19][28]/P0001  , \wishbone_bd_ram_mem3_reg[19][29]/P0001  , \wishbone_bd_ram_mem3_reg[19][30]/P0001  , \wishbone_bd_ram_mem3_reg[19][31]/P0001  , \wishbone_bd_ram_mem3_reg[1][24]/P0001  , \wishbone_bd_ram_mem3_reg[1][25]/P0001  , \wishbone_bd_ram_mem3_reg[1][26]/P0001  , \wishbone_bd_ram_mem3_reg[1][27]/P0001  , \wishbone_bd_ram_mem3_reg[1][28]/P0001  , \wishbone_bd_ram_mem3_reg[1][29]/P0001  , \wishbone_bd_ram_mem3_reg[1][30]/P0001  , \wishbone_bd_ram_mem3_reg[1][31]/P0001  , \wishbone_bd_ram_mem3_reg[200][24]/P0001  , \wishbone_bd_ram_mem3_reg[200][25]/P0001  , \wishbone_bd_ram_mem3_reg[200][26]/P0001  , \wishbone_bd_ram_mem3_reg[200][27]/P0001  , \wishbone_bd_ram_mem3_reg[200][28]/P0001  , \wishbone_bd_ram_mem3_reg[200][29]/P0001  , \wishbone_bd_ram_mem3_reg[200][30]/P0001  , \wishbone_bd_ram_mem3_reg[200][31]/P0001  , \wishbone_bd_ram_mem3_reg[201][24]/P0001  , \wishbone_bd_ram_mem3_reg[201][25]/P0001  , \wishbone_bd_ram_mem3_reg[201][26]/P0001  , \wishbone_bd_ram_mem3_reg[201][27]/P0001  , \wishbone_bd_ram_mem3_reg[201][28]/P0001  , \wishbone_bd_ram_mem3_reg[201][29]/P0001  , \wishbone_bd_ram_mem3_reg[201][30]/P0001  , \wishbone_bd_ram_mem3_reg[201][31]/P0001  , \wishbone_bd_ram_mem3_reg[202][24]/P0001  , \wishbone_bd_ram_mem3_reg[202][25]/P0001  , \wishbone_bd_ram_mem3_reg[202][26]/P0001  , \wishbone_bd_ram_mem3_reg[202][27]/P0001  , \wishbone_bd_ram_mem3_reg[202][28]/P0001  , \wishbone_bd_ram_mem3_reg[202][29]/P0001  , \wishbone_bd_ram_mem3_reg[202][30]/P0001  , \wishbone_bd_ram_mem3_reg[202][31]/P0001  , \wishbone_bd_ram_mem3_reg[203][24]/P0001  , \wishbone_bd_ram_mem3_reg[203][25]/P0001  , \wishbone_bd_ram_mem3_reg[203][26]/P0001  , \wishbone_bd_ram_mem3_reg[203][27]/P0001  , \wishbone_bd_ram_mem3_reg[203][28]/P0001  , \wishbone_bd_ram_mem3_reg[203][29]/P0001  , \wishbone_bd_ram_mem3_reg[203][30]/P0001  , \wishbone_bd_ram_mem3_reg[203][31]/P0001  , \wishbone_bd_ram_mem3_reg[204][24]/P0001  , \wishbone_bd_ram_mem3_reg[204][25]/P0001  , \wishbone_bd_ram_mem3_reg[204][26]/P0001  , \wishbone_bd_ram_mem3_reg[204][27]/P0001  , \wishbone_bd_ram_mem3_reg[204][28]/P0001  , \wishbone_bd_ram_mem3_reg[204][29]/P0001  , \wishbone_bd_ram_mem3_reg[204][30]/P0001  , \wishbone_bd_ram_mem3_reg[204][31]/P0001  , \wishbone_bd_ram_mem3_reg[205][24]/P0001  , \wishbone_bd_ram_mem3_reg[205][25]/P0001  , \wishbone_bd_ram_mem3_reg[205][26]/P0001  , \wishbone_bd_ram_mem3_reg[205][27]/P0001  , \wishbone_bd_ram_mem3_reg[205][28]/P0001  , \wishbone_bd_ram_mem3_reg[205][29]/P0001  , \wishbone_bd_ram_mem3_reg[205][30]/P0001  , \wishbone_bd_ram_mem3_reg[205][31]/P0001  , \wishbone_bd_ram_mem3_reg[206][24]/P0001  , \wishbone_bd_ram_mem3_reg[206][25]/P0001  , \wishbone_bd_ram_mem3_reg[206][26]/P0001  , \wishbone_bd_ram_mem3_reg[206][27]/P0001  , \wishbone_bd_ram_mem3_reg[206][28]/P0001  , \wishbone_bd_ram_mem3_reg[206][29]/P0001  , \wishbone_bd_ram_mem3_reg[206][30]/P0001  , \wishbone_bd_ram_mem3_reg[206][31]/P0001  , \wishbone_bd_ram_mem3_reg[207][24]/P0001  , \wishbone_bd_ram_mem3_reg[207][25]/P0001  , \wishbone_bd_ram_mem3_reg[207][26]/P0001  , \wishbone_bd_ram_mem3_reg[207][27]/P0001  , \wishbone_bd_ram_mem3_reg[207][28]/P0001  , \wishbone_bd_ram_mem3_reg[207][29]/P0001  , \wishbone_bd_ram_mem3_reg[207][30]/P0001  , \wishbone_bd_ram_mem3_reg[207][31]/P0001  , \wishbone_bd_ram_mem3_reg[208][24]/P0001  , \wishbone_bd_ram_mem3_reg[208][25]/P0001  , \wishbone_bd_ram_mem3_reg[208][26]/P0001  , \wishbone_bd_ram_mem3_reg[208][27]/P0001  , \wishbone_bd_ram_mem3_reg[208][28]/P0001  , \wishbone_bd_ram_mem3_reg[208][29]/P0001  , \wishbone_bd_ram_mem3_reg[208][30]/P0001  , \wishbone_bd_ram_mem3_reg[208][31]/P0001  , \wishbone_bd_ram_mem3_reg[209][24]/P0001  , \wishbone_bd_ram_mem3_reg[209][25]/P0001  , \wishbone_bd_ram_mem3_reg[209][26]/P0001  , \wishbone_bd_ram_mem3_reg[209][27]/P0001  , \wishbone_bd_ram_mem3_reg[209][28]/P0001  , \wishbone_bd_ram_mem3_reg[209][29]/P0001  , \wishbone_bd_ram_mem3_reg[209][30]/P0001  , \wishbone_bd_ram_mem3_reg[209][31]/P0001  , \wishbone_bd_ram_mem3_reg[20][24]/P0001  , \wishbone_bd_ram_mem3_reg[20][25]/P0001  , \wishbone_bd_ram_mem3_reg[20][26]/P0001  , \wishbone_bd_ram_mem3_reg[20][27]/P0001  , \wishbone_bd_ram_mem3_reg[20][28]/P0001  , \wishbone_bd_ram_mem3_reg[20][29]/P0001  , \wishbone_bd_ram_mem3_reg[20][30]/P0001  , \wishbone_bd_ram_mem3_reg[20][31]/P0001  , \wishbone_bd_ram_mem3_reg[210][24]/P0001  , \wishbone_bd_ram_mem3_reg[210][25]/P0001  , \wishbone_bd_ram_mem3_reg[210][26]/P0001  , \wishbone_bd_ram_mem3_reg[210][27]/P0001  , \wishbone_bd_ram_mem3_reg[210][28]/P0001  , \wishbone_bd_ram_mem3_reg[210][29]/P0001  , \wishbone_bd_ram_mem3_reg[210][30]/P0001  , \wishbone_bd_ram_mem3_reg[210][31]/P0001  , \wishbone_bd_ram_mem3_reg[211][24]/P0001  , \wishbone_bd_ram_mem3_reg[211][25]/P0001  , \wishbone_bd_ram_mem3_reg[211][26]/P0001  , \wishbone_bd_ram_mem3_reg[211][27]/P0001  , \wishbone_bd_ram_mem3_reg[211][28]/P0001  , \wishbone_bd_ram_mem3_reg[211][29]/P0001  , \wishbone_bd_ram_mem3_reg[211][30]/P0001  , \wishbone_bd_ram_mem3_reg[211][31]/P0001  , \wishbone_bd_ram_mem3_reg[212][24]/P0001  , \wishbone_bd_ram_mem3_reg[212][25]/P0001  , \wishbone_bd_ram_mem3_reg[212][26]/P0001  , \wishbone_bd_ram_mem3_reg[212][27]/P0001  , \wishbone_bd_ram_mem3_reg[212][28]/P0001  , \wishbone_bd_ram_mem3_reg[212][29]/P0001  , \wishbone_bd_ram_mem3_reg[212][30]/P0001  , \wishbone_bd_ram_mem3_reg[212][31]/P0001  , \wishbone_bd_ram_mem3_reg[213][24]/P0001  , \wishbone_bd_ram_mem3_reg[213][25]/P0001  , \wishbone_bd_ram_mem3_reg[213][26]/P0001  , \wishbone_bd_ram_mem3_reg[213][27]/P0001  , \wishbone_bd_ram_mem3_reg[213][28]/P0001  , \wishbone_bd_ram_mem3_reg[213][29]/P0001  , \wishbone_bd_ram_mem3_reg[213][30]/P0001  , \wishbone_bd_ram_mem3_reg[213][31]/P0001  , \wishbone_bd_ram_mem3_reg[214][24]/P0001  , \wishbone_bd_ram_mem3_reg[214][25]/P0001  , \wishbone_bd_ram_mem3_reg[214][26]/P0001  , \wishbone_bd_ram_mem3_reg[214][27]/P0001  , \wishbone_bd_ram_mem3_reg[214][28]/P0001  , \wishbone_bd_ram_mem3_reg[214][29]/P0001  , \wishbone_bd_ram_mem3_reg[214][30]/P0001  , \wishbone_bd_ram_mem3_reg[214][31]/P0001  , \wishbone_bd_ram_mem3_reg[215][24]/P0001  , \wishbone_bd_ram_mem3_reg[215][25]/P0001  , \wishbone_bd_ram_mem3_reg[215][26]/P0001  , \wishbone_bd_ram_mem3_reg[215][27]/P0001  , \wishbone_bd_ram_mem3_reg[215][28]/P0001  , \wishbone_bd_ram_mem3_reg[215][29]/P0001  , \wishbone_bd_ram_mem3_reg[215][30]/P0001  , \wishbone_bd_ram_mem3_reg[215][31]/P0001  , \wishbone_bd_ram_mem3_reg[216][24]/P0001  , \wishbone_bd_ram_mem3_reg[216][25]/P0001  , \wishbone_bd_ram_mem3_reg[216][26]/P0001  , \wishbone_bd_ram_mem3_reg[216][27]/P0001  , \wishbone_bd_ram_mem3_reg[216][28]/P0001  , \wishbone_bd_ram_mem3_reg[216][29]/P0001  , \wishbone_bd_ram_mem3_reg[216][30]/P0001  , \wishbone_bd_ram_mem3_reg[216][31]/P0001  , \wishbone_bd_ram_mem3_reg[217][24]/P0001  , \wishbone_bd_ram_mem3_reg[217][25]/P0001  , \wishbone_bd_ram_mem3_reg[217][26]/P0001  , \wishbone_bd_ram_mem3_reg[217][27]/P0001  , \wishbone_bd_ram_mem3_reg[217][28]/P0001  , \wishbone_bd_ram_mem3_reg[217][29]/P0001  , \wishbone_bd_ram_mem3_reg[217][30]/P0001  , \wishbone_bd_ram_mem3_reg[217][31]/P0001  , \wishbone_bd_ram_mem3_reg[218][24]/P0001  , \wishbone_bd_ram_mem3_reg[218][25]/P0001  , \wishbone_bd_ram_mem3_reg[218][26]/P0001  , \wishbone_bd_ram_mem3_reg[218][27]/P0001  , \wishbone_bd_ram_mem3_reg[218][28]/P0001  , \wishbone_bd_ram_mem3_reg[218][29]/P0001  , \wishbone_bd_ram_mem3_reg[218][30]/P0001  , \wishbone_bd_ram_mem3_reg[218][31]/P0001  , \wishbone_bd_ram_mem3_reg[219][24]/P0001  , \wishbone_bd_ram_mem3_reg[219][25]/P0001  , \wishbone_bd_ram_mem3_reg[219][26]/P0001  , \wishbone_bd_ram_mem3_reg[219][27]/P0001  , \wishbone_bd_ram_mem3_reg[219][28]/P0001  , \wishbone_bd_ram_mem3_reg[219][29]/P0001  , \wishbone_bd_ram_mem3_reg[219][30]/P0001  , \wishbone_bd_ram_mem3_reg[219][31]/P0001  , \wishbone_bd_ram_mem3_reg[21][24]/P0001  , \wishbone_bd_ram_mem3_reg[21][25]/P0001  , \wishbone_bd_ram_mem3_reg[21][26]/P0001  , \wishbone_bd_ram_mem3_reg[21][27]/P0001  , \wishbone_bd_ram_mem3_reg[21][28]/P0001  , \wishbone_bd_ram_mem3_reg[21][29]/P0001  , \wishbone_bd_ram_mem3_reg[21][30]/P0001  , \wishbone_bd_ram_mem3_reg[21][31]/P0001  , \wishbone_bd_ram_mem3_reg[220][24]/P0001  , \wishbone_bd_ram_mem3_reg[220][25]/P0001  , \wishbone_bd_ram_mem3_reg[220][26]/P0001  , \wishbone_bd_ram_mem3_reg[220][27]/P0001  , \wishbone_bd_ram_mem3_reg[220][28]/P0001  , \wishbone_bd_ram_mem3_reg[220][29]/P0001  , \wishbone_bd_ram_mem3_reg[220][30]/P0001  , \wishbone_bd_ram_mem3_reg[220][31]/P0001  , \wishbone_bd_ram_mem3_reg[221][24]/P0001  , \wishbone_bd_ram_mem3_reg[221][25]/P0001  , \wishbone_bd_ram_mem3_reg[221][26]/P0001  , \wishbone_bd_ram_mem3_reg[221][27]/P0001  , \wishbone_bd_ram_mem3_reg[221][28]/P0001  , \wishbone_bd_ram_mem3_reg[221][29]/P0001  , \wishbone_bd_ram_mem3_reg[221][30]/P0001  , \wishbone_bd_ram_mem3_reg[221][31]/P0001  , \wishbone_bd_ram_mem3_reg[222][24]/P0001  , \wishbone_bd_ram_mem3_reg[222][25]/P0001  , \wishbone_bd_ram_mem3_reg[222][26]/P0001  , \wishbone_bd_ram_mem3_reg[222][27]/P0001  , \wishbone_bd_ram_mem3_reg[222][28]/P0001  , \wishbone_bd_ram_mem3_reg[222][29]/P0001  , \wishbone_bd_ram_mem3_reg[222][30]/P0001  , \wishbone_bd_ram_mem3_reg[222][31]/P0001  , \wishbone_bd_ram_mem3_reg[223][24]/P0001  , \wishbone_bd_ram_mem3_reg[223][25]/P0001  , \wishbone_bd_ram_mem3_reg[223][26]/P0001  , \wishbone_bd_ram_mem3_reg[223][27]/P0001  , \wishbone_bd_ram_mem3_reg[223][28]/P0001  , \wishbone_bd_ram_mem3_reg[223][29]/P0001  , \wishbone_bd_ram_mem3_reg[223][30]/P0001  , \wishbone_bd_ram_mem3_reg[223][31]/P0001  , \wishbone_bd_ram_mem3_reg[224][24]/P0001  , \wishbone_bd_ram_mem3_reg[224][25]/P0001  , \wishbone_bd_ram_mem3_reg[224][26]/P0001  , \wishbone_bd_ram_mem3_reg[224][27]/P0001  , \wishbone_bd_ram_mem3_reg[224][28]/P0001  , \wishbone_bd_ram_mem3_reg[224][29]/P0001  , \wishbone_bd_ram_mem3_reg[224][30]/P0001  , \wishbone_bd_ram_mem3_reg[224][31]/P0001  , \wishbone_bd_ram_mem3_reg[225][24]/P0001  , \wishbone_bd_ram_mem3_reg[225][25]/P0001  , \wishbone_bd_ram_mem3_reg[225][26]/P0001  , \wishbone_bd_ram_mem3_reg[225][27]/P0001  , \wishbone_bd_ram_mem3_reg[225][28]/P0001  , \wishbone_bd_ram_mem3_reg[225][29]/P0001  , \wishbone_bd_ram_mem3_reg[225][30]/P0001  , \wishbone_bd_ram_mem3_reg[225][31]/P0001  , \wishbone_bd_ram_mem3_reg[226][24]/P0001  , \wishbone_bd_ram_mem3_reg[226][25]/P0001  , \wishbone_bd_ram_mem3_reg[226][26]/P0001  , \wishbone_bd_ram_mem3_reg[226][27]/P0001  , \wishbone_bd_ram_mem3_reg[226][28]/P0001  , \wishbone_bd_ram_mem3_reg[226][29]/P0001  , \wishbone_bd_ram_mem3_reg[226][30]/P0001  , \wishbone_bd_ram_mem3_reg[226][31]/P0001  , \wishbone_bd_ram_mem3_reg[227][24]/P0001  , \wishbone_bd_ram_mem3_reg[227][25]/P0001  , \wishbone_bd_ram_mem3_reg[227][26]/P0001  , \wishbone_bd_ram_mem3_reg[227][27]/P0001  , \wishbone_bd_ram_mem3_reg[227][28]/P0001  , \wishbone_bd_ram_mem3_reg[227][29]/P0001  , \wishbone_bd_ram_mem3_reg[227][30]/P0001  , \wishbone_bd_ram_mem3_reg[227][31]/P0001  , \wishbone_bd_ram_mem3_reg[228][24]/P0001  , \wishbone_bd_ram_mem3_reg[228][25]/P0001  , \wishbone_bd_ram_mem3_reg[228][26]/P0001  , \wishbone_bd_ram_mem3_reg[228][27]/P0001  , \wishbone_bd_ram_mem3_reg[228][28]/P0001  , \wishbone_bd_ram_mem3_reg[228][29]/P0001  , \wishbone_bd_ram_mem3_reg[228][30]/P0001  , \wishbone_bd_ram_mem3_reg[228][31]/P0001  , \wishbone_bd_ram_mem3_reg[229][24]/P0001  , \wishbone_bd_ram_mem3_reg[229][25]/P0001  , \wishbone_bd_ram_mem3_reg[229][26]/P0001  , \wishbone_bd_ram_mem3_reg[229][27]/P0001  , \wishbone_bd_ram_mem3_reg[229][28]/P0001  , \wishbone_bd_ram_mem3_reg[229][29]/P0001  , \wishbone_bd_ram_mem3_reg[229][30]/P0001  , \wishbone_bd_ram_mem3_reg[229][31]/P0001  , \wishbone_bd_ram_mem3_reg[22][24]/P0001  , \wishbone_bd_ram_mem3_reg[22][25]/P0001  , \wishbone_bd_ram_mem3_reg[22][26]/P0001  , \wishbone_bd_ram_mem3_reg[22][27]/P0001  , \wishbone_bd_ram_mem3_reg[22][28]/P0001  , \wishbone_bd_ram_mem3_reg[22][29]/P0001  , \wishbone_bd_ram_mem3_reg[22][30]/P0001  , \wishbone_bd_ram_mem3_reg[22][31]/P0001  , \wishbone_bd_ram_mem3_reg[230][24]/P0001  , \wishbone_bd_ram_mem3_reg[230][25]/P0001  , \wishbone_bd_ram_mem3_reg[230][26]/P0001  , \wishbone_bd_ram_mem3_reg[230][27]/P0001  , \wishbone_bd_ram_mem3_reg[230][28]/P0001  , \wishbone_bd_ram_mem3_reg[230][29]/P0001  , \wishbone_bd_ram_mem3_reg[230][30]/P0001  , \wishbone_bd_ram_mem3_reg[230][31]/P0001  , \wishbone_bd_ram_mem3_reg[231][24]/P0001  , \wishbone_bd_ram_mem3_reg[231][25]/P0001  , \wishbone_bd_ram_mem3_reg[231][26]/P0001  , \wishbone_bd_ram_mem3_reg[231][27]/P0001  , \wishbone_bd_ram_mem3_reg[231][28]/P0001  , \wishbone_bd_ram_mem3_reg[231][29]/P0001  , \wishbone_bd_ram_mem3_reg[231][30]/P0001  , \wishbone_bd_ram_mem3_reg[231][31]/P0001  , \wishbone_bd_ram_mem3_reg[232][24]/P0001  , \wishbone_bd_ram_mem3_reg[232][25]/P0001  , \wishbone_bd_ram_mem3_reg[232][26]/P0001  , \wishbone_bd_ram_mem3_reg[232][27]/P0001  , \wishbone_bd_ram_mem3_reg[232][28]/P0001  , \wishbone_bd_ram_mem3_reg[232][29]/P0001  , \wishbone_bd_ram_mem3_reg[232][30]/P0001  , \wishbone_bd_ram_mem3_reg[232][31]/P0001  , \wishbone_bd_ram_mem3_reg[233][24]/P0001  , \wishbone_bd_ram_mem3_reg[233][25]/P0001  , \wishbone_bd_ram_mem3_reg[233][26]/P0001  , \wishbone_bd_ram_mem3_reg[233][27]/P0001  , \wishbone_bd_ram_mem3_reg[233][28]/P0001  , \wishbone_bd_ram_mem3_reg[233][29]/P0001  , \wishbone_bd_ram_mem3_reg[233][30]/P0001  , \wishbone_bd_ram_mem3_reg[233][31]/P0001  , \wishbone_bd_ram_mem3_reg[234][24]/P0001  , \wishbone_bd_ram_mem3_reg[234][25]/P0001  , \wishbone_bd_ram_mem3_reg[234][26]/P0001  , \wishbone_bd_ram_mem3_reg[234][27]/P0001  , \wishbone_bd_ram_mem3_reg[234][28]/P0001  , \wishbone_bd_ram_mem3_reg[234][29]/P0001  , \wishbone_bd_ram_mem3_reg[234][30]/P0001  , \wishbone_bd_ram_mem3_reg[234][31]/P0001  , \wishbone_bd_ram_mem3_reg[235][24]/P0001  , \wishbone_bd_ram_mem3_reg[235][25]/P0001  , \wishbone_bd_ram_mem3_reg[235][26]/P0001  , \wishbone_bd_ram_mem3_reg[235][27]/P0001  , \wishbone_bd_ram_mem3_reg[235][28]/P0001  , \wishbone_bd_ram_mem3_reg[235][29]/P0001  , \wishbone_bd_ram_mem3_reg[235][30]/P0001  , \wishbone_bd_ram_mem3_reg[235][31]/P0001  , \wishbone_bd_ram_mem3_reg[236][24]/P0001  , \wishbone_bd_ram_mem3_reg[236][25]/P0001  , \wishbone_bd_ram_mem3_reg[236][26]/P0001  , \wishbone_bd_ram_mem3_reg[236][27]/P0001  , \wishbone_bd_ram_mem3_reg[236][28]/P0001  , \wishbone_bd_ram_mem3_reg[236][29]/P0001  , \wishbone_bd_ram_mem3_reg[236][30]/P0001  , \wishbone_bd_ram_mem3_reg[236][31]/P0001  , \wishbone_bd_ram_mem3_reg[237][24]/P0001  , \wishbone_bd_ram_mem3_reg[237][25]/P0001  , \wishbone_bd_ram_mem3_reg[237][26]/P0001  , \wishbone_bd_ram_mem3_reg[237][27]/P0001  , \wishbone_bd_ram_mem3_reg[237][28]/P0001  , \wishbone_bd_ram_mem3_reg[237][29]/P0001  , \wishbone_bd_ram_mem3_reg[237][30]/P0001  , \wishbone_bd_ram_mem3_reg[237][31]/P0001  , \wishbone_bd_ram_mem3_reg[238][24]/P0001  , \wishbone_bd_ram_mem3_reg[238][25]/P0001  , \wishbone_bd_ram_mem3_reg[238][26]/P0001  , \wishbone_bd_ram_mem3_reg[238][27]/P0001  , \wishbone_bd_ram_mem3_reg[238][28]/P0001  , \wishbone_bd_ram_mem3_reg[238][29]/P0001  , \wishbone_bd_ram_mem3_reg[238][30]/P0001  , \wishbone_bd_ram_mem3_reg[238][31]/P0001  , \wishbone_bd_ram_mem3_reg[239][24]/P0001  , \wishbone_bd_ram_mem3_reg[239][25]/P0001  , \wishbone_bd_ram_mem3_reg[239][26]/P0001  , \wishbone_bd_ram_mem3_reg[239][27]/P0001  , \wishbone_bd_ram_mem3_reg[239][28]/P0001  , \wishbone_bd_ram_mem3_reg[239][29]/P0001  , \wishbone_bd_ram_mem3_reg[239][30]/P0001  , \wishbone_bd_ram_mem3_reg[239][31]/P0001  , \wishbone_bd_ram_mem3_reg[23][24]/P0001  , \wishbone_bd_ram_mem3_reg[23][25]/P0001  , \wishbone_bd_ram_mem3_reg[23][26]/P0001  , \wishbone_bd_ram_mem3_reg[23][27]/P0001  , \wishbone_bd_ram_mem3_reg[23][28]/P0001  , \wishbone_bd_ram_mem3_reg[23][29]/P0001  , \wishbone_bd_ram_mem3_reg[23][30]/P0001  , \wishbone_bd_ram_mem3_reg[23][31]/P0001  , \wishbone_bd_ram_mem3_reg[240][24]/P0001  , \wishbone_bd_ram_mem3_reg[240][25]/P0001  , \wishbone_bd_ram_mem3_reg[240][26]/P0001  , \wishbone_bd_ram_mem3_reg[240][27]/P0001  , \wishbone_bd_ram_mem3_reg[240][28]/P0001  , \wishbone_bd_ram_mem3_reg[240][29]/P0001  , \wishbone_bd_ram_mem3_reg[240][30]/P0001  , \wishbone_bd_ram_mem3_reg[240][31]/P0001  , \wishbone_bd_ram_mem3_reg[241][24]/P0001  , \wishbone_bd_ram_mem3_reg[241][25]/P0001  , \wishbone_bd_ram_mem3_reg[241][26]/P0001  , \wishbone_bd_ram_mem3_reg[241][27]/P0001  , \wishbone_bd_ram_mem3_reg[241][28]/P0001  , \wishbone_bd_ram_mem3_reg[241][29]/P0001  , \wishbone_bd_ram_mem3_reg[241][30]/P0001  , \wishbone_bd_ram_mem3_reg[241][31]/P0001  , \wishbone_bd_ram_mem3_reg[242][24]/P0001  , \wishbone_bd_ram_mem3_reg[242][25]/P0001  , \wishbone_bd_ram_mem3_reg[242][26]/P0001  , \wishbone_bd_ram_mem3_reg[242][27]/P0001  , \wishbone_bd_ram_mem3_reg[242][28]/P0001  , \wishbone_bd_ram_mem3_reg[242][29]/P0001  , \wishbone_bd_ram_mem3_reg[242][30]/P0001  , \wishbone_bd_ram_mem3_reg[242][31]/P0001  , \wishbone_bd_ram_mem3_reg[243][24]/P0001  , \wishbone_bd_ram_mem3_reg[243][25]/P0001  , \wishbone_bd_ram_mem3_reg[243][26]/P0001  , \wishbone_bd_ram_mem3_reg[243][27]/P0001  , \wishbone_bd_ram_mem3_reg[243][28]/P0001  , \wishbone_bd_ram_mem3_reg[243][29]/P0001  , \wishbone_bd_ram_mem3_reg[243][30]/P0001  , \wishbone_bd_ram_mem3_reg[243][31]/P0001  , \wishbone_bd_ram_mem3_reg[244][24]/P0001  , \wishbone_bd_ram_mem3_reg[244][25]/P0001  , \wishbone_bd_ram_mem3_reg[244][26]/P0001  , \wishbone_bd_ram_mem3_reg[244][27]/P0001  , \wishbone_bd_ram_mem3_reg[244][28]/P0001  , \wishbone_bd_ram_mem3_reg[244][29]/P0001  , \wishbone_bd_ram_mem3_reg[244][30]/P0001  , \wishbone_bd_ram_mem3_reg[244][31]/P0001  , \wishbone_bd_ram_mem3_reg[245][24]/P0001  , \wishbone_bd_ram_mem3_reg[245][25]/P0001  , \wishbone_bd_ram_mem3_reg[245][26]/P0001  , \wishbone_bd_ram_mem3_reg[245][27]/P0001  , \wishbone_bd_ram_mem3_reg[245][28]/P0001  , \wishbone_bd_ram_mem3_reg[245][29]/P0001  , \wishbone_bd_ram_mem3_reg[245][30]/P0001  , \wishbone_bd_ram_mem3_reg[245][31]/P0001  , \wishbone_bd_ram_mem3_reg[246][24]/P0001  , \wishbone_bd_ram_mem3_reg[246][25]/P0001  , \wishbone_bd_ram_mem3_reg[246][26]/P0001  , \wishbone_bd_ram_mem3_reg[246][27]/P0001  , \wishbone_bd_ram_mem3_reg[246][28]/P0001  , \wishbone_bd_ram_mem3_reg[246][29]/P0001  , \wishbone_bd_ram_mem3_reg[246][30]/P0001  , \wishbone_bd_ram_mem3_reg[246][31]/P0001  , \wishbone_bd_ram_mem3_reg[247][24]/P0001  , \wishbone_bd_ram_mem3_reg[247][25]/P0001  , \wishbone_bd_ram_mem3_reg[247][26]/P0001  , \wishbone_bd_ram_mem3_reg[247][27]/P0001  , \wishbone_bd_ram_mem3_reg[247][28]/P0001  , \wishbone_bd_ram_mem3_reg[247][29]/P0001  , \wishbone_bd_ram_mem3_reg[247][30]/P0001  , \wishbone_bd_ram_mem3_reg[247][31]/P0001  , \wishbone_bd_ram_mem3_reg[248][24]/P0001  , \wishbone_bd_ram_mem3_reg[248][25]/P0001  , \wishbone_bd_ram_mem3_reg[248][26]/P0001  , \wishbone_bd_ram_mem3_reg[248][27]/P0001  , \wishbone_bd_ram_mem3_reg[248][28]/P0001  , \wishbone_bd_ram_mem3_reg[248][29]/P0001  , \wishbone_bd_ram_mem3_reg[248][30]/P0001  , \wishbone_bd_ram_mem3_reg[248][31]/P0001  , \wishbone_bd_ram_mem3_reg[249][24]/P0001  , \wishbone_bd_ram_mem3_reg[249][25]/P0001  , \wishbone_bd_ram_mem3_reg[249][26]/P0001  , \wishbone_bd_ram_mem3_reg[249][27]/P0001  , \wishbone_bd_ram_mem3_reg[249][28]/P0001  , \wishbone_bd_ram_mem3_reg[249][29]/P0001  , \wishbone_bd_ram_mem3_reg[249][30]/P0001  , \wishbone_bd_ram_mem3_reg[249][31]/P0001  , \wishbone_bd_ram_mem3_reg[24][24]/P0001  , \wishbone_bd_ram_mem3_reg[24][25]/P0001  , \wishbone_bd_ram_mem3_reg[24][26]/P0001  , \wishbone_bd_ram_mem3_reg[24][27]/P0001  , \wishbone_bd_ram_mem3_reg[24][28]/P0001  , \wishbone_bd_ram_mem3_reg[24][29]/P0001  , \wishbone_bd_ram_mem3_reg[24][30]/P0001  , \wishbone_bd_ram_mem3_reg[24][31]/P0001  , \wishbone_bd_ram_mem3_reg[250][24]/P0001  , \wishbone_bd_ram_mem3_reg[250][25]/P0001  , \wishbone_bd_ram_mem3_reg[250][26]/P0001  , \wishbone_bd_ram_mem3_reg[250][27]/P0001  , \wishbone_bd_ram_mem3_reg[250][28]/P0001  , \wishbone_bd_ram_mem3_reg[250][29]/P0001  , \wishbone_bd_ram_mem3_reg[250][30]/P0001  , \wishbone_bd_ram_mem3_reg[250][31]/P0001  , \wishbone_bd_ram_mem3_reg[251][24]/P0001  , \wishbone_bd_ram_mem3_reg[251][25]/P0001  , \wishbone_bd_ram_mem3_reg[251][26]/P0001  , \wishbone_bd_ram_mem3_reg[251][27]/P0001  , \wishbone_bd_ram_mem3_reg[251][28]/P0001  , \wishbone_bd_ram_mem3_reg[251][29]/P0001  , \wishbone_bd_ram_mem3_reg[251][30]/P0001  , \wishbone_bd_ram_mem3_reg[251][31]/P0001  , \wishbone_bd_ram_mem3_reg[252][24]/P0001  , \wishbone_bd_ram_mem3_reg[252][25]/P0001  , \wishbone_bd_ram_mem3_reg[252][26]/P0001  , \wishbone_bd_ram_mem3_reg[252][27]/P0001  , \wishbone_bd_ram_mem3_reg[252][28]/P0001  , \wishbone_bd_ram_mem3_reg[252][29]/P0001  , \wishbone_bd_ram_mem3_reg[252][30]/P0001  , \wishbone_bd_ram_mem3_reg[252][31]/P0001  , \wishbone_bd_ram_mem3_reg[253][24]/P0001  , \wishbone_bd_ram_mem3_reg[253][25]/P0001  , \wishbone_bd_ram_mem3_reg[253][26]/P0001  , \wishbone_bd_ram_mem3_reg[253][27]/P0001  , \wishbone_bd_ram_mem3_reg[253][28]/P0001  , \wishbone_bd_ram_mem3_reg[253][29]/P0001  , \wishbone_bd_ram_mem3_reg[253][30]/P0001  , \wishbone_bd_ram_mem3_reg[253][31]/P0001  , \wishbone_bd_ram_mem3_reg[254][24]/P0001  , \wishbone_bd_ram_mem3_reg[254][25]/P0001  , \wishbone_bd_ram_mem3_reg[254][26]/P0001  , \wishbone_bd_ram_mem3_reg[254][27]/P0001  , \wishbone_bd_ram_mem3_reg[254][28]/P0001  , \wishbone_bd_ram_mem3_reg[254][29]/P0001  , \wishbone_bd_ram_mem3_reg[254][30]/P0001  , \wishbone_bd_ram_mem3_reg[254][31]/P0001  , \wishbone_bd_ram_mem3_reg[255][24]/P0001  , \wishbone_bd_ram_mem3_reg[255][25]/P0001  , \wishbone_bd_ram_mem3_reg[255][26]/P0001  , \wishbone_bd_ram_mem3_reg[255][27]/P0001  , \wishbone_bd_ram_mem3_reg[255][28]/P0001  , \wishbone_bd_ram_mem3_reg[255][29]/P0001  , \wishbone_bd_ram_mem3_reg[255][30]/P0001  , \wishbone_bd_ram_mem3_reg[255][31]/P0001  , \wishbone_bd_ram_mem3_reg[25][24]/P0001  , \wishbone_bd_ram_mem3_reg[25][25]/P0001  , \wishbone_bd_ram_mem3_reg[25][26]/P0001  , \wishbone_bd_ram_mem3_reg[25][27]/P0001  , \wishbone_bd_ram_mem3_reg[25][28]/P0001  , \wishbone_bd_ram_mem3_reg[25][29]/P0001  , \wishbone_bd_ram_mem3_reg[25][30]/P0001  , \wishbone_bd_ram_mem3_reg[25][31]/P0001  , \wishbone_bd_ram_mem3_reg[26][24]/P0001  , \wishbone_bd_ram_mem3_reg[26][25]/P0001  , \wishbone_bd_ram_mem3_reg[26][26]/P0001  , \wishbone_bd_ram_mem3_reg[26][27]/P0001  , \wishbone_bd_ram_mem3_reg[26][28]/P0001  , \wishbone_bd_ram_mem3_reg[26][29]/P0001  , \wishbone_bd_ram_mem3_reg[26][30]/P0001  , \wishbone_bd_ram_mem3_reg[26][31]/P0001  , \wishbone_bd_ram_mem3_reg[27][24]/P0001  , \wishbone_bd_ram_mem3_reg[27][25]/P0001  , \wishbone_bd_ram_mem3_reg[27][26]/P0001  , \wishbone_bd_ram_mem3_reg[27][27]/P0001  , \wishbone_bd_ram_mem3_reg[27][28]/P0001  , \wishbone_bd_ram_mem3_reg[27][29]/P0001  , \wishbone_bd_ram_mem3_reg[27][30]/P0001  , \wishbone_bd_ram_mem3_reg[27][31]/P0001  , \wishbone_bd_ram_mem3_reg[28][24]/P0001  , \wishbone_bd_ram_mem3_reg[28][25]/P0001  , \wishbone_bd_ram_mem3_reg[28][26]/P0001  , \wishbone_bd_ram_mem3_reg[28][27]/P0001  , \wishbone_bd_ram_mem3_reg[28][28]/P0001  , \wishbone_bd_ram_mem3_reg[28][29]/P0001  , \wishbone_bd_ram_mem3_reg[28][30]/P0001  , \wishbone_bd_ram_mem3_reg[28][31]/P0001  , \wishbone_bd_ram_mem3_reg[29][24]/P0001  , \wishbone_bd_ram_mem3_reg[29][25]/P0001  , \wishbone_bd_ram_mem3_reg[29][26]/P0001  , \wishbone_bd_ram_mem3_reg[29][27]/P0001  , \wishbone_bd_ram_mem3_reg[29][28]/P0001  , \wishbone_bd_ram_mem3_reg[29][29]/P0001  , \wishbone_bd_ram_mem3_reg[29][30]/P0001  , \wishbone_bd_ram_mem3_reg[29][31]/P0001  , \wishbone_bd_ram_mem3_reg[2][24]/P0001  , \wishbone_bd_ram_mem3_reg[2][25]/P0001  , \wishbone_bd_ram_mem3_reg[2][26]/P0001  , \wishbone_bd_ram_mem3_reg[2][27]/P0001  , \wishbone_bd_ram_mem3_reg[2][28]/P0001  , \wishbone_bd_ram_mem3_reg[2][29]/P0001  , \wishbone_bd_ram_mem3_reg[2][30]/P0001  , \wishbone_bd_ram_mem3_reg[2][31]/P0001  , \wishbone_bd_ram_mem3_reg[30][24]/P0001  , \wishbone_bd_ram_mem3_reg[30][25]/P0001  , \wishbone_bd_ram_mem3_reg[30][26]/P0001  , \wishbone_bd_ram_mem3_reg[30][27]/P0001  , \wishbone_bd_ram_mem3_reg[30][28]/P0001  , \wishbone_bd_ram_mem3_reg[30][29]/P0001  , \wishbone_bd_ram_mem3_reg[30][30]/P0001  , \wishbone_bd_ram_mem3_reg[30][31]/P0001  , \wishbone_bd_ram_mem3_reg[31][24]/P0001  , \wishbone_bd_ram_mem3_reg[31][25]/P0001  , \wishbone_bd_ram_mem3_reg[31][26]/P0001  , \wishbone_bd_ram_mem3_reg[31][27]/P0001  , \wishbone_bd_ram_mem3_reg[31][28]/P0001  , \wishbone_bd_ram_mem3_reg[31][29]/P0001  , \wishbone_bd_ram_mem3_reg[31][30]/P0001  , \wishbone_bd_ram_mem3_reg[31][31]/P0001  , \wishbone_bd_ram_mem3_reg[32][24]/P0001  , \wishbone_bd_ram_mem3_reg[32][25]/P0001  , \wishbone_bd_ram_mem3_reg[32][26]/P0001  , \wishbone_bd_ram_mem3_reg[32][27]/P0001  , \wishbone_bd_ram_mem3_reg[32][28]/P0001  , \wishbone_bd_ram_mem3_reg[32][29]/P0001  , \wishbone_bd_ram_mem3_reg[32][30]/P0001  , \wishbone_bd_ram_mem3_reg[32][31]/P0001  , \wishbone_bd_ram_mem3_reg[33][24]/P0001  , \wishbone_bd_ram_mem3_reg[33][25]/P0001  , \wishbone_bd_ram_mem3_reg[33][26]/P0001  , \wishbone_bd_ram_mem3_reg[33][27]/P0001  , \wishbone_bd_ram_mem3_reg[33][28]/P0001  , \wishbone_bd_ram_mem3_reg[33][29]/P0001  , \wishbone_bd_ram_mem3_reg[33][30]/P0001  , \wishbone_bd_ram_mem3_reg[33][31]/P0001  , \wishbone_bd_ram_mem3_reg[34][24]/P0001  , \wishbone_bd_ram_mem3_reg[34][25]/P0001  , \wishbone_bd_ram_mem3_reg[34][26]/P0001  , \wishbone_bd_ram_mem3_reg[34][27]/P0001  , \wishbone_bd_ram_mem3_reg[34][28]/P0001  , \wishbone_bd_ram_mem3_reg[34][29]/P0001  , \wishbone_bd_ram_mem3_reg[34][30]/P0001  , \wishbone_bd_ram_mem3_reg[34][31]/P0001  , \wishbone_bd_ram_mem3_reg[35][24]/P0001  , \wishbone_bd_ram_mem3_reg[35][25]/P0001  , \wishbone_bd_ram_mem3_reg[35][26]/P0001  , \wishbone_bd_ram_mem3_reg[35][27]/P0001  , \wishbone_bd_ram_mem3_reg[35][28]/P0001  , \wishbone_bd_ram_mem3_reg[35][29]/P0001  , \wishbone_bd_ram_mem3_reg[35][30]/P0001  , \wishbone_bd_ram_mem3_reg[35][31]/P0001  , \wishbone_bd_ram_mem3_reg[36][24]/P0001  , \wishbone_bd_ram_mem3_reg[36][25]/P0001  , \wishbone_bd_ram_mem3_reg[36][26]/P0001  , \wishbone_bd_ram_mem3_reg[36][27]/P0001  , \wishbone_bd_ram_mem3_reg[36][28]/P0001  , \wishbone_bd_ram_mem3_reg[36][29]/P0001  , \wishbone_bd_ram_mem3_reg[36][30]/P0001  , \wishbone_bd_ram_mem3_reg[36][31]/P0001  , \wishbone_bd_ram_mem3_reg[37][24]/P0001  , \wishbone_bd_ram_mem3_reg[37][25]/P0001  , \wishbone_bd_ram_mem3_reg[37][26]/P0001  , \wishbone_bd_ram_mem3_reg[37][27]/P0001  , \wishbone_bd_ram_mem3_reg[37][28]/P0001  , \wishbone_bd_ram_mem3_reg[37][29]/P0001  , \wishbone_bd_ram_mem3_reg[37][30]/P0001  , \wishbone_bd_ram_mem3_reg[37][31]/P0001  , \wishbone_bd_ram_mem3_reg[38][24]/P0001  , \wishbone_bd_ram_mem3_reg[38][25]/P0001  , \wishbone_bd_ram_mem3_reg[38][26]/P0001  , \wishbone_bd_ram_mem3_reg[38][27]/P0001  , \wishbone_bd_ram_mem3_reg[38][28]/P0001  , \wishbone_bd_ram_mem3_reg[38][29]/P0001  , \wishbone_bd_ram_mem3_reg[38][30]/P0001  , \wishbone_bd_ram_mem3_reg[38][31]/P0001  , \wishbone_bd_ram_mem3_reg[39][24]/P0001  , \wishbone_bd_ram_mem3_reg[39][25]/P0001  , \wishbone_bd_ram_mem3_reg[39][26]/P0001  , \wishbone_bd_ram_mem3_reg[39][27]/P0001  , \wishbone_bd_ram_mem3_reg[39][28]/P0001  , \wishbone_bd_ram_mem3_reg[39][29]/P0001  , \wishbone_bd_ram_mem3_reg[39][30]/P0001  , \wishbone_bd_ram_mem3_reg[39][31]/P0001  , \wishbone_bd_ram_mem3_reg[3][24]/P0001  , \wishbone_bd_ram_mem3_reg[3][25]/P0001  , \wishbone_bd_ram_mem3_reg[3][26]/P0001  , \wishbone_bd_ram_mem3_reg[3][27]/P0001  , \wishbone_bd_ram_mem3_reg[3][28]/P0001  , \wishbone_bd_ram_mem3_reg[3][29]/P0001  , \wishbone_bd_ram_mem3_reg[3][30]/P0001  , \wishbone_bd_ram_mem3_reg[3][31]/P0001  , \wishbone_bd_ram_mem3_reg[40][24]/P0001  , \wishbone_bd_ram_mem3_reg[40][25]/P0001  , \wishbone_bd_ram_mem3_reg[40][26]/P0001  , \wishbone_bd_ram_mem3_reg[40][27]/P0001  , \wishbone_bd_ram_mem3_reg[40][28]/P0001  , \wishbone_bd_ram_mem3_reg[40][29]/P0001  , \wishbone_bd_ram_mem3_reg[40][30]/P0001  , \wishbone_bd_ram_mem3_reg[40][31]/P0001  , \wishbone_bd_ram_mem3_reg[41][24]/P0001  , \wishbone_bd_ram_mem3_reg[41][25]/P0001  , \wishbone_bd_ram_mem3_reg[41][26]/P0001  , \wishbone_bd_ram_mem3_reg[41][27]/P0001  , \wishbone_bd_ram_mem3_reg[41][28]/P0001  , \wishbone_bd_ram_mem3_reg[41][29]/P0001  , \wishbone_bd_ram_mem3_reg[41][30]/P0001  , \wishbone_bd_ram_mem3_reg[41][31]/P0001  , \wishbone_bd_ram_mem3_reg[42][24]/P0001  , \wishbone_bd_ram_mem3_reg[42][25]/P0001  , \wishbone_bd_ram_mem3_reg[42][26]/P0001  , \wishbone_bd_ram_mem3_reg[42][27]/P0001  , \wishbone_bd_ram_mem3_reg[42][28]/P0001  , \wishbone_bd_ram_mem3_reg[42][29]/P0001  , \wishbone_bd_ram_mem3_reg[42][30]/P0001  , \wishbone_bd_ram_mem3_reg[42][31]/P0001  , \wishbone_bd_ram_mem3_reg[43][24]/P0001  , \wishbone_bd_ram_mem3_reg[43][25]/P0001  , \wishbone_bd_ram_mem3_reg[43][26]/P0001  , \wishbone_bd_ram_mem3_reg[43][27]/P0001  , \wishbone_bd_ram_mem3_reg[43][28]/P0001  , \wishbone_bd_ram_mem3_reg[43][29]/P0001  , \wishbone_bd_ram_mem3_reg[43][30]/P0001  , \wishbone_bd_ram_mem3_reg[43][31]/P0001  , \wishbone_bd_ram_mem3_reg[44][24]/P0001  , \wishbone_bd_ram_mem3_reg[44][25]/P0001  , \wishbone_bd_ram_mem3_reg[44][26]/P0001  , \wishbone_bd_ram_mem3_reg[44][27]/P0001  , \wishbone_bd_ram_mem3_reg[44][28]/P0001  , \wishbone_bd_ram_mem3_reg[44][29]/P0001  , \wishbone_bd_ram_mem3_reg[44][30]/P0001  , \wishbone_bd_ram_mem3_reg[44][31]/P0001  , \wishbone_bd_ram_mem3_reg[45][24]/P0001  , \wishbone_bd_ram_mem3_reg[45][25]/P0001  , \wishbone_bd_ram_mem3_reg[45][26]/P0001  , \wishbone_bd_ram_mem3_reg[45][27]/P0001  , \wishbone_bd_ram_mem3_reg[45][28]/P0001  , \wishbone_bd_ram_mem3_reg[45][29]/P0001  , \wishbone_bd_ram_mem3_reg[45][30]/P0001  , \wishbone_bd_ram_mem3_reg[45][31]/P0001  , \wishbone_bd_ram_mem3_reg[46][24]/P0001  , \wishbone_bd_ram_mem3_reg[46][25]/P0001  , \wishbone_bd_ram_mem3_reg[46][26]/P0001  , \wishbone_bd_ram_mem3_reg[46][27]/P0001  , \wishbone_bd_ram_mem3_reg[46][28]/P0001  , \wishbone_bd_ram_mem3_reg[46][29]/P0001  , \wishbone_bd_ram_mem3_reg[46][30]/P0001  , \wishbone_bd_ram_mem3_reg[46][31]/P0001  , \wishbone_bd_ram_mem3_reg[47][24]/P0001  , \wishbone_bd_ram_mem3_reg[47][25]/P0001  , \wishbone_bd_ram_mem3_reg[47][26]/P0001  , \wishbone_bd_ram_mem3_reg[47][27]/P0001  , \wishbone_bd_ram_mem3_reg[47][28]/P0001  , \wishbone_bd_ram_mem3_reg[47][29]/P0001  , \wishbone_bd_ram_mem3_reg[47][30]/P0001  , \wishbone_bd_ram_mem3_reg[47][31]/P0001  , \wishbone_bd_ram_mem3_reg[48][24]/P0001  , \wishbone_bd_ram_mem3_reg[48][25]/P0001  , \wishbone_bd_ram_mem3_reg[48][26]/P0001  , \wishbone_bd_ram_mem3_reg[48][27]/P0001  , \wishbone_bd_ram_mem3_reg[48][28]/P0001  , \wishbone_bd_ram_mem3_reg[48][29]/P0001  , \wishbone_bd_ram_mem3_reg[48][30]/P0001  , \wishbone_bd_ram_mem3_reg[48][31]/P0001  , \wishbone_bd_ram_mem3_reg[49][24]/P0001  , \wishbone_bd_ram_mem3_reg[49][25]/P0001  , \wishbone_bd_ram_mem3_reg[49][26]/P0001  , \wishbone_bd_ram_mem3_reg[49][27]/P0001  , \wishbone_bd_ram_mem3_reg[49][28]/P0001  , \wishbone_bd_ram_mem3_reg[49][29]/P0001  , \wishbone_bd_ram_mem3_reg[49][30]/P0001  , \wishbone_bd_ram_mem3_reg[49][31]/P0001  , \wishbone_bd_ram_mem3_reg[4][24]/P0001  , \wishbone_bd_ram_mem3_reg[4][25]/P0001  , \wishbone_bd_ram_mem3_reg[4][26]/P0001  , \wishbone_bd_ram_mem3_reg[4][27]/P0001  , \wishbone_bd_ram_mem3_reg[4][28]/P0001  , \wishbone_bd_ram_mem3_reg[4][29]/P0001  , \wishbone_bd_ram_mem3_reg[4][30]/P0001  , \wishbone_bd_ram_mem3_reg[4][31]/P0001  , \wishbone_bd_ram_mem3_reg[50][24]/P0001  , \wishbone_bd_ram_mem3_reg[50][25]/P0001  , \wishbone_bd_ram_mem3_reg[50][26]/P0001  , \wishbone_bd_ram_mem3_reg[50][27]/P0001  , \wishbone_bd_ram_mem3_reg[50][28]/P0001  , \wishbone_bd_ram_mem3_reg[50][29]/P0001  , \wishbone_bd_ram_mem3_reg[50][30]/P0001  , \wishbone_bd_ram_mem3_reg[50][31]/P0001  , \wishbone_bd_ram_mem3_reg[51][24]/P0001  , \wishbone_bd_ram_mem3_reg[51][25]/P0001  , \wishbone_bd_ram_mem3_reg[51][26]/P0001  , \wishbone_bd_ram_mem3_reg[51][27]/P0001  , \wishbone_bd_ram_mem3_reg[51][28]/P0001  , \wishbone_bd_ram_mem3_reg[51][29]/P0001  , \wishbone_bd_ram_mem3_reg[51][30]/P0001  , \wishbone_bd_ram_mem3_reg[51][31]/P0001  , \wishbone_bd_ram_mem3_reg[52][24]/P0001  , \wishbone_bd_ram_mem3_reg[52][25]/P0001  , \wishbone_bd_ram_mem3_reg[52][26]/P0001  , \wishbone_bd_ram_mem3_reg[52][27]/P0001  , \wishbone_bd_ram_mem3_reg[52][28]/P0001  , \wishbone_bd_ram_mem3_reg[52][29]/P0001  , \wishbone_bd_ram_mem3_reg[52][30]/P0001  , \wishbone_bd_ram_mem3_reg[52][31]/P0001  , \wishbone_bd_ram_mem3_reg[53][24]/P0001  , \wishbone_bd_ram_mem3_reg[53][25]/P0001  , \wishbone_bd_ram_mem3_reg[53][26]/P0001  , \wishbone_bd_ram_mem3_reg[53][27]/P0001  , \wishbone_bd_ram_mem3_reg[53][28]/P0001  , \wishbone_bd_ram_mem3_reg[53][29]/P0001  , \wishbone_bd_ram_mem3_reg[53][30]/P0001  , \wishbone_bd_ram_mem3_reg[53][31]/P0001  , \wishbone_bd_ram_mem3_reg[54][24]/P0001  , \wishbone_bd_ram_mem3_reg[54][25]/P0001  , \wishbone_bd_ram_mem3_reg[54][26]/P0001  , \wishbone_bd_ram_mem3_reg[54][27]/P0001  , \wishbone_bd_ram_mem3_reg[54][28]/P0001  , \wishbone_bd_ram_mem3_reg[54][29]/P0001  , \wishbone_bd_ram_mem3_reg[54][30]/P0001  , \wishbone_bd_ram_mem3_reg[54][31]/P0001  , \wishbone_bd_ram_mem3_reg[55][24]/P0001  , \wishbone_bd_ram_mem3_reg[55][25]/P0001  , \wishbone_bd_ram_mem3_reg[55][26]/P0001  , \wishbone_bd_ram_mem3_reg[55][27]/P0001  , \wishbone_bd_ram_mem3_reg[55][28]/P0001  , \wishbone_bd_ram_mem3_reg[55][29]/P0001  , \wishbone_bd_ram_mem3_reg[55][30]/P0001  , \wishbone_bd_ram_mem3_reg[55][31]/P0001  , \wishbone_bd_ram_mem3_reg[56][24]/P0001  , \wishbone_bd_ram_mem3_reg[56][25]/P0001  , \wishbone_bd_ram_mem3_reg[56][26]/P0001  , \wishbone_bd_ram_mem3_reg[56][27]/P0001  , \wishbone_bd_ram_mem3_reg[56][28]/P0001  , \wishbone_bd_ram_mem3_reg[56][29]/P0001  , \wishbone_bd_ram_mem3_reg[56][30]/P0001  , \wishbone_bd_ram_mem3_reg[56][31]/P0001  , \wishbone_bd_ram_mem3_reg[57][24]/P0001  , \wishbone_bd_ram_mem3_reg[57][25]/P0001  , \wishbone_bd_ram_mem3_reg[57][26]/P0001  , \wishbone_bd_ram_mem3_reg[57][27]/P0001  , \wishbone_bd_ram_mem3_reg[57][28]/P0001  , \wishbone_bd_ram_mem3_reg[57][29]/P0001  , \wishbone_bd_ram_mem3_reg[57][30]/P0001  , \wishbone_bd_ram_mem3_reg[57][31]/P0001  , \wishbone_bd_ram_mem3_reg[58][24]/P0001  , \wishbone_bd_ram_mem3_reg[58][25]/P0001  , \wishbone_bd_ram_mem3_reg[58][26]/P0001  , \wishbone_bd_ram_mem3_reg[58][27]/P0001  , \wishbone_bd_ram_mem3_reg[58][28]/P0001  , \wishbone_bd_ram_mem3_reg[58][29]/P0001  , \wishbone_bd_ram_mem3_reg[58][30]/P0001  , \wishbone_bd_ram_mem3_reg[58][31]/P0001  , \wishbone_bd_ram_mem3_reg[59][24]/P0001  , \wishbone_bd_ram_mem3_reg[59][25]/P0001  , \wishbone_bd_ram_mem3_reg[59][26]/P0001  , \wishbone_bd_ram_mem3_reg[59][27]/P0001  , \wishbone_bd_ram_mem3_reg[59][28]/P0001  , \wishbone_bd_ram_mem3_reg[59][29]/P0001  , \wishbone_bd_ram_mem3_reg[59][30]/P0001  , \wishbone_bd_ram_mem3_reg[59][31]/P0001  , \wishbone_bd_ram_mem3_reg[5][24]/P0001  , \wishbone_bd_ram_mem3_reg[5][25]/P0001  , \wishbone_bd_ram_mem3_reg[5][26]/P0001  , \wishbone_bd_ram_mem3_reg[5][27]/P0001  , \wishbone_bd_ram_mem3_reg[5][28]/P0001  , \wishbone_bd_ram_mem3_reg[5][29]/P0001  , \wishbone_bd_ram_mem3_reg[5][30]/P0001  , \wishbone_bd_ram_mem3_reg[5][31]/P0001  , \wishbone_bd_ram_mem3_reg[60][24]/P0001  , \wishbone_bd_ram_mem3_reg[60][25]/P0001  , \wishbone_bd_ram_mem3_reg[60][26]/P0001  , \wishbone_bd_ram_mem3_reg[60][27]/P0001  , \wishbone_bd_ram_mem3_reg[60][28]/P0001  , \wishbone_bd_ram_mem3_reg[60][29]/P0001  , \wishbone_bd_ram_mem3_reg[60][30]/P0001  , \wishbone_bd_ram_mem3_reg[60][31]/P0001  , \wishbone_bd_ram_mem3_reg[61][24]/P0001  , \wishbone_bd_ram_mem3_reg[61][25]/P0001  , \wishbone_bd_ram_mem3_reg[61][26]/P0001  , \wishbone_bd_ram_mem3_reg[61][27]/P0001  , \wishbone_bd_ram_mem3_reg[61][28]/P0001  , \wishbone_bd_ram_mem3_reg[61][29]/P0001  , \wishbone_bd_ram_mem3_reg[61][30]/P0001  , \wishbone_bd_ram_mem3_reg[61][31]/P0001  , \wishbone_bd_ram_mem3_reg[62][24]/P0001  , \wishbone_bd_ram_mem3_reg[62][25]/P0001  , \wishbone_bd_ram_mem3_reg[62][26]/P0001  , \wishbone_bd_ram_mem3_reg[62][27]/P0001  , \wishbone_bd_ram_mem3_reg[62][28]/P0001  , \wishbone_bd_ram_mem3_reg[62][29]/P0001  , \wishbone_bd_ram_mem3_reg[62][30]/P0001  , \wishbone_bd_ram_mem3_reg[62][31]/P0001  , \wishbone_bd_ram_mem3_reg[63][24]/P0001  , \wishbone_bd_ram_mem3_reg[63][25]/P0001  , \wishbone_bd_ram_mem3_reg[63][26]/P0001  , \wishbone_bd_ram_mem3_reg[63][27]/P0001  , \wishbone_bd_ram_mem3_reg[63][28]/P0001  , \wishbone_bd_ram_mem3_reg[63][29]/P0001  , \wishbone_bd_ram_mem3_reg[63][30]/P0001  , \wishbone_bd_ram_mem3_reg[63][31]/P0001  , \wishbone_bd_ram_mem3_reg[64][24]/P0001  , \wishbone_bd_ram_mem3_reg[64][25]/P0001  , \wishbone_bd_ram_mem3_reg[64][26]/P0001  , \wishbone_bd_ram_mem3_reg[64][27]/P0001  , \wishbone_bd_ram_mem3_reg[64][28]/P0001  , \wishbone_bd_ram_mem3_reg[64][29]/P0001  , \wishbone_bd_ram_mem3_reg[64][30]/P0001  , \wishbone_bd_ram_mem3_reg[64][31]/P0001  , \wishbone_bd_ram_mem3_reg[65][24]/P0001  , \wishbone_bd_ram_mem3_reg[65][25]/P0001  , \wishbone_bd_ram_mem3_reg[65][26]/P0001  , \wishbone_bd_ram_mem3_reg[65][27]/P0001  , \wishbone_bd_ram_mem3_reg[65][28]/P0001  , \wishbone_bd_ram_mem3_reg[65][29]/P0001  , \wishbone_bd_ram_mem3_reg[65][30]/P0001  , \wishbone_bd_ram_mem3_reg[65][31]/P0001  , \wishbone_bd_ram_mem3_reg[66][24]/P0001  , \wishbone_bd_ram_mem3_reg[66][25]/P0001  , \wishbone_bd_ram_mem3_reg[66][26]/P0001  , \wishbone_bd_ram_mem3_reg[66][27]/P0001  , \wishbone_bd_ram_mem3_reg[66][28]/P0001  , \wishbone_bd_ram_mem3_reg[66][29]/P0001  , \wishbone_bd_ram_mem3_reg[66][30]/P0001  , \wishbone_bd_ram_mem3_reg[66][31]/P0001  , \wishbone_bd_ram_mem3_reg[67][24]/P0001  , \wishbone_bd_ram_mem3_reg[67][25]/P0001  , \wishbone_bd_ram_mem3_reg[67][26]/P0001  , \wishbone_bd_ram_mem3_reg[67][27]/P0001  , \wishbone_bd_ram_mem3_reg[67][28]/P0001  , \wishbone_bd_ram_mem3_reg[67][29]/P0001  , \wishbone_bd_ram_mem3_reg[67][30]/P0001  , \wishbone_bd_ram_mem3_reg[67][31]/P0001  , \wishbone_bd_ram_mem3_reg[68][24]/P0001  , \wishbone_bd_ram_mem3_reg[68][25]/P0001  , \wishbone_bd_ram_mem3_reg[68][26]/P0001  , \wishbone_bd_ram_mem3_reg[68][27]/P0001  , \wishbone_bd_ram_mem3_reg[68][28]/P0001  , \wishbone_bd_ram_mem3_reg[68][29]/P0001  , \wishbone_bd_ram_mem3_reg[68][30]/P0001  , \wishbone_bd_ram_mem3_reg[68][31]/P0001  , \wishbone_bd_ram_mem3_reg[69][24]/P0001  , \wishbone_bd_ram_mem3_reg[69][25]/P0001  , \wishbone_bd_ram_mem3_reg[69][26]/P0001  , \wishbone_bd_ram_mem3_reg[69][27]/P0001  , \wishbone_bd_ram_mem3_reg[69][28]/P0001  , \wishbone_bd_ram_mem3_reg[69][29]/P0001  , \wishbone_bd_ram_mem3_reg[69][30]/P0001  , \wishbone_bd_ram_mem3_reg[69][31]/P0001  , \wishbone_bd_ram_mem3_reg[6][24]/P0001  , \wishbone_bd_ram_mem3_reg[6][25]/P0001  , \wishbone_bd_ram_mem3_reg[6][26]/P0001  , \wishbone_bd_ram_mem3_reg[6][27]/P0001  , \wishbone_bd_ram_mem3_reg[6][28]/P0001  , \wishbone_bd_ram_mem3_reg[6][29]/P0001  , \wishbone_bd_ram_mem3_reg[6][30]/P0001  , \wishbone_bd_ram_mem3_reg[6][31]/P0001  , \wishbone_bd_ram_mem3_reg[70][24]/P0001  , \wishbone_bd_ram_mem3_reg[70][25]/P0001  , \wishbone_bd_ram_mem3_reg[70][26]/P0001  , \wishbone_bd_ram_mem3_reg[70][27]/P0001  , \wishbone_bd_ram_mem3_reg[70][28]/P0001  , \wishbone_bd_ram_mem3_reg[70][29]/P0001  , \wishbone_bd_ram_mem3_reg[70][30]/P0001  , \wishbone_bd_ram_mem3_reg[70][31]/P0001  , \wishbone_bd_ram_mem3_reg[71][24]/P0001  , \wishbone_bd_ram_mem3_reg[71][25]/P0001  , \wishbone_bd_ram_mem3_reg[71][26]/P0001  , \wishbone_bd_ram_mem3_reg[71][27]/P0001  , \wishbone_bd_ram_mem3_reg[71][28]/P0001  , \wishbone_bd_ram_mem3_reg[71][29]/P0001  , \wishbone_bd_ram_mem3_reg[71][30]/P0001  , \wishbone_bd_ram_mem3_reg[71][31]/P0001  , \wishbone_bd_ram_mem3_reg[72][24]/P0001  , \wishbone_bd_ram_mem3_reg[72][25]/P0001  , \wishbone_bd_ram_mem3_reg[72][26]/P0001  , \wishbone_bd_ram_mem3_reg[72][27]/P0001  , \wishbone_bd_ram_mem3_reg[72][28]/P0001  , \wishbone_bd_ram_mem3_reg[72][29]/P0001  , \wishbone_bd_ram_mem3_reg[72][30]/P0001  , \wishbone_bd_ram_mem3_reg[72][31]/P0001  , \wishbone_bd_ram_mem3_reg[73][24]/P0001  , \wishbone_bd_ram_mem3_reg[73][25]/P0001  , \wishbone_bd_ram_mem3_reg[73][26]/P0001  , \wishbone_bd_ram_mem3_reg[73][27]/P0001  , \wishbone_bd_ram_mem3_reg[73][28]/P0001  , \wishbone_bd_ram_mem3_reg[73][29]/P0001  , \wishbone_bd_ram_mem3_reg[73][30]/P0001  , \wishbone_bd_ram_mem3_reg[73][31]/P0001  , \wishbone_bd_ram_mem3_reg[74][24]/P0001  , \wishbone_bd_ram_mem3_reg[74][25]/P0001  , \wishbone_bd_ram_mem3_reg[74][26]/P0001  , \wishbone_bd_ram_mem3_reg[74][27]/P0001  , \wishbone_bd_ram_mem3_reg[74][28]/P0001  , \wishbone_bd_ram_mem3_reg[74][29]/P0001  , \wishbone_bd_ram_mem3_reg[74][30]/P0001  , \wishbone_bd_ram_mem3_reg[74][31]/P0001  , \wishbone_bd_ram_mem3_reg[75][24]/P0001  , \wishbone_bd_ram_mem3_reg[75][25]/P0001  , \wishbone_bd_ram_mem3_reg[75][26]/P0001  , \wishbone_bd_ram_mem3_reg[75][27]/P0001  , \wishbone_bd_ram_mem3_reg[75][28]/P0001  , \wishbone_bd_ram_mem3_reg[75][29]/P0001  , \wishbone_bd_ram_mem3_reg[75][30]/P0001  , \wishbone_bd_ram_mem3_reg[75][31]/P0001  , \wishbone_bd_ram_mem3_reg[76][24]/P0001  , \wishbone_bd_ram_mem3_reg[76][25]/P0001  , \wishbone_bd_ram_mem3_reg[76][26]/P0001  , \wishbone_bd_ram_mem3_reg[76][27]/P0001  , \wishbone_bd_ram_mem3_reg[76][28]/P0001  , \wishbone_bd_ram_mem3_reg[76][29]/P0001  , \wishbone_bd_ram_mem3_reg[76][30]/P0001  , \wishbone_bd_ram_mem3_reg[76][31]/P0001  , \wishbone_bd_ram_mem3_reg[77][24]/P0001  , \wishbone_bd_ram_mem3_reg[77][25]/P0001  , \wishbone_bd_ram_mem3_reg[77][26]/P0001  , \wishbone_bd_ram_mem3_reg[77][27]/P0001  , \wishbone_bd_ram_mem3_reg[77][28]/P0001  , \wishbone_bd_ram_mem3_reg[77][29]/P0001  , \wishbone_bd_ram_mem3_reg[77][30]/P0001  , \wishbone_bd_ram_mem3_reg[77][31]/P0001  , \wishbone_bd_ram_mem3_reg[78][24]/P0001  , \wishbone_bd_ram_mem3_reg[78][25]/P0001  , \wishbone_bd_ram_mem3_reg[78][26]/P0001  , \wishbone_bd_ram_mem3_reg[78][27]/P0001  , \wishbone_bd_ram_mem3_reg[78][28]/P0001  , \wishbone_bd_ram_mem3_reg[78][29]/P0001  , \wishbone_bd_ram_mem3_reg[78][30]/P0001  , \wishbone_bd_ram_mem3_reg[78][31]/P0001  , \wishbone_bd_ram_mem3_reg[79][24]/P0001  , \wishbone_bd_ram_mem3_reg[79][25]/P0001  , \wishbone_bd_ram_mem3_reg[79][26]/P0001  , \wishbone_bd_ram_mem3_reg[79][27]/P0001  , \wishbone_bd_ram_mem3_reg[79][28]/P0001  , \wishbone_bd_ram_mem3_reg[79][29]/P0001  , \wishbone_bd_ram_mem3_reg[79][30]/P0001  , \wishbone_bd_ram_mem3_reg[79][31]/P0001  , \wishbone_bd_ram_mem3_reg[7][24]/P0001  , \wishbone_bd_ram_mem3_reg[7][25]/P0001  , \wishbone_bd_ram_mem3_reg[7][26]/P0001  , \wishbone_bd_ram_mem3_reg[7][27]/P0001  , \wishbone_bd_ram_mem3_reg[7][28]/P0001  , \wishbone_bd_ram_mem3_reg[7][29]/P0001  , \wishbone_bd_ram_mem3_reg[7][30]/P0001  , \wishbone_bd_ram_mem3_reg[7][31]/P0001  , \wishbone_bd_ram_mem3_reg[80][24]/P0001  , \wishbone_bd_ram_mem3_reg[80][25]/P0001  , \wishbone_bd_ram_mem3_reg[80][26]/P0001  , \wishbone_bd_ram_mem3_reg[80][27]/P0001  , \wishbone_bd_ram_mem3_reg[80][28]/P0001  , \wishbone_bd_ram_mem3_reg[80][29]/P0001  , \wishbone_bd_ram_mem3_reg[80][30]/P0001  , \wishbone_bd_ram_mem3_reg[80][31]/P0001  , \wishbone_bd_ram_mem3_reg[81][24]/P0001  , \wishbone_bd_ram_mem3_reg[81][25]/P0001  , \wishbone_bd_ram_mem3_reg[81][26]/P0001  , \wishbone_bd_ram_mem3_reg[81][27]/P0001  , \wishbone_bd_ram_mem3_reg[81][28]/P0001  , \wishbone_bd_ram_mem3_reg[81][29]/P0001  , \wishbone_bd_ram_mem3_reg[81][30]/P0001  , \wishbone_bd_ram_mem3_reg[81][31]/P0001  , \wishbone_bd_ram_mem3_reg[82][24]/P0001  , \wishbone_bd_ram_mem3_reg[82][25]/P0001  , \wishbone_bd_ram_mem3_reg[82][26]/P0001  , \wishbone_bd_ram_mem3_reg[82][27]/P0001  , \wishbone_bd_ram_mem3_reg[82][28]/P0001  , \wishbone_bd_ram_mem3_reg[82][29]/P0001  , \wishbone_bd_ram_mem3_reg[82][30]/P0001  , \wishbone_bd_ram_mem3_reg[82][31]/P0001  , \wishbone_bd_ram_mem3_reg[83][24]/P0001  , \wishbone_bd_ram_mem3_reg[83][25]/P0001  , \wishbone_bd_ram_mem3_reg[83][26]/P0001  , \wishbone_bd_ram_mem3_reg[83][27]/P0001  , \wishbone_bd_ram_mem3_reg[83][28]/P0001  , \wishbone_bd_ram_mem3_reg[83][29]/P0001  , \wishbone_bd_ram_mem3_reg[83][30]/P0001  , \wishbone_bd_ram_mem3_reg[83][31]/P0001  , \wishbone_bd_ram_mem3_reg[84][24]/P0001  , \wishbone_bd_ram_mem3_reg[84][25]/P0001  , \wishbone_bd_ram_mem3_reg[84][26]/P0001  , \wishbone_bd_ram_mem3_reg[84][27]/P0001  , \wishbone_bd_ram_mem3_reg[84][28]/P0001  , \wishbone_bd_ram_mem3_reg[84][29]/P0001  , \wishbone_bd_ram_mem3_reg[84][30]/P0001  , \wishbone_bd_ram_mem3_reg[84][31]/P0001  , \wishbone_bd_ram_mem3_reg[85][24]/P0001  , \wishbone_bd_ram_mem3_reg[85][25]/P0001  , \wishbone_bd_ram_mem3_reg[85][26]/P0001  , \wishbone_bd_ram_mem3_reg[85][27]/P0001  , \wishbone_bd_ram_mem3_reg[85][28]/P0001  , \wishbone_bd_ram_mem3_reg[85][29]/P0001  , \wishbone_bd_ram_mem3_reg[85][30]/P0001  , \wishbone_bd_ram_mem3_reg[85][31]/P0001  , \wishbone_bd_ram_mem3_reg[86][24]/P0001  , \wishbone_bd_ram_mem3_reg[86][25]/P0001  , \wishbone_bd_ram_mem3_reg[86][26]/P0001  , \wishbone_bd_ram_mem3_reg[86][27]/P0001  , \wishbone_bd_ram_mem3_reg[86][28]/P0001  , \wishbone_bd_ram_mem3_reg[86][29]/P0001  , \wishbone_bd_ram_mem3_reg[86][30]/P0001  , \wishbone_bd_ram_mem3_reg[86][31]/P0001  , \wishbone_bd_ram_mem3_reg[87][24]/P0001  , \wishbone_bd_ram_mem3_reg[87][25]/P0001  , \wishbone_bd_ram_mem3_reg[87][26]/P0001  , \wishbone_bd_ram_mem3_reg[87][27]/P0001  , \wishbone_bd_ram_mem3_reg[87][28]/P0001  , \wishbone_bd_ram_mem3_reg[87][29]/P0001  , \wishbone_bd_ram_mem3_reg[87][30]/P0001  , \wishbone_bd_ram_mem3_reg[87][31]/P0001  , \wishbone_bd_ram_mem3_reg[88][24]/P0001  , \wishbone_bd_ram_mem3_reg[88][25]/P0001  , \wishbone_bd_ram_mem3_reg[88][26]/P0001  , \wishbone_bd_ram_mem3_reg[88][27]/P0001  , \wishbone_bd_ram_mem3_reg[88][28]/P0001  , \wishbone_bd_ram_mem3_reg[88][29]/P0001  , \wishbone_bd_ram_mem3_reg[88][30]/P0001  , \wishbone_bd_ram_mem3_reg[88][31]/P0001  , \wishbone_bd_ram_mem3_reg[89][24]/P0001  , \wishbone_bd_ram_mem3_reg[89][25]/P0001  , \wishbone_bd_ram_mem3_reg[89][26]/P0001  , \wishbone_bd_ram_mem3_reg[89][27]/P0001  , \wishbone_bd_ram_mem3_reg[89][28]/P0001  , \wishbone_bd_ram_mem3_reg[89][29]/P0001  , \wishbone_bd_ram_mem3_reg[89][30]/P0001  , \wishbone_bd_ram_mem3_reg[89][31]/P0001  , \wishbone_bd_ram_mem3_reg[8][24]/P0001  , \wishbone_bd_ram_mem3_reg[8][25]/P0001  , \wishbone_bd_ram_mem3_reg[8][26]/P0001  , \wishbone_bd_ram_mem3_reg[8][27]/P0001  , \wishbone_bd_ram_mem3_reg[8][28]/P0001  , \wishbone_bd_ram_mem3_reg[8][29]/P0001  , \wishbone_bd_ram_mem3_reg[8][30]/P0001  , \wishbone_bd_ram_mem3_reg[8][31]/P0001  , \wishbone_bd_ram_mem3_reg[90][24]/P0001  , \wishbone_bd_ram_mem3_reg[90][25]/P0001  , \wishbone_bd_ram_mem3_reg[90][26]/P0001  , \wishbone_bd_ram_mem3_reg[90][27]/P0001  , \wishbone_bd_ram_mem3_reg[90][28]/P0001  , \wishbone_bd_ram_mem3_reg[90][29]/P0001  , \wishbone_bd_ram_mem3_reg[90][30]/P0001  , \wishbone_bd_ram_mem3_reg[90][31]/P0001  , \wishbone_bd_ram_mem3_reg[91][24]/P0001  , \wishbone_bd_ram_mem3_reg[91][25]/P0001  , \wishbone_bd_ram_mem3_reg[91][26]/P0001  , \wishbone_bd_ram_mem3_reg[91][27]/P0001  , \wishbone_bd_ram_mem3_reg[91][28]/P0001  , \wishbone_bd_ram_mem3_reg[91][29]/P0001  , \wishbone_bd_ram_mem3_reg[91][30]/P0001  , \wishbone_bd_ram_mem3_reg[91][31]/P0001  , \wishbone_bd_ram_mem3_reg[92][24]/P0001  , \wishbone_bd_ram_mem3_reg[92][25]/P0001  , \wishbone_bd_ram_mem3_reg[92][26]/P0001  , \wishbone_bd_ram_mem3_reg[92][27]/P0001  , \wishbone_bd_ram_mem3_reg[92][28]/P0001  , \wishbone_bd_ram_mem3_reg[92][29]/P0001  , \wishbone_bd_ram_mem3_reg[92][30]/P0001  , \wishbone_bd_ram_mem3_reg[92][31]/P0001  , \wishbone_bd_ram_mem3_reg[93][24]/P0001  , \wishbone_bd_ram_mem3_reg[93][25]/P0001  , \wishbone_bd_ram_mem3_reg[93][26]/P0001  , \wishbone_bd_ram_mem3_reg[93][27]/P0001  , \wishbone_bd_ram_mem3_reg[93][28]/P0001  , \wishbone_bd_ram_mem3_reg[93][29]/P0001  , \wishbone_bd_ram_mem3_reg[93][30]/P0001  , \wishbone_bd_ram_mem3_reg[93][31]/P0001  , \wishbone_bd_ram_mem3_reg[94][24]/P0001  , \wishbone_bd_ram_mem3_reg[94][25]/P0001  , \wishbone_bd_ram_mem3_reg[94][26]/P0001  , \wishbone_bd_ram_mem3_reg[94][27]/P0001  , \wishbone_bd_ram_mem3_reg[94][28]/P0001  , \wishbone_bd_ram_mem3_reg[94][29]/P0001  , \wishbone_bd_ram_mem3_reg[94][30]/P0001  , \wishbone_bd_ram_mem3_reg[94][31]/P0001  , \wishbone_bd_ram_mem3_reg[95][24]/P0001  , \wishbone_bd_ram_mem3_reg[95][25]/P0001  , \wishbone_bd_ram_mem3_reg[95][26]/P0001  , \wishbone_bd_ram_mem3_reg[95][27]/P0001  , \wishbone_bd_ram_mem3_reg[95][28]/P0001  , \wishbone_bd_ram_mem3_reg[95][29]/P0001  , \wishbone_bd_ram_mem3_reg[95][30]/P0001  , \wishbone_bd_ram_mem3_reg[95][31]/P0001  , \wishbone_bd_ram_mem3_reg[96][24]/P0001  , \wishbone_bd_ram_mem3_reg[96][25]/P0001  , \wishbone_bd_ram_mem3_reg[96][26]/P0001  , \wishbone_bd_ram_mem3_reg[96][27]/P0001  , \wishbone_bd_ram_mem3_reg[96][28]/P0001  , \wishbone_bd_ram_mem3_reg[96][29]/P0001  , \wishbone_bd_ram_mem3_reg[96][30]/P0001  , \wishbone_bd_ram_mem3_reg[96][31]/P0001  , \wishbone_bd_ram_mem3_reg[97][24]/P0001  , \wishbone_bd_ram_mem3_reg[97][25]/P0001  , \wishbone_bd_ram_mem3_reg[97][26]/P0001  , \wishbone_bd_ram_mem3_reg[97][27]/P0001  , \wishbone_bd_ram_mem3_reg[97][28]/P0001  , \wishbone_bd_ram_mem3_reg[97][29]/P0001  , \wishbone_bd_ram_mem3_reg[97][30]/P0001  , \wishbone_bd_ram_mem3_reg[97][31]/P0001  , \wishbone_bd_ram_mem3_reg[98][24]/P0001  , \wishbone_bd_ram_mem3_reg[98][25]/P0001  , \wishbone_bd_ram_mem3_reg[98][26]/P0001  , \wishbone_bd_ram_mem3_reg[98][27]/P0001  , \wishbone_bd_ram_mem3_reg[98][28]/P0001  , \wishbone_bd_ram_mem3_reg[98][29]/P0001  , \wishbone_bd_ram_mem3_reg[98][30]/P0001  , \wishbone_bd_ram_mem3_reg[98][31]/P0001  , \wishbone_bd_ram_mem3_reg[99][24]/P0001  , \wishbone_bd_ram_mem3_reg[99][25]/P0001  , \wishbone_bd_ram_mem3_reg[99][26]/P0001  , \wishbone_bd_ram_mem3_reg[99][27]/P0001  , \wishbone_bd_ram_mem3_reg[99][28]/P0001  , \wishbone_bd_ram_mem3_reg[99][29]/P0001  , \wishbone_bd_ram_mem3_reg[99][30]/P0001  , \wishbone_bd_ram_mem3_reg[99][31]/P0001  , \wishbone_bd_ram_mem3_reg[9][24]/P0001  , \wishbone_bd_ram_mem3_reg[9][25]/P0001  , \wishbone_bd_ram_mem3_reg[9][26]/P0001  , \wishbone_bd_ram_mem3_reg[9][27]/P0001  , \wishbone_bd_ram_mem3_reg[9][28]/P0001  , \wishbone_bd_ram_mem3_reg[9][29]/P0001  , \wishbone_bd_ram_mem3_reg[9][30]/P0001  , \wishbone_bd_ram_mem3_reg[9][31]/P0001  , \wishbone_bd_ram_raddr_reg[0]/P0001  , \wishbone_bd_ram_raddr_reg[1]/NET0131  , \wishbone_bd_ram_raddr_reg[2]/NET0131  , \wishbone_bd_ram_raddr_reg[3]/P0001  , \wishbone_bd_ram_raddr_reg[4]/NET0131  , \wishbone_bd_ram_raddr_reg[5]/NET0131  , \wishbone_bd_ram_raddr_reg[6]/NET0131  , \wishbone_bd_ram_raddr_reg[7]/NET0131  , \wishbone_cyc_cleared_reg/NET0131  , \wishbone_r_RxEn_q_reg/NET0131  , \wishbone_r_TxEn_q_reg/NET0131  , \wishbone_ram_addr_reg[0]/NET0131  , \wishbone_ram_addr_reg[1]/NET0131  , \wishbone_ram_addr_reg[2]/NET0131  , \wishbone_ram_addr_reg[3]/NET0131  , \wishbone_ram_addr_reg[4]/NET0131  , \wishbone_ram_addr_reg[5]/NET0131  , \wishbone_ram_addr_reg[6]/NET0131  , \wishbone_ram_addr_reg[7]/NET0131  , \wishbone_ram_di_reg[0]/NET0131  , \wishbone_ram_di_reg[10]/NET0131  , \wishbone_ram_di_reg[11]/NET0131  , \wishbone_ram_di_reg[12]/NET0131  , \wishbone_ram_di_reg[13]/NET0131  , \wishbone_ram_di_reg[14]/NET0131  , \wishbone_ram_di_reg[15]/NET0131  , \wishbone_ram_di_reg[16]/NET0131  , \wishbone_ram_di_reg[17]/NET0131  , \wishbone_ram_di_reg[18]/NET0131  , \wishbone_ram_di_reg[19]/NET0131  , \wishbone_ram_di_reg[1]/NET0131  , \wishbone_ram_di_reg[20]/NET0131  , \wishbone_ram_di_reg[21]/NET0131  , \wishbone_ram_di_reg[22]/NET0131  , \wishbone_ram_di_reg[23]/NET0131  , \wishbone_ram_di_reg[24]/NET0131  , \wishbone_ram_di_reg[25]/NET0131  , \wishbone_ram_di_reg[26]/NET0131  , \wishbone_ram_di_reg[27]/NET0131  , \wishbone_ram_di_reg[28]/NET0131  , \wishbone_ram_di_reg[29]/NET0131  , \wishbone_ram_di_reg[2]/NET0131  , \wishbone_ram_di_reg[30]/NET0131  , \wishbone_ram_di_reg[31]/NET0131  , \wishbone_ram_di_reg[3]/NET0131  , \wishbone_ram_di_reg[4]/NET0131  , \wishbone_ram_di_reg[5]/NET0131  , \wishbone_ram_di_reg[6]/NET0131  , \wishbone_ram_di_reg[7]/NET0131  , \wishbone_ram_di_reg[8]/NET0131  , \wishbone_ram_di_reg[9]/NET0131  , \wishbone_rx_burst_cnt_reg[0]/NET0131  , \wishbone_rx_burst_cnt_reg[1]/NET0131  , \wishbone_rx_burst_cnt_reg[2]/NET0131  , \wishbone_rx_burst_en_reg/NET0131  , \wishbone_rx_fifo_cnt_reg[0]/NET0131  , \wishbone_rx_fifo_cnt_reg[1]/NET0131  , \wishbone_rx_fifo_cnt_reg[2]/NET0131  , \wishbone_rx_fifo_cnt_reg[3]/NET0131  , \wishbone_rx_fifo_cnt_reg[4]/NET0131  , \wishbone_rx_fifo_fifo_reg[0][0]/P0001  , \wishbone_rx_fifo_fifo_reg[0][10]/P0001  , \wishbone_rx_fifo_fifo_reg[0][11]/P0001  , \wishbone_rx_fifo_fifo_reg[0][12]/P0001  , \wishbone_rx_fifo_fifo_reg[0][13]/P0001  , \wishbone_rx_fifo_fifo_reg[0][14]/P0001  , \wishbone_rx_fifo_fifo_reg[0][15]/P0001  , \wishbone_rx_fifo_fifo_reg[0][16]/P0001  , \wishbone_rx_fifo_fifo_reg[0][17]/P0001  , \wishbone_rx_fifo_fifo_reg[0][18]/P0001  , \wishbone_rx_fifo_fifo_reg[0][19]/P0001  , \wishbone_rx_fifo_fifo_reg[0][1]/P0001  , \wishbone_rx_fifo_fifo_reg[0][20]/P0001  , \wishbone_rx_fifo_fifo_reg[0][21]/P0001  , \wishbone_rx_fifo_fifo_reg[0][22]/P0001  , \wishbone_rx_fifo_fifo_reg[0][23]/P0001  , \wishbone_rx_fifo_fifo_reg[0][24]/P0001  , \wishbone_rx_fifo_fifo_reg[0][25]/P0001  , \wishbone_rx_fifo_fifo_reg[0][26]/P0001  , \wishbone_rx_fifo_fifo_reg[0][27]/P0001  , \wishbone_rx_fifo_fifo_reg[0][28]/P0001  , \wishbone_rx_fifo_fifo_reg[0][29]/P0001  , \wishbone_rx_fifo_fifo_reg[0][2]/P0001  , \wishbone_rx_fifo_fifo_reg[0][30]/P0001  , \wishbone_rx_fifo_fifo_reg[0][31]/P0001  , \wishbone_rx_fifo_fifo_reg[0][3]/P0001  , \wishbone_rx_fifo_fifo_reg[0][4]/P0001  , \wishbone_rx_fifo_fifo_reg[0][5]/P0001  , \wishbone_rx_fifo_fifo_reg[0][6]/P0001  , \wishbone_rx_fifo_fifo_reg[0][7]/P0001  , \wishbone_rx_fifo_fifo_reg[0][8]/P0001  , \wishbone_rx_fifo_fifo_reg[0][9]/P0001  , \wishbone_rx_fifo_fifo_reg[10][0]/P0001  , \wishbone_rx_fifo_fifo_reg[10][10]/P0001  , \wishbone_rx_fifo_fifo_reg[10][11]/P0001  , \wishbone_rx_fifo_fifo_reg[10][12]/P0001  , \wishbone_rx_fifo_fifo_reg[10][13]/P0001  , \wishbone_rx_fifo_fifo_reg[10][14]/P0001  , \wishbone_rx_fifo_fifo_reg[10][15]/P0001  , \wishbone_rx_fifo_fifo_reg[10][16]/P0001  , \wishbone_rx_fifo_fifo_reg[10][17]/P0001  , \wishbone_rx_fifo_fifo_reg[10][18]/P0001  , \wishbone_rx_fifo_fifo_reg[10][19]/P0001  , \wishbone_rx_fifo_fifo_reg[10][1]/P0001  , \wishbone_rx_fifo_fifo_reg[10][20]/P0001  , \wishbone_rx_fifo_fifo_reg[10][21]/P0001  , \wishbone_rx_fifo_fifo_reg[10][22]/P0001  , \wishbone_rx_fifo_fifo_reg[10][23]/P0001  , \wishbone_rx_fifo_fifo_reg[10][24]/P0001  , \wishbone_rx_fifo_fifo_reg[10][25]/P0001  , \wishbone_rx_fifo_fifo_reg[10][26]/P0001  , \wishbone_rx_fifo_fifo_reg[10][27]/P0001  , \wishbone_rx_fifo_fifo_reg[10][28]/P0001  , \wishbone_rx_fifo_fifo_reg[10][29]/P0001  , \wishbone_rx_fifo_fifo_reg[10][2]/P0001  , \wishbone_rx_fifo_fifo_reg[10][30]/P0001  , \wishbone_rx_fifo_fifo_reg[10][31]/P0001  , \wishbone_rx_fifo_fifo_reg[10][3]/P0001  , \wishbone_rx_fifo_fifo_reg[10][4]/P0001  , \wishbone_rx_fifo_fifo_reg[10][5]/P0001  , \wishbone_rx_fifo_fifo_reg[10][6]/P0001  , \wishbone_rx_fifo_fifo_reg[10][7]/P0001  , \wishbone_rx_fifo_fifo_reg[10][8]/P0001  , \wishbone_rx_fifo_fifo_reg[10][9]/P0001  , \wishbone_rx_fifo_fifo_reg[11][0]/P0001  , \wishbone_rx_fifo_fifo_reg[11][10]/P0001  , \wishbone_rx_fifo_fifo_reg[11][11]/P0001  , \wishbone_rx_fifo_fifo_reg[11][12]/P0001  , \wishbone_rx_fifo_fifo_reg[11][13]/P0001  , \wishbone_rx_fifo_fifo_reg[11][14]/P0001  , \wishbone_rx_fifo_fifo_reg[11][15]/P0001  , \wishbone_rx_fifo_fifo_reg[11][16]/P0001  , \wishbone_rx_fifo_fifo_reg[11][17]/P0001  , \wishbone_rx_fifo_fifo_reg[11][18]/P0001  , \wishbone_rx_fifo_fifo_reg[11][19]/P0001  , \wishbone_rx_fifo_fifo_reg[11][1]/P0001  , \wishbone_rx_fifo_fifo_reg[11][20]/P0001  , \wishbone_rx_fifo_fifo_reg[11][21]/P0001  , \wishbone_rx_fifo_fifo_reg[11][22]/P0001  , \wishbone_rx_fifo_fifo_reg[11][23]/P0001  , \wishbone_rx_fifo_fifo_reg[11][24]/P0001  , \wishbone_rx_fifo_fifo_reg[11][25]/P0001  , \wishbone_rx_fifo_fifo_reg[11][26]/P0001  , \wishbone_rx_fifo_fifo_reg[11][27]/P0001  , \wishbone_rx_fifo_fifo_reg[11][28]/P0001  , \wishbone_rx_fifo_fifo_reg[11][29]/P0001  , \wishbone_rx_fifo_fifo_reg[11][2]/P0001  , \wishbone_rx_fifo_fifo_reg[11][30]/P0001  , \wishbone_rx_fifo_fifo_reg[11][31]/P0001  , \wishbone_rx_fifo_fifo_reg[11][3]/P0001  , \wishbone_rx_fifo_fifo_reg[11][4]/P0001  , \wishbone_rx_fifo_fifo_reg[11][5]/P0001  , \wishbone_rx_fifo_fifo_reg[11][6]/P0001  , \wishbone_rx_fifo_fifo_reg[11][7]/P0001  , \wishbone_rx_fifo_fifo_reg[11][8]/P0001  , \wishbone_rx_fifo_fifo_reg[11][9]/P0001  , \wishbone_rx_fifo_fifo_reg[12][0]/P0001  , \wishbone_rx_fifo_fifo_reg[12][10]/P0001  , \wishbone_rx_fifo_fifo_reg[12][11]/P0001  , \wishbone_rx_fifo_fifo_reg[12][12]/P0001  , \wishbone_rx_fifo_fifo_reg[12][13]/P0001  , \wishbone_rx_fifo_fifo_reg[12][14]/P0001  , \wishbone_rx_fifo_fifo_reg[12][15]/P0001  , \wishbone_rx_fifo_fifo_reg[12][16]/P0001  , \wishbone_rx_fifo_fifo_reg[12][17]/P0001  , \wishbone_rx_fifo_fifo_reg[12][18]/P0001  , \wishbone_rx_fifo_fifo_reg[12][19]/P0001  , \wishbone_rx_fifo_fifo_reg[12][1]/P0001  , \wishbone_rx_fifo_fifo_reg[12][20]/P0001  , \wishbone_rx_fifo_fifo_reg[12][21]/P0001  , \wishbone_rx_fifo_fifo_reg[12][22]/P0001  , \wishbone_rx_fifo_fifo_reg[12][23]/P0001  , \wishbone_rx_fifo_fifo_reg[12][24]/P0001  , \wishbone_rx_fifo_fifo_reg[12][25]/P0001  , \wishbone_rx_fifo_fifo_reg[12][26]/P0001  , \wishbone_rx_fifo_fifo_reg[12][27]/P0001  , \wishbone_rx_fifo_fifo_reg[12][28]/P0001  , \wishbone_rx_fifo_fifo_reg[12][29]/P0001  , \wishbone_rx_fifo_fifo_reg[12][2]/P0001  , \wishbone_rx_fifo_fifo_reg[12][30]/P0001  , \wishbone_rx_fifo_fifo_reg[12][31]/P0001  , \wishbone_rx_fifo_fifo_reg[12][3]/P0001  , \wishbone_rx_fifo_fifo_reg[12][4]/P0001  , \wishbone_rx_fifo_fifo_reg[12][5]/P0001  , \wishbone_rx_fifo_fifo_reg[12][6]/P0001  , \wishbone_rx_fifo_fifo_reg[12][7]/P0001  , \wishbone_rx_fifo_fifo_reg[12][8]/P0001  , \wishbone_rx_fifo_fifo_reg[12][9]/P0001  , \wishbone_rx_fifo_fifo_reg[13][0]/P0001  , \wishbone_rx_fifo_fifo_reg[13][10]/P0001  , \wishbone_rx_fifo_fifo_reg[13][11]/P0001  , \wishbone_rx_fifo_fifo_reg[13][12]/P0001  , \wishbone_rx_fifo_fifo_reg[13][13]/P0001  , \wishbone_rx_fifo_fifo_reg[13][14]/P0001  , \wishbone_rx_fifo_fifo_reg[13][15]/P0001  , \wishbone_rx_fifo_fifo_reg[13][16]/P0001  , \wishbone_rx_fifo_fifo_reg[13][17]/P0001  , \wishbone_rx_fifo_fifo_reg[13][18]/P0001  , \wishbone_rx_fifo_fifo_reg[13][19]/P0001  , \wishbone_rx_fifo_fifo_reg[13][1]/P0001  , \wishbone_rx_fifo_fifo_reg[13][20]/P0001  , \wishbone_rx_fifo_fifo_reg[13][21]/P0001  , \wishbone_rx_fifo_fifo_reg[13][22]/P0001  , \wishbone_rx_fifo_fifo_reg[13][23]/P0001  , \wishbone_rx_fifo_fifo_reg[13][24]/P0001  , \wishbone_rx_fifo_fifo_reg[13][25]/P0001  , \wishbone_rx_fifo_fifo_reg[13][26]/P0001  , \wishbone_rx_fifo_fifo_reg[13][27]/P0001  , \wishbone_rx_fifo_fifo_reg[13][28]/P0001  , \wishbone_rx_fifo_fifo_reg[13][29]/P0001  , \wishbone_rx_fifo_fifo_reg[13][2]/P0001  , \wishbone_rx_fifo_fifo_reg[13][30]/P0001  , \wishbone_rx_fifo_fifo_reg[13][31]/P0001  , \wishbone_rx_fifo_fifo_reg[13][3]/P0001  , \wishbone_rx_fifo_fifo_reg[13][4]/P0001  , \wishbone_rx_fifo_fifo_reg[13][5]/P0001  , \wishbone_rx_fifo_fifo_reg[13][6]/P0001  , \wishbone_rx_fifo_fifo_reg[13][7]/P0001  , \wishbone_rx_fifo_fifo_reg[13][8]/P0001  , \wishbone_rx_fifo_fifo_reg[13][9]/P0001  , \wishbone_rx_fifo_fifo_reg[14][0]/P0001  , \wishbone_rx_fifo_fifo_reg[14][10]/P0001  , \wishbone_rx_fifo_fifo_reg[14][11]/P0001  , \wishbone_rx_fifo_fifo_reg[14][12]/P0001  , \wishbone_rx_fifo_fifo_reg[14][13]/P0001  , \wishbone_rx_fifo_fifo_reg[14][14]/P0001  , \wishbone_rx_fifo_fifo_reg[14][15]/P0001  , \wishbone_rx_fifo_fifo_reg[14][16]/P0001  , \wishbone_rx_fifo_fifo_reg[14][17]/P0001  , \wishbone_rx_fifo_fifo_reg[14][18]/P0001  , \wishbone_rx_fifo_fifo_reg[14][19]/P0001  , \wishbone_rx_fifo_fifo_reg[14][1]/P0001  , \wishbone_rx_fifo_fifo_reg[14][20]/P0001  , \wishbone_rx_fifo_fifo_reg[14][21]/P0001  , \wishbone_rx_fifo_fifo_reg[14][22]/P0001  , \wishbone_rx_fifo_fifo_reg[14][23]/P0001  , \wishbone_rx_fifo_fifo_reg[14][24]/P0001  , \wishbone_rx_fifo_fifo_reg[14][25]/P0001  , \wishbone_rx_fifo_fifo_reg[14][26]/P0001  , \wishbone_rx_fifo_fifo_reg[14][27]/P0001  , \wishbone_rx_fifo_fifo_reg[14][28]/P0001  , \wishbone_rx_fifo_fifo_reg[14][29]/P0001  , \wishbone_rx_fifo_fifo_reg[14][2]/P0001  , \wishbone_rx_fifo_fifo_reg[14][30]/P0001  , \wishbone_rx_fifo_fifo_reg[14][31]/P0001  , \wishbone_rx_fifo_fifo_reg[14][3]/P0001  , \wishbone_rx_fifo_fifo_reg[14][4]/P0001  , \wishbone_rx_fifo_fifo_reg[14][5]/P0001  , \wishbone_rx_fifo_fifo_reg[14][6]/P0001  , \wishbone_rx_fifo_fifo_reg[14][7]/P0001  , \wishbone_rx_fifo_fifo_reg[14][8]/P0001  , \wishbone_rx_fifo_fifo_reg[14][9]/P0001  , \wishbone_rx_fifo_fifo_reg[15][0]/P0001  , \wishbone_rx_fifo_fifo_reg[15][10]/P0001  , \wishbone_rx_fifo_fifo_reg[15][11]/P0001  , \wishbone_rx_fifo_fifo_reg[15][12]/P0001  , \wishbone_rx_fifo_fifo_reg[15][13]/P0001  , \wishbone_rx_fifo_fifo_reg[15][14]/P0001  , \wishbone_rx_fifo_fifo_reg[15][15]/P0001  , \wishbone_rx_fifo_fifo_reg[15][16]/P0001  , \wishbone_rx_fifo_fifo_reg[15][17]/P0001  , \wishbone_rx_fifo_fifo_reg[15][18]/P0001  , \wishbone_rx_fifo_fifo_reg[15][19]/P0001  , \wishbone_rx_fifo_fifo_reg[15][1]/P0001  , \wishbone_rx_fifo_fifo_reg[15][20]/P0001  , \wishbone_rx_fifo_fifo_reg[15][21]/P0001  , \wishbone_rx_fifo_fifo_reg[15][22]/P0001  , \wishbone_rx_fifo_fifo_reg[15][23]/P0001  , \wishbone_rx_fifo_fifo_reg[15][24]/P0001  , \wishbone_rx_fifo_fifo_reg[15][25]/P0001  , \wishbone_rx_fifo_fifo_reg[15][26]/P0001  , \wishbone_rx_fifo_fifo_reg[15][27]/P0001  , \wishbone_rx_fifo_fifo_reg[15][28]/P0001  , \wishbone_rx_fifo_fifo_reg[15][29]/P0001  , \wishbone_rx_fifo_fifo_reg[15][2]/P0001  , \wishbone_rx_fifo_fifo_reg[15][30]/P0001  , \wishbone_rx_fifo_fifo_reg[15][31]/P0001  , \wishbone_rx_fifo_fifo_reg[15][3]/P0001  , \wishbone_rx_fifo_fifo_reg[15][4]/P0001  , \wishbone_rx_fifo_fifo_reg[15][5]/P0001  , \wishbone_rx_fifo_fifo_reg[15][6]/P0001  , \wishbone_rx_fifo_fifo_reg[15][7]/P0001  , \wishbone_rx_fifo_fifo_reg[15][8]/P0001  , \wishbone_rx_fifo_fifo_reg[15][9]/P0001  , \wishbone_rx_fifo_fifo_reg[1][0]/P0001  , \wishbone_rx_fifo_fifo_reg[1][10]/P0001  , \wishbone_rx_fifo_fifo_reg[1][11]/P0001  , \wishbone_rx_fifo_fifo_reg[1][12]/P0001  , \wishbone_rx_fifo_fifo_reg[1][13]/P0001  , \wishbone_rx_fifo_fifo_reg[1][14]/P0001  , \wishbone_rx_fifo_fifo_reg[1][15]/P0001  , \wishbone_rx_fifo_fifo_reg[1][16]/P0001  , \wishbone_rx_fifo_fifo_reg[1][17]/P0001  , \wishbone_rx_fifo_fifo_reg[1][18]/P0001  , \wishbone_rx_fifo_fifo_reg[1][19]/P0001  , \wishbone_rx_fifo_fifo_reg[1][1]/P0001  , \wishbone_rx_fifo_fifo_reg[1][20]/P0001  , \wishbone_rx_fifo_fifo_reg[1][21]/P0001  , \wishbone_rx_fifo_fifo_reg[1][22]/P0001  , \wishbone_rx_fifo_fifo_reg[1][23]/P0001  , \wishbone_rx_fifo_fifo_reg[1][24]/P0001  , \wishbone_rx_fifo_fifo_reg[1][25]/P0001  , \wishbone_rx_fifo_fifo_reg[1][26]/P0001  , \wishbone_rx_fifo_fifo_reg[1][27]/P0001  , \wishbone_rx_fifo_fifo_reg[1][28]/P0001  , \wishbone_rx_fifo_fifo_reg[1][29]/P0001  , \wishbone_rx_fifo_fifo_reg[1][2]/P0001  , \wishbone_rx_fifo_fifo_reg[1][30]/P0001  , \wishbone_rx_fifo_fifo_reg[1][31]/P0001  , \wishbone_rx_fifo_fifo_reg[1][3]/P0001  , \wishbone_rx_fifo_fifo_reg[1][4]/P0001  , \wishbone_rx_fifo_fifo_reg[1][5]/P0001  , \wishbone_rx_fifo_fifo_reg[1][6]/P0001  , \wishbone_rx_fifo_fifo_reg[1][7]/P0001  , \wishbone_rx_fifo_fifo_reg[1][8]/P0001  , \wishbone_rx_fifo_fifo_reg[1][9]/P0001  , \wishbone_rx_fifo_fifo_reg[2][0]/P0001  , \wishbone_rx_fifo_fifo_reg[2][10]/P0001  , \wishbone_rx_fifo_fifo_reg[2][11]/P0001  , \wishbone_rx_fifo_fifo_reg[2][12]/P0001  , \wishbone_rx_fifo_fifo_reg[2][13]/P0001  , \wishbone_rx_fifo_fifo_reg[2][14]/P0001  , \wishbone_rx_fifo_fifo_reg[2][15]/P0001  , \wishbone_rx_fifo_fifo_reg[2][16]/P0001  , \wishbone_rx_fifo_fifo_reg[2][17]/P0001  , \wishbone_rx_fifo_fifo_reg[2][18]/P0001  , \wishbone_rx_fifo_fifo_reg[2][19]/P0001  , \wishbone_rx_fifo_fifo_reg[2][1]/P0001  , \wishbone_rx_fifo_fifo_reg[2][20]/P0001  , \wishbone_rx_fifo_fifo_reg[2][21]/P0001  , \wishbone_rx_fifo_fifo_reg[2][22]/P0001  , \wishbone_rx_fifo_fifo_reg[2][23]/P0001  , \wishbone_rx_fifo_fifo_reg[2][24]/P0001  , \wishbone_rx_fifo_fifo_reg[2][25]/P0001  , \wishbone_rx_fifo_fifo_reg[2][26]/P0001  , \wishbone_rx_fifo_fifo_reg[2][27]/P0001  , \wishbone_rx_fifo_fifo_reg[2][28]/P0001  , \wishbone_rx_fifo_fifo_reg[2][29]/P0001  , \wishbone_rx_fifo_fifo_reg[2][2]/P0001  , \wishbone_rx_fifo_fifo_reg[2][30]/P0001  , \wishbone_rx_fifo_fifo_reg[2][31]/P0001  , \wishbone_rx_fifo_fifo_reg[2][3]/P0001  , \wishbone_rx_fifo_fifo_reg[2][4]/P0001  , \wishbone_rx_fifo_fifo_reg[2][5]/P0001  , \wishbone_rx_fifo_fifo_reg[2][6]/P0001  , \wishbone_rx_fifo_fifo_reg[2][7]/P0001  , \wishbone_rx_fifo_fifo_reg[2][8]/P0001  , \wishbone_rx_fifo_fifo_reg[2][9]/P0001  , \wishbone_rx_fifo_fifo_reg[3][0]/P0001  , \wishbone_rx_fifo_fifo_reg[3][10]/P0001  , \wishbone_rx_fifo_fifo_reg[3][11]/P0001  , \wishbone_rx_fifo_fifo_reg[3][12]/P0001  , \wishbone_rx_fifo_fifo_reg[3][13]/P0001  , \wishbone_rx_fifo_fifo_reg[3][14]/P0001  , \wishbone_rx_fifo_fifo_reg[3][15]/P0001  , \wishbone_rx_fifo_fifo_reg[3][16]/P0001  , \wishbone_rx_fifo_fifo_reg[3][17]/P0001  , \wishbone_rx_fifo_fifo_reg[3][18]/P0001  , \wishbone_rx_fifo_fifo_reg[3][19]/P0001  , \wishbone_rx_fifo_fifo_reg[3][1]/P0001  , \wishbone_rx_fifo_fifo_reg[3][20]/P0001  , \wishbone_rx_fifo_fifo_reg[3][21]/P0001  , \wishbone_rx_fifo_fifo_reg[3][22]/P0001  , \wishbone_rx_fifo_fifo_reg[3][23]/P0001  , \wishbone_rx_fifo_fifo_reg[3][24]/P0001  , \wishbone_rx_fifo_fifo_reg[3][25]/P0001  , \wishbone_rx_fifo_fifo_reg[3][26]/P0001  , \wishbone_rx_fifo_fifo_reg[3][27]/P0001  , \wishbone_rx_fifo_fifo_reg[3][28]/P0001  , \wishbone_rx_fifo_fifo_reg[3][29]/P0001  , \wishbone_rx_fifo_fifo_reg[3][2]/P0001  , \wishbone_rx_fifo_fifo_reg[3][30]/P0001  , \wishbone_rx_fifo_fifo_reg[3][31]/P0001  , \wishbone_rx_fifo_fifo_reg[3][3]/P0001  , \wishbone_rx_fifo_fifo_reg[3][4]/P0001  , \wishbone_rx_fifo_fifo_reg[3][5]/P0001  , \wishbone_rx_fifo_fifo_reg[3][6]/P0001  , \wishbone_rx_fifo_fifo_reg[3][7]/P0001  , \wishbone_rx_fifo_fifo_reg[3][8]/P0001  , \wishbone_rx_fifo_fifo_reg[3][9]/P0001  , \wishbone_rx_fifo_fifo_reg[4][0]/P0001  , \wishbone_rx_fifo_fifo_reg[4][10]/P0001  , \wishbone_rx_fifo_fifo_reg[4][11]/P0001  , \wishbone_rx_fifo_fifo_reg[4][12]/P0001  , \wishbone_rx_fifo_fifo_reg[4][13]/P0001  , \wishbone_rx_fifo_fifo_reg[4][14]/P0001  , \wishbone_rx_fifo_fifo_reg[4][15]/P0001  , \wishbone_rx_fifo_fifo_reg[4][16]/P0001  , \wishbone_rx_fifo_fifo_reg[4][17]/P0001  , \wishbone_rx_fifo_fifo_reg[4][18]/P0001  , \wishbone_rx_fifo_fifo_reg[4][19]/P0001  , \wishbone_rx_fifo_fifo_reg[4][1]/P0001  , \wishbone_rx_fifo_fifo_reg[4][20]/P0001  , \wishbone_rx_fifo_fifo_reg[4][21]/P0001  , \wishbone_rx_fifo_fifo_reg[4][22]/P0001  , \wishbone_rx_fifo_fifo_reg[4][23]/P0001  , \wishbone_rx_fifo_fifo_reg[4][24]/P0001  , \wishbone_rx_fifo_fifo_reg[4][25]/P0001  , \wishbone_rx_fifo_fifo_reg[4][26]/P0001  , \wishbone_rx_fifo_fifo_reg[4][27]/P0001  , \wishbone_rx_fifo_fifo_reg[4][28]/P0001  , \wishbone_rx_fifo_fifo_reg[4][29]/P0001  , \wishbone_rx_fifo_fifo_reg[4][2]/P0001  , \wishbone_rx_fifo_fifo_reg[4][30]/P0001  , \wishbone_rx_fifo_fifo_reg[4][31]/P0001  , \wishbone_rx_fifo_fifo_reg[4][3]/P0001  , \wishbone_rx_fifo_fifo_reg[4][4]/P0001  , \wishbone_rx_fifo_fifo_reg[4][5]/P0001  , \wishbone_rx_fifo_fifo_reg[4][6]/P0001  , \wishbone_rx_fifo_fifo_reg[4][7]/P0001  , \wishbone_rx_fifo_fifo_reg[4][8]/P0001  , \wishbone_rx_fifo_fifo_reg[4][9]/P0001  , \wishbone_rx_fifo_fifo_reg[5][0]/P0001  , \wishbone_rx_fifo_fifo_reg[5][10]/P0001  , \wishbone_rx_fifo_fifo_reg[5][11]/P0001  , \wishbone_rx_fifo_fifo_reg[5][12]/P0001  , \wishbone_rx_fifo_fifo_reg[5][13]/P0001  , \wishbone_rx_fifo_fifo_reg[5][14]/P0001  , \wishbone_rx_fifo_fifo_reg[5][15]/P0001  , \wishbone_rx_fifo_fifo_reg[5][16]/P0001  , \wishbone_rx_fifo_fifo_reg[5][17]/P0001  , \wishbone_rx_fifo_fifo_reg[5][18]/P0001  , \wishbone_rx_fifo_fifo_reg[5][19]/P0001  , \wishbone_rx_fifo_fifo_reg[5][1]/P0001  , \wishbone_rx_fifo_fifo_reg[5][20]/P0001  , \wishbone_rx_fifo_fifo_reg[5][21]/P0001  , \wishbone_rx_fifo_fifo_reg[5][22]/P0001  , \wishbone_rx_fifo_fifo_reg[5][23]/P0001  , \wishbone_rx_fifo_fifo_reg[5][24]/P0001  , \wishbone_rx_fifo_fifo_reg[5][25]/P0001  , \wishbone_rx_fifo_fifo_reg[5][26]/P0001  , \wishbone_rx_fifo_fifo_reg[5][27]/P0001  , \wishbone_rx_fifo_fifo_reg[5][28]/P0001  , \wishbone_rx_fifo_fifo_reg[5][29]/P0001  , \wishbone_rx_fifo_fifo_reg[5][2]/P0001  , \wishbone_rx_fifo_fifo_reg[5][30]/P0001  , \wishbone_rx_fifo_fifo_reg[5][31]/P0001  , \wishbone_rx_fifo_fifo_reg[5][3]/P0001  , \wishbone_rx_fifo_fifo_reg[5][4]/P0001  , \wishbone_rx_fifo_fifo_reg[5][5]/P0001  , \wishbone_rx_fifo_fifo_reg[5][6]/P0001  , \wishbone_rx_fifo_fifo_reg[5][7]/P0001  , \wishbone_rx_fifo_fifo_reg[5][8]/P0001  , \wishbone_rx_fifo_fifo_reg[5][9]/P0001  , \wishbone_rx_fifo_fifo_reg[6][0]/P0001  , \wishbone_rx_fifo_fifo_reg[6][10]/P0001  , \wishbone_rx_fifo_fifo_reg[6][11]/P0001  , \wishbone_rx_fifo_fifo_reg[6][12]/P0001  , \wishbone_rx_fifo_fifo_reg[6][13]/P0001  , \wishbone_rx_fifo_fifo_reg[6][14]/P0001  , \wishbone_rx_fifo_fifo_reg[6][15]/P0001  , \wishbone_rx_fifo_fifo_reg[6][16]/P0001  , \wishbone_rx_fifo_fifo_reg[6][17]/P0001  , \wishbone_rx_fifo_fifo_reg[6][18]/P0001  , \wishbone_rx_fifo_fifo_reg[6][19]/P0001  , \wishbone_rx_fifo_fifo_reg[6][1]/P0001  , \wishbone_rx_fifo_fifo_reg[6][20]/P0001  , \wishbone_rx_fifo_fifo_reg[6][21]/P0001  , \wishbone_rx_fifo_fifo_reg[6][22]/P0001  , \wishbone_rx_fifo_fifo_reg[6][23]/P0001  , \wishbone_rx_fifo_fifo_reg[6][24]/P0001  , \wishbone_rx_fifo_fifo_reg[6][25]/P0001  , \wishbone_rx_fifo_fifo_reg[6][26]/P0001  , \wishbone_rx_fifo_fifo_reg[6][27]/P0001  , \wishbone_rx_fifo_fifo_reg[6][28]/P0001  , \wishbone_rx_fifo_fifo_reg[6][29]/P0001  , \wishbone_rx_fifo_fifo_reg[6][2]/P0001  , \wishbone_rx_fifo_fifo_reg[6][30]/P0001  , \wishbone_rx_fifo_fifo_reg[6][31]/P0001  , \wishbone_rx_fifo_fifo_reg[6][3]/P0001  , \wishbone_rx_fifo_fifo_reg[6][4]/P0001  , \wishbone_rx_fifo_fifo_reg[6][5]/P0001  , \wishbone_rx_fifo_fifo_reg[6][6]/P0001  , \wishbone_rx_fifo_fifo_reg[6][7]/P0001  , \wishbone_rx_fifo_fifo_reg[6][8]/P0001  , \wishbone_rx_fifo_fifo_reg[6][9]/P0001  , \wishbone_rx_fifo_fifo_reg[7][0]/P0001  , \wishbone_rx_fifo_fifo_reg[7][10]/P0001  , \wishbone_rx_fifo_fifo_reg[7][11]/P0001  , \wishbone_rx_fifo_fifo_reg[7][12]/P0001  , \wishbone_rx_fifo_fifo_reg[7][13]/P0001  , \wishbone_rx_fifo_fifo_reg[7][14]/P0001  , \wishbone_rx_fifo_fifo_reg[7][15]/P0001  , \wishbone_rx_fifo_fifo_reg[7][16]/P0001  , \wishbone_rx_fifo_fifo_reg[7][17]/P0001  , \wishbone_rx_fifo_fifo_reg[7][18]/P0001  , \wishbone_rx_fifo_fifo_reg[7][19]/P0001  , \wishbone_rx_fifo_fifo_reg[7][1]/P0001  , \wishbone_rx_fifo_fifo_reg[7][20]/P0001  , \wishbone_rx_fifo_fifo_reg[7][21]/P0001  , \wishbone_rx_fifo_fifo_reg[7][22]/P0001  , \wishbone_rx_fifo_fifo_reg[7][23]/P0001  , \wishbone_rx_fifo_fifo_reg[7][24]/P0001  , \wishbone_rx_fifo_fifo_reg[7][25]/P0001  , \wishbone_rx_fifo_fifo_reg[7][26]/P0001  , \wishbone_rx_fifo_fifo_reg[7][27]/P0001  , \wishbone_rx_fifo_fifo_reg[7][28]/P0001  , \wishbone_rx_fifo_fifo_reg[7][29]/P0001  , \wishbone_rx_fifo_fifo_reg[7][2]/P0001  , \wishbone_rx_fifo_fifo_reg[7][30]/P0001  , \wishbone_rx_fifo_fifo_reg[7][31]/P0001  , \wishbone_rx_fifo_fifo_reg[7][3]/P0001  , \wishbone_rx_fifo_fifo_reg[7][4]/P0001  , \wishbone_rx_fifo_fifo_reg[7][5]/P0001  , \wishbone_rx_fifo_fifo_reg[7][6]/P0001  , \wishbone_rx_fifo_fifo_reg[7][7]/P0001  , \wishbone_rx_fifo_fifo_reg[7][8]/P0001  , \wishbone_rx_fifo_fifo_reg[7][9]/P0001  , \wishbone_rx_fifo_fifo_reg[8][0]/P0001  , \wishbone_rx_fifo_fifo_reg[8][10]/P0001  , \wishbone_rx_fifo_fifo_reg[8][11]/P0001  , \wishbone_rx_fifo_fifo_reg[8][12]/P0001  , \wishbone_rx_fifo_fifo_reg[8][13]/P0001  , \wishbone_rx_fifo_fifo_reg[8][14]/P0001  , \wishbone_rx_fifo_fifo_reg[8][15]/P0001  , \wishbone_rx_fifo_fifo_reg[8][16]/P0001  , \wishbone_rx_fifo_fifo_reg[8][17]/P0001  , \wishbone_rx_fifo_fifo_reg[8][18]/P0001  , \wishbone_rx_fifo_fifo_reg[8][19]/P0001  , \wishbone_rx_fifo_fifo_reg[8][1]/P0001  , \wishbone_rx_fifo_fifo_reg[8][20]/P0001  , \wishbone_rx_fifo_fifo_reg[8][21]/P0001  , \wishbone_rx_fifo_fifo_reg[8][22]/P0001  , \wishbone_rx_fifo_fifo_reg[8][23]/P0001  , \wishbone_rx_fifo_fifo_reg[8][24]/P0001  , \wishbone_rx_fifo_fifo_reg[8][25]/P0001  , \wishbone_rx_fifo_fifo_reg[8][26]/P0001  , \wishbone_rx_fifo_fifo_reg[8][27]/P0001  , \wishbone_rx_fifo_fifo_reg[8][28]/P0001  , \wishbone_rx_fifo_fifo_reg[8][29]/P0001  , \wishbone_rx_fifo_fifo_reg[8][2]/P0001  , \wishbone_rx_fifo_fifo_reg[8][30]/P0001  , \wishbone_rx_fifo_fifo_reg[8][31]/P0001  , \wishbone_rx_fifo_fifo_reg[8][3]/P0001  , \wishbone_rx_fifo_fifo_reg[8][4]/P0001  , \wishbone_rx_fifo_fifo_reg[8][5]/P0001  , \wishbone_rx_fifo_fifo_reg[8][6]/P0001  , \wishbone_rx_fifo_fifo_reg[8][7]/P0001  , \wishbone_rx_fifo_fifo_reg[8][8]/P0001  , \wishbone_rx_fifo_fifo_reg[8][9]/P0001  , \wishbone_rx_fifo_fifo_reg[9][0]/P0001  , \wishbone_rx_fifo_fifo_reg[9][10]/P0001  , \wishbone_rx_fifo_fifo_reg[9][11]/P0001  , \wishbone_rx_fifo_fifo_reg[9][12]/P0001  , \wishbone_rx_fifo_fifo_reg[9][13]/P0001  , \wishbone_rx_fifo_fifo_reg[9][14]/P0001  , \wishbone_rx_fifo_fifo_reg[9][15]/P0001  , \wishbone_rx_fifo_fifo_reg[9][16]/P0001  , \wishbone_rx_fifo_fifo_reg[9][17]/P0001  , \wishbone_rx_fifo_fifo_reg[9][18]/P0001  , \wishbone_rx_fifo_fifo_reg[9][19]/P0001  , \wishbone_rx_fifo_fifo_reg[9][1]/P0001  , \wishbone_rx_fifo_fifo_reg[9][20]/P0001  , \wishbone_rx_fifo_fifo_reg[9][21]/P0001  , \wishbone_rx_fifo_fifo_reg[9][22]/P0001  , \wishbone_rx_fifo_fifo_reg[9][23]/P0001  , \wishbone_rx_fifo_fifo_reg[9][24]/P0001  , \wishbone_rx_fifo_fifo_reg[9][25]/P0001  , \wishbone_rx_fifo_fifo_reg[9][26]/P0001  , \wishbone_rx_fifo_fifo_reg[9][27]/P0001  , \wishbone_rx_fifo_fifo_reg[9][28]/P0001  , \wishbone_rx_fifo_fifo_reg[9][29]/P0001  , \wishbone_rx_fifo_fifo_reg[9][2]/P0001  , \wishbone_rx_fifo_fifo_reg[9][30]/P0001  , \wishbone_rx_fifo_fifo_reg[9][31]/P0001  , \wishbone_rx_fifo_fifo_reg[9][3]/P0001  , \wishbone_rx_fifo_fifo_reg[9][4]/P0001  , \wishbone_rx_fifo_fifo_reg[9][5]/P0001  , \wishbone_rx_fifo_fifo_reg[9][6]/P0001  , \wishbone_rx_fifo_fifo_reg[9][7]/P0001  , \wishbone_rx_fifo_fifo_reg[9][8]/P0001  , \wishbone_rx_fifo_fifo_reg[9][9]/P0001  , \wishbone_rx_fifo_read_pointer_reg[0]/NET0131  , \wishbone_rx_fifo_read_pointer_reg[1]/NET0131  , \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  , \wishbone_rx_fifo_read_pointer_reg[3]/NET0131  , \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  , \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  , \wishbone_rx_fifo_write_pointer_reg[2]/NET0131  , \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  , \wishbone_tx_burst_cnt_reg[0]/NET0131  , \wishbone_tx_burst_cnt_reg[1]/NET0131  , \wishbone_tx_burst_cnt_reg[2]/NET0131  , \wishbone_tx_burst_en_reg/NET0131  , \wishbone_tx_fifo_cnt_reg[0]/NET0131  , \wishbone_tx_fifo_cnt_reg[1]/NET0131  , \wishbone_tx_fifo_cnt_reg[2]/NET0131  , \wishbone_tx_fifo_cnt_reg[3]/NET0131  , \wishbone_tx_fifo_cnt_reg[4]/NET0131  , \wishbone_tx_fifo_data_out_reg[0]/P0001  , \wishbone_tx_fifo_data_out_reg[10]/P0001  , \wishbone_tx_fifo_data_out_reg[11]/P0001  , \wishbone_tx_fifo_data_out_reg[12]/P0001  , \wishbone_tx_fifo_data_out_reg[13]/P0001  , \wishbone_tx_fifo_data_out_reg[14]/P0001  , \wishbone_tx_fifo_data_out_reg[15]/P0001  , \wishbone_tx_fifo_data_out_reg[16]/P0001  , \wishbone_tx_fifo_data_out_reg[17]/P0001  , \wishbone_tx_fifo_data_out_reg[18]/P0001  , \wishbone_tx_fifo_data_out_reg[19]/P0001  , \wishbone_tx_fifo_data_out_reg[1]/P0001  , \wishbone_tx_fifo_data_out_reg[20]/P0001  , \wishbone_tx_fifo_data_out_reg[21]/P0001  , \wishbone_tx_fifo_data_out_reg[22]/P0001  , \wishbone_tx_fifo_data_out_reg[23]/P0001  , \wishbone_tx_fifo_data_out_reg[24]/P0001  , \wishbone_tx_fifo_data_out_reg[25]/P0001  , \wishbone_tx_fifo_data_out_reg[26]/P0001  , \wishbone_tx_fifo_data_out_reg[27]/P0001  , \wishbone_tx_fifo_data_out_reg[28]/P0001  , \wishbone_tx_fifo_data_out_reg[29]/P0001  , \wishbone_tx_fifo_data_out_reg[2]/P0001  , \wishbone_tx_fifo_data_out_reg[30]/P0001  , \wishbone_tx_fifo_data_out_reg[31]/P0001  , \wishbone_tx_fifo_data_out_reg[3]/P0001  , \wishbone_tx_fifo_data_out_reg[4]/P0001  , \wishbone_tx_fifo_data_out_reg[5]/P0001  , \wishbone_tx_fifo_data_out_reg[6]/P0001  , \wishbone_tx_fifo_data_out_reg[7]/P0001  , \wishbone_tx_fifo_data_out_reg[8]/P0001  , \wishbone_tx_fifo_data_out_reg[9]/P0001  , \wishbone_tx_fifo_fifo_reg[0][0]/P0001  , \wishbone_tx_fifo_fifo_reg[0][10]/P0001  , \wishbone_tx_fifo_fifo_reg[0][11]/P0001  , \wishbone_tx_fifo_fifo_reg[0][12]/P0001  , \wishbone_tx_fifo_fifo_reg[0][13]/P0001  , \wishbone_tx_fifo_fifo_reg[0][14]/P0001  , \wishbone_tx_fifo_fifo_reg[0][15]/P0001  , \wishbone_tx_fifo_fifo_reg[0][16]/P0001  , \wishbone_tx_fifo_fifo_reg[0][17]/P0001  , \wishbone_tx_fifo_fifo_reg[0][18]/P0001  , \wishbone_tx_fifo_fifo_reg[0][19]/P0001  , \wishbone_tx_fifo_fifo_reg[0][1]/P0001  , \wishbone_tx_fifo_fifo_reg[0][20]/P0001  , \wishbone_tx_fifo_fifo_reg[0][21]/P0001  , \wishbone_tx_fifo_fifo_reg[0][22]/P0001  , \wishbone_tx_fifo_fifo_reg[0][23]/P0001  , \wishbone_tx_fifo_fifo_reg[0][24]/P0001  , \wishbone_tx_fifo_fifo_reg[0][25]/P0001  , \wishbone_tx_fifo_fifo_reg[0][26]/P0001  , \wishbone_tx_fifo_fifo_reg[0][27]/P0001  , \wishbone_tx_fifo_fifo_reg[0][28]/P0001  , \wishbone_tx_fifo_fifo_reg[0][29]/P0001  , \wishbone_tx_fifo_fifo_reg[0][2]/P0001  , \wishbone_tx_fifo_fifo_reg[0][30]/P0001  , \wishbone_tx_fifo_fifo_reg[0][31]/P0001  , \wishbone_tx_fifo_fifo_reg[0][3]/P0001  , \wishbone_tx_fifo_fifo_reg[0][4]/P0001  , \wishbone_tx_fifo_fifo_reg[0][5]/P0001  , \wishbone_tx_fifo_fifo_reg[0][6]/P0001  , \wishbone_tx_fifo_fifo_reg[0][7]/P0001  , \wishbone_tx_fifo_fifo_reg[0][8]/P0001  , \wishbone_tx_fifo_fifo_reg[0][9]/P0001  , \wishbone_tx_fifo_fifo_reg[10][0]/P0001  , \wishbone_tx_fifo_fifo_reg[10][10]/P0001  , \wishbone_tx_fifo_fifo_reg[10][11]/P0001  , \wishbone_tx_fifo_fifo_reg[10][12]/P0001  , \wishbone_tx_fifo_fifo_reg[10][13]/P0001  , \wishbone_tx_fifo_fifo_reg[10][14]/P0001  , \wishbone_tx_fifo_fifo_reg[10][15]/P0001  , \wishbone_tx_fifo_fifo_reg[10][16]/P0001  , \wishbone_tx_fifo_fifo_reg[10][17]/P0001  , \wishbone_tx_fifo_fifo_reg[10][18]/P0001  , \wishbone_tx_fifo_fifo_reg[10][19]/P0001  , \wishbone_tx_fifo_fifo_reg[10][1]/P0001  , \wishbone_tx_fifo_fifo_reg[10][20]/P0001  , \wishbone_tx_fifo_fifo_reg[10][21]/P0001  , \wishbone_tx_fifo_fifo_reg[10][22]/P0001  , \wishbone_tx_fifo_fifo_reg[10][23]/P0001  , \wishbone_tx_fifo_fifo_reg[10][24]/P0001  , \wishbone_tx_fifo_fifo_reg[10][25]/P0001  , \wishbone_tx_fifo_fifo_reg[10][26]/P0001  , \wishbone_tx_fifo_fifo_reg[10][27]/P0001  , \wishbone_tx_fifo_fifo_reg[10][28]/P0001  , \wishbone_tx_fifo_fifo_reg[10][29]/P0001  , \wishbone_tx_fifo_fifo_reg[10][2]/P0001  , \wishbone_tx_fifo_fifo_reg[10][30]/P0001  , \wishbone_tx_fifo_fifo_reg[10][31]/P0001  , \wishbone_tx_fifo_fifo_reg[10][3]/P0001  , \wishbone_tx_fifo_fifo_reg[10][4]/P0001  , \wishbone_tx_fifo_fifo_reg[10][5]/P0001  , \wishbone_tx_fifo_fifo_reg[10][6]/P0001  , \wishbone_tx_fifo_fifo_reg[10][7]/P0001  , \wishbone_tx_fifo_fifo_reg[10][8]/P0001  , \wishbone_tx_fifo_fifo_reg[10][9]/P0001  , \wishbone_tx_fifo_fifo_reg[11][0]/P0001  , \wishbone_tx_fifo_fifo_reg[11][10]/P0001  , \wishbone_tx_fifo_fifo_reg[11][11]/P0001  , \wishbone_tx_fifo_fifo_reg[11][12]/P0001  , \wishbone_tx_fifo_fifo_reg[11][13]/P0001  , \wishbone_tx_fifo_fifo_reg[11][14]/P0001  , \wishbone_tx_fifo_fifo_reg[11][15]/P0001  , \wishbone_tx_fifo_fifo_reg[11][16]/P0001  , \wishbone_tx_fifo_fifo_reg[11][17]/P0001  , \wishbone_tx_fifo_fifo_reg[11][18]/P0001  , \wishbone_tx_fifo_fifo_reg[11][19]/P0001  , \wishbone_tx_fifo_fifo_reg[11][1]/P0001  , \wishbone_tx_fifo_fifo_reg[11][20]/P0001  , \wishbone_tx_fifo_fifo_reg[11][21]/P0001  , \wishbone_tx_fifo_fifo_reg[11][22]/P0001  , \wishbone_tx_fifo_fifo_reg[11][23]/P0001  , \wishbone_tx_fifo_fifo_reg[11][24]/P0001  , \wishbone_tx_fifo_fifo_reg[11][25]/P0001  , \wishbone_tx_fifo_fifo_reg[11][26]/P0001  , \wishbone_tx_fifo_fifo_reg[11][27]/P0001  , \wishbone_tx_fifo_fifo_reg[11][28]/P0001  , \wishbone_tx_fifo_fifo_reg[11][29]/P0001  , \wishbone_tx_fifo_fifo_reg[11][2]/P0001  , \wishbone_tx_fifo_fifo_reg[11][30]/P0001  , \wishbone_tx_fifo_fifo_reg[11][31]/P0001  , \wishbone_tx_fifo_fifo_reg[11][3]/P0001  , \wishbone_tx_fifo_fifo_reg[11][4]/P0001  , \wishbone_tx_fifo_fifo_reg[11][5]/P0001  , \wishbone_tx_fifo_fifo_reg[11][6]/P0001  , \wishbone_tx_fifo_fifo_reg[11][7]/P0001  , \wishbone_tx_fifo_fifo_reg[11][8]/P0001  , \wishbone_tx_fifo_fifo_reg[11][9]/P0001  , \wishbone_tx_fifo_fifo_reg[12][0]/P0001  , \wishbone_tx_fifo_fifo_reg[12][10]/P0001  , \wishbone_tx_fifo_fifo_reg[12][11]/P0001  , \wishbone_tx_fifo_fifo_reg[12][12]/P0001  , \wishbone_tx_fifo_fifo_reg[12][13]/P0001  , \wishbone_tx_fifo_fifo_reg[12][14]/P0001  , \wishbone_tx_fifo_fifo_reg[12][15]/P0001  , \wishbone_tx_fifo_fifo_reg[12][16]/P0001  , \wishbone_tx_fifo_fifo_reg[12][17]/P0001  , \wishbone_tx_fifo_fifo_reg[12][18]/P0001  , \wishbone_tx_fifo_fifo_reg[12][19]/P0001  , \wishbone_tx_fifo_fifo_reg[12][1]/P0001  , \wishbone_tx_fifo_fifo_reg[12][20]/P0001  , \wishbone_tx_fifo_fifo_reg[12][21]/P0001  , \wishbone_tx_fifo_fifo_reg[12][22]/P0001  , \wishbone_tx_fifo_fifo_reg[12][23]/P0001  , \wishbone_tx_fifo_fifo_reg[12][24]/P0001  , \wishbone_tx_fifo_fifo_reg[12][25]/P0001  , \wishbone_tx_fifo_fifo_reg[12][26]/P0001  , \wishbone_tx_fifo_fifo_reg[12][27]/P0001  , \wishbone_tx_fifo_fifo_reg[12][28]/P0001  , \wishbone_tx_fifo_fifo_reg[12][29]/P0001  , \wishbone_tx_fifo_fifo_reg[12][2]/P0001  , \wishbone_tx_fifo_fifo_reg[12][30]/P0001  , \wishbone_tx_fifo_fifo_reg[12][31]/P0001  , \wishbone_tx_fifo_fifo_reg[12][3]/P0001  , \wishbone_tx_fifo_fifo_reg[12][4]/P0001  , \wishbone_tx_fifo_fifo_reg[12][5]/P0001  , \wishbone_tx_fifo_fifo_reg[12][6]/P0001  , \wishbone_tx_fifo_fifo_reg[12][7]/P0001  , \wishbone_tx_fifo_fifo_reg[12][8]/P0001  , \wishbone_tx_fifo_fifo_reg[12][9]/P0001  , \wishbone_tx_fifo_fifo_reg[13][0]/P0001  , \wishbone_tx_fifo_fifo_reg[13][10]/P0001  , \wishbone_tx_fifo_fifo_reg[13][11]/P0001  , \wishbone_tx_fifo_fifo_reg[13][12]/P0001  , \wishbone_tx_fifo_fifo_reg[13][13]/P0001  , \wishbone_tx_fifo_fifo_reg[13][14]/P0001  , \wishbone_tx_fifo_fifo_reg[13][15]/P0001  , \wishbone_tx_fifo_fifo_reg[13][16]/P0001  , \wishbone_tx_fifo_fifo_reg[13][17]/P0001  , \wishbone_tx_fifo_fifo_reg[13][18]/P0001  , \wishbone_tx_fifo_fifo_reg[13][19]/P0001  , \wishbone_tx_fifo_fifo_reg[13][1]/P0001  , \wishbone_tx_fifo_fifo_reg[13][20]/P0001  , \wishbone_tx_fifo_fifo_reg[13][21]/P0001  , \wishbone_tx_fifo_fifo_reg[13][22]/P0001  , \wishbone_tx_fifo_fifo_reg[13][23]/P0001  , \wishbone_tx_fifo_fifo_reg[13][24]/P0001  , \wishbone_tx_fifo_fifo_reg[13][25]/P0001  , \wishbone_tx_fifo_fifo_reg[13][26]/P0001  , \wishbone_tx_fifo_fifo_reg[13][27]/P0001  , \wishbone_tx_fifo_fifo_reg[13][28]/P0001  , \wishbone_tx_fifo_fifo_reg[13][29]/P0001  , \wishbone_tx_fifo_fifo_reg[13][2]/P0001  , \wishbone_tx_fifo_fifo_reg[13][30]/P0001  , \wishbone_tx_fifo_fifo_reg[13][31]/P0001  , \wishbone_tx_fifo_fifo_reg[13][3]/P0001  , \wishbone_tx_fifo_fifo_reg[13][4]/P0001  , \wishbone_tx_fifo_fifo_reg[13][5]/P0001  , \wishbone_tx_fifo_fifo_reg[13][6]/P0001  , \wishbone_tx_fifo_fifo_reg[13][7]/P0001  , \wishbone_tx_fifo_fifo_reg[13][8]/P0001  , \wishbone_tx_fifo_fifo_reg[13][9]/P0001  , \wishbone_tx_fifo_fifo_reg[14][0]/P0001  , \wishbone_tx_fifo_fifo_reg[14][10]/P0001  , \wishbone_tx_fifo_fifo_reg[14][11]/P0001  , \wishbone_tx_fifo_fifo_reg[14][12]/P0001  , \wishbone_tx_fifo_fifo_reg[14][13]/P0001  , \wishbone_tx_fifo_fifo_reg[14][14]/P0001  , \wishbone_tx_fifo_fifo_reg[14][15]/P0001  , \wishbone_tx_fifo_fifo_reg[14][16]/P0001  , \wishbone_tx_fifo_fifo_reg[14][17]/P0001  , \wishbone_tx_fifo_fifo_reg[14][18]/P0001  , \wishbone_tx_fifo_fifo_reg[14][19]/P0001  , \wishbone_tx_fifo_fifo_reg[14][1]/P0001  , \wishbone_tx_fifo_fifo_reg[14][20]/P0001  , \wishbone_tx_fifo_fifo_reg[14][21]/P0001  , \wishbone_tx_fifo_fifo_reg[14][22]/P0001  , \wishbone_tx_fifo_fifo_reg[14][23]/P0001  , \wishbone_tx_fifo_fifo_reg[14][24]/P0001  , \wishbone_tx_fifo_fifo_reg[14][25]/P0001  , \wishbone_tx_fifo_fifo_reg[14][26]/P0001  , \wishbone_tx_fifo_fifo_reg[14][27]/P0001  , \wishbone_tx_fifo_fifo_reg[14][28]/P0001  , \wishbone_tx_fifo_fifo_reg[14][29]/P0001  , \wishbone_tx_fifo_fifo_reg[14][2]/P0001  , \wishbone_tx_fifo_fifo_reg[14][30]/P0001  , \wishbone_tx_fifo_fifo_reg[14][31]/P0001  , \wishbone_tx_fifo_fifo_reg[14][3]/P0001  , \wishbone_tx_fifo_fifo_reg[14][4]/P0001  , \wishbone_tx_fifo_fifo_reg[14][5]/P0001  , \wishbone_tx_fifo_fifo_reg[14][6]/P0001  , \wishbone_tx_fifo_fifo_reg[14][7]/P0001  , \wishbone_tx_fifo_fifo_reg[14][8]/P0001  , \wishbone_tx_fifo_fifo_reg[14][9]/P0001  , \wishbone_tx_fifo_fifo_reg[15][0]/P0001  , \wishbone_tx_fifo_fifo_reg[15][10]/P0001  , \wishbone_tx_fifo_fifo_reg[15][11]/P0001  , \wishbone_tx_fifo_fifo_reg[15][12]/P0001  , \wishbone_tx_fifo_fifo_reg[15][13]/P0001  , \wishbone_tx_fifo_fifo_reg[15][14]/P0001  , \wishbone_tx_fifo_fifo_reg[15][15]/P0001  , \wishbone_tx_fifo_fifo_reg[15][16]/P0001  , \wishbone_tx_fifo_fifo_reg[15][17]/P0001  , \wishbone_tx_fifo_fifo_reg[15][18]/P0001  , \wishbone_tx_fifo_fifo_reg[15][19]/P0001  , \wishbone_tx_fifo_fifo_reg[15][1]/P0001  , \wishbone_tx_fifo_fifo_reg[15][20]/P0001  , \wishbone_tx_fifo_fifo_reg[15][21]/P0001  , \wishbone_tx_fifo_fifo_reg[15][22]/P0001  , \wishbone_tx_fifo_fifo_reg[15][23]/P0001  , \wishbone_tx_fifo_fifo_reg[15][24]/P0001  , \wishbone_tx_fifo_fifo_reg[15][25]/P0001  , \wishbone_tx_fifo_fifo_reg[15][26]/P0001  , \wishbone_tx_fifo_fifo_reg[15][27]/P0001  , \wishbone_tx_fifo_fifo_reg[15][28]/P0001  , \wishbone_tx_fifo_fifo_reg[15][29]/P0001  , \wishbone_tx_fifo_fifo_reg[15][2]/P0001  , \wishbone_tx_fifo_fifo_reg[15][30]/P0001  , \wishbone_tx_fifo_fifo_reg[15][31]/P0001  , \wishbone_tx_fifo_fifo_reg[15][3]/P0001  , \wishbone_tx_fifo_fifo_reg[15][4]/P0001  , \wishbone_tx_fifo_fifo_reg[15][5]/P0001  , \wishbone_tx_fifo_fifo_reg[15][6]/P0001  , \wishbone_tx_fifo_fifo_reg[15][7]/P0001  , \wishbone_tx_fifo_fifo_reg[15][8]/P0001  , \wishbone_tx_fifo_fifo_reg[15][9]/P0001  , \wishbone_tx_fifo_fifo_reg[1][0]/P0001  , \wishbone_tx_fifo_fifo_reg[1][10]/P0001  , \wishbone_tx_fifo_fifo_reg[1][11]/P0001  , \wishbone_tx_fifo_fifo_reg[1][12]/P0001  , \wishbone_tx_fifo_fifo_reg[1][13]/P0001  , \wishbone_tx_fifo_fifo_reg[1][14]/P0001  , \wishbone_tx_fifo_fifo_reg[1][15]/P0001  , \wishbone_tx_fifo_fifo_reg[1][16]/P0001  , \wishbone_tx_fifo_fifo_reg[1][17]/P0001  , \wishbone_tx_fifo_fifo_reg[1][18]/P0001  , \wishbone_tx_fifo_fifo_reg[1][19]/P0001  , \wishbone_tx_fifo_fifo_reg[1][1]/P0001  , \wishbone_tx_fifo_fifo_reg[1][20]/P0001  , \wishbone_tx_fifo_fifo_reg[1][21]/P0001  , \wishbone_tx_fifo_fifo_reg[1][22]/P0001  , \wishbone_tx_fifo_fifo_reg[1][23]/P0001  , \wishbone_tx_fifo_fifo_reg[1][24]/P0001  , \wishbone_tx_fifo_fifo_reg[1][25]/P0001  , \wishbone_tx_fifo_fifo_reg[1][26]/P0001  , \wishbone_tx_fifo_fifo_reg[1][27]/P0001  , \wishbone_tx_fifo_fifo_reg[1][28]/P0001  , \wishbone_tx_fifo_fifo_reg[1][29]/P0001  , \wishbone_tx_fifo_fifo_reg[1][2]/P0001  , \wishbone_tx_fifo_fifo_reg[1][30]/P0001  , \wishbone_tx_fifo_fifo_reg[1][31]/P0001  , \wishbone_tx_fifo_fifo_reg[1][3]/P0001  , \wishbone_tx_fifo_fifo_reg[1][4]/P0001  , \wishbone_tx_fifo_fifo_reg[1][5]/P0001  , \wishbone_tx_fifo_fifo_reg[1][6]/P0001  , \wishbone_tx_fifo_fifo_reg[1][7]/P0001  , \wishbone_tx_fifo_fifo_reg[1][8]/P0001  , \wishbone_tx_fifo_fifo_reg[1][9]/P0001  , \wishbone_tx_fifo_fifo_reg[2][0]/P0001  , \wishbone_tx_fifo_fifo_reg[2][10]/P0001  , \wishbone_tx_fifo_fifo_reg[2][11]/P0001  , \wishbone_tx_fifo_fifo_reg[2][12]/P0001  , \wishbone_tx_fifo_fifo_reg[2][13]/P0001  , \wishbone_tx_fifo_fifo_reg[2][14]/P0001  , \wishbone_tx_fifo_fifo_reg[2][15]/P0001  , \wishbone_tx_fifo_fifo_reg[2][16]/P0001  , \wishbone_tx_fifo_fifo_reg[2][17]/P0001  , \wishbone_tx_fifo_fifo_reg[2][18]/P0001  , \wishbone_tx_fifo_fifo_reg[2][19]/P0001  , \wishbone_tx_fifo_fifo_reg[2][1]/P0001  , \wishbone_tx_fifo_fifo_reg[2][20]/P0001  , \wishbone_tx_fifo_fifo_reg[2][21]/P0001  , \wishbone_tx_fifo_fifo_reg[2][22]/P0001  , \wishbone_tx_fifo_fifo_reg[2][23]/P0001  , \wishbone_tx_fifo_fifo_reg[2][24]/P0001  , \wishbone_tx_fifo_fifo_reg[2][25]/P0001  , \wishbone_tx_fifo_fifo_reg[2][26]/P0001  , \wishbone_tx_fifo_fifo_reg[2][27]/P0001  , \wishbone_tx_fifo_fifo_reg[2][28]/P0001  , \wishbone_tx_fifo_fifo_reg[2][29]/P0001  , \wishbone_tx_fifo_fifo_reg[2][2]/P0001  , \wishbone_tx_fifo_fifo_reg[2][30]/P0001  , \wishbone_tx_fifo_fifo_reg[2][31]/P0001  , \wishbone_tx_fifo_fifo_reg[2][3]/P0001  , \wishbone_tx_fifo_fifo_reg[2][4]/P0001  , \wishbone_tx_fifo_fifo_reg[2][5]/P0001  , \wishbone_tx_fifo_fifo_reg[2][6]/P0001  , \wishbone_tx_fifo_fifo_reg[2][7]/P0001  , \wishbone_tx_fifo_fifo_reg[2][8]/P0001  , \wishbone_tx_fifo_fifo_reg[2][9]/P0001  , \wishbone_tx_fifo_fifo_reg[3][0]/P0001  , \wishbone_tx_fifo_fifo_reg[3][10]/P0001  , \wishbone_tx_fifo_fifo_reg[3][11]/P0001  , \wishbone_tx_fifo_fifo_reg[3][12]/P0001  , \wishbone_tx_fifo_fifo_reg[3][13]/P0001  , \wishbone_tx_fifo_fifo_reg[3][14]/P0001  , \wishbone_tx_fifo_fifo_reg[3][15]/P0001  , \wishbone_tx_fifo_fifo_reg[3][16]/P0001  , \wishbone_tx_fifo_fifo_reg[3][17]/P0001  , \wishbone_tx_fifo_fifo_reg[3][18]/P0001  , \wishbone_tx_fifo_fifo_reg[3][19]/P0001  , \wishbone_tx_fifo_fifo_reg[3][1]/P0001  , \wishbone_tx_fifo_fifo_reg[3][20]/P0001  , \wishbone_tx_fifo_fifo_reg[3][21]/P0001  , \wishbone_tx_fifo_fifo_reg[3][22]/P0001  , \wishbone_tx_fifo_fifo_reg[3][23]/P0001  , \wishbone_tx_fifo_fifo_reg[3][24]/P0001  , \wishbone_tx_fifo_fifo_reg[3][25]/P0001  , \wishbone_tx_fifo_fifo_reg[3][26]/P0001  , \wishbone_tx_fifo_fifo_reg[3][27]/P0001  , \wishbone_tx_fifo_fifo_reg[3][28]/P0001  , \wishbone_tx_fifo_fifo_reg[3][29]/P0001  , \wishbone_tx_fifo_fifo_reg[3][2]/P0001  , \wishbone_tx_fifo_fifo_reg[3][30]/P0001  , \wishbone_tx_fifo_fifo_reg[3][31]/P0001  , \wishbone_tx_fifo_fifo_reg[3][3]/P0001  , \wishbone_tx_fifo_fifo_reg[3][4]/P0001  , \wishbone_tx_fifo_fifo_reg[3][5]/P0001  , \wishbone_tx_fifo_fifo_reg[3][6]/P0001  , \wishbone_tx_fifo_fifo_reg[3][7]/P0001  , \wishbone_tx_fifo_fifo_reg[3][8]/P0001  , \wishbone_tx_fifo_fifo_reg[3][9]/P0001  , \wishbone_tx_fifo_fifo_reg[4][0]/P0001  , \wishbone_tx_fifo_fifo_reg[4][10]/P0001  , \wishbone_tx_fifo_fifo_reg[4][11]/P0001  , \wishbone_tx_fifo_fifo_reg[4][12]/P0001  , \wishbone_tx_fifo_fifo_reg[4][13]/P0001  , \wishbone_tx_fifo_fifo_reg[4][14]/P0001  , \wishbone_tx_fifo_fifo_reg[4][15]/P0001  , \wishbone_tx_fifo_fifo_reg[4][16]/P0001  , \wishbone_tx_fifo_fifo_reg[4][17]/P0001  , \wishbone_tx_fifo_fifo_reg[4][18]/P0001  , \wishbone_tx_fifo_fifo_reg[4][19]/P0001  , \wishbone_tx_fifo_fifo_reg[4][1]/P0001  , \wishbone_tx_fifo_fifo_reg[4][20]/P0001  , \wishbone_tx_fifo_fifo_reg[4][21]/P0001  , \wishbone_tx_fifo_fifo_reg[4][22]/P0001  , \wishbone_tx_fifo_fifo_reg[4][23]/P0001  , \wishbone_tx_fifo_fifo_reg[4][24]/P0001  , \wishbone_tx_fifo_fifo_reg[4][25]/P0001  , \wishbone_tx_fifo_fifo_reg[4][26]/P0001  , \wishbone_tx_fifo_fifo_reg[4][27]/P0001  , \wishbone_tx_fifo_fifo_reg[4][28]/P0001  , \wishbone_tx_fifo_fifo_reg[4][29]/P0001  , \wishbone_tx_fifo_fifo_reg[4][2]/P0001  , \wishbone_tx_fifo_fifo_reg[4][30]/P0001  , \wishbone_tx_fifo_fifo_reg[4][31]/P0001  , \wishbone_tx_fifo_fifo_reg[4][3]/P0001  , \wishbone_tx_fifo_fifo_reg[4][4]/P0001  , \wishbone_tx_fifo_fifo_reg[4][5]/P0001  , \wishbone_tx_fifo_fifo_reg[4][6]/P0001  , \wishbone_tx_fifo_fifo_reg[4][7]/P0001  , \wishbone_tx_fifo_fifo_reg[4][8]/P0001  , \wishbone_tx_fifo_fifo_reg[4][9]/P0001  , \wishbone_tx_fifo_fifo_reg[5][0]/P0001  , \wishbone_tx_fifo_fifo_reg[5][10]/P0001  , \wishbone_tx_fifo_fifo_reg[5][11]/P0001  , \wishbone_tx_fifo_fifo_reg[5][12]/P0001  , \wishbone_tx_fifo_fifo_reg[5][13]/P0001  , \wishbone_tx_fifo_fifo_reg[5][14]/P0001  , \wishbone_tx_fifo_fifo_reg[5][15]/P0001  , \wishbone_tx_fifo_fifo_reg[5][16]/P0001  , \wishbone_tx_fifo_fifo_reg[5][17]/P0001  , \wishbone_tx_fifo_fifo_reg[5][18]/P0001  , \wishbone_tx_fifo_fifo_reg[5][19]/P0001  , \wishbone_tx_fifo_fifo_reg[5][1]/P0001  , \wishbone_tx_fifo_fifo_reg[5][20]/P0001  , \wishbone_tx_fifo_fifo_reg[5][21]/P0001  , \wishbone_tx_fifo_fifo_reg[5][22]/P0001  , \wishbone_tx_fifo_fifo_reg[5][23]/P0001  , \wishbone_tx_fifo_fifo_reg[5][24]/P0001  , \wishbone_tx_fifo_fifo_reg[5][25]/P0001  , \wishbone_tx_fifo_fifo_reg[5][26]/P0001  , \wishbone_tx_fifo_fifo_reg[5][27]/P0001  , \wishbone_tx_fifo_fifo_reg[5][28]/P0001  , \wishbone_tx_fifo_fifo_reg[5][29]/P0001  , \wishbone_tx_fifo_fifo_reg[5][2]/P0001  , \wishbone_tx_fifo_fifo_reg[5][30]/P0001  , \wishbone_tx_fifo_fifo_reg[5][31]/P0001  , \wishbone_tx_fifo_fifo_reg[5][3]/P0001  , \wishbone_tx_fifo_fifo_reg[5][4]/P0001  , \wishbone_tx_fifo_fifo_reg[5][5]/P0001  , \wishbone_tx_fifo_fifo_reg[5][6]/P0001  , \wishbone_tx_fifo_fifo_reg[5][7]/P0001  , \wishbone_tx_fifo_fifo_reg[5][8]/P0001  , \wishbone_tx_fifo_fifo_reg[5][9]/P0001  , \wishbone_tx_fifo_fifo_reg[6][0]/P0001  , \wishbone_tx_fifo_fifo_reg[6][10]/P0001  , \wishbone_tx_fifo_fifo_reg[6][11]/P0001  , \wishbone_tx_fifo_fifo_reg[6][12]/P0001  , \wishbone_tx_fifo_fifo_reg[6][13]/P0001  , \wishbone_tx_fifo_fifo_reg[6][14]/P0001  , \wishbone_tx_fifo_fifo_reg[6][15]/P0001  , \wishbone_tx_fifo_fifo_reg[6][16]/P0001  , \wishbone_tx_fifo_fifo_reg[6][17]/P0001  , \wishbone_tx_fifo_fifo_reg[6][18]/P0001  , \wishbone_tx_fifo_fifo_reg[6][19]/P0001  , \wishbone_tx_fifo_fifo_reg[6][1]/P0001  , \wishbone_tx_fifo_fifo_reg[6][20]/P0001  , \wishbone_tx_fifo_fifo_reg[6][21]/P0001  , \wishbone_tx_fifo_fifo_reg[6][22]/P0001  , \wishbone_tx_fifo_fifo_reg[6][23]/P0001  , \wishbone_tx_fifo_fifo_reg[6][24]/P0001  , \wishbone_tx_fifo_fifo_reg[6][25]/P0001  , \wishbone_tx_fifo_fifo_reg[6][26]/P0001  , \wishbone_tx_fifo_fifo_reg[6][27]/P0001  , \wishbone_tx_fifo_fifo_reg[6][28]/P0001  , \wishbone_tx_fifo_fifo_reg[6][29]/P0001  , \wishbone_tx_fifo_fifo_reg[6][2]/P0001  , \wishbone_tx_fifo_fifo_reg[6][30]/P0001  , \wishbone_tx_fifo_fifo_reg[6][31]/P0001  , \wishbone_tx_fifo_fifo_reg[6][3]/P0001  , \wishbone_tx_fifo_fifo_reg[6][4]/P0001  , \wishbone_tx_fifo_fifo_reg[6][5]/P0001  , \wishbone_tx_fifo_fifo_reg[6][6]/P0001  , \wishbone_tx_fifo_fifo_reg[6][7]/P0001  , \wishbone_tx_fifo_fifo_reg[6][8]/P0001  , \wishbone_tx_fifo_fifo_reg[6][9]/P0001  , \wishbone_tx_fifo_fifo_reg[7][0]/P0001  , \wishbone_tx_fifo_fifo_reg[7][10]/P0001  , \wishbone_tx_fifo_fifo_reg[7][11]/P0001  , \wishbone_tx_fifo_fifo_reg[7][12]/P0001  , \wishbone_tx_fifo_fifo_reg[7][13]/P0001  , \wishbone_tx_fifo_fifo_reg[7][14]/P0001  , \wishbone_tx_fifo_fifo_reg[7][15]/P0001  , \wishbone_tx_fifo_fifo_reg[7][16]/P0001  , \wishbone_tx_fifo_fifo_reg[7][17]/P0001  , \wishbone_tx_fifo_fifo_reg[7][18]/P0001  , \wishbone_tx_fifo_fifo_reg[7][19]/P0001  , \wishbone_tx_fifo_fifo_reg[7][1]/P0001  , \wishbone_tx_fifo_fifo_reg[7][20]/P0001  , \wishbone_tx_fifo_fifo_reg[7][21]/P0001  , \wishbone_tx_fifo_fifo_reg[7][22]/P0001  , \wishbone_tx_fifo_fifo_reg[7][23]/P0001  , \wishbone_tx_fifo_fifo_reg[7][24]/P0001  , \wishbone_tx_fifo_fifo_reg[7][25]/P0001  , \wishbone_tx_fifo_fifo_reg[7][26]/P0001  , \wishbone_tx_fifo_fifo_reg[7][27]/P0001  , \wishbone_tx_fifo_fifo_reg[7][28]/P0001  , \wishbone_tx_fifo_fifo_reg[7][29]/P0001  , \wishbone_tx_fifo_fifo_reg[7][2]/P0001  , \wishbone_tx_fifo_fifo_reg[7][30]/P0001  , \wishbone_tx_fifo_fifo_reg[7][31]/P0001  , \wishbone_tx_fifo_fifo_reg[7][3]/P0001  , \wishbone_tx_fifo_fifo_reg[7][4]/P0001  , \wishbone_tx_fifo_fifo_reg[7][5]/P0001  , \wishbone_tx_fifo_fifo_reg[7][6]/P0001  , \wishbone_tx_fifo_fifo_reg[7][7]/P0001  , \wishbone_tx_fifo_fifo_reg[7][8]/P0001  , \wishbone_tx_fifo_fifo_reg[7][9]/P0001  , \wishbone_tx_fifo_fifo_reg[8][0]/P0001  , \wishbone_tx_fifo_fifo_reg[8][10]/P0001  , \wishbone_tx_fifo_fifo_reg[8][11]/P0001  , \wishbone_tx_fifo_fifo_reg[8][12]/P0001  , \wishbone_tx_fifo_fifo_reg[8][13]/P0001  , \wishbone_tx_fifo_fifo_reg[8][14]/P0001  , \wishbone_tx_fifo_fifo_reg[8][15]/P0001  , \wishbone_tx_fifo_fifo_reg[8][16]/P0001  , \wishbone_tx_fifo_fifo_reg[8][17]/P0001  , \wishbone_tx_fifo_fifo_reg[8][18]/P0001  , \wishbone_tx_fifo_fifo_reg[8][19]/P0001  , \wishbone_tx_fifo_fifo_reg[8][1]/P0001  , \wishbone_tx_fifo_fifo_reg[8][20]/P0001  , \wishbone_tx_fifo_fifo_reg[8][21]/P0001  , \wishbone_tx_fifo_fifo_reg[8][22]/P0001  , \wishbone_tx_fifo_fifo_reg[8][23]/P0001  , \wishbone_tx_fifo_fifo_reg[8][24]/P0001  , \wishbone_tx_fifo_fifo_reg[8][25]/P0001  , \wishbone_tx_fifo_fifo_reg[8][26]/P0001  , \wishbone_tx_fifo_fifo_reg[8][27]/P0001  , \wishbone_tx_fifo_fifo_reg[8][28]/P0001  , \wishbone_tx_fifo_fifo_reg[8][29]/P0001  , \wishbone_tx_fifo_fifo_reg[8][2]/P0001  , \wishbone_tx_fifo_fifo_reg[8][30]/P0001  , \wishbone_tx_fifo_fifo_reg[8][31]/P0001  , \wishbone_tx_fifo_fifo_reg[8][3]/P0001  , \wishbone_tx_fifo_fifo_reg[8][4]/P0001  , \wishbone_tx_fifo_fifo_reg[8][5]/P0001  , \wishbone_tx_fifo_fifo_reg[8][6]/P0001  , \wishbone_tx_fifo_fifo_reg[8][7]/P0001  , \wishbone_tx_fifo_fifo_reg[8][8]/P0001  , \wishbone_tx_fifo_fifo_reg[8][9]/P0001  , \wishbone_tx_fifo_fifo_reg[9][0]/P0001  , \wishbone_tx_fifo_fifo_reg[9][10]/P0001  , \wishbone_tx_fifo_fifo_reg[9][11]/P0001  , \wishbone_tx_fifo_fifo_reg[9][12]/P0001  , \wishbone_tx_fifo_fifo_reg[9][13]/P0001  , \wishbone_tx_fifo_fifo_reg[9][14]/P0001  , \wishbone_tx_fifo_fifo_reg[9][15]/P0001  , \wishbone_tx_fifo_fifo_reg[9][16]/P0001  , \wishbone_tx_fifo_fifo_reg[9][17]/P0001  , \wishbone_tx_fifo_fifo_reg[9][18]/P0001  , \wishbone_tx_fifo_fifo_reg[9][19]/P0001  , \wishbone_tx_fifo_fifo_reg[9][1]/P0001  , \wishbone_tx_fifo_fifo_reg[9][20]/P0001  , \wishbone_tx_fifo_fifo_reg[9][21]/P0001  , \wishbone_tx_fifo_fifo_reg[9][22]/P0001  , \wishbone_tx_fifo_fifo_reg[9][23]/P0001  , \wishbone_tx_fifo_fifo_reg[9][24]/P0001  , \wishbone_tx_fifo_fifo_reg[9][25]/P0001  , \wishbone_tx_fifo_fifo_reg[9][26]/P0001  , \wishbone_tx_fifo_fifo_reg[9][27]/P0001  , \wishbone_tx_fifo_fifo_reg[9][28]/P0001  , \wishbone_tx_fifo_fifo_reg[9][29]/P0001  , \wishbone_tx_fifo_fifo_reg[9][2]/P0001  , \wishbone_tx_fifo_fifo_reg[9][30]/P0001  , \wishbone_tx_fifo_fifo_reg[9][31]/P0001  , \wishbone_tx_fifo_fifo_reg[9][3]/P0001  , \wishbone_tx_fifo_fifo_reg[9][4]/P0001  , \wishbone_tx_fifo_fifo_reg[9][5]/P0001  , \wishbone_tx_fifo_fifo_reg[9][6]/P0001  , \wishbone_tx_fifo_fifo_reg[9][7]/P0001  , \wishbone_tx_fifo_fifo_reg[9][8]/P0001  , \wishbone_tx_fifo_fifo_reg[9][9]/P0001  , \wishbone_tx_fifo_read_pointer_reg[0]/NET0131  , \wishbone_tx_fifo_read_pointer_reg[1]/NET0131  , \wishbone_tx_fifo_read_pointer_reg[2]/NET0131  , \wishbone_tx_fifo_read_pointer_reg[3]/NET0131  , \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  , \wishbone_tx_fifo_write_pointer_reg[1]/NET0131  , \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  , \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  , \_al_n1  , \g215539/_0_  , \g215543/_0_  , \g215547/_0_  , \g215551/_0_  , \g215552/_0_  , \g215578/_0_  , \g215587/_1_  , \g215589/_1_  , \g215591/_1_  , \g215593/_1_  , \g215595/_1_  , \g215597/_1_  , \g215599/_1_  , \g215601/_1_  , \g215603/_1_  , \g215605/_1_  , \g215607/_1_  , \g215609/_1_  , \g215611/_1_  , \g215613/_1_  , \g215615/_1_  , \g215617/_1_  , \g215618/_0_  , \g215619/_0_  , \g215620/_0_  , \g215632/_1_  , \g215634/_0_  , \g215635/_0_  , \g215636/_0_  , \g215637/_0_  , \g215638/_0_  , \g215639/_0_  , \g215655/_1_  , \g215657/_1_  , \g215659/_1_  , \g215661/_1_  , \g215662/_0_  , \g215663/_0_  , \g215664/_0_  , \g215665/_0_  , \g215668/_0_  , \g215674/_0_  , \g215677/_0_  , \g215686/_0_  , \g215695/_0_  , \g215696/_0_  , \g215702/_1__syn_2  , \g215705/_0_  , \g215706/_0_  , \g215716/_0_  , \g215717/_0_  , \g215718/_0_  , \g215726/_0_  , \g215727/_0_  , \g215728/_0_  , \g215760/_0_  , \g215764/_0_  , \g215765/_0_  , \g215766/_0_  , \g215767/_3_  , \g215768/_3_  , \g215769/_3_  , \g215770/_3_  , \g215771/_3_  , \g215772/_3_  , \g215773/_3_  , \g215774/_3_  , \g215775/_3_  , \g215776/_3_  , \g215777/_3_  , \g215778/_3_  , \g215779/_3_  , \g215780/_3_  , \g215790/_0_  , \g215791/_0_  , \g215792/_0_  , \g215793/_0_  , \g215801/_0_  , \g215802/_0_  , \g215803/_0_  , \g215804/_0_  , \g215812/_0_  , \g215813/_0_  , \g215821/_0_  , \g215823/_0_  , \g215831/_0_  , \g215832/_0_  , \g215833/_0_  , \g215845/_0_  , \g215846/_0_  , \g215847/_0_  , \g215872/_0_  , \g215873/_0_  , \g215874/_0_  , \g215904/_0_  , \g215905/_0_  , \g215906/_0_  , \g215907/_0_  , \g215908/_0_  , \g215909/_0_  , \g215910/_0_  , \g215911/_0_  , \g215912/_0_  , \g215913/_0_  , \g215914/_0_  , \g215915/_0_  , \g215916/_0_  , \g215917/_0_  , \g215918/_0_  , \g215919/_0_  , \g215920/_0_  , \g215923/_0_  , \g215926/_0_  , \g215941/_0_  , \g215942/_0_  , \g215943/_0_  , \g215944/_0_  , \g215945/_0_  , \g215946/_0_  , \g215947/_0_  , \g215948/_0_  , \g215949/_0_  , \g215950/_0_  , \g215951/_0_  , \g215952/_0_  , \g215953/_0_  , \g215954/_0_  , \g215955/_0_  , \g215956/_0_  , \g215957/_0_  , \g215959/_00_  , \g215960/_0_  , \g215962/_0_  , \g215964/_0_  , \g215966/_0_  , \g215972/_0_  , \g216035/_0_  , \g216037/_0_  , \g216038/_0_  , \g216039/_0_  , \g216040/_0_  , \g216041/_0_  , \g216042/_0_  , \g216046/_0_  , \g216048/_0_  , \g216057/_0_  , \g216263/_0_  , \g216264/_0_  , \g216265/_0_  , \g216266/_0_  , \g216267/_0_  , \g216268/_0_  , \g216269/_0_  , \g216270/_0_  , \g216271/_0_  , \g216272/_0_  , \g216273/_0_  , \g216284/_0_  , \g216289/_0_  , \g216290/_0_  , \g216292/_0_  , \g216296/_0_  , \g216297/_0_  , \g216300/_0_  , \g216301/_0_  , \g216302/_0_  , \g216303/_0_  , \g216304/_0_  , \g216305/_0_  , \g216306/_0_  , \g216307/_0_  , \g216310/_3_  , \g216311/_3_  , \g216314/u3_syn_7  , \g216322/_3_  , \g216323/_3_  , \g216324/_3_  , \g216325/_3_  , \g216326/_3_  , \g216327/_3_  , \g216328/_3_  , \g216329/_3_  , \g216369/_0_  , \g216370/_0_  , \g216371/_0_  , \g216372/_0_  , \g216373/_0_  , \g216374/_0_  , \g216375/_0_  , \g216376/_0_  , \g216379/_0_  , \g216380/_0_  , \g216381/_0_  , \g216385/_0_  , \g216389/_0_  , \g216390/_0_  , \g216402/_0_  , \g216404/_0_  , \g216405/_0_  , \g216406/_0_  , \g216407/_0_  , \g216408/_0_  , \g216409/_0_  , \g216410/_0_  , \g216411/_0_  , \g216412/_0_  , \g216413/_0_  , \g216414/_0_  , \g216415/_0_  , \g216416/_0_  , \g216417/_0_  , \g216418/_0_  , \g216419/_0_  , \g216420/_0_  , \g216421/_0_  , \g216422/_0_  , \g216423/_0_  , \g216424/_0_  , \g216425/_0_  , \g216426/_0_  , \g216427/_0_  , \g216428/_0_  , \g216429/_0_  , \g216430/_0_  , \g216431/_0_  , \g216432/_0_  , \g216433/_0_  , \g216434/_0_  , \g216435/_0_  , \g216436/_0_  , \g216437/_0_  , \g216438/_0_  , \g216439/_3_  , \g216447/_3_  , \g216448/_3_  , \g216452/_0_  , \g216453/_0_  , \g216454/_0_  , \g216455/_0_  , \g216456/_0_  , \g216457/_0_  , \g216458/_3_  , \g216459/_3_  , \g216461/_3_  , \g216462/_3_  , \g216463/_3_  , \g216464/_3_  , \g216465/_3_  , \g216466/_0_  , \g216467/_3_  , \g216468/_3_  , \g216469/_3_  , \g216470/_3_  , \g216471/_3_  , \g216473/_3_  , \g216474/_3_  , \g216475/_3_  , \g216476/_3_  , \g216477/_3_  , \g216478/_0_  , \g216479/_3_  , \g216480/_3_  , \g216481/_3_  , \g216492/_0_  , \g216494/_0_  , \g216495/_3_  , \g216496/_3_  , \g216498/_3_  , \g216499/_3_  , \g216500/_3_  , \g216513/_3_  , \g216514/_3_  , \g216515/_3_  , \g216516/_3_  , \g216517/_3_  , \g216518/_3_  , \g216519/_3_  , \g216520/_3_  , \g216521/_3_  , \g216522/_3_  , \g216523/_3_  , \g216524/_3_  , \g216525/_3_  , \g216526/_3_  , \g216527/_3_  , \g216528/_3_  , \g216529/_3_  , \g216530/_3_  , \g216531/_3_  , \g216532/_3_  , \g216533/_3_  , \g216534/_3_  , \g216535/_3_  , \g216536/_3_  , \g216537/_3_  , \g216538/_3_  , \g216555/_3_  , \g216556/_3_  , \g216557/_3_  , \g216560/_3_  , \g216561/_3_  , \g216562/_3_  , \g216563/_3_  , \g216564/_3_  , \g216565/_3_  , \g216566/_3_  , \g216567/_3_  , \g216568/_3_  , \g216569/_3_  , \g216570/_3_  , \g216571/_3_  , \g216575/_3_  , \g216576/_3_  , \g216577/_3_  , \g216578/_3_  , \g216579/_3_  , \g216580/_3_  , \g216581/_3_  , \g216582/_3_  , \g216583/_3_  , \g216586/_3_  , \g216587/_3_  , \g216588/_3_  , \g216589/_3_  , \g216590/_3_  , \g216591/_3_  , \g216592/_3_  , \g216593/_3_  , \g216594/_3_  , \g216595/_3_  , \g216600/_3_  , \g216683/_0_  , \g216689/_0_  , \g216693/_0_  , \g216694/_0_  , \g216727/_0_  , \g216728/_0_  , \g216729/_0_  , \g216732/_0_  , \g216733/_0_  , \g216734/_0_  , \g216735/_0_  , \g216736/_0_  , \g216737/_0_  , \g216738/_0_  , \g216739/_0_  , \g216740/_0_  , \g216741/_0_  , \g216742/_0_  , \g216743/_0_  , \g216744/_0_  , \g216745/_0_  , \g216746/_0_  , \g216748/_0_  , \g216751/_0_  , \g216754/_0_  , \g216762/_0_  , \g216934/_2_  , \g216952/_0_  , \g216955/_0_  , \g216969/_0_  , \g216979/_0_  , \g216984/_0_  , \g216996/_0_  , \g217002/_0_  , \g217014/_0_  , \g217015/_0_  , \g217016/_0_  , \g217017/_0_  , \g217018/_0_  , \g217019/_0_  , \g217023/_0_  , \g217116/_0_  , \g217146/_3_  , \g217149/_0_  , \g217151/_0_  , \g217160/_0_  , \g217167/_0_  , \g217168/_0_  , \g217169/_0_  , \g217170/_0_  , \g217171/_0_  , \g217172/_0_  , \g217173/_0_  , \g217174/_0_  , \g217175/_0_  , \g217176/_0_  , \g217177/_0_  , \g217178/_0_  , \g217179/_0_  , \g217180/_0_  , \g217181/_0_  , \g217182/_0_  , \g217183/_0_  , \g217187/_0_  , \g217188/_0_  , \g217189/_0_  , \g217193/_0_  , \g217194/_0_  , \g217195/_0_  , \g217196/_0_  , \g217202/_0_  , \g217205/_0_  , \g217206/_0_  , \g217207/_0_  , \g217208/_0_  , \g217209/_0_  , \g217210/_0_  , \g217211/_0_  , \g217212/_0_  , \g217213/_0_  , \g217214/_0_  , \g217215/_0_  , \g217216/_0_  , \g217217/_0_  , \g217218/_0_  , \g217219/_0_  , \g217220/_0_  , \g217223/_0_  , \g217231/_0_  , \g217237/_0_  , \g217238/_0_  , \g217242/_0_  , \g217243/_0_  , \g217250/_3_  , \g217251/_3_  , \g217252/_3_  , \g217253/_3_  , \g217254/_3_  , \g217255/_3_  , \g217256/_3_  , \g217257/_3_  , \g217258/_3_  , \g217259/_3_  , \g217260/_3_  , \g217261/_3_  , \g217262/_3_  , \g217263/_3_  , \g217264/_3_  , \g217265/_3_  , \g217266/_3_  , \g217267/_3_  , \g217268/_3_  , \g217269/_3_  , \g217270/_3_  , \g217271/_3_  , \g217272/_3_  , \g217273/_3_  , \g217274/_3_  , \g217275/_3_  , \g217276/_3_  , \g217277/_3_  , \g217278/_3_  , \g217279/_3_  , \g217280/_3_  , \g217281/_3_  , \g217282/_3_  , \g217283/_3_  , \g217284/_3_  , \g217285/_3_  , \g217286/_3_  , \g217287/_3_  , \g217288/_3_  , \g217289/_3_  , \g217290/_3_  , \g217291/_3_  , \g217292/_3_  , \g217293/_3_  , \g217294/_3_  , \g217295/_3_  , \g217296/_3_  , \g217297/_3_  , \g217298/_3_  , \g217299/_3_  , \g217300/_3_  , \g217301/_3_  , \g217302/_3_  , \g217303/_3_  , \g217304/_3_  , \g217305/_3_  , \g217306/_3_  , \g217307/_3_  , \g217308/_3_  , \g217309/_3_  , \g217310/_3_  , \g217311/_3_  , \g217312/_3_  , \g217313/_3_  , \g217318/_0_  , \g217662/_0_  , \g217663/_0_  , \g217682/_0_  , \g217697/_0_  , \g217698/_0_  , \g217699/_0_  , \g217700/_0_  , \g217701/_0_  , \g217705/_0_  , \g217711/_0_  , \g217747/_0_  , \g217753/_00_  , \g217775/_0_  , \g217781/_0_  , \g217784/_0_  , \g217785/_0_  , \g217786/_0_  , \g217787/_0_  , \g217788/_0_  , \g217790/_0_  , \g217815/_0_  , \g217817/_0_  , \g218145/_0_  , \g218148/_0_  , \g218150/_0_  , \g218167/_0_  , \g218168/_0_  , \g218234/_0_  , \g218235/_0_  , \g218236/_0_  , \g218238/_0_  , \g218242/_0_  , \g218332/_0_  , \g218335/_0_  , \g218336/_0_  , \g218337/_0_  , \g218338/_0_  , \g218339/_0_  , \g218340/_0_  , \g218341/_0_  , \g218342/_0_  , \g218343/_0_  , \g218344/_0_  , \g218345/_0_  , \g218346/_0_  , \g218347/_0_  , \g218348/_0_  , \g218349/_0_  , \g218350/_0_  , \g218351/_0_  , \g218352/_0_  , \g218353/_0_  , \g218354/_0_  , \g218355/_0_  , \g218356/_0_  , \g218357/_0_  , \g218358/_0_  , \g218359/_0_  , \g218360/_0_  , \g218398/_3_  , \g218430/_0_  , \g218440/_0_  , \g218452/u3_syn_4  , \g218495/u3_syn_4  , \g218517/u3_syn_4  , \g218554/u3_syn_4  , \g218575/u3_syn_4  , \g218600/u3_syn_4  , \g218621/u3_syn_4  , \g218638/u3_syn_4  , \g218659/u3_syn_4  , \g218673/u3_syn_4  , \g218707/u3_syn_4  , \g218735/_3_  , \g219186/_0_  , \g219187/_0_  , \g219188/_0_  , \g219189/_0_  , \g219190/_0_  , \g219196/_0_  , \g219198/_0_  , \g219199/_0_  , \g219200/_0_  , \g219308/_0_  , \g219314/_0_  , \g219326/_0_  , \g219328/_0_  , \g219348/_0_  , \g219351/_0_  , \g219363/_0_  , \g219364/_0_  , \g219365/_0_  , \g219366/_0_  , \g219367/_0_  , \g219368/_0_  , \g219369/_0_  , \g219376/_0_  , \g219381/_0_  , \g219382/_0_  , \g219384/_0_  , \g219385/_0_  , \g219391/_0_  , \g219394/_0_  , \g219395/_0_  , \g219396/_0_  , \g219397/_0_  , \g219398/_0_  , \g219399/_0_  , \g219400/_0_  , \g219401/_0_  , \g219402/_0_  , \g219403/_0_  , \g219404/_0_  , \g219405/_0_  , \g219406/_0_  , \g219407/_0_  , \g219408/_0_  , \g219409/_0_  , \g219410/_0_  , \g219411/_0_  , \g219412/_0_  , \g219413/_0_  , \g219414/_0_  , \g219415/_0_  , \g219416/_0_  , \g219417/_0_  , \g219418/_0_  , \g219419/_0_  , \g219420/_0_  , \g219421/_0_  , \g219422/_0_  , \g219423/_0_  , \g219424/_0_  , \g219425/_0_  , \g219426/_0_  , \g219427/_0_  , \g219428/_0_  , \g219429/_0_  , \g219430/_0_  , \g219431/_0_  , \g219432/_0_  , \g219433/_0_  , \g219434/_0_  , \g219435/_0_  , \g219436/_0_  , \g219437/_0_  , \g219438/_0_  , \g219439/_0_  , \g219440/_0_  , \g219441/_0_  , \g219442/_0_  , \g219443/_0_  , \g219444/_0_  , \g219445/_0_  , \g219446/_0_  , \g219447/_0_  , \g219449/_0_  , \g219450/_0_  , \g219451/_0_  , \g219452/_0_  , \g219453/_0_  , \g219454/_0_  , \g219455/_0_  , \g219456/_0_  , \g219457/_0_  , \g219458/_0_  , \g219464/u3_syn_7  , \g219496/u3_syn_4  , \g219512/u3_syn_4  , \g219526/u3_syn_4  , \g219549/u3_syn_4  , \g219571/u3_syn_4  , \g219588/u3_syn_4  , \g219603/u3_syn_4  , \g219621/u3_syn_4  , \g219636/_3_  , \g219652/u3_syn_4  , \g219676/_3_  , \g219686/_0_  , \g219689/_0_  , \g219694/_3_  , \g220062/_0_  , \g220068/_0_  , \g220069/_0_  , \g220072/_0_  , \g220084/_0_  , \g220149/_0_  , \g220162/_0_  , \g220317/_0_  , \g220360/_2_  , \g220368/_2_  , \g220369/_0_  , \g220370/_0_  , \g220371/_0_  , \g220372/_0_  , \g220376/_0_  , \g220390/_0_  , \g220395/_0_  , \g220499/_0_  , \g220500/_0_  , \g220501/_0_  , \g220502/_0_  , \g220503/_0_  , \g220504/_0_  , \g220505/_0_  , \g220506/_0_  , \g220507/_0_  , \g220508/_0_  , \g220509/_0_  , \g220510/_0_  , \g220511/_0_  , \g220512/_0_  , \g220513/_0_  , \g220514/_0_  , \g220515/_0_  , \g220516/_0_  , \g220517/_0_  , \g220518/_0_  , \g220519/_0_  , \g220520/_0_  , \g220521/_0_  , \g220522/_0_  , \g220523/_0_  , \g220524/_0_  , \g220525/_0_  , \g220526/_0_  , \g220527/_0_  , \g220528/_0_  , \g220529/_0_  , \g220530/_0_  , \g220531/_0_  , \g220532/_0_  , \g220533/_0_  , \g220534/_0_  , \g220535/_0_  , \g220557/_0_  , \g220558/_0_  , \g220559/_0_  , \g220560/_0_  , \g220561/_0_  , \g220562/_0_  , \g220563/_0_  , \g220564/_0_  , \g220565/_0_  , \g220566/_0_  , \g220567/_0_  , \g220568/_0_  , \g220569/_0_  , \g220570/_0_  , \g220571/_0_  , \g220572/_0_  , \g220573/_0_  , \g220574/_0_  , \g220575/_0_  , \g220576/_0_  , \g220577/_0_  , \g220578/_0_  , \g220579/_0_  , \g220580/_0_  , \g220581/_0_  , \g220582/_0_  , \g220583/_0_  , \g220584/_0_  , \g220585/_0_  , \g220586/_0_  , \g220587/_0_  , \g220588/_0_  , \g220589/_0_  , \g220590/_0_  , \g220591/_0_  , \g220592/_0_  , \g220593/_0_  , \g220594/_0_  , \g220595/_0_  , \g220596/_0_  , \g220597/_0_  , \g220598/_0_  , \g220599/_0_  , \g220600/_0_  , \g220601/_0_  , \g220602/_0_  , \g220603/_0_  , \g220604/_0_  , \g220605/_0_  , \g220606/_0_  , \g220607/_0_  , \g220608/_0_  , \g220609/_0_  , \g220610/_0_  , \g220611/_0_  , \g220612/_0_  , \g220613/_0_  , \g220614/_0_  , \g220615/_0_  , \g220616/_0_  , \g220617/_0_  , \g220618/_0_  , \g220619/_0_  , \g220620/_0_  , \g220621/_0_  , \g220622/_0_  , \g220623/_0_  , \g220624/_0_  , \g220625/_0_  , \g220626/_0_  , \g220627/_0_  , \g220628/_0_  , \g220629/_0_  , \g220630/_0_  , \g220631/_0_  , \g220632/_0_  , \g220633/_0_  , \g220634/_0_  , \g220635/_0_  , \g220636/_0_  , \g220637/_0_  , \g220638/_0_  , \g220639/_0_  , \g220640/_0_  , \g220641/_0_  , \g220642/_0_  , \g220643/_0_  , \g220644/_0_  , \g220645/_0_  , \g220646/_0_  , \g220647/_0_  , \g220648/_0_  , \g220649/_0_  , \g220650/_0_  , \g220651/_0_  , \g220652/_0_  , \g220653/_0_  , \g220654/_0_  , \g220655/_0_  , \g220656/_0_  , \g220657/_0_  , \g220658/_0_  , \g220659/_0_  , \g220660/_0_  , \g220661/_0_  , \g220662/_0_  , \g220663/_0_  , \g220664/_0_  , \g220665/_0_  , \g220666/_0_  , \g220674/_0_  , \g220679/u3_syn_7  , \g220711/u3_syn_4  , \g220726/u3_syn_4  , \g220739/u3_syn_4  , \g220751/u3_syn_4  , \g220759/u3_syn_4  , \g220773/u3_syn_4  , \g220782/u3_syn_4  , \g220805/u3_syn_4  , \g220828/u3_syn_4  , \g220921/_0_  , \g220930/u3_syn_4  , \g220949/_3_  , \g220994/_3_  , \g221207/_0_  , \g221213/_0_  , \g221223/_0_  , \g221224/_0_  , \g221225/_0_  , \g221226/_0_  , \g221231/_0_  , \g221232/_0_  , \g221234/_0_  , \g221235/_0_  , \g221246/_2_  , \g221249/_2_  , \g221265/_0_  , \g221287/_0_  , \g221325/_0_  , \g221326/_0_  , \g221447/_0_  , \g221449/_0_  , \g221452/_0_  , \g221469/_0_  , \g221473/_0_  , \g221503/_0_  , \g221510/_0_  , \g221512/_0_  , \g221516/_0_  , \g221517/_0_  , \g221524/_0_  , \g221530/_0_  , \g221592/_0_  , \g221593/_0_  , \g221634/u3_syn_4  , \g221669/u3_syn_4  , \g221789/u3_syn_4  , \g221813/u3_syn_4  , \g221829/u3_syn_4  , \g221861/u3_syn_4  , \g221876/_0_  , \g221935/_0_  , \g221944/_3_  , \g230200/_0_  , \g230201/_0_  , \g230205/_0_  , \g230295/_0_  , \g230297/_0_  , \g230298/_0_  , \g230300/_0_  , \g230302/_0_  , \g230303/_0_  , \g230343/_0_  , \g230368/_0_  , \g230511/_0_  , \g230531/_0_  , \g230635/_2_  , \g230661/_0_  , \g230715/_1__syn_2  , \g230731/_0_  , \g230766/_0_  , \g230784/_0_  , \g230785/_0_  , \g230786/_0_  , \g230787/_0_  , \g230797/_0_  , \g230798/_0_  , \g230803/_0_  , \g230804/_00_  , \g230805/_00_  , \g230806/_00_  , \g230807/_00_  , \g230808/_00_  , \g230809/_00_  , \g230815/_0_  , \g230816/_2_  , \g230817/_2_  , \g230829/_0_  , \g230834/_0_  , \g230835/_0_  , \g230836/_0_  , \g230837/_0_  , \g230844/_0_  , \g230863/_3_  , \g230864/_3_  , \g230870/_0_  , \g230988/_3_  , \g231010/_3_  , \g231016/_3_  , \g231042/_3_  , \g231471/_0_  , \g231472/_0_  , \g231476/_3_  , \g231480/_3_  , \g231484/_3_  , \g231504/_0_  , \g231532/_0_  , \g231542/_0_  , \g231560/_1_  , \g231578/_1_  , \g231580/_0_  , \g231590/_1__syn_2  , \g231615/_0_  , \g231623/_1_  , \g231634/_2_  , \g231635/_0_  , \g231638/_2_  , \g231640/_0_  , \g231653/_2_  , \g231787/_0_  , \g231931/_0_  , \g231939/_3_  , \g231940/_0_  , \g231951/_0_  , \g231955/_0_  , \g231956/_0_  , \g231959/_2_  , \g231960/_0_  , \g231964/_0_  , \g231965/_0_  , \g231975/_0_  , \g231986/_1_  , \g231987/_1_  , \g231989/_1_  , \g231990/_1_  , \g231991/_0_  , \g231992/_0_  , \g231995/_0_  , \g231998/_0_  , \g231999/_0_  , \g232002/_3_  , \g232035/u3_syn_4  , \g232038/u3_syn_4  , \g232046/u3_syn_4  , \g232054/u3_syn_4  , \g232062/u3_syn_4  , \g232070/u3_syn_4  , \g232078/u3_syn_4  , \g232079/u3_syn_4  , \g232087/u3_syn_4  , \g232096/u3_syn_4  , \g232104/u3_syn_4  , \g232112/u3_syn_4  , \g232120/u3_syn_4  , \g232128/u3_syn_4  , \g232136/u3_syn_4  , \g232144/u3_syn_4  , \g232152/u3_syn_4  , \g232161/u3_syn_4  , \g232169/u3_syn_4  , \g232177/u3_syn_4  , \g232185/u3_syn_4  , \g232186/u3_syn_4  , \g232194/u3_syn_4  , \g232202/u3_syn_4  , \g232210/u3_syn_4  , \g232218/u3_syn_4  , \g232226/u3_syn_4  , \g232234/u3_syn_4  , \g232242/u3_syn_4  , \g232251/u3_syn_4  , \g232259/u3_syn_4  , \g232267/u3_syn_4  , \g232275/u3_syn_4  , \g232283/u3_syn_4  , \g232291/u3_syn_4  , \g232299/u3_syn_4  , \g232307/u3_syn_4  , \g232315/u3_syn_4  , \g232324/u3_syn_4  , \g232332/u3_syn_4  , \g232341/u3_syn_4  , \g232349/u3_syn_4  , \g232357/u3_syn_4  , \g232366/u3_syn_4  , \g232374/u3_syn_4  , \g232382/u3_syn_4  , \g232390/u3_syn_4  , \g232398/u3_syn_4  , \g232406/u3_syn_4  , \g232414/u3_syn_4  , \g232422/u3_syn_4  , \g232427/u3_syn_4  , \g232431/u3_syn_4  , \g232439/u3_syn_4  , \g232444/u3_syn_4  , \g232452/u3_syn_4  , \g232461/u3_syn_4  , \g232471/u3_syn_4  , \g232479/u3_syn_4  , \g232487/u3_syn_4  , \g232495/u3_syn_4  , \g232503/u3_syn_4  , \g232506/u3_syn_4  , \g232514/u3_syn_4  , \g232527/u3_syn_4  , \g232530/u3_syn_4  , \g232536/u3_syn_4  , \g232544/u3_syn_4  , \g232551/u3_syn_4  , \g232557/u3_syn_4  , \g232568/u3_syn_4  , \g232576/u3_syn_4  , \g232585/u3_syn_4  , \g232593/u3_syn_4  , \g232597/u3_syn_4  , \g232609/u3_syn_4  , \g232617/u3_syn_4  , \g232625/u3_syn_4  , \g232633/u3_syn_4  , \g232641/u3_syn_4  , \g232649/u3_syn_4  , \g232657/u3_syn_4  , \g232665/u3_syn_4  , \g232673/u3_syn_4  , \g232681/u3_syn_4  , \g232689/u3_syn_4  , \g232697/u3_syn_4  , \g232705/u3_syn_4  , \g232713/u3_syn_4  , \g232717/u3_syn_4  , \g232729/u3_syn_4  , \g232737/u3_syn_4  , \g232745/u3_syn_4  , \g232749/u3_syn_4  , \g232761/u3_syn_4  , \g232768/u3_syn_4  , \g232777/u3_syn_4  , \g232785/u3_syn_4  , \g232793/u3_syn_4  , \g232801/u3_syn_4  , \g232809/u3_syn_4  , \g232815/u3_syn_4  , \g232823/u3_syn_4  , \g232833/u3_syn_4  , \g232841/u3_syn_4  , \g232846/u3_syn_4  , \g232851/u3_syn_4  , \g232865/u3_syn_4  , \g232873/u3_syn_4  , \g232881/u3_syn_4  , \g232882/u3_syn_4  , \g232895/u3_syn_4  , \g232904/u3_syn_4  , \g232913/u3_syn_4  , \g232921/u3_syn_4  , \g232928/u3_syn_4  , \g232934/u3_syn_4  , \g232945/u3_syn_4  , \g232953/u3_syn_4  , \g232954/u3_syn_4  , \g232969/u3_syn_4  , \g232977/u3_syn_4  , \g232981/u3_syn_4  , \g232993/u3_syn_4  , \g232995/u3_syn_4  , \g233009/u3_syn_4  , \g233017/u3_syn_4  , \g233025/u3_syn_4  , \g233033/u3_syn_4  , \g233041/u3_syn_4  , \g233047/u3_syn_4  , \g233057/u3_syn_4  , \g233065/u3_syn_4  , \g233073/u3_syn_4  , \g233081/u3_syn_4  , \g233087/u3_syn_4  , \g233097/u3_syn_4  , \g233105/u3_syn_4  , \g233113/u3_syn_4  , \g233121/u3_syn_4  , \g233128/u3_syn_4  , \g233134/u3_syn_4  , \g233144/u3_syn_4  , \g233153/u3_syn_4  , \g233161/u3_syn_4  , \g233169/u3_syn_4  , \g233177/u3_syn_4  , \g233185/u3_syn_4  , \g233193/u3_syn_4  , \g233201/u3_syn_4  , \g233209/u3_syn_4  , \g233217/u3_syn_4  , \g233219/u3_syn_4  , \g233229/u3_syn_4  , \g233241/u3_syn_4  , \g233249/u3_syn_4  , \g233257/u3_syn_4  , \g233265/u3_syn_4  , \g233273/u3_syn_4  , \g233281/u3_syn_4  , \g233289/u3_syn_4  , \g233297/u3_syn_4  , \g233305/u3_syn_4  , \g233313/u3_syn_4  , \g233321/u3_syn_4  , \g233329/u3_syn_4  , \g233337/u3_syn_4  , \g233345/u3_syn_4  , \g233353/u3_syn_4  , \g233361/u3_syn_4  , \g233369/u3_syn_4  , \g233377/u3_syn_4  , \g233382/u3_syn_4  , \g233392/u3_syn_4  , \g233394/u3_syn_4  , \g233409/u3_syn_4  , \g233417/u3_syn_4  , \g233425/u3_syn_4  , \g233433/u3_syn_4  , \g233441/u3_syn_4  , \g233449/u3_syn_4  , \g233453/u3_syn_4  , \g233465/u3_syn_4  , \g233473/u3_syn_4  , \g233481/u3_syn_4  , \g233489/u3_syn_4  , \g233497/u3_syn_4  , \g233505/u3_syn_4  , \g233513/u3_syn_4  , \g233516/u3_syn_4  , \g233529/u3_syn_4  , \g233531/u3_syn_4  , \g233546/u3_syn_4  , \g233554/u3_syn_4  , \g233562/u3_syn_4  , \g233570/u3_syn_4  , \g233578/u3_syn_4  , \g233586/u3_syn_4  , \g233594/u3_syn_4  , \g233602/u3_syn_4  , \g233603/u3_syn_4  , \g233618/u3_syn_4  , \g233626/u3_syn_4  , \g233634/u3_syn_4  , \g233642/u3_syn_4  , \g233650/u3_syn_4  , \g233658/u3_syn_4  , \g233666/u3_syn_4  , \g233674/u3_syn_4  , \g233682/u3_syn_4  , \g233690/u3_syn_4  , \g233698/u3_syn_4  , \g233706/u3_syn_4  , \g233714/u3_syn_4  , \g233722/u3_syn_4  , \g233730/u3_syn_4  , \g233738/u3_syn_4  , \g233746/u3_syn_4  , \g233754/u3_syn_4  , \g233762/u3_syn_4  , \g233770/u3_syn_4  , \g233778/u3_syn_4  , \g233783/u3_syn_4  , \g233794/u3_syn_4  , \g233802/u3_syn_4  , \g233806/u3_syn_4  , \g233818/u3_syn_4  , \g233826/u3_syn_4  , \g233828/u3_syn_4  , \g233838/u3_syn_4  , \g233850/u3_syn_4  , \g233858/u3_syn_4  , \g233860/u3_syn_4  , \g233870/u3_syn_4  , \g233881/u3_syn_4  , \g233890/u3_syn_4  , \g233899/u3_syn_4  , \g233908/u3_syn_4  , \g233917/u3_syn_4  , \g233919/u3_syn_4  , \g233927/u3_syn_4  , \g233935/u3_syn_4  , \g233943/u3_syn_4  , \g233945/u3_syn_4  , \g233953/u3_syn_4  , \g233961/u3_syn_4  , \g233969/u3_syn_4  , \g233977/u3_syn_4  , \g233985/u3_syn_4  , \g233993/u3_syn_4  , \g234001/u3_syn_4  , \g234008/u3_syn_4  , \g234009/u3_syn_4  , \g234024/u3_syn_4  , \g234032/u3_syn_4  , \g234038/u3_syn_4  , \g234056/u3_syn_4  , \g234063/u3_syn_4  , \g234071/u3_syn_4  , \g234079/u3_syn_4  , \g234098/u3_syn_4  , \g234106/u3_syn_4  , \g234114/u3_syn_4  , \g234122/u3_syn_4  , \g234130/u3_syn_4  , \g234138/u3_syn_4  , \g234145/u3_syn_4  , \g234156/u3_syn_4  , \g234162/u3_syn_4  , \g234171/u3_syn_4  , \g234183/u3_syn_4  , \g234248/u3_syn_4  , \g234265/u3_syn_4  , \g234273/u3_syn_4  , \g234281/u3_syn_4  , \g234289/u3_syn_4  , \g234297/u3_syn_4  , \g234306/u3_syn_4  , \g234314/u3_syn_4  , \g234322/u3_syn_4  , \g234331/u3_syn_4  , \g234339/u3_syn_4  , \g234347/u3_syn_4  , \g234355/u3_syn_4  , \g234363/u3_syn_4  , \g234371/u3_syn_4  , \g234379/u3_syn_4  , \g234387/u3_syn_4  , \g234395/u3_syn_4  , \g234403/u3_syn_4  , \g234411/u3_syn_4  , \g234419/u3_syn_4  , \g234427/u3_syn_4  , \g234435/u3_syn_4  , \g234443/u3_syn_4  , \g234451/u3_syn_4  , \g234459/u3_syn_4  , \g234467/u3_syn_4  , \g234475/u3_syn_4  , \g234483/u3_syn_4  , \g234491/u3_syn_4  , \g234499/u3_syn_4  , \g234507/u3_syn_4  , \g234515/u3_syn_4  , \g234523/u3_syn_4  , \g234531/u3_syn_4  , \g234539/u3_syn_4  , \g234547/u3_syn_4  , \g234555/u3_syn_4  , \g234563/u3_syn_4  , \g234571/u3_syn_4  , \g234579/u3_syn_4  , \g234587/u3_syn_4  , \g234595/u3_syn_4  , \g234604/u3_syn_4  , \g234612/u3_syn_4  , \g234620/u3_syn_4  , \g234628/u3_syn_4  , \g234636/u3_syn_4  , \g234644/u3_syn_4  , \g234652/u3_syn_4  , \g234660/u3_syn_4  , \g234668/u3_syn_4  , \g234676/u3_syn_4  , \g234684/u3_syn_4  , \g234692/u3_syn_4  , \g234700/u3_syn_4  , \g234708/u3_syn_4  , \g234716/u3_syn_4  , \g234725/u3_syn_4  , \g234733/u3_syn_4  , \g234741/u3_syn_4  , \g234749/u3_syn_4  , \g234757/u3_syn_4  , \g234765/u3_syn_4  , \g234773/u3_syn_4  , \g234781/u3_syn_4  , \g234789/u3_syn_4  , \g234798/u3_syn_4  , \g234806/u3_syn_4  , \g234814/u3_syn_4  , \g234822/u3_syn_4  , \g234830/u3_syn_4  , \g234838/u3_syn_4  , \g235911/u3_syn_4  , \g235912/u3_syn_4  , \g235920/u3_syn_4  , \g235928/u3_syn_4  , \g235936/u3_syn_4  , \g235944/u3_syn_4  , \g235952/u3_syn_4  , \g235960/u3_syn_4  , \g235968/u3_syn_4  , \g235976/u3_syn_4  , \g235984/u3_syn_4  , \g235992/u3_syn_4  , \g236000/u3_syn_4  , \g236008/u3_syn_4  , \g236016/u3_syn_4  , \g236021/u3_syn_4  , \g236025/u3_syn_4  , \g236033/u3_syn_4  , \g236041/u3_syn_4  , \g236049/u3_syn_4  , \g236057/u3_syn_4  , \g236065/u3_syn_4  , \g236073/u3_syn_4  , \g236081/u3_syn_4  , \g236089/u3_syn_4  , \g236097/u3_syn_4  , \g236105/u3_syn_4  , \g236113/u3_syn_4  , \g236121/u3_syn_4  , \g236129/u3_syn_4  , \g236137/u3_syn_4  , \g236145/u3_syn_4  , \g236153/u3_syn_4  , \g236161/u3_syn_4  , \g236169/u3_syn_4  , \g236177/u3_syn_4  , \g236185/u3_syn_4  , \g236193/u3_syn_4  , \g236196/u3_syn_4  , \g236198/u3_syn_4  , \g236203/u3_syn_4  , \g236211/u3_syn_4  , \g236219/u3_syn_4  , \g236220/u3_syn_4  , \g236229/u3_syn_4  , \g236232/u3_syn_4  , \g236238/u3_syn_4  , \g236246/u3_syn_4  , \g236255/u3_syn_4  , \g236263/u3_syn_4  , \g236271/u3_syn_4  , \g236275/u3_syn_4  , \g236280/u3_syn_4  , \g236288/u3_syn_4  , \g236296/u3_syn_4  , \g236304/u3_syn_4  , \g236305/u3_syn_4  , \g236306/u3_syn_4  , \g236315/u3_syn_4  , \g236323/u3_syn_4  , \g236331/u3_syn_4  , \g236334/u3_syn_4  , \g236340/u3_syn_4  , \g236348/u3_syn_4  , \g236357/u3_syn_4  , \g236359/u3_syn_4  , \g236367/u3_syn_4  , \g236374/u3_syn_4  , \g236376/u3_syn_4  , \g236377/u3_syn_4  , \g236385/u3_syn_4  , \g236393/u3_syn_4  , \g236402/u3_syn_4  , \g236410/u3_syn_4  , \g236419/u3_syn_4  , \g236427/u3_syn_4  , \g236433/u3_syn_4  , \g236436/u3_syn_4  , \g236444/u3_syn_4  , \g236452/u3_syn_4  , \g236460/u3_syn_4  , \g236468/u3_syn_4  , \g236476/u3_syn_4  , \g236484/u3_syn_4  , \g236492/u3_syn_4  , \g236500/u3_syn_4  , \g236508/u3_syn_4  , \g236516/u3_syn_4  , \g236518/u3_syn_4  , \g236525/u3_syn_4  , \g236533/u3_syn_4  , \g236542/u3_syn_4  , \g236550/u3_syn_4  , \g236559/u3_syn_4  , \g236567/u3_syn_4  , \g236575/u3_syn_4  , \g236583/u3_syn_4  , \g236591/u3_syn_4  , \g236599/u3_syn_4  , \g236607/u3_syn_4  , \g236608/u3_syn_4  , \g236616/u3_syn_4  , \g236624/u3_syn_4  , \g236632/u3_syn_4  , \g236640/u3_syn_4  , \g236647/u3_syn_4  , \g236649/u3_syn_4  , \g236659/u3_syn_4  , \g236671/u3_syn_4  , \g236677/u3_syn_4  , \g236688/u3_syn_4  , \g236696/u3_syn_4  , \g236705/u3_syn_4  , \g236712/u3_syn_4  , \g236718/u3_syn_4  , \g236729/u3_syn_4  , \g236732/u3_syn_4  , \g236745/u3_syn_4  , \g236753/u3_syn_4  , \g236761/u3_syn_4  , \g236769/u3_syn_4  , \g236777/u3_syn_4  , \g236779/u3_syn_4  , \g236788/u3_syn_4  , \g236800/u3_syn_4  , \g236802/u3_syn_4  , \g236805/u3_syn_4  , \g236813/u3_syn_4  , \g236825/u3_syn_4  , \g236829/u3_syn_4  , \g236837/u3_syn_4  , \g236849/u3_syn_4  , \g236854/u3_syn_4  , \g236860/u3_syn_4  , \g236872/u3_syn_4  , \g236878/u3_syn_4  , \g236884/u3_syn_4  , \g236896/u3_syn_4  , \g236903/u3_syn_4  , \g236908/u3_syn_4  , \g236920/u3_syn_4  , \g236930/u3_syn_4  , \g236939/u3_syn_4  , \g236947/u3_syn_4  , \g236949/u3_syn_4  , \g236956/u3_syn_4  , \g236962/u3_syn_4  , \g236965/u3_syn_4  , \g236980/u3_syn_4  , \g236988/u3_syn_4  , \g236989/u3_syn_4  , \g237004/u3_syn_4  , \g237005/u3_syn_4  , \g237020/u3_syn_4  , \g237021/u3_syn_4  , \g237033/u3_syn_4  , \g237044/u3_syn_4  , \g237045/u3_syn_4  , \g237056/u3_syn_4  , \g237068/u3_syn_4  , \g237076/u3_syn_4  , \g237084/u3_syn_4  , \g237092/u3_syn_4  , \g237095/u3_syn_4  , \g237107/u3_syn_4  , \g237110/u3_syn_4  , \g237119/u3_syn_4  , \g237131/u3_syn_4  , \g237135/u3_syn_4  , \g237148/u3_syn_4  , \g237152/u3_syn_4  , \g237165/u3_syn_4  , \g237168/u3_syn_4  , \g237180/u3_syn_4  , \g237185/u3_syn_4  , \g237192/u3_syn_4  , \g237204/u3_syn_4  , \g237209/u3_syn_4  , \g237215/u3_syn_4  , \g237229/u3_syn_4  , \g237231/u3_syn_4  , \g237245/u3_syn_4  , \g237251/u3_syn_4  , \g237260/u3_syn_4  , \g237262/u3_syn_4  , \g237277/u3_syn_4  , \g237281/u3_syn_4  , \g237293/u3_syn_4  , \g237294/u3_syn_4  , \g237310/u3_syn_4  , \g237311/u3_syn_4  , \g237323/u3_syn_4  , \g237334/u3_syn_4  , \g237342/u3_syn_4  , \g237350/u3_syn_4  , \g237353/u3_syn_4  , \g237359/u3_syn_4  , \g237367/u3_syn_4  , \g237368/u3_syn_4  , \g237378/u3_syn_4  , \g237391/u3_syn_4  , \g237392/u3_syn_4  , \g237403/u3_syn_4  , \g237415/u3_syn_4  , \g237417/u3_syn_4  , \g237431/u3_syn_4  , \g237439/u3_syn_4  , \g237440/u3_syn_4  , \g237454/u3_syn_4  , \g237457/u3_syn_4  , \g237472/u3_syn_4  , \g237480/u3_syn_4  , \g237488/u3_syn_4  , \g237496/u3_syn_4  , \g237499/u3_syn_4  , \g237512/u3_syn_4  , \g237515/u3_syn_4  , \g237525/u3_syn_4  , \g237529/u3_syn_4  , \g237535/u3_syn_4  , \g237541/u3_syn_4  , \g237553/u3_syn_4  , \g237561/u3_syn_4  , \g237569/u3_syn_4  , \g237575/u3_syn_4  , \g237578/u3_syn_4  , \g237581/u3_syn_4  , \g237591/u3_syn_4  , \g237602/u3_syn_4  , \g237610/u3_syn_4  , \g237617/u3_syn_4  , \g237623/u3_syn_4  , \g237633/u3_syn_4  , \g237635/u3_syn_4  , \g237648/u3_syn_4  , \g237658/u3_syn_4  , \g237659/u3_syn_4  , \g237660/u3_syn_4  , \g237668/u3_syn_4  , \g237675/u3_syn_4  , \g237684/u3_syn_4  , \g237692/u3_syn_4  , \g237693/u3_syn_4  , \g237705/u3_syn_4  , \g237716/u3_syn_4  , \g237717/u3_syn_4  , \g237729/u3_syn_4  , \g237740/u3_syn_4  , \g237741/u3_syn_4  , \g237756/u3_syn_4  , \g237764/u3_syn_4  , \g237768/u3_syn_4  , \g237780/u3_syn_4  , \g237782/u3_syn_4  , \g237792/u3_syn_4  , \g237804/u3_syn_4  , \g237812/u3_syn_4  , \g237820/u3_syn_4  , \g237828/u3_syn_4  , \g237836/u3_syn_4  , \g237844/u3_syn_4  , \g237852/u3_syn_4  , \g237860/u3_syn_4  , \g237868/u3_syn_4  , \g237876/u3_syn_4  , \g237884/u3_syn_4  , \g237888/u3_syn_4  , \g237895/u3_syn_4  , \g237907/u3_syn_4  , \g237916/u3_syn_4  , \g237924/u3_syn_4  , \g237931/u3_syn_4  , \g237940/u3_syn_4  , \g237949/u3_syn_4  , \g237950/u3_syn_4  , \g237955/u3_syn_4  , \g237961/u3_syn_4  , \g237965/u3_syn_4  , \g237975/u3_syn_4  , \g237983/u3_syn_4  , \g237989/u3_syn_4  , \g237999/u3_syn_4  , \g238007/u3_syn_4  , \g238015/u3_syn_4  , \g238017/u3_syn_4  , \g238033/u3_syn_4  , \g238035/u3_syn_4  , \g238049/u3_syn_4  , \g238057/u3_syn_4  , \g238065/u3_syn_4  , \g238072/u3_syn_4  , \g238081/u3_syn_4  , \g238082/u3_syn_4  , \g238097/u3_syn_4  , \g238105/u3_syn_4  , \g238113/u3_syn_4  , \g238114/u3_syn_4  , \g238129/u3_syn_4  , \g238137/u3_syn_4  , \g238145/u3_syn_4  , \g238153/u3_syn_4  , \g238161/u3_syn_4  , \g238163/u3_syn_4  , \g238177/u3_syn_4  , \g238179/u3_syn_4  , \g238194/u3_syn_4  , \g238197/u3_syn_4  , \g238209/u3_syn_4  , \g238213/u3_syn_4  , \g238225/u3_syn_4  , \g238229/u3_syn_4  , \g238237/u3_syn_4  , \g238250/u3_syn_4  , \g238257/u3_syn_4  , \g238263/u3_syn_4  , \g238269/u3_syn_4  , \g238282/u3_syn_4  , \g238285/u3_syn_4  , \g238298/u3_syn_4  , \g238301/u3_syn_4  , \g238314/u3_syn_4  , \g238316/u3_syn_4  , \g238329/u3_syn_4  , \g238338/u3_syn_4  , \g238346/u3_syn_4  , \g238351/u3_syn_4  , \g238356/u3_syn_4  , \g238368/u3_syn_4  , \g238378/u3_syn_4  , \g238386/u3_syn_4  , \g238394/u3_syn_4  , \g238402/u3_syn_4  , \g238409/u3_syn_4  , \g238412/u3_syn_4  , \g238427/u3_syn_4  , \g238429/u3_syn_4  , \g238443/u3_syn_4  , \g238448/u3_syn_4  , \g238457/u3_syn_4  , \g238460/u3_syn_4  , \g238472/u3_syn_4  , \g238484/u3_syn_4  , \g238492/u3_syn_4  , \g238500/u3_syn_4  , \g238505/u3_syn_4  , \g238516/u3_syn_4  , \g238524/u3_syn_4  , \g238532/u3_syn_4  , \g238534/u3_syn_4  , \g238544/u3_syn_4  , \g238549/u3_syn_4  , \g238550/u3_syn_4  , \g238565/u3_syn_4  , \g238566/u3_syn_4  , \g238582/u3_syn_4  , \g238583/u3_syn_4  , \g238594/u3_syn_4  , \g238606/u3_syn_4  , \g238614/u3_syn_4  , \g238615/u3_syn_4  , \g238619/u3_syn_4  , \g238631/u3_syn_4  , \g238639/u3_syn_4  , \g238647/u3_syn_4  , \g238649/u3_syn_4  , \g238659/u3_syn_4  , \g238670/u3_syn_4  , \g238671/u3_syn_4  , \g238680/u3_syn_4  , \g238688/u3_syn_4  , \g238691/u3_syn_4  , \g238696/u3_syn_4  , \g238705/u3_syn_4  , \g238708/u3_syn_4  , \g238721/u3_syn_4  , \g238724/u3_syn_4  , \g238736/u3_syn_4  , \g238745/u3_syn_4  , \g238753/u3_syn_4  , \g238757/u3_syn_4  , \g238764/u3_syn_4  , \g238776/u3_syn_4  , \g238781/u3_syn_4  , \g238787/u3_syn_4  , \g238799/u3_syn_4  , \g238807/u3_syn_4  , \g238811/u3_syn_4  , \g238824/u3_syn_4  , \g238830/u3_syn_4  , \g238841/u3_syn_4  , \g238843/u3_syn_4  , \g238855/u3_syn_4  , \g238859/u3_syn_4  , \g238863/u3_syn_4  , \g238868/u3_syn_4  , \g238880/u3_syn_4  , \g238888/u3_syn_4  , \g238892/u3_syn_4  , \g238903/u3_syn_4  , \g238911/u3_syn_4  , \g238915/u3_syn_4  , \g238927/u3_syn_4  , \g238937/u3_syn_4  , \g238945/u3_syn_4  , \g238953/u3_syn_4  , \g238961/u3_syn_4  , \g238970/u3_syn_4  , \g238971/u3_syn_4  , \g238983/u3_syn_4  , \g238994/u3_syn_4  , \g239002/u3_syn_4  , \g239009/u3_syn_4  , \g239015/u3_syn_4  , \g239025/u3_syn_4  , \g239030/u3_syn_4  , \g239041/u3_syn_4  , \g239048/u3_syn_4  , \g239053/u3_syn_4  , \g239065/u3_syn_4  , \g239073/u3_syn_4  , \g239081/u3_syn_4  , \g239082/u3_syn_4  , \g239093/u3_syn_4  , \g239105/u3_syn_4  , \g239108/u3_syn_4  , \g239117/u3_syn_4  , \g239129/u3_syn_4  , \g239137/u3_syn_4  , \g239139/u3_syn_4  , \g239148/u3_syn_4  , \g239160/u3_syn_4  , \g239162/u3_syn_4  , \g239172/u3_syn_4  , \g239184/u3_syn_4  , \g239187/u3_syn_4  , \g239189/u3_syn_4  , \g239201/u3_syn_4  , \g239208/u3_syn_4  , \g239217/u3_syn_4  , \g239219/u3_syn_4  , \g239226/u3_syn_4  , \g239234/u3_syn_4  , \g239242/u3_syn_4  , \g239246/u3_syn_4  , \g239257/u3_syn_4  , \g239258/u3_syn_4  , \g239263/u3_syn_4  , \g239275/u3_syn_4  , \g239277/u3_syn_4  , \g239291/u3_syn_4  , \g239296/u3_syn_4  , \g239308/u3_syn_4  , \g239311/u3_syn_4  , \g239322/u3_syn_4  , \g239329/u3_syn_4  , \g239338/u3_syn_4  , \g239339/u3_syn_4  , \g239346/u3_syn_4  , \g239351/u3_syn_4  , \g239363/u3_syn_4  , \g239370/u3_syn_4  , \g239375/u3_syn_4  , \g239387/u3_syn_4  , \g239395/u3_syn_4  , \g239418/u3_syn_4  , \g239439/u3_syn_4  , \g239442/u3_syn_4  , \g239454/u3_syn_4  , \g239464/u3_syn_4  , \g239470/u3_syn_4  , \g239481/u3_syn_4  , \g239487/u3_syn_4  , \g239497/u3_syn_4  , \g239520/u3_syn_4  , \g239532/u3_syn_4  , \g239543/u3_syn_4  , \g239551/u3_syn_4  , \g239552/u3_syn_4  , \g239567/u3_syn_4  , \g239575/u3_syn_4  , \g239579/u3_syn_4  , \g239592/u3_syn_4  , \g239594/u3_syn_4  , \g239608/u3_syn_4  , \g239626/u3_syn_4  , \g239634/u3_syn_4  , \g239646/u3_syn_4  , \g239649/u3_syn_4  , \g239657/u3_syn_4  , \g239670/u3_syn_4  , \g239673/u3_syn_4  , \g239686/u3_syn_4  , \g239694/u3_syn_4  , \g239695/u3_syn_4  , \g239701/u3_syn_4  , \g239705/u3_syn_4  , \g239709/u3_syn_4  , \g239715/u3_syn_4  , \g239717/u3_syn_4  , \g239726/u3_syn_4  , \g239734/u3_syn_4  , \g239735/u3_syn_4  , \g239743/u3_syn_4  , \g239760/u3_syn_4  , \g239768/u3_syn_4  , \g239776/u3_syn_4  , \g239784/u3_syn_4  , \g239793/u3_syn_4  , \g239801/u3_syn_4  , \g239817/u3_syn_4  , \g239818/u3_syn_4  , \g239848/u3_syn_4  , \g239856/u3_syn_4  , \g239872/u3_syn_4  , \g239880/u3_syn_4  , \g239888/u3_syn_4  , \g239896/u3_syn_4  , \g239904/u3_syn_4  , \g239912/u3_syn_4  , \g239920/u3_syn_4  , \g239928/u3_syn_4  , \g239936/u3_syn_4  , \g239951/u3_syn_4  , \g239963/u3_syn_4  , \g239979/u3_syn_4  , \g239986/u3_syn_4  , \g239999/u3_syn_4  , \g240000/u3_syn_4  , \g240008/u3_syn_4  , \g240012/u3_syn_4  , \g240018/u3_syn_4  , \g240026/u3_syn_4  , \g240034/u3_syn_4  , \g240042/u3_syn_4  , \g240050/u3_syn_4  , \g240074/u3_syn_4  , \g240091/u3_syn_4  , \g240122/u3_syn_4  , \g240147/u3_syn_4  , \g240209/u3_syn_4  , \g240219/u3_syn_4  , \g240259/u3_syn_4  , \g240334/u3_syn_4  , \g240406/u3_syn_4  , \g240416/u3_syn_4  , \g240424/u3_syn_4  , \g240432/u3_syn_4  , \g240440/u3_syn_4  , \g240448/u3_syn_4  , \g240456/u3_syn_4  , \g240464/u3_syn_4  , \g240472/u3_syn_4  , \g240480/u3_syn_4  , \g240488/u3_syn_4  , \g240496/u3_syn_4  , \g240504/u3_syn_4  , \g240512/u3_syn_4  , \g240520/u3_syn_4  , \g240530/u3_syn_4  , \g240538/u3_syn_4  , \g240547/u3_syn_4  , \g240555/u3_syn_4  , \g240563/u3_syn_4  , \g240571/u3_syn_4  , \g240579/u3_syn_4  , \g240587/u3_syn_4  , \g240595/u3_syn_4  , \g240603/u3_syn_4  , \g240611/u3_syn_4  , \g240619/u3_syn_4  , \g240627/u3_syn_4  , \g240635/u3_syn_4  , \g240643/u3_syn_4  , \g240651/u3_syn_4  , \g240659/u3_syn_4  , \g240667/u3_syn_4  , \g240675/u3_syn_4  , \g240683/u3_syn_4  , \g240691/u3_syn_4  , \g240699/u3_syn_4  , \g240707/u3_syn_4  , \g240715/u3_syn_4  , \g240723/u3_syn_4  , \g240731/u3_syn_4  , \g240739/u3_syn_4  , \g240747/u3_syn_4  , \g240755/u3_syn_4  , \g240763/u3_syn_4  , \g240771/u3_syn_4  , \g240779/u3_syn_4  , \g240787/u3_syn_4  , \g240795/u3_syn_4  , \g240803/u3_syn_4  , \g240811/u3_syn_4  , \g240819/u3_syn_4  , \g240827/u3_syn_4  , \g240835/u3_syn_4  , \g240843/u3_syn_4  , \g240851/u3_syn_4  , \g240859/u3_syn_4  , \g240867/u3_syn_4  , \g240875/u3_syn_4  , \g240883/u3_syn_4  , \g240891/u3_syn_4  , \g240899/u3_syn_4  , \g240907/u3_syn_4  , \g240915/u3_syn_4  , \g240923/u3_syn_4  , \g240931/u3_syn_4  , \g240939/u3_syn_4  , \g240947/u3_syn_4  , \g240955/u3_syn_4  , \g240963/u3_syn_4  , \g240971/u3_syn_4  , \g240979/u3_syn_4  , \g240987/u3_syn_4  , \g240995/u3_syn_4  , \g241003/u3_syn_4  , \g241011/u3_syn_4  , \g241019/u3_syn_4  , \g241027/u3_syn_4  , \g241036/u3_syn_4  , \g241044/u3_syn_4  , \g241052/u3_syn_4  , \g241060/u3_syn_4  , \g241068/u3_syn_4  , \g241076/u3_syn_4  , \g241084/u3_syn_4  , \g241092/u3_syn_4  , \g241100/u3_syn_4  , \g241108/u3_syn_4  , \g241116/u3_syn_4  , \g241124/u3_syn_4  , \g241132/u3_syn_4  , \g241140/u3_syn_4  , \g241148/u3_syn_4  , \g241156/u3_syn_4  , \g241164/u3_syn_4  , \g241172/u3_syn_4  , \g241180/u3_syn_4  , \g241188/u3_syn_4  , \g241196/u3_syn_4  , \g241205/u3_syn_4  , \g241213/u3_syn_4  , \g241221/u3_syn_4  , \g241229/u3_syn_4  , \g241237/u3_syn_4  , \g241245/u3_syn_4  , \g241253/u3_syn_4  , \g241261/u3_syn_4  , \g241269/u3_syn_4  , \g241277/u3_syn_4  , \g241285/u3_syn_4  , \g241293/u3_syn_4  , \g241301/u3_syn_4  , \g241309/u3_syn_4  , \g241317/u3_syn_4  , \g241325/u3_syn_4  , \g241333/u3_syn_4  , \g241341/u3_syn_4  , \g241349/u3_syn_4  , \g241358/u3_syn_4  , \g241366/u3_syn_4  , \g241374/u3_syn_4  , \g241382/u3_syn_4  , \g241390/u3_syn_4  , \g241398/u3_syn_4  , \g241406/u3_syn_4  , \g241415/u3_syn_4  , \g241424/u3_syn_4  , \g241433/u3_syn_4  , \g241441/u3_syn_4  , \g241449/u3_syn_4  , \g241459/u3_syn_4  , \g241470/u3_syn_4  , \g241480/u3_syn_4  , \g241489/u3_syn_4  , \g241497/u3_syn_4  , \g241505/u3_syn_4  , \g241513/u3_syn_4  , \g241545/_3_  , \g241580/_00_  , \g241737/_0_  , \g241752/_0_  , \g241755/_0_  , \g241767/_2__syn_2  , \g241781/_1__syn_2  , \g241782/_0_  , \g241803/_1__syn_2  , \g241805/_0_  , \g241812/_1__syn_2  , \g241814/_1__syn_2  , \g241816/_1__syn_2  , \g241819/_1__syn_2  , \g241822/_1__syn_2  , \g241823/_0_  , \g241833/_1__syn_2  , \g241843/_1__syn_2  , \g241844/_1__syn_2  , \g241848/_1__syn_2  , \g241855/_1__syn_2  , \g241868/_1__syn_2  , \g242013/_1__syn_2  , \g242015/_1__syn_2  , \g242017/_1__syn_2  , \g242021/_1__syn_2  , \g242039/_1__syn_2  , \g242081/_0_  , \g242086/_0_  , \g242101/_3_  , \g242116/_0_  , \g242135/_2_  , \g242147/_0_  , \g242158/_0_  , \g242196/_0_  , \g242202/_0_  , \g242203/_0_  , \g242204/_0_  , \g242212/_0_  , \g242226/_01_  , \g242281/_0_  , \g242407/_0_  , \g242410/_0_  , \g242426/_0_  , \g242438/_2_  , \g242466/_0_  , \g242530/_0_  , \g242532/_0_  , \g243397/_0_  , \g245925/_0_  , \g245932/_0_  , \g245933/_0_  , \g245986/_3_  , \g250157/_3_  , \g250202/_0_  , \g250246/_1_  , \g250248/_0_  , \g250250/_0_  , \g250305/_0_  , \g250323/_0_  , \g250373/_0_  , \g250377/_0_  , \g250412/_0_  , \g250413/_0_  , \g250418/_0_  , \g250419/_0_  , \g250421/_0_  , \g250433/_0_  , \g250448/_3_  , \g250567/_3_  , \g258965/_0_  , \g259006/_0_  , \g259471/_0_  , \g259473/_2_  , \g260557/_0_  , \g261035/_0_  , \g261095/_3_  , \g261207/_2__syn_2  , \g261754/_0_  , \g262017/_0_  , \g262045/_0_  , \g262046/_0_  , \g262100/_3_  , \g263539/_1_  , \g263574/_0_  , \g263858/_0_  , \g264104/_1_  , \g264107/_1_  , \g264117/_0_  , \g264282/_0_  , \g264511/_0_  , \g264541/_0_  , \g264562/_0_  , \g264618/_0_  , \g264660/_0_  , \g264681/_3_  , \g264727/_0_  , \g265013/_0_  , \g265084/_0_  , \g265378/_0_  , \g265413/_0_  , \g265446/_0_  , \g265486/_0_  , \g265524/_3_  , \g265528/_3_  , \g265548/_3_  , \g265579/_0_  , \g265768/_0_  , \g265801/_0_  , \g265819/_1_  , \g265853/_0_  , \g265933/_0_  , \g266022/_0_  , \g266183/_1_  , \g281909/_0_  , \g281965/_1_  , \g282284/_1_  , \g282639/_1_  , \g283047/_0_  , \g283157/_1_  , \g283184/_0_  , \g283334/_3_  , int_o_pad , \m_wb_adr_o[0]_pad  , \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2  , \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3  , \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3  , \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3  , \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3  , \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3  , \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3  , \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3  );
  input \CarrierSense_Tx2_reg/NET0131  ;
  input \Collision_Tx1_reg/NET0131  ;
  input \Collision_Tx2_reg/NET0131  ;
  input \RstTxPauseRq_reg/NET0131  ;
  input \RxAbortRst_reg/NET0131  ;
  input \RxAbort_latch_reg/NET0131  ;
  input \RxAbort_wb_reg/NET0131  ;
  input \RxEnSync_reg/NET0131  ;
  input \TPauseRq_reg/NET0131  ;
  input \TxPauseRq_sync2_reg/NET0131  ;
  input \TxPauseRq_sync3_reg/NET0131  ;
  input \WillSendControlFrame_sync2_reg/NET0131  ;
  input \WillSendControlFrame_sync3_reg/NET0131  ;
  input \WillTransmit_q2_reg/P0001  ;
  input \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131  ;
  input \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131  ;
  input \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131  ;
  input \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_IPGR1_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_IPGT_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_IPGT_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_IPGT_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_IPGT_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_IPGT_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_IPGT_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_IPGT_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131  ;
  input \ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MODER_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_MODER_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_MODER_2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  ;
  input \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  ;
  input \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131  ;
  input \ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131  ;
  input \ethreg1_ResetRxCIrq_sync2_reg/NET0131  ;
  input \ethreg1_ResetRxCIrq_sync3_reg/NET0131  ;
  input \ethreg1_ResetTxCIrq_sync2_reg/NET0131  ;
  input \ethreg1_SetRxCIrq_reg/NET0131  ;
  input \ethreg1_SetRxCIrq_rxclk_reg/NET0131  ;
  input \ethreg1_SetRxCIrq_sync2_reg/NET0131  ;
  input \ethreg1_SetRxCIrq_sync3_reg/NET0131  ;
  input \ethreg1_SetTxCIrq_reg/NET0131  ;
  input \ethreg1_SetTxCIrq_sync2_reg/NET0131  ;
  input \ethreg1_SetTxCIrq_sync3_reg/NET0131  ;
  input \ethreg1_SetTxCIrq_txclk_reg/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131  ;
  input \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131  ;
  input \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131  ;
  input \ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131  ;
  input \ethreg1_irq_busy_reg/NET0131  ;
  input \ethreg1_irq_rxb_reg/NET0131  ;
  input \ethreg1_irq_rxc_reg/NET0131  ;
  input \ethreg1_irq_rxe_reg/NET0131  ;
  input \ethreg1_irq_txb_reg/NET0131  ;
  input \ethreg1_irq_txc_reg/NET0131  ;
  input \ethreg1_irq_txe_reg/NET0131  ;
  input m_wb_ack_i_pad ;
  input \m_wb_adr_o[10]_pad  ;
  input \m_wb_adr_o[11]_pad  ;
  input \m_wb_adr_o[12]_pad  ;
  input \m_wb_adr_o[13]_pad  ;
  input \m_wb_adr_o[14]_pad  ;
  input \m_wb_adr_o[15]_pad  ;
  input \m_wb_adr_o[16]_pad  ;
  input \m_wb_adr_o[17]_pad  ;
  input \m_wb_adr_o[18]_pad  ;
  input \m_wb_adr_o[19]_pad  ;
  input \m_wb_adr_o[20]_pad  ;
  input \m_wb_adr_o[21]_pad  ;
  input \m_wb_adr_o[22]_pad  ;
  input \m_wb_adr_o[23]_pad  ;
  input \m_wb_adr_o[24]_pad  ;
  input \m_wb_adr_o[25]_pad  ;
  input \m_wb_adr_o[26]_pad  ;
  input \m_wb_adr_o[27]_pad  ;
  input \m_wb_adr_o[28]_pad  ;
  input \m_wb_adr_o[29]_pad  ;
  input \m_wb_adr_o[2]_pad  ;
  input \m_wb_adr_o[30]_pad  ;
  input \m_wb_adr_o[31]_pad  ;
  input \m_wb_adr_o[3]_pad  ;
  input \m_wb_adr_o[4]_pad  ;
  input \m_wb_adr_o[5]_pad  ;
  input \m_wb_adr_o[6]_pad  ;
  input \m_wb_adr_o[7]_pad  ;
  input \m_wb_adr_o[8]_pad  ;
  input \m_wb_adr_o[9]_pad  ;
  input \m_wb_dat_i[10]_pad  ;
  input \m_wb_dat_i[11]_pad  ;
  input \m_wb_dat_i[12]_pad  ;
  input \m_wb_dat_i[13]_pad  ;
  input \m_wb_dat_i[14]_pad  ;
  input \m_wb_dat_i[15]_pad  ;
  input \m_wb_dat_i[16]_pad  ;
  input \m_wb_dat_i[17]_pad  ;
  input \m_wb_dat_i[18]_pad  ;
  input \m_wb_dat_i[19]_pad  ;
  input \m_wb_dat_i[1]_pad  ;
  input \m_wb_dat_i[20]_pad  ;
  input \m_wb_dat_i[22]_pad  ;
  input \m_wb_dat_i[23]_pad  ;
  input \m_wb_dat_i[24]_pad  ;
  input \m_wb_dat_i[25]_pad  ;
  input \m_wb_dat_i[26]_pad  ;
  input \m_wb_dat_i[27]_pad  ;
  input \m_wb_dat_i[28]_pad  ;
  input \m_wb_dat_i[29]_pad  ;
  input \m_wb_dat_i[2]_pad  ;
  input \m_wb_dat_i[30]_pad  ;
  input \m_wb_dat_i[31]_pad  ;
  input \m_wb_dat_i[3]_pad  ;
  input \m_wb_dat_i[4]_pad  ;
  input \m_wb_dat_i[5]_pad  ;
  input \m_wb_dat_i[6]_pad  ;
  input \m_wb_dat_i[7]_pad  ;
  input \m_wb_dat_i[8]_pad  ;
  input m_wb_err_i_pad ;
  input \m_wb_sel_o[0]_pad  ;
  input \m_wb_sel_o[1]_pad  ;
  input \m_wb_sel_o[2]_pad  ;
  input \m_wb_sel_o[3]_pad  ;
  input m_wb_stb_o_pad ;
  input m_wb_we_o_pad ;
  input \maccontrol1_MuxedAbort_reg/NET0131  ;
  input \maccontrol1_MuxedDone_reg/NET0131  ;
  input \maccontrol1_TxAbortInLatched_reg/NET0131  ;
  input \maccontrol1_TxDoneInLatched_reg/NET0131  ;
  input \maccontrol1_TxUsedDataOutDetected_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_AddressOK_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131  ;
  input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131  ;
  input \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  ;
  input \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  ;
  input \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  ;
  input \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
  input \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  ;
  input \maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_Divider2_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131  ;
  input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131  ;
  input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131  ;
  input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131  ;
  input \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131  ;
  input \maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  ;
  input \maccontrol1_receivecontrol1_Pause_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131  ;
  input \maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131  ;
  input \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  ;
  input \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131  ;
  input \maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131  ;
  input \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  ;
  input \maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131  ;
  input \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131  ;
  input \maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131  ;
  input \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131  ;
  input \maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001  ;
  input \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131  ;
  input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131  ;
  input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  ;
  input \maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131  ;
  input \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131  ;
  input \maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001  ;
  input \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  ;
  input \maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131  ;
  input \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131  ;
  input \macstatus1_CarrierSenseLost_reg/NET0131  ;
  input \macstatus1_DeferLatched_reg/NET0131  ;
  input \macstatus1_DribbleNibble_reg/NET0131  ;
  input \macstatus1_InvalidSymbol_reg/NET0131  ;
  input \macstatus1_LatchedCrcError_reg/NET0131  ;
  input \macstatus1_LatchedMRxErr_reg/NET0131  ;
  input \macstatus1_LateCollLatched_reg/P0002  ;
  input \macstatus1_LoadRxStatus_reg/NET0131  ;
  input \macstatus1_ReceiveEnd_reg/NET0131  ;
  input \macstatus1_ReceivedPacketTooBig_reg/NET0131  ;
  input \macstatus1_RetryCntLatched_reg[0]/P0002  ;
  input \macstatus1_RetryCntLatched_reg[1]/P0002  ;
  input \macstatus1_RetryCntLatched_reg[2]/P0002  ;
  input \macstatus1_RetryCntLatched_reg[3]/P0002  ;
  input \macstatus1_RetryLimit_reg/P0002  ;
  input \macstatus1_RxColWindow_reg/NET0131  ;
  input \macstatus1_RxLateCollision_reg/NET0131  ;
  input \macstatus1_ShortFrame_reg/NET0131  ;
  input mcoll_pad_i_pad ;
  input md_pad_i_pad ;
  input mdc_pad_o_pad ;
  input \miim1_BitCounter_reg[0]/NET0131  ;
  input \miim1_BitCounter_reg[1]/NET0131  ;
  input \miim1_BitCounter_reg[2]/NET0131  ;
  input \miim1_BitCounter_reg[3]/NET0131  ;
  input \miim1_BitCounter_reg[4]/NET0131  ;
  input \miim1_BitCounter_reg[5]/NET0131  ;
  input \miim1_BitCounter_reg[6]/NET0131  ;
  input \miim1_EndBusy_reg/NET0131  ;
  input \miim1_InProgress_q1_reg/NET0131  ;
  input \miim1_InProgress_q2_reg/NET0131  ;
  input \miim1_InProgress_q3_reg/NET0131  ;
  input \miim1_InProgress_reg/NET0131  ;
  input \miim1_LatchByte0_d_reg/NET0131  ;
  input \miim1_LatchByte1_d_reg/NET0131  ;
  input \miim1_LatchByte_reg[0]/NET0131  ;
  input \miim1_LatchByte_reg[1]/NET0131  ;
  input \miim1_Nvalid_reg/NET0131  ;
  input \miim1_RStatStart_q1_reg/NET0131  ;
  input \miim1_RStatStart_q2_reg/NET0131  ;
  input \miim1_RStatStart_reg/NET0131  ;
  input \miim1_RStat_q2_reg/NET0131  ;
  input \miim1_RStat_q3_reg/NET0131  ;
  input \miim1_ScanStat_q2_reg/NET0131  ;
  input \miim1_SyncStatMdcEn_reg/NET0131  ;
  input \miim1_WCtrlDataStart_q1_reg/NET0131  ;
  input \miim1_WCtrlDataStart_q2_reg/NET0131  ;
  input \miim1_WCtrlDataStart_q_reg/NET0131  ;
  input \miim1_WCtrlDataStart_reg/NET0131  ;
  input \miim1_WCtrlData_q2_reg/NET0131  ;
  input \miim1_WCtrlData_q3_reg/NET0131  ;
  input \miim1_WriteOp_reg/NET0131  ;
  input \miim1_clkgen_Counter_reg[0]/NET0131  ;
  input \miim1_clkgen_Counter_reg[1]/NET0131  ;
  input \miim1_clkgen_Counter_reg[2]/NET0131  ;
  input \miim1_clkgen_Counter_reg[3]/NET0131  ;
  input \miim1_clkgen_Counter_reg[4]/NET0131  ;
  input \miim1_clkgen_Counter_reg[5]/NET0131  ;
  input \miim1_clkgen_Counter_reg[6]/NET0131  ;
  input \miim1_outctrl_Mdo_2d_reg/NET0131  ;
  input \miim1_shftrg_LinkFail_reg/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[0]/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[1]/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[2]/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[3]/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[4]/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[5]/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[6]/NET0131  ;
  input \miim1_shftrg_ShiftReg_reg[7]/NET0131  ;
  input \mrxd_pad_i[0]_pad  ;
  input \mrxd_pad_i[1]_pad  ;
  input \mrxd_pad_i[2]_pad  ;
  input \mrxd_pad_i[3]_pad  ;
  input mrxdv_pad_i_pad ;
  input mrxerr_pad_i_pad ;
  input \mtxd_pad_o[0]_pad  ;
  input \mtxd_pad_o[1]_pad  ;
  input \mtxd_pad_o[2]_pad  ;
  input \mtxd_pad_o[3]_pad  ;
  input mtxen_pad_o_pad ;
  input mtxerr_pad_o_pad ;
  input \rxethmac1_Broadcast_reg/NET0131  ;
  input \rxethmac1_CrcHashGood_reg/P0001  ;
  input \rxethmac1_CrcHash_reg[0]/P0001  ;
  input \rxethmac1_CrcHash_reg[1]/P0001  ;
  input \rxethmac1_CrcHash_reg[2]/P0001  ;
  input \rxethmac1_CrcHash_reg[3]/P0001  ;
  input \rxethmac1_CrcHash_reg[4]/P0001  ;
  input \rxethmac1_CrcHash_reg[5]/P0001  ;
  input \rxethmac1_DelayData_reg/NET0131  ;
  input \rxethmac1_LatchedByte_reg[0]/NET0131  ;
  input \rxethmac1_LatchedByte_reg[1]/NET0131  ;
  input \rxethmac1_LatchedByte_reg[2]/NET0131  ;
  input \rxethmac1_LatchedByte_reg[3]/NET0131  ;
  input \rxethmac1_LatchedByte_reg[4]/NET0131  ;
  input \rxethmac1_LatchedByte_reg[5]/NET0131  ;
  input \rxethmac1_LatchedByte_reg[6]/NET0131  ;
  input \rxethmac1_LatchedByte_reg[7]/NET0131  ;
  input \rxethmac1_Multicast_reg/NET0131  ;
  input \rxethmac1_RxData_d_reg[0]/NET0131  ;
  input \rxethmac1_RxData_d_reg[1]/NET0131  ;
  input \rxethmac1_RxData_d_reg[2]/NET0131  ;
  input \rxethmac1_RxData_d_reg[3]/NET0131  ;
  input \rxethmac1_RxData_d_reg[4]/NET0131  ;
  input \rxethmac1_RxData_d_reg[5]/NET0131  ;
  input \rxethmac1_RxData_d_reg[6]/NET0131  ;
  input \rxethmac1_RxData_d_reg[7]/NET0131  ;
  input \rxethmac1_RxData_reg[0]/NET0131  ;
  input \rxethmac1_RxData_reg[1]/NET0131  ;
  input \rxethmac1_RxData_reg[2]/NET0131  ;
  input \rxethmac1_RxData_reg[3]/NET0131  ;
  input \rxethmac1_RxData_reg[4]/NET0131  ;
  input \rxethmac1_RxData_reg[5]/NET0131  ;
  input \rxethmac1_RxData_reg[6]/NET0131  ;
  input \rxethmac1_RxData_reg[7]/NET0131  ;
  input \rxethmac1_RxEndFrm_d_reg/NET0131  ;
  input \rxethmac1_RxEndFrm_reg/NET0131  ;
  input \rxethmac1_RxStartFrm_reg/NET0131  ;
  input \rxethmac1_RxValid_reg/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[0]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[10]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[11]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[12]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[13]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[14]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[15]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[16]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[17]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[18]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[19]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[1]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[20]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[21]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[22]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[23]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[24]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[25]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[26]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[27]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[28]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[29]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[2]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[30]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[31]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[3]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[4]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[5]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[6]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[7]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[8]/NET0131  ;
  input \rxethmac1_crcrx_Crc_reg[9]/NET0131  ;
  input \rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131  ;
  input \rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131  ;
  input \rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131  ;
  input \rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  input \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  input \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  ;
  input \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  ;
  input \rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  ;
  input \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  ;
  input \rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131  ;
  input \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  ;
  input \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  ;
  input \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131  ;
  input \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131  ;
  input \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  input \rxethmac1_rxstatem1_StateData1_reg/NET0131  ;
  input \rxethmac1_rxstatem1_StateDrop_reg/NET0131  ;
  input \rxethmac1_rxstatem1_StateIdle_reg/NET0131  ;
  input \rxethmac1_rxstatem1_StatePreamble_reg/NET0131  ;
  input \rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  input \txethmac1_ColWindow_reg/NET0131  ;
  input \txethmac1_PacketFinished_q_reg/NET0131  ;
  input \txethmac1_RetryCnt_reg[0]/NET0131  ;
  input \txethmac1_RetryCnt_reg[1]/NET0131  ;
  input \txethmac1_RetryCnt_reg[2]/NET0131  ;
  input \txethmac1_RetryCnt_reg[3]/NET0131  ;
  input \txethmac1_StatusLatch_reg/NET0131  ;
  input \txethmac1_StopExcessiveDeferOccured_reg/NET0131  ;
  input \txethmac1_TxAbort_reg/NET0131  ;
  input \txethmac1_TxDone_reg/NET0131  ;
  input \txethmac1_TxRetry_reg/NET0131  ;
  input \txethmac1_TxUsedData_reg/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[0]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[1]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[2]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[3]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[4]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[5]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[6]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[7]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[8]/NET0131  ;
  input \txethmac1_random1_RandomLatched_reg[9]/NET0131  ;
  input \txethmac1_random1_x_reg[1]/NET0131  ;
  input \txethmac1_random1_x_reg[2]/NET0131  ;
  input \txethmac1_random1_x_reg[3]/NET0131  ;
  input \txethmac1_random1_x_reg[4]/NET0131  ;
  input \txethmac1_random1_x_reg[5]/NET0131  ;
  input \txethmac1_random1_x_reg[6]/NET0131  ;
  input \txethmac1_random1_x_reg[7]/NET0131  ;
  input \txethmac1_random1_x_reg[8]/NET0131  ;
  input \txethmac1_random1_x_reg[9]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  ;
  input \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
  input \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  ;
  input \txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131  ;
  input \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[14]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[15]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  ;
  input \txethmac1_txcounters1_NibCnt_reg[9]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[0]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[10]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[11]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[12]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[13]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[14]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[15]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[16]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[17]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[18]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[19]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[1]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[20]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[21]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[22]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[23]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[24]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[25]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[26]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[27]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[28]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[29]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[2]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[30]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[31]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[3]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[4]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[5]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[6]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[7]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[8]/NET0131  ;
  input \txethmac1_txcrc_Crc_reg[9]/NET0131  ;
  input \txethmac1_txstatem1_Rule1_reg/NET0131  ;
  input \txethmac1_txstatem1_StateBackOff_reg/NET0131  ;
  input \txethmac1_txstatem1_StateData_reg[0]/NET0131  ;
  input \txethmac1_txstatem1_StateData_reg[1]/NET0131  ;
  input \txethmac1_txstatem1_StateDefer_reg/NET0131  ;
  input \txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  input \txethmac1_txstatem1_StateIPG_reg/NET0131  ;
  input \txethmac1_txstatem1_StateIdle_reg/NET0131  ;
  input \txethmac1_txstatem1_StateJam_q_reg/NET0131  ;
  input \txethmac1_txstatem1_StateJam_reg/NET0131  ;
  input \txethmac1_txstatem1_StatePAD_reg/NET0131  ;
  input \txethmac1_txstatem1_StatePreamble_reg/NET0131  ;
  input wb_ack_o_pad ;
  input \wb_adr_i[10]_pad  ;
  input \wb_adr_i[11]_pad  ;
  input \wb_adr_i[2]_pad  ;
  input \wb_adr_i[3]_pad  ;
  input \wb_adr_i[4]_pad  ;
  input \wb_adr_i[5]_pad  ;
  input \wb_adr_i[6]_pad  ;
  input \wb_adr_i[7]_pad  ;
  input \wb_adr_i[8]_pad  ;
  input \wb_adr_i[9]_pad  ;
  input wb_cyc_i_pad ;
  input \wb_dat_i[0]_pad  ;
  input \wb_dat_i[10]_pad  ;
  input \wb_dat_i[11]_pad  ;
  input \wb_dat_i[12]_pad  ;
  input \wb_dat_i[13]_pad  ;
  input \wb_dat_i[14]_pad  ;
  input \wb_dat_i[15]_pad  ;
  input \wb_dat_i[16]_pad  ;
  input \wb_dat_i[17]_pad  ;
  input \wb_dat_i[18]_pad  ;
  input \wb_dat_i[19]_pad  ;
  input \wb_dat_i[1]_pad  ;
  input \wb_dat_i[20]_pad  ;
  input \wb_dat_i[21]_pad  ;
  input \wb_dat_i[22]_pad  ;
  input \wb_dat_i[23]_pad  ;
  input \wb_dat_i[24]_pad  ;
  input \wb_dat_i[25]_pad  ;
  input \wb_dat_i[26]_pad  ;
  input \wb_dat_i[27]_pad  ;
  input \wb_dat_i[28]_pad  ;
  input \wb_dat_i[29]_pad  ;
  input \wb_dat_i[2]_pad  ;
  input \wb_dat_i[30]_pad  ;
  input \wb_dat_i[31]_pad  ;
  input \wb_dat_i[3]_pad  ;
  input \wb_dat_i[4]_pad  ;
  input \wb_dat_i[5]_pad  ;
  input \wb_dat_i[6]_pad  ;
  input \wb_dat_i[7]_pad  ;
  input \wb_dat_i[8]_pad  ;
  input \wb_dat_i[9]_pad  ;
  input wb_err_o_pad ;
  input wb_rst_i_pad ;
  input \wb_sel_i[0]_pad  ;
  input \wb_sel_i[1]_pad  ;
  input \wb_sel_i[2]_pad  ;
  input \wb_sel_i[3]_pad  ;
  input wb_stb_i_pad ;
  input wb_we_i_pad ;
  input \wishbone_BDRead_reg/NET0131  ;
  input \wishbone_BDWrite_reg[0]/NET0131  ;
  input \wishbone_BDWrite_reg[1]/NET0131  ;
  input \wishbone_BDWrite_reg[2]/NET0131  ;
  input \wishbone_BDWrite_reg[3]/NET0131  ;
  input \wishbone_BlockReadTxDataFromMemory_reg/NET0131  ;
  input \wishbone_BlockingIncrementTxPointer_reg/NET0131  ;
  input \wishbone_BlockingTxBDRead_reg/NET0131  ;
  input \wishbone_BlockingTxStatusWrite_reg/NET0131  ;
  input \wishbone_BlockingTxStatusWrite_sync2_reg/NET0131  ;
  input \wishbone_BlockingTxStatusWrite_sync3_reg/NET0131  ;
  input \wishbone_Busy_IRQ_rck_reg/NET0131  ;
  input \wishbone_Busy_IRQ_sync2_reg/P0001  ;
  input \wishbone_Busy_IRQ_sync3_reg/P0001  ;
  input \wishbone_Busy_IRQ_syncb2_reg/P0001  ;
  input \wishbone_Flop_reg/NET0131  ;
  input \wishbone_IncrTxPointer_reg/NET0131  ;
  input \wishbone_LastByteIn_reg/NET0131  ;
  input \wishbone_LastWord_reg/NET0131  ;
  input \wishbone_LatchValidBytes_q_reg/NET0131  ;
  input \wishbone_LatchValidBytes_reg/NET0131  ;
  input \wishbone_LatchedRxLength_reg[0]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[10]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[11]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[12]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[13]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[14]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[15]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[1]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[2]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[3]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[4]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[5]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[6]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[7]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[8]/NET0131  ;
  input \wishbone_LatchedRxLength_reg[9]/NET0131  ;
  input \wishbone_LatchedRxStartFrm_reg/NET0131  ;
  input \wishbone_LatchedTxLength_reg[0]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[10]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[11]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[12]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[13]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[14]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[15]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[1]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[2]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[3]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[4]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[5]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[6]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[7]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[8]/NET0131  ;
  input \wishbone_LatchedTxLength_reg[9]/NET0131  ;
  input \wishbone_MasterWbRX_reg/NET0131  ;
  input \wishbone_MasterWbTX_reg/NET0131  ;
  input \wishbone_ReadTxDataFromFifo_sync2_reg/NET0131  ;
  input \wishbone_ReadTxDataFromFifo_sync3_reg/NET0131  ;
  input \wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131  ;
  input \wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131  ;
  input \wishbone_ReadTxDataFromFifo_tck_reg/NET0131  ;
  input \wishbone_ReadTxDataFromMemory_reg/NET0131  ;
  input \wishbone_RxAbortLatched_reg/NET0131  ;
  input \wishbone_RxAbortSync2_reg/NET0131  ;
  input \wishbone_RxAbortSync3_reg/NET0131  ;
  input \wishbone_RxAbortSync4_reg/NET0131  ;
  input \wishbone_RxAbortSyncb2_reg/NET0131  ;
  input \wishbone_RxBDAddress_reg[1]/NET0131  ;
  input \wishbone_RxBDAddress_reg[2]/NET0131  ;
  input \wishbone_RxBDAddress_reg[3]/NET0131  ;
  input \wishbone_RxBDAddress_reg[4]/NET0131  ;
  input \wishbone_RxBDAddress_reg[5]/NET0131  ;
  input \wishbone_RxBDAddress_reg[6]/NET0131  ;
  input \wishbone_RxBDAddress_reg[7]/NET0131  ;
  input \wishbone_RxBDRead_reg/NET0131  ;
  input \wishbone_RxBDReady_reg/NET0131  ;
  input \wishbone_RxB_IRQ_reg/NET0131  ;
  input \wishbone_RxByteCnt_reg[0]/NET0131  ;
  input \wishbone_RxByteCnt_reg[1]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[10]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[11]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[12]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[13]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[14]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[15]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[16]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[17]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[18]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[19]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[20]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[21]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[22]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[23]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[24]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[25]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[26]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[27]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[28]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[29]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[30]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[31]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[8]/NET0131  ;
  input \wishbone_RxDataLatched1_reg[9]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[0]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[10]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[11]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[12]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[13]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[14]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[15]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[16]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[17]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[18]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[19]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[1]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[20]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[21]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[22]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[23]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[24]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[25]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[26]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[27]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[28]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[29]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[2]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[30]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[31]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[3]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[4]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[5]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[6]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[7]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[8]/NET0131  ;
  input \wishbone_RxDataLatched2_reg[9]/NET0131  ;
  input \wishbone_RxE_IRQ_reg/NET0131  ;
  input \wishbone_RxEn_needed_reg/NET0131  ;
  input \wishbone_RxEn_q_reg/NET0131  ;
  input \wishbone_RxEn_reg/NET0131  ;
  input \wishbone_RxEnableWindow_reg/NET0131  ;
  input \wishbone_RxOverrun_reg/NET0131  ;
  input \wishbone_RxPointerLSB_rst_reg[0]/NET0131  ;
  input \wishbone_RxPointerLSB_rst_reg[1]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[10]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[11]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[12]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[13]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[14]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[15]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[16]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[17]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[18]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[19]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[20]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[21]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[22]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[23]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[24]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[25]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[26]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[27]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[28]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[29]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[2]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[30]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[31]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[3]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[4]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[5]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[6]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[7]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[8]/NET0131  ;
  input \wishbone_RxPointerMSB_reg[9]/NET0131  ;
  input \wishbone_RxPointerRead_reg/NET0131  ;
  input \wishbone_RxReady_reg/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[0]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[1]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[2]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[3]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[4]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[5]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[6]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[7]/NET0131  ;
  input \wishbone_RxStatusInLatched_reg[8]/NET0131  ;
  input \wishbone_RxStatusWriteLatched_reg/NET0131  ;
  input \wishbone_RxStatusWriteLatched_sync2_reg/NET0131  ;
  input \wishbone_RxStatusWriteLatched_syncb2_reg/NET0131  ;
  input \wishbone_RxStatus_reg[13]/NET0131  ;
  input \wishbone_RxStatus_reg[14]/NET0131  ;
  input \wishbone_RxValidBytes_reg[0]/NET0131  ;
  input \wishbone_RxValidBytes_reg[1]/NET0131  ;
  input \wishbone_ShiftEndedSync1_reg/NET0131  ;
  input \wishbone_ShiftEndedSync2_reg/NET0131  ;
  input \wishbone_ShiftEndedSync3_reg/NET0131  ;
  input \wishbone_ShiftEndedSync_c1_reg/NET0131  ;
  input \wishbone_ShiftEndedSync_c2_reg/NET0131  ;
  input \wishbone_ShiftEnded_rck_reg/NET0131  ;
  input \wishbone_ShiftEnded_reg/NET0131  ;
  input \wishbone_ShiftWillEnd_reg/NET0131  ;
  input \wishbone_StartOccured_reg/NET0131  ;
  input \wishbone_SyncRxStartFrm_q2_reg/NET0131  ;
  input \wishbone_SyncRxStartFrm_q_reg/NET0131  ;
  input \wishbone_TxAbortPacketBlocked_reg/NET0131  ;
  input \wishbone_TxAbortPacket_NotCleared_reg/NET0131  ;
  input \wishbone_TxAbortPacket_reg/NET0131  ;
  input \wishbone_TxAbort_q_reg/NET0131  ;
  input \wishbone_TxAbort_wb_q_reg/NET0131  ;
  input \wishbone_TxAbort_wb_reg/NET0131  ;
  input \wishbone_TxBDAddress_reg[1]/NET0131  ;
  input \wishbone_TxBDAddress_reg[2]/NET0131  ;
  input \wishbone_TxBDAddress_reg[3]/NET0131  ;
  input \wishbone_TxBDAddress_reg[4]/NET0131  ;
  input \wishbone_TxBDAddress_reg[5]/NET0131  ;
  input \wishbone_TxBDAddress_reg[6]/NET0131  ;
  input \wishbone_TxBDAddress_reg[7]/NET0131  ;
  input \wishbone_TxBDRead_reg/NET0131  ;
  input \wishbone_TxBDReady_reg/NET0131  ;
  input \wishbone_TxB_IRQ_reg/NET0131  ;
  input \wishbone_TxByteCnt_reg[0]/NET0131  ;
  input \wishbone_TxByteCnt_reg[1]/NET0131  ;
  input \wishbone_TxDataLatched_reg[0]/NET0131  ;
  input \wishbone_TxDataLatched_reg[10]/NET0131  ;
  input \wishbone_TxDataLatched_reg[11]/NET0131  ;
  input \wishbone_TxDataLatched_reg[12]/NET0131  ;
  input \wishbone_TxDataLatched_reg[13]/NET0131  ;
  input \wishbone_TxDataLatched_reg[14]/NET0131  ;
  input \wishbone_TxDataLatched_reg[15]/NET0131  ;
  input \wishbone_TxDataLatched_reg[16]/NET0131  ;
  input \wishbone_TxDataLatched_reg[17]/NET0131  ;
  input \wishbone_TxDataLatched_reg[18]/NET0131  ;
  input \wishbone_TxDataLatched_reg[19]/NET0131  ;
  input \wishbone_TxDataLatched_reg[1]/NET0131  ;
  input \wishbone_TxDataLatched_reg[20]/NET0131  ;
  input \wishbone_TxDataLatched_reg[21]/NET0131  ;
  input \wishbone_TxDataLatched_reg[22]/NET0131  ;
  input \wishbone_TxDataLatched_reg[23]/NET0131  ;
  input \wishbone_TxDataLatched_reg[24]/NET0131  ;
  input \wishbone_TxDataLatched_reg[25]/NET0131  ;
  input \wishbone_TxDataLatched_reg[26]/NET0131  ;
  input \wishbone_TxDataLatched_reg[27]/NET0131  ;
  input \wishbone_TxDataLatched_reg[28]/NET0131  ;
  input \wishbone_TxDataLatched_reg[29]/NET0131  ;
  input \wishbone_TxDataLatched_reg[2]/NET0131  ;
  input \wishbone_TxDataLatched_reg[30]/NET0131  ;
  input \wishbone_TxDataLatched_reg[31]/NET0131  ;
  input \wishbone_TxDataLatched_reg[3]/NET0131  ;
  input \wishbone_TxDataLatched_reg[4]/NET0131  ;
  input \wishbone_TxDataLatched_reg[5]/NET0131  ;
  input \wishbone_TxDataLatched_reg[6]/NET0131  ;
  input \wishbone_TxDataLatched_reg[7]/NET0131  ;
  input \wishbone_TxDataLatched_reg[8]/NET0131  ;
  input \wishbone_TxDataLatched_reg[9]/NET0131  ;
  input \wishbone_TxData_reg[0]/NET0131  ;
  input \wishbone_TxData_reg[1]/NET0131  ;
  input \wishbone_TxData_reg[2]/NET0131  ;
  input \wishbone_TxData_reg[3]/NET0131  ;
  input \wishbone_TxData_reg[4]/NET0131  ;
  input \wishbone_TxData_reg[5]/NET0131  ;
  input \wishbone_TxData_reg[6]/NET0131  ;
  input \wishbone_TxData_reg[7]/NET0131  ;
  input \wishbone_TxDonePacketBlocked_reg/NET0131  ;
  input \wishbone_TxDonePacket_NotCleared_reg/NET0131  ;
  input \wishbone_TxDonePacket_reg/NET0131  ;
  input \wishbone_TxDone_wb_q_reg/NET0131  ;
  input \wishbone_TxDone_wb_reg/NET0131  ;
  input \wishbone_TxE_IRQ_reg/NET0131  ;
  input \wishbone_TxEn_needed_reg/NET0131  ;
  input \wishbone_TxEn_q_reg/NET0131  ;
  input \wishbone_TxEn_reg/NET0131  ;
  input \wishbone_TxEndFrm_reg/NET0131  ;
  input \wishbone_TxEndFrm_wb_reg/NET0131  ;
  input \wishbone_TxLength_reg[0]/NET0131  ;
  input \wishbone_TxLength_reg[10]/NET0131  ;
  input \wishbone_TxLength_reg[11]/NET0131  ;
  input \wishbone_TxLength_reg[12]/NET0131  ;
  input \wishbone_TxLength_reg[13]/NET0131  ;
  input \wishbone_TxLength_reg[14]/NET0131  ;
  input \wishbone_TxLength_reg[15]/NET0131  ;
  input \wishbone_TxLength_reg[1]/NET0131  ;
  input \wishbone_TxLength_reg[2]/NET0131  ;
  input \wishbone_TxLength_reg[3]/NET0131  ;
  input \wishbone_TxLength_reg[4]/NET0131  ;
  input \wishbone_TxLength_reg[5]/NET0131  ;
  input \wishbone_TxLength_reg[6]/NET0131  ;
  input \wishbone_TxLength_reg[7]/NET0131  ;
  input \wishbone_TxLength_reg[8]/NET0131  ;
  input \wishbone_TxLength_reg[9]/NET0131  ;
  input \wishbone_TxPointerLSB_reg[0]/NET0131  ;
  input \wishbone_TxPointerLSB_reg[1]/NET0131  ;
  input \wishbone_TxPointerLSB_rst_reg[0]/NET0131  ;
  input \wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[10]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[11]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[12]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[13]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[14]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[15]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[16]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[17]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[18]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[19]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[20]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[21]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[22]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[23]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[24]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[25]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[26]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[27]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[28]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[29]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[2]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[30]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[31]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[3]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[4]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[5]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[6]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[7]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[8]/NET0131  ;
  input \wishbone_TxPointerMSB_reg[9]/NET0131  ;
  input \wishbone_TxPointerRead_reg/NET0131  ;
  input \wishbone_TxRetryPacketBlocked_reg/NET0131  ;
  input \wishbone_TxRetryPacket_NotCleared_reg/NET0131  ;
  input \wishbone_TxRetryPacket_reg/NET0131  ;
  input \wishbone_TxRetry_q_reg/NET0131  ;
  input \wishbone_TxRetry_wb_q_reg/NET0131  ;
  input \wishbone_TxRetry_wb_reg/NET0131  ;
  input \wishbone_TxStartFrm_reg/NET0131  ;
  input \wishbone_TxStartFrm_sync2_reg/NET0131  ;
  input \wishbone_TxStartFrm_syncb2_reg/NET0131  ;
  input \wishbone_TxStartFrm_wb_reg/NET0131  ;
  input \wishbone_TxStatus_reg[11]/NET0131  ;
  input \wishbone_TxStatus_reg[12]/NET0131  ;
  input \wishbone_TxStatus_reg[13]/NET0131  ;
  input \wishbone_TxStatus_reg[14]/NET0131  ;
  input \wishbone_TxUnderRun_reg/NET0131  ;
  input \wishbone_TxUnderRun_sync1_reg/NET0131  ;
  input \wishbone_TxUnderRun_wb_reg/NET0131  ;
  input \wishbone_TxUsedData_q_reg/NET0131  ;
  input \wishbone_TxValidBytesLatched_reg[0]/NET0131  ;
  input \wishbone_TxValidBytesLatched_reg[1]/NET0131  ;
  input \wishbone_WB_ACK_O_reg/P0001  ;
  input \wishbone_WbEn_q_reg/NET0131  ;
  input \wishbone_WbEn_reg/NET0131  ;
  input \wishbone_WriteRxDataToFifoSync2_reg/NET0131  ;
  input \wishbone_WriteRxDataToFifoSync3_reg/NET0131  ;
  input \wishbone_WriteRxDataToFifo_reg/NET0131  ;
  input \wishbone_bd_ram_mem0_reg[0][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[0][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[0][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[0][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[0][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[0][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[0][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[0][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[100][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[101][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[102][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[103][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[104][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[105][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[106][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[107][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[108][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[109][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[10][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[110][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[111][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[112][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[113][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[114][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[115][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[116][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[117][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[118][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[119][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[11][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[120][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[121][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[122][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[123][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[124][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[125][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[126][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[127][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[128][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[129][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[12][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[130][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[131][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[132][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[133][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[134][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[135][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[136][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[137][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[138][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[139][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[13][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[140][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[141][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[142][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[143][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[144][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[145][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[146][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[147][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[148][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[149][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[14][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[150][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[151][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[152][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[153][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[154][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[155][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[156][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[157][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[158][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[159][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[15][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[160][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[161][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[162][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[163][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[164][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[165][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[166][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[167][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[168][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[169][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[16][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[170][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[171][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[172][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[173][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[174][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[175][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[176][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[177][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[178][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[179][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[17][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[180][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[181][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[182][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[183][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[184][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[185][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[186][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[187][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[188][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[189][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[18][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[190][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[191][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[192][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[193][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[194][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[195][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[196][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[197][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[198][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[199][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[19][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[1][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[200][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[201][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[202][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[203][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[204][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[205][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[206][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[207][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[208][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[209][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[20][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[210][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[211][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[212][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[213][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[214][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[215][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[216][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[217][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[218][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[219][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[21][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[220][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[221][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[222][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[223][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[224][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[225][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[226][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[227][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[228][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[229][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[22][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[230][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[231][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[232][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[233][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[234][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[235][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[236][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[237][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[238][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[239][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[23][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[240][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[241][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[242][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[243][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[244][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[245][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[246][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[247][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[248][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[249][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[24][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[250][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[251][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[252][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[253][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[254][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[255][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[25][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[26][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[27][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[28][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[29][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[2][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[30][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[31][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[32][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[33][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[34][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[35][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[36][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[37][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[38][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[39][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[3][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[40][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[41][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[42][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[43][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[44][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[45][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[46][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[47][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[48][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[49][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[4][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[50][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[51][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[52][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[53][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[54][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[55][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[56][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[57][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[58][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[59][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[5][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[60][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[61][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[62][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[63][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[64][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[65][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[66][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[67][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[68][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[69][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[6][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[70][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[71][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[72][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[73][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[74][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[75][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[76][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[77][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[78][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[79][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[7][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[80][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[81][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[82][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[83][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[84][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[85][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[86][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[87][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[88][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[89][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[8][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[90][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[91][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[92][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[93][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[94][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[95][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[96][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[97][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[98][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[99][7]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][0]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][1]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][2]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][3]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][4]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][5]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][6]/P0001  ;
  input \wishbone_bd_ram_mem0_reg[9][7]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[0][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[100][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[101][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[102][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[103][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[104][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[105][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[106][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[107][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[108][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[109][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[10][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[110][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[111][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[112][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[113][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[114][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[115][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[116][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[117][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[118][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[119][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[11][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[120][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[121][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[122][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[123][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[124][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[125][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[126][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[127][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[128][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[129][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[12][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[130][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[131][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[132][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[133][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[134][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[135][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[136][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[137][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[138][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[139][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[13][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[140][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[141][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[142][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[143][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[144][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[145][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[146][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[147][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[148][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[149][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[14][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[150][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[151][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[152][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[153][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[154][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[155][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[156][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[157][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[158][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[159][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[15][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[160][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[161][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[162][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[163][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[164][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[165][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[166][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[167][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[168][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[169][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[16][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[170][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[171][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[172][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[173][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[174][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[175][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[176][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[177][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[178][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[179][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[17][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[180][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[181][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[182][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[183][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[184][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[185][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[186][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[187][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[188][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[189][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[18][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[190][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[191][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[192][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[193][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[194][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[195][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[196][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[197][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[198][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[199][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[19][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[1][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[200][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[201][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[202][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[203][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[204][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[205][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[206][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[207][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[208][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[209][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[20][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[210][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[211][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[212][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[213][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[214][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[215][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[216][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[217][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[218][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[219][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[21][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[220][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[221][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[222][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[223][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[224][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[225][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[226][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[227][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[228][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[229][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[22][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[230][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[231][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[232][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[233][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[234][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[235][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[236][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[237][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[238][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[239][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[23][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[240][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[241][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[242][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[243][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[244][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[245][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[246][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[247][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[248][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[249][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[24][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[250][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[251][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[252][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[253][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[254][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[255][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[25][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[26][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[27][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[28][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[29][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[2][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[30][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[31][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[32][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[33][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[34][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[35][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[36][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[37][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[38][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[39][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[3][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[40][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[41][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[42][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[43][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[44][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[45][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[46][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[47][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[48][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[49][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[4][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[50][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[51][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[52][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[53][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[54][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[55][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[56][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[57][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[58][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[59][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[5][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[60][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[61][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[62][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[63][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[64][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[65][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[66][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[67][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[68][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[69][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[6][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[70][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[71][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[72][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[73][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[74][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[75][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[76][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[77][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[78][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[79][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[7][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[80][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[81][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[82][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[83][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[84][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[85][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[86][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[87][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[88][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[89][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[8][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[90][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[91][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[92][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[93][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[94][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[95][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[96][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[97][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[98][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[99][9]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][10]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][11]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][12]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][13]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][14]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][15]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][8]/P0001  ;
  input \wishbone_bd_ram_mem1_reg[9][9]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[0][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[100][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[101][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[102][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[103][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[104][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[105][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[106][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[107][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[108][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[109][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[10][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[110][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[111][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[112][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[113][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[114][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[115][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[116][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[117][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[118][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[119][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[11][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[120][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[121][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[122][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[123][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[124][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[125][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[126][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[127][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[128][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[129][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[12][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[130][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[131][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[132][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[133][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[134][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[135][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[136][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[137][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[138][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[139][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[13][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[140][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[141][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[142][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[143][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[144][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[145][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[146][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[147][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[148][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[149][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[14][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[150][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[151][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[152][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[153][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[154][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[155][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[156][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[157][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[158][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[159][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[15][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[160][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[161][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[162][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[163][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[164][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[165][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[166][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[167][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[168][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[169][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[16][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[170][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[171][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[172][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[173][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[174][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[175][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[176][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[177][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[178][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[179][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[17][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[180][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[181][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[182][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[183][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[184][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[185][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[186][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[187][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[188][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[189][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[18][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[190][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[191][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[192][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[193][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[194][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[195][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[196][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[197][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[198][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[199][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[19][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[1][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[200][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[201][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[202][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[203][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[204][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[205][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[206][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[207][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[208][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[209][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[20][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[210][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[211][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[212][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[213][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[214][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[215][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[216][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[217][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[218][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[219][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[21][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[220][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[221][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[222][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[223][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[224][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[225][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[226][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[227][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[228][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[229][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[22][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[230][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[231][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[232][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[233][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[234][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[235][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[236][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[237][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[238][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[239][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[23][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[240][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[241][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[242][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[243][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[244][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[245][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[246][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[247][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[248][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[249][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[24][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[250][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[251][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[252][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[253][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[254][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[255][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[25][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[26][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[27][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[28][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[29][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[2][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[30][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[31][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[32][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[33][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[34][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[35][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[36][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[37][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[38][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[39][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[3][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[40][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[41][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[42][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[43][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[44][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[45][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[46][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[47][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[48][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[49][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[4][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[50][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[51][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[52][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[53][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[54][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[55][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[56][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[57][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[58][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[59][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[5][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[60][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[61][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[62][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[63][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[64][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[65][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[66][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[67][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[68][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[69][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[6][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[70][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[71][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[72][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[73][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[74][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[75][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[76][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[77][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[78][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[79][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[7][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[80][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[81][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[82][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[83][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[84][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[85][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[86][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[87][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[88][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[89][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[8][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[90][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[91][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[92][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[93][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[94][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[95][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[96][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[97][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[98][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[99][23]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][16]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][17]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][18]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][19]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][20]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][21]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][22]/P0001  ;
  input \wishbone_bd_ram_mem2_reg[9][23]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[0][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[100][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[101][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[102][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[103][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[104][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[105][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[106][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[107][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[108][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[109][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[10][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[110][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[111][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[112][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[113][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[114][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[115][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[116][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[117][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[118][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[119][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[11][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[120][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[121][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[122][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[123][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[124][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[125][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[126][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[127][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[128][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[129][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[12][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[130][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[131][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[132][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[133][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[134][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[135][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[136][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[137][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[138][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[139][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[13][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[140][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[141][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[142][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[143][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[144][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[145][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[146][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[147][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[148][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[149][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[14][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[150][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[151][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[152][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[153][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[154][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[155][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[156][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[157][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[158][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[159][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[15][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[160][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[161][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[162][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[163][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[164][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[165][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[166][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[167][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[168][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[169][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[16][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[170][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[171][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[172][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[173][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[174][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[175][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[176][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[177][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[178][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[179][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[17][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[180][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[181][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[182][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[183][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[184][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[185][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[186][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[187][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[188][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[189][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[18][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[190][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[191][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[192][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[193][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[194][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[195][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[196][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[197][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[198][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[199][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[19][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[1][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[200][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[201][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[202][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[203][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[204][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[205][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[206][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[207][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[208][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[209][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[20][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[210][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[211][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[212][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[213][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[214][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[215][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[216][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[217][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[218][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[219][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[21][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[220][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[221][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[222][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[223][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[224][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[225][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[226][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[227][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[228][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[229][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[22][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[230][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[231][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[232][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[233][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[234][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[235][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[236][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[237][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[238][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[239][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[23][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[240][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[241][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[242][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[243][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[244][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[245][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[246][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[247][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[248][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[249][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[24][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[250][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[251][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[252][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[253][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[254][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[255][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[25][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[26][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[27][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[28][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[29][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[2][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[30][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[31][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[32][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[33][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[34][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[35][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[36][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[37][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[38][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[39][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[3][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[40][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[41][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[42][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[43][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[44][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[45][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[46][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[47][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[48][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[49][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[4][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[50][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[51][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[52][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[53][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[54][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[55][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[56][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[57][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[58][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[59][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[5][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[60][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[61][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[62][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[63][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[64][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[65][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[66][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[67][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[68][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[69][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[6][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[70][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[71][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[72][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[73][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[74][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[75][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[76][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[77][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[78][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[79][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[7][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[80][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[81][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[82][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[83][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[84][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[85][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[86][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[87][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[88][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[89][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[8][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[90][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[91][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[92][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[93][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[94][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[95][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[96][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[97][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[98][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[99][31]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][24]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][25]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][26]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][27]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][28]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][29]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][30]/P0001  ;
  input \wishbone_bd_ram_mem3_reg[9][31]/P0001  ;
  input \wishbone_bd_ram_raddr_reg[0]/P0001  ;
  input \wishbone_bd_ram_raddr_reg[1]/NET0131  ;
  input \wishbone_bd_ram_raddr_reg[2]/NET0131  ;
  input \wishbone_bd_ram_raddr_reg[3]/P0001  ;
  input \wishbone_bd_ram_raddr_reg[4]/NET0131  ;
  input \wishbone_bd_ram_raddr_reg[5]/NET0131  ;
  input \wishbone_bd_ram_raddr_reg[6]/NET0131  ;
  input \wishbone_bd_ram_raddr_reg[7]/NET0131  ;
  input \wishbone_cyc_cleared_reg/NET0131  ;
  input \wishbone_r_RxEn_q_reg/NET0131  ;
  input \wishbone_r_TxEn_q_reg/NET0131  ;
  input \wishbone_ram_addr_reg[0]/NET0131  ;
  input \wishbone_ram_addr_reg[1]/NET0131  ;
  input \wishbone_ram_addr_reg[2]/NET0131  ;
  input \wishbone_ram_addr_reg[3]/NET0131  ;
  input \wishbone_ram_addr_reg[4]/NET0131  ;
  input \wishbone_ram_addr_reg[5]/NET0131  ;
  input \wishbone_ram_addr_reg[6]/NET0131  ;
  input \wishbone_ram_addr_reg[7]/NET0131  ;
  input \wishbone_ram_di_reg[0]/NET0131  ;
  input \wishbone_ram_di_reg[10]/NET0131  ;
  input \wishbone_ram_di_reg[11]/NET0131  ;
  input \wishbone_ram_di_reg[12]/NET0131  ;
  input \wishbone_ram_di_reg[13]/NET0131  ;
  input \wishbone_ram_di_reg[14]/NET0131  ;
  input \wishbone_ram_di_reg[15]/NET0131  ;
  input \wishbone_ram_di_reg[16]/NET0131  ;
  input \wishbone_ram_di_reg[17]/NET0131  ;
  input \wishbone_ram_di_reg[18]/NET0131  ;
  input \wishbone_ram_di_reg[19]/NET0131  ;
  input \wishbone_ram_di_reg[1]/NET0131  ;
  input \wishbone_ram_di_reg[20]/NET0131  ;
  input \wishbone_ram_di_reg[21]/NET0131  ;
  input \wishbone_ram_di_reg[22]/NET0131  ;
  input \wishbone_ram_di_reg[23]/NET0131  ;
  input \wishbone_ram_di_reg[24]/NET0131  ;
  input \wishbone_ram_di_reg[25]/NET0131  ;
  input \wishbone_ram_di_reg[26]/NET0131  ;
  input \wishbone_ram_di_reg[27]/NET0131  ;
  input \wishbone_ram_di_reg[28]/NET0131  ;
  input \wishbone_ram_di_reg[29]/NET0131  ;
  input \wishbone_ram_di_reg[2]/NET0131  ;
  input \wishbone_ram_di_reg[30]/NET0131  ;
  input \wishbone_ram_di_reg[31]/NET0131  ;
  input \wishbone_ram_di_reg[3]/NET0131  ;
  input \wishbone_ram_di_reg[4]/NET0131  ;
  input \wishbone_ram_di_reg[5]/NET0131  ;
  input \wishbone_ram_di_reg[6]/NET0131  ;
  input \wishbone_ram_di_reg[7]/NET0131  ;
  input \wishbone_ram_di_reg[8]/NET0131  ;
  input \wishbone_ram_di_reg[9]/NET0131  ;
  input \wishbone_rx_burst_cnt_reg[0]/NET0131  ;
  input \wishbone_rx_burst_cnt_reg[1]/NET0131  ;
  input \wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  input \wishbone_rx_burst_en_reg/NET0131  ;
  input \wishbone_rx_fifo_cnt_reg[0]/NET0131  ;
  input \wishbone_rx_fifo_cnt_reg[1]/NET0131  ;
  input \wishbone_rx_fifo_cnt_reg[2]/NET0131  ;
  input \wishbone_rx_fifo_cnt_reg[3]/NET0131  ;
  input \wishbone_rx_fifo_cnt_reg[4]/NET0131  ;
  input \wishbone_rx_fifo_fifo_reg[0][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[0][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[10][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[11][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[12][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[13][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[14][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[15][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[1][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[2][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[3][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[4][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[5][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[6][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[7][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[8][9]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][0]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][10]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][11]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][12]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][13]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][14]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][15]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][16]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][17]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][18]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][19]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][1]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][20]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][21]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][22]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][23]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][24]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][25]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][26]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][27]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][28]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][29]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][2]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][30]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][31]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][3]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][4]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][5]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][6]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][7]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][8]/P0001  ;
  input \wishbone_rx_fifo_fifo_reg[9][9]/P0001  ;
  input \wishbone_rx_fifo_read_pointer_reg[0]/NET0131  ;
  input \wishbone_rx_fifo_read_pointer_reg[1]/NET0131  ;
  input \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  ;
  input \wishbone_rx_fifo_read_pointer_reg[3]/NET0131  ;
  input \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  ;
  input \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  input \wishbone_rx_fifo_write_pointer_reg[2]/NET0131  ;
  input \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
  input \wishbone_tx_burst_cnt_reg[0]/NET0131  ;
  input \wishbone_tx_burst_cnt_reg[1]/NET0131  ;
  input \wishbone_tx_burst_cnt_reg[2]/NET0131  ;
  input \wishbone_tx_burst_en_reg/NET0131  ;
  input \wishbone_tx_fifo_cnt_reg[0]/NET0131  ;
  input \wishbone_tx_fifo_cnt_reg[1]/NET0131  ;
  input \wishbone_tx_fifo_cnt_reg[2]/NET0131  ;
  input \wishbone_tx_fifo_cnt_reg[3]/NET0131  ;
  input \wishbone_tx_fifo_cnt_reg[4]/NET0131  ;
  input \wishbone_tx_fifo_data_out_reg[0]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[10]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[11]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[12]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[13]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[14]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[15]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[16]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[17]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[18]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[19]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[1]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[20]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[21]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[22]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[23]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[24]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[25]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[26]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[27]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[28]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[29]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[2]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[30]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[31]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[3]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[4]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[5]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[6]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[7]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[8]/P0001  ;
  input \wishbone_tx_fifo_data_out_reg[9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[0][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[10][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[11][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[12][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[13][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[14][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[15][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[1][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[2][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[3][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[4][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[5][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[6][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[7][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[8][9]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][0]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][10]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][11]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][12]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][13]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][14]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][15]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][16]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][17]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][18]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][19]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][1]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][20]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][21]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][22]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][23]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][24]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][25]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][26]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][27]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][28]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][29]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][2]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][30]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][31]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][3]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][4]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][5]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][6]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][7]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][8]/P0001  ;
  input \wishbone_tx_fifo_fifo_reg[9][9]/P0001  ;
  input \wishbone_tx_fifo_read_pointer_reg[0]/NET0131  ;
  input \wishbone_tx_fifo_read_pointer_reg[1]/NET0131  ;
  input \wishbone_tx_fifo_read_pointer_reg[2]/NET0131  ;
  input \wishbone_tx_fifo_read_pointer_reg[3]/NET0131  ;
  input \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  ;
  input \wishbone_tx_fifo_write_pointer_reg[1]/NET0131  ;
  input \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  ;
  input \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
  output \_al_n1  ;
  output \g215539/_0_  ;
  output \g215543/_0_  ;
  output \g215547/_0_  ;
  output \g215551/_0_  ;
  output \g215552/_0_  ;
  output \g215578/_0_  ;
  output \g215587/_1_  ;
  output \g215589/_1_  ;
  output \g215591/_1_  ;
  output \g215593/_1_  ;
  output \g215595/_1_  ;
  output \g215597/_1_  ;
  output \g215599/_1_  ;
  output \g215601/_1_  ;
  output \g215603/_1_  ;
  output \g215605/_1_  ;
  output \g215607/_1_  ;
  output \g215609/_1_  ;
  output \g215611/_1_  ;
  output \g215613/_1_  ;
  output \g215615/_1_  ;
  output \g215617/_1_  ;
  output \g215618/_0_  ;
  output \g215619/_0_  ;
  output \g215620/_0_  ;
  output \g215632/_1_  ;
  output \g215634/_0_  ;
  output \g215635/_0_  ;
  output \g215636/_0_  ;
  output \g215637/_0_  ;
  output \g215638/_0_  ;
  output \g215639/_0_  ;
  output \g215655/_1_  ;
  output \g215657/_1_  ;
  output \g215659/_1_  ;
  output \g215661/_1_  ;
  output \g215662/_0_  ;
  output \g215663/_0_  ;
  output \g215664/_0_  ;
  output \g215665/_0_  ;
  output \g215668/_0_  ;
  output \g215674/_0_  ;
  output \g215677/_0_  ;
  output \g215686/_0_  ;
  output \g215695/_0_  ;
  output \g215696/_0_  ;
  output \g215702/_1__syn_2  ;
  output \g215705/_0_  ;
  output \g215706/_0_  ;
  output \g215716/_0_  ;
  output \g215717/_0_  ;
  output \g215718/_0_  ;
  output \g215726/_0_  ;
  output \g215727/_0_  ;
  output \g215728/_0_  ;
  output \g215760/_0_  ;
  output \g215764/_0_  ;
  output \g215765/_0_  ;
  output \g215766/_0_  ;
  output \g215767/_3_  ;
  output \g215768/_3_  ;
  output \g215769/_3_  ;
  output \g215770/_3_  ;
  output \g215771/_3_  ;
  output \g215772/_3_  ;
  output \g215773/_3_  ;
  output \g215774/_3_  ;
  output \g215775/_3_  ;
  output \g215776/_3_  ;
  output \g215777/_3_  ;
  output \g215778/_3_  ;
  output \g215779/_3_  ;
  output \g215780/_3_  ;
  output \g215790/_0_  ;
  output \g215791/_0_  ;
  output \g215792/_0_  ;
  output \g215793/_0_  ;
  output \g215801/_0_  ;
  output \g215802/_0_  ;
  output \g215803/_0_  ;
  output \g215804/_0_  ;
  output \g215812/_0_  ;
  output \g215813/_0_  ;
  output \g215821/_0_  ;
  output \g215823/_0_  ;
  output \g215831/_0_  ;
  output \g215832/_0_  ;
  output \g215833/_0_  ;
  output \g215845/_0_  ;
  output \g215846/_0_  ;
  output \g215847/_0_  ;
  output \g215872/_0_  ;
  output \g215873/_0_  ;
  output \g215874/_0_  ;
  output \g215904/_0_  ;
  output \g215905/_0_  ;
  output \g215906/_0_  ;
  output \g215907/_0_  ;
  output \g215908/_0_  ;
  output \g215909/_0_  ;
  output \g215910/_0_  ;
  output \g215911/_0_  ;
  output \g215912/_0_  ;
  output \g215913/_0_  ;
  output \g215914/_0_  ;
  output \g215915/_0_  ;
  output \g215916/_0_  ;
  output \g215917/_0_  ;
  output \g215918/_0_  ;
  output \g215919/_0_  ;
  output \g215920/_0_  ;
  output \g215923/_0_  ;
  output \g215926/_0_  ;
  output \g215941/_0_  ;
  output \g215942/_0_  ;
  output \g215943/_0_  ;
  output \g215944/_0_  ;
  output \g215945/_0_  ;
  output \g215946/_0_  ;
  output \g215947/_0_  ;
  output \g215948/_0_  ;
  output \g215949/_0_  ;
  output \g215950/_0_  ;
  output \g215951/_0_  ;
  output \g215952/_0_  ;
  output \g215953/_0_  ;
  output \g215954/_0_  ;
  output \g215955/_0_  ;
  output \g215956/_0_  ;
  output \g215957/_0_  ;
  output \g215959/_00_  ;
  output \g215960/_0_  ;
  output \g215962/_0_  ;
  output \g215964/_0_  ;
  output \g215966/_0_  ;
  output \g215972/_0_  ;
  output \g216035/_0_  ;
  output \g216037/_0_  ;
  output \g216038/_0_  ;
  output \g216039/_0_  ;
  output \g216040/_0_  ;
  output \g216041/_0_  ;
  output \g216042/_0_  ;
  output \g216046/_0_  ;
  output \g216048/_0_  ;
  output \g216057/_0_  ;
  output \g216263/_0_  ;
  output \g216264/_0_  ;
  output \g216265/_0_  ;
  output \g216266/_0_  ;
  output \g216267/_0_  ;
  output \g216268/_0_  ;
  output \g216269/_0_  ;
  output \g216270/_0_  ;
  output \g216271/_0_  ;
  output \g216272/_0_  ;
  output \g216273/_0_  ;
  output \g216284/_0_  ;
  output \g216289/_0_  ;
  output \g216290/_0_  ;
  output \g216292/_0_  ;
  output \g216296/_0_  ;
  output \g216297/_0_  ;
  output \g216300/_0_  ;
  output \g216301/_0_  ;
  output \g216302/_0_  ;
  output \g216303/_0_  ;
  output \g216304/_0_  ;
  output \g216305/_0_  ;
  output \g216306/_0_  ;
  output \g216307/_0_  ;
  output \g216310/_3_  ;
  output \g216311/_3_  ;
  output \g216314/u3_syn_7  ;
  output \g216322/_3_  ;
  output \g216323/_3_  ;
  output \g216324/_3_  ;
  output \g216325/_3_  ;
  output \g216326/_3_  ;
  output \g216327/_3_  ;
  output \g216328/_3_  ;
  output \g216329/_3_  ;
  output \g216369/_0_  ;
  output \g216370/_0_  ;
  output \g216371/_0_  ;
  output \g216372/_0_  ;
  output \g216373/_0_  ;
  output \g216374/_0_  ;
  output \g216375/_0_  ;
  output \g216376/_0_  ;
  output \g216379/_0_  ;
  output \g216380/_0_  ;
  output \g216381/_0_  ;
  output \g216385/_0_  ;
  output \g216389/_0_  ;
  output \g216390/_0_  ;
  output \g216402/_0_  ;
  output \g216404/_0_  ;
  output \g216405/_0_  ;
  output \g216406/_0_  ;
  output \g216407/_0_  ;
  output \g216408/_0_  ;
  output \g216409/_0_  ;
  output \g216410/_0_  ;
  output \g216411/_0_  ;
  output \g216412/_0_  ;
  output \g216413/_0_  ;
  output \g216414/_0_  ;
  output \g216415/_0_  ;
  output \g216416/_0_  ;
  output \g216417/_0_  ;
  output \g216418/_0_  ;
  output \g216419/_0_  ;
  output \g216420/_0_  ;
  output \g216421/_0_  ;
  output \g216422/_0_  ;
  output \g216423/_0_  ;
  output \g216424/_0_  ;
  output \g216425/_0_  ;
  output \g216426/_0_  ;
  output \g216427/_0_  ;
  output \g216428/_0_  ;
  output \g216429/_0_  ;
  output \g216430/_0_  ;
  output \g216431/_0_  ;
  output \g216432/_0_  ;
  output \g216433/_0_  ;
  output \g216434/_0_  ;
  output \g216435/_0_  ;
  output \g216436/_0_  ;
  output \g216437/_0_  ;
  output \g216438/_0_  ;
  output \g216439/_3_  ;
  output \g216447/_3_  ;
  output \g216448/_3_  ;
  output \g216452/_0_  ;
  output \g216453/_0_  ;
  output \g216454/_0_  ;
  output \g216455/_0_  ;
  output \g216456/_0_  ;
  output \g216457/_0_  ;
  output \g216458/_3_  ;
  output \g216459/_3_  ;
  output \g216461/_3_  ;
  output \g216462/_3_  ;
  output \g216463/_3_  ;
  output \g216464/_3_  ;
  output \g216465/_3_  ;
  output \g216466/_0_  ;
  output \g216467/_3_  ;
  output \g216468/_3_  ;
  output \g216469/_3_  ;
  output \g216470/_3_  ;
  output \g216471/_3_  ;
  output \g216473/_3_  ;
  output \g216474/_3_  ;
  output \g216475/_3_  ;
  output \g216476/_3_  ;
  output \g216477/_3_  ;
  output \g216478/_0_  ;
  output \g216479/_3_  ;
  output \g216480/_3_  ;
  output \g216481/_3_  ;
  output \g216492/_0_  ;
  output \g216494/_0_  ;
  output \g216495/_3_  ;
  output \g216496/_3_  ;
  output \g216498/_3_  ;
  output \g216499/_3_  ;
  output \g216500/_3_  ;
  output \g216513/_3_  ;
  output \g216514/_3_  ;
  output \g216515/_3_  ;
  output \g216516/_3_  ;
  output \g216517/_3_  ;
  output \g216518/_3_  ;
  output \g216519/_3_  ;
  output \g216520/_3_  ;
  output \g216521/_3_  ;
  output \g216522/_3_  ;
  output \g216523/_3_  ;
  output \g216524/_3_  ;
  output \g216525/_3_  ;
  output \g216526/_3_  ;
  output \g216527/_3_  ;
  output \g216528/_3_  ;
  output \g216529/_3_  ;
  output \g216530/_3_  ;
  output \g216531/_3_  ;
  output \g216532/_3_  ;
  output \g216533/_3_  ;
  output \g216534/_3_  ;
  output \g216535/_3_  ;
  output \g216536/_3_  ;
  output \g216537/_3_  ;
  output \g216538/_3_  ;
  output \g216555/_3_  ;
  output \g216556/_3_  ;
  output \g216557/_3_  ;
  output \g216560/_3_  ;
  output \g216561/_3_  ;
  output \g216562/_3_  ;
  output \g216563/_3_  ;
  output \g216564/_3_  ;
  output \g216565/_3_  ;
  output \g216566/_3_  ;
  output \g216567/_3_  ;
  output \g216568/_3_  ;
  output \g216569/_3_  ;
  output \g216570/_3_  ;
  output \g216571/_3_  ;
  output \g216575/_3_  ;
  output \g216576/_3_  ;
  output \g216577/_3_  ;
  output \g216578/_3_  ;
  output \g216579/_3_  ;
  output \g216580/_3_  ;
  output \g216581/_3_  ;
  output \g216582/_3_  ;
  output \g216583/_3_  ;
  output \g216586/_3_  ;
  output \g216587/_3_  ;
  output \g216588/_3_  ;
  output \g216589/_3_  ;
  output \g216590/_3_  ;
  output \g216591/_3_  ;
  output \g216592/_3_  ;
  output \g216593/_3_  ;
  output \g216594/_3_  ;
  output \g216595/_3_  ;
  output \g216600/_3_  ;
  output \g216683/_0_  ;
  output \g216689/_0_  ;
  output \g216693/_0_  ;
  output \g216694/_0_  ;
  output \g216727/_0_  ;
  output \g216728/_0_  ;
  output \g216729/_0_  ;
  output \g216732/_0_  ;
  output \g216733/_0_  ;
  output \g216734/_0_  ;
  output \g216735/_0_  ;
  output \g216736/_0_  ;
  output \g216737/_0_  ;
  output \g216738/_0_  ;
  output \g216739/_0_  ;
  output \g216740/_0_  ;
  output \g216741/_0_  ;
  output \g216742/_0_  ;
  output \g216743/_0_  ;
  output \g216744/_0_  ;
  output \g216745/_0_  ;
  output \g216746/_0_  ;
  output \g216748/_0_  ;
  output \g216751/_0_  ;
  output \g216754/_0_  ;
  output \g216762/_0_  ;
  output \g216934/_2_  ;
  output \g216952/_0_  ;
  output \g216955/_0_  ;
  output \g216969/_0_  ;
  output \g216979/_0_  ;
  output \g216984/_0_  ;
  output \g216996/_0_  ;
  output \g217002/_0_  ;
  output \g217014/_0_  ;
  output \g217015/_0_  ;
  output \g217016/_0_  ;
  output \g217017/_0_  ;
  output \g217018/_0_  ;
  output \g217019/_0_  ;
  output \g217023/_0_  ;
  output \g217116/_0_  ;
  output \g217146/_3_  ;
  output \g217149/_0_  ;
  output \g217151/_0_  ;
  output \g217160/_0_  ;
  output \g217167/_0_  ;
  output \g217168/_0_  ;
  output \g217169/_0_  ;
  output \g217170/_0_  ;
  output \g217171/_0_  ;
  output \g217172/_0_  ;
  output \g217173/_0_  ;
  output \g217174/_0_  ;
  output \g217175/_0_  ;
  output \g217176/_0_  ;
  output \g217177/_0_  ;
  output \g217178/_0_  ;
  output \g217179/_0_  ;
  output \g217180/_0_  ;
  output \g217181/_0_  ;
  output \g217182/_0_  ;
  output \g217183/_0_  ;
  output \g217187/_0_  ;
  output \g217188/_0_  ;
  output \g217189/_0_  ;
  output \g217193/_0_  ;
  output \g217194/_0_  ;
  output \g217195/_0_  ;
  output \g217196/_0_  ;
  output \g217202/_0_  ;
  output \g217205/_0_  ;
  output \g217206/_0_  ;
  output \g217207/_0_  ;
  output \g217208/_0_  ;
  output \g217209/_0_  ;
  output \g217210/_0_  ;
  output \g217211/_0_  ;
  output \g217212/_0_  ;
  output \g217213/_0_  ;
  output \g217214/_0_  ;
  output \g217215/_0_  ;
  output \g217216/_0_  ;
  output \g217217/_0_  ;
  output \g217218/_0_  ;
  output \g217219/_0_  ;
  output \g217220/_0_  ;
  output \g217223/_0_  ;
  output \g217231/_0_  ;
  output \g217237/_0_  ;
  output \g217238/_0_  ;
  output \g217242/_0_  ;
  output \g217243/_0_  ;
  output \g217250/_3_  ;
  output \g217251/_3_  ;
  output \g217252/_3_  ;
  output \g217253/_3_  ;
  output \g217254/_3_  ;
  output \g217255/_3_  ;
  output \g217256/_3_  ;
  output \g217257/_3_  ;
  output \g217258/_3_  ;
  output \g217259/_3_  ;
  output \g217260/_3_  ;
  output \g217261/_3_  ;
  output \g217262/_3_  ;
  output \g217263/_3_  ;
  output \g217264/_3_  ;
  output \g217265/_3_  ;
  output \g217266/_3_  ;
  output \g217267/_3_  ;
  output \g217268/_3_  ;
  output \g217269/_3_  ;
  output \g217270/_3_  ;
  output \g217271/_3_  ;
  output \g217272/_3_  ;
  output \g217273/_3_  ;
  output \g217274/_3_  ;
  output \g217275/_3_  ;
  output \g217276/_3_  ;
  output \g217277/_3_  ;
  output \g217278/_3_  ;
  output \g217279/_3_  ;
  output \g217280/_3_  ;
  output \g217281/_3_  ;
  output \g217282/_3_  ;
  output \g217283/_3_  ;
  output \g217284/_3_  ;
  output \g217285/_3_  ;
  output \g217286/_3_  ;
  output \g217287/_3_  ;
  output \g217288/_3_  ;
  output \g217289/_3_  ;
  output \g217290/_3_  ;
  output \g217291/_3_  ;
  output \g217292/_3_  ;
  output \g217293/_3_  ;
  output \g217294/_3_  ;
  output \g217295/_3_  ;
  output \g217296/_3_  ;
  output \g217297/_3_  ;
  output \g217298/_3_  ;
  output \g217299/_3_  ;
  output \g217300/_3_  ;
  output \g217301/_3_  ;
  output \g217302/_3_  ;
  output \g217303/_3_  ;
  output \g217304/_3_  ;
  output \g217305/_3_  ;
  output \g217306/_3_  ;
  output \g217307/_3_  ;
  output \g217308/_3_  ;
  output \g217309/_3_  ;
  output \g217310/_3_  ;
  output \g217311/_3_  ;
  output \g217312/_3_  ;
  output \g217313/_3_  ;
  output \g217318/_0_  ;
  output \g217662/_0_  ;
  output \g217663/_0_  ;
  output \g217682/_0_  ;
  output \g217697/_0_  ;
  output \g217698/_0_  ;
  output \g217699/_0_  ;
  output \g217700/_0_  ;
  output \g217701/_0_  ;
  output \g217705/_0_  ;
  output \g217711/_0_  ;
  output \g217747/_0_  ;
  output \g217753/_00_  ;
  output \g217775/_0_  ;
  output \g217781/_0_  ;
  output \g217784/_0_  ;
  output \g217785/_0_  ;
  output \g217786/_0_  ;
  output \g217787/_0_  ;
  output \g217788/_0_  ;
  output \g217790/_0_  ;
  output \g217815/_0_  ;
  output \g217817/_0_  ;
  output \g218145/_0_  ;
  output \g218148/_0_  ;
  output \g218150/_0_  ;
  output \g218167/_0_  ;
  output \g218168/_0_  ;
  output \g218234/_0_  ;
  output \g218235/_0_  ;
  output \g218236/_0_  ;
  output \g218238/_0_  ;
  output \g218242/_0_  ;
  output \g218332/_0_  ;
  output \g218335/_0_  ;
  output \g218336/_0_  ;
  output \g218337/_0_  ;
  output \g218338/_0_  ;
  output \g218339/_0_  ;
  output \g218340/_0_  ;
  output \g218341/_0_  ;
  output \g218342/_0_  ;
  output \g218343/_0_  ;
  output \g218344/_0_  ;
  output \g218345/_0_  ;
  output \g218346/_0_  ;
  output \g218347/_0_  ;
  output \g218348/_0_  ;
  output \g218349/_0_  ;
  output \g218350/_0_  ;
  output \g218351/_0_  ;
  output \g218352/_0_  ;
  output \g218353/_0_  ;
  output \g218354/_0_  ;
  output \g218355/_0_  ;
  output \g218356/_0_  ;
  output \g218357/_0_  ;
  output \g218358/_0_  ;
  output \g218359/_0_  ;
  output \g218360/_0_  ;
  output \g218398/_3_  ;
  output \g218430/_0_  ;
  output \g218440/_0_  ;
  output \g218452/u3_syn_4  ;
  output \g218495/u3_syn_4  ;
  output \g218517/u3_syn_4  ;
  output \g218554/u3_syn_4  ;
  output \g218575/u3_syn_4  ;
  output \g218600/u3_syn_4  ;
  output \g218621/u3_syn_4  ;
  output \g218638/u3_syn_4  ;
  output \g218659/u3_syn_4  ;
  output \g218673/u3_syn_4  ;
  output \g218707/u3_syn_4  ;
  output \g218735/_3_  ;
  output \g219186/_0_  ;
  output \g219187/_0_  ;
  output \g219188/_0_  ;
  output \g219189/_0_  ;
  output \g219190/_0_  ;
  output \g219196/_0_  ;
  output \g219198/_0_  ;
  output \g219199/_0_  ;
  output \g219200/_0_  ;
  output \g219308/_0_  ;
  output \g219314/_0_  ;
  output \g219326/_0_  ;
  output \g219328/_0_  ;
  output \g219348/_0_  ;
  output \g219351/_0_  ;
  output \g219363/_0_  ;
  output \g219364/_0_  ;
  output \g219365/_0_  ;
  output \g219366/_0_  ;
  output \g219367/_0_  ;
  output \g219368/_0_  ;
  output \g219369/_0_  ;
  output \g219376/_0_  ;
  output \g219381/_0_  ;
  output \g219382/_0_  ;
  output \g219384/_0_  ;
  output \g219385/_0_  ;
  output \g219391/_0_  ;
  output \g219394/_0_  ;
  output \g219395/_0_  ;
  output \g219396/_0_  ;
  output \g219397/_0_  ;
  output \g219398/_0_  ;
  output \g219399/_0_  ;
  output \g219400/_0_  ;
  output \g219401/_0_  ;
  output \g219402/_0_  ;
  output \g219403/_0_  ;
  output \g219404/_0_  ;
  output \g219405/_0_  ;
  output \g219406/_0_  ;
  output \g219407/_0_  ;
  output \g219408/_0_  ;
  output \g219409/_0_  ;
  output \g219410/_0_  ;
  output \g219411/_0_  ;
  output \g219412/_0_  ;
  output \g219413/_0_  ;
  output \g219414/_0_  ;
  output \g219415/_0_  ;
  output \g219416/_0_  ;
  output \g219417/_0_  ;
  output \g219418/_0_  ;
  output \g219419/_0_  ;
  output \g219420/_0_  ;
  output \g219421/_0_  ;
  output \g219422/_0_  ;
  output \g219423/_0_  ;
  output \g219424/_0_  ;
  output \g219425/_0_  ;
  output \g219426/_0_  ;
  output \g219427/_0_  ;
  output \g219428/_0_  ;
  output \g219429/_0_  ;
  output \g219430/_0_  ;
  output \g219431/_0_  ;
  output \g219432/_0_  ;
  output \g219433/_0_  ;
  output \g219434/_0_  ;
  output \g219435/_0_  ;
  output \g219436/_0_  ;
  output \g219437/_0_  ;
  output \g219438/_0_  ;
  output \g219439/_0_  ;
  output \g219440/_0_  ;
  output \g219441/_0_  ;
  output \g219442/_0_  ;
  output \g219443/_0_  ;
  output \g219444/_0_  ;
  output \g219445/_0_  ;
  output \g219446/_0_  ;
  output \g219447/_0_  ;
  output \g219449/_0_  ;
  output \g219450/_0_  ;
  output \g219451/_0_  ;
  output \g219452/_0_  ;
  output \g219453/_0_  ;
  output \g219454/_0_  ;
  output \g219455/_0_  ;
  output \g219456/_0_  ;
  output \g219457/_0_  ;
  output \g219458/_0_  ;
  output \g219464/u3_syn_7  ;
  output \g219496/u3_syn_4  ;
  output \g219512/u3_syn_4  ;
  output \g219526/u3_syn_4  ;
  output \g219549/u3_syn_4  ;
  output \g219571/u3_syn_4  ;
  output \g219588/u3_syn_4  ;
  output \g219603/u3_syn_4  ;
  output \g219621/u3_syn_4  ;
  output \g219636/_3_  ;
  output \g219652/u3_syn_4  ;
  output \g219676/_3_  ;
  output \g219686/_0_  ;
  output \g219689/_0_  ;
  output \g219694/_3_  ;
  output \g220062/_0_  ;
  output \g220068/_0_  ;
  output \g220069/_0_  ;
  output \g220072/_0_  ;
  output \g220084/_0_  ;
  output \g220149/_0_  ;
  output \g220162/_0_  ;
  output \g220317/_0_  ;
  output \g220360/_2_  ;
  output \g220368/_2_  ;
  output \g220369/_0_  ;
  output \g220370/_0_  ;
  output \g220371/_0_  ;
  output \g220372/_0_  ;
  output \g220376/_0_  ;
  output \g220390/_0_  ;
  output \g220395/_0_  ;
  output \g220499/_0_  ;
  output \g220500/_0_  ;
  output \g220501/_0_  ;
  output \g220502/_0_  ;
  output \g220503/_0_  ;
  output \g220504/_0_  ;
  output \g220505/_0_  ;
  output \g220506/_0_  ;
  output \g220507/_0_  ;
  output \g220508/_0_  ;
  output \g220509/_0_  ;
  output \g220510/_0_  ;
  output \g220511/_0_  ;
  output \g220512/_0_  ;
  output \g220513/_0_  ;
  output \g220514/_0_  ;
  output \g220515/_0_  ;
  output \g220516/_0_  ;
  output \g220517/_0_  ;
  output \g220518/_0_  ;
  output \g220519/_0_  ;
  output \g220520/_0_  ;
  output \g220521/_0_  ;
  output \g220522/_0_  ;
  output \g220523/_0_  ;
  output \g220524/_0_  ;
  output \g220525/_0_  ;
  output \g220526/_0_  ;
  output \g220527/_0_  ;
  output \g220528/_0_  ;
  output \g220529/_0_  ;
  output \g220530/_0_  ;
  output \g220531/_0_  ;
  output \g220532/_0_  ;
  output \g220533/_0_  ;
  output \g220534/_0_  ;
  output \g220535/_0_  ;
  output \g220557/_0_  ;
  output \g220558/_0_  ;
  output \g220559/_0_  ;
  output \g220560/_0_  ;
  output \g220561/_0_  ;
  output \g220562/_0_  ;
  output \g220563/_0_  ;
  output \g220564/_0_  ;
  output \g220565/_0_  ;
  output \g220566/_0_  ;
  output \g220567/_0_  ;
  output \g220568/_0_  ;
  output \g220569/_0_  ;
  output \g220570/_0_  ;
  output \g220571/_0_  ;
  output \g220572/_0_  ;
  output \g220573/_0_  ;
  output \g220574/_0_  ;
  output \g220575/_0_  ;
  output \g220576/_0_  ;
  output \g220577/_0_  ;
  output \g220578/_0_  ;
  output \g220579/_0_  ;
  output \g220580/_0_  ;
  output \g220581/_0_  ;
  output \g220582/_0_  ;
  output \g220583/_0_  ;
  output \g220584/_0_  ;
  output \g220585/_0_  ;
  output \g220586/_0_  ;
  output \g220587/_0_  ;
  output \g220588/_0_  ;
  output \g220589/_0_  ;
  output \g220590/_0_  ;
  output \g220591/_0_  ;
  output \g220592/_0_  ;
  output \g220593/_0_  ;
  output \g220594/_0_  ;
  output \g220595/_0_  ;
  output \g220596/_0_  ;
  output \g220597/_0_  ;
  output \g220598/_0_  ;
  output \g220599/_0_  ;
  output \g220600/_0_  ;
  output \g220601/_0_  ;
  output \g220602/_0_  ;
  output \g220603/_0_  ;
  output \g220604/_0_  ;
  output \g220605/_0_  ;
  output \g220606/_0_  ;
  output \g220607/_0_  ;
  output \g220608/_0_  ;
  output \g220609/_0_  ;
  output \g220610/_0_  ;
  output \g220611/_0_  ;
  output \g220612/_0_  ;
  output \g220613/_0_  ;
  output \g220614/_0_  ;
  output \g220615/_0_  ;
  output \g220616/_0_  ;
  output \g220617/_0_  ;
  output \g220618/_0_  ;
  output \g220619/_0_  ;
  output \g220620/_0_  ;
  output \g220621/_0_  ;
  output \g220622/_0_  ;
  output \g220623/_0_  ;
  output \g220624/_0_  ;
  output \g220625/_0_  ;
  output \g220626/_0_  ;
  output \g220627/_0_  ;
  output \g220628/_0_  ;
  output \g220629/_0_  ;
  output \g220630/_0_  ;
  output \g220631/_0_  ;
  output \g220632/_0_  ;
  output \g220633/_0_  ;
  output \g220634/_0_  ;
  output \g220635/_0_  ;
  output \g220636/_0_  ;
  output \g220637/_0_  ;
  output \g220638/_0_  ;
  output \g220639/_0_  ;
  output \g220640/_0_  ;
  output \g220641/_0_  ;
  output \g220642/_0_  ;
  output \g220643/_0_  ;
  output \g220644/_0_  ;
  output \g220645/_0_  ;
  output \g220646/_0_  ;
  output \g220647/_0_  ;
  output \g220648/_0_  ;
  output \g220649/_0_  ;
  output \g220650/_0_  ;
  output \g220651/_0_  ;
  output \g220652/_0_  ;
  output \g220653/_0_  ;
  output \g220654/_0_  ;
  output \g220655/_0_  ;
  output \g220656/_0_  ;
  output \g220657/_0_  ;
  output \g220658/_0_  ;
  output \g220659/_0_  ;
  output \g220660/_0_  ;
  output \g220661/_0_  ;
  output \g220662/_0_  ;
  output \g220663/_0_  ;
  output \g220664/_0_  ;
  output \g220665/_0_  ;
  output \g220666/_0_  ;
  output \g220674/_0_  ;
  output \g220679/u3_syn_7  ;
  output \g220711/u3_syn_4  ;
  output \g220726/u3_syn_4  ;
  output \g220739/u3_syn_4  ;
  output \g220751/u3_syn_4  ;
  output \g220759/u3_syn_4  ;
  output \g220773/u3_syn_4  ;
  output \g220782/u3_syn_4  ;
  output \g220805/u3_syn_4  ;
  output \g220828/u3_syn_4  ;
  output \g220921/_0_  ;
  output \g220930/u3_syn_4  ;
  output \g220949/_3_  ;
  output \g220994/_3_  ;
  output \g221207/_0_  ;
  output \g221213/_0_  ;
  output \g221223/_0_  ;
  output \g221224/_0_  ;
  output \g221225/_0_  ;
  output \g221226/_0_  ;
  output \g221231/_0_  ;
  output \g221232/_0_  ;
  output \g221234/_0_  ;
  output \g221235/_0_  ;
  output \g221246/_2_  ;
  output \g221249/_2_  ;
  output \g221265/_0_  ;
  output \g221287/_0_  ;
  output \g221325/_0_  ;
  output \g221326/_0_  ;
  output \g221447/_0_  ;
  output \g221449/_0_  ;
  output \g221452/_0_  ;
  output \g221469/_0_  ;
  output \g221473/_0_  ;
  output \g221503/_0_  ;
  output \g221510/_0_  ;
  output \g221512/_0_  ;
  output \g221516/_0_  ;
  output \g221517/_0_  ;
  output \g221524/_0_  ;
  output \g221530/_0_  ;
  output \g221592/_0_  ;
  output \g221593/_0_  ;
  output \g221634/u3_syn_4  ;
  output \g221669/u3_syn_4  ;
  output \g221789/u3_syn_4  ;
  output \g221813/u3_syn_4  ;
  output \g221829/u3_syn_4  ;
  output \g221861/u3_syn_4  ;
  output \g221876/_0_  ;
  output \g221935/_0_  ;
  output \g221944/_3_  ;
  output \g230200/_0_  ;
  output \g230201/_0_  ;
  output \g230205/_0_  ;
  output \g230295/_0_  ;
  output \g230297/_0_  ;
  output \g230298/_0_  ;
  output \g230300/_0_  ;
  output \g230302/_0_  ;
  output \g230303/_0_  ;
  output \g230343/_0_  ;
  output \g230368/_0_  ;
  output \g230511/_0_  ;
  output \g230531/_0_  ;
  output \g230635/_2_  ;
  output \g230661/_0_  ;
  output \g230715/_1__syn_2  ;
  output \g230731/_0_  ;
  output \g230766/_0_  ;
  output \g230784/_0_  ;
  output \g230785/_0_  ;
  output \g230786/_0_  ;
  output \g230787/_0_  ;
  output \g230797/_0_  ;
  output \g230798/_0_  ;
  output \g230803/_0_  ;
  output \g230804/_00_  ;
  output \g230805/_00_  ;
  output \g230806/_00_  ;
  output \g230807/_00_  ;
  output \g230808/_00_  ;
  output \g230809/_00_  ;
  output \g230815/_0_  ;
  output \g230816/_2_  ;
  output \g230817/_2_  ;
  output \g230829/_0_  ;
  output \g230834/_0_  ;
  output \g230835/_0_  ;
  output \g230836/_0_  ;
  output \g230837/_0_  ;
  output \g230844/_0_  ;
  output \g230863/_3_  ;
  output \g230864/_3_  ;
  output \g230870/_0_  ;
  output \g230988/_3_  ;
  output \g231010/_3_  ;
  output \g231016/_3_  ;
  output \g231042/_3_  ;
  output \g231471/_0_  ;
  output \g231472/_0_  ;
  output \g231476/_3_  ;
  output \g231480/_3_  ;
  output \g231484/_3_  ;
  output \g231504/_0_  ;
  output \g231532/_0_  ;
  output \g231542/_0_  ;
  output \g231560/_1_  ;
  output \g231578/_1_  ;
  output \g231580/_0_  ;
  output \g231590/_1__syn_2  ;
  output \g231615/_0_  ;
  output \g231623/_1_  ;
  output \g231634/_2_  ;
  output \g231635/_0_  ;
  output \g231638/_2_  ;
  output \g231640/_0_  ;
  output \g231653/_2_  ;
  output \g231787/_0_  ;
  output \g231931/_0_  ;
  output \g231939/_3_  ;
  output \g231940/_0_  ;
  output \g231951/_0_  ;
  output \g231955/_0_  ;
  output \g231956/_0_  ;
  output \g231959/_2_  ;
  output \g231960/_0_  ;
  output \g231964/_0_  ;
  output \g231965/_0_  ;
  output \g231975/_0_  ;
  output \g231986/_1_  ;
  output \g231987/_1_  ;
  output \g231989/_1_  ;
  output \g231990/_1_  ;
  output \g231991/_0_  ;
  output \g231992/_0_  ;
  output \g231995/_0_  ;
  output \g231998/_0_  ;
  output \g231999/_0_  ;
  output \g232002/_3_  ;
  output \g232035/u3_syn_4  ;
  output \g232038/u3_syn_4  ;
  output \g232046/u3_syn_4  ;
  output \g232054/u3_syn_4  ;
  output \g232062/u3_syn_4  ;
  output \g232070/u3_syn_4  ;
  output \g232078/u3_syn_4  ;
  output \g232079/u3_syn_4  ;
  output \g232087/u3_syn_4  ;
  output \g232096/u3_syn_4  ;
  output \g232104/u3_syn_4  ;
  output \g232112/u3_syn_4  ;
  output \g232120/u3_syn_4  ;
  output \g232128/u3_syn_4  ;
  output \g232136/u3_syn_4  ;
  output \g232144/u3_syn_4  ;
  output \g232152/u3_syn_4  ;
  output \g232161/u3_syn_4  ;
  output \g232169/u3_syn_4  ;
  output \g232177/u3_syn_4  ;
  output \g232185/u3_syn_4  ;
  output \g232186/u3_syn_4  ;
  output \g232194/u3_syn_4  ;
  output \g232202/u3_syn_4  ;
  output \g232210/u3_syn_4  ;
  output \g232218/u3_syn_4  ;
  output \g232226/u3_syn_4  ;
  output \g232234/u3_syn_4  ;
  output \g232242/u3_syn_4  ;
  output \g232251/u3_syn_4  ;
  output \g232259/u3_syn_4  ;
  output \g232267/u3_syn_4  ;
  output \g232275/u3_syn_4  ;
  output \g232283/u3_syn_4  ;
  output \g232291/u3_syn_4  ;
  output \g232299/u3_syn_4  ;
  output \g232307/u3_syn_4  ;
  output \g232315/u3_syn_4  ;
  output \g232324/u3_syn_4  ;
  output \g232332/u3_syn_4  ;
  output \g232341/u3_syn_4  ;
  output \g232349/u3_syn_4  ;
  output \g232357/u3_syn_4  ;
  output \g232366/u3_syn_4  ;
  output \g232374/u3_syn_4  ;
  output \g232382/u3_syn_4  ;
  output \g232390/u3_syn_4  ;
  output \g232398/u3_syn_4  ;
  output \g232406/u3_syn_4  ;
  output \g232414/u3_syn_4  ;
  output \g232422/u3_syn_4  ;
  output \g232427/u3_syn_4  ;
  output \g232431/u3_syn_4  ;
  output \g232439/u3_syn_4  ;
  output \g232444/u3_syn_4  ;
  output \g232452/u3_syn_4  ;
  output \g232461/u3_syn_4  ;
  output \g232471/u3_syn_4  ;
  output \g232479/u3_syn_4  ;
  output \g232487/u3_syn_4  ;
  output \g232495/u3_syn_4  ;
  output \g232503/u3_syn_4  ;
  output \g232506/u3_syn_4  ;
  output \g232514/u3_syn_4  ;
  output \g232527/u3_syn_4  ;
  output \g232530/u3_syn_4  ;
  output \g232536/u3_syn_4  ;
  output \g232544/u3_syn_4  ;
  output \g232551/u3_syn_4  ;
  output \g232557/u3_syn_4  ;
  output \g232568/u3_syn_4  ;
  output \g232576/u3_syn_4  ;
  output \g232585/u3_syn_4  ;
  output \g232593/u3_syn_4  ;
  output \g232597/u3_syn_4  ;
  output \g232609/u3_syn_4  ;
  output \g232617/u3_syn_4  ;
  output \g232625/u3_syn_4  ;
  output \g232633/u3_syn_4  ;
  output \g232641/u3_syn_4  ;
  output \g232649/u3_syn_4  ;
  output \g232657/u3_syn_4  ;
  output \g232665/u3_syn_4  ;
  output \g232673/u3_syn_4  ;
  output \g232681/u3_syn_4  ;
  output \g232689/u3_syn_4  ;
  output \g232697/u3_syn_4  ;
  output \g232705/u3_syn_4  ;
  output \g232713/u3_syn_4  ;
  output \g232717/u3_syn_4  ;
  output \g232729/u3_syn_4  ;
  output \g232737/u3_syn_4  ;
  output \g232745/u3_syn_4  ;
  output \g232749/u3_syn_4  ;
  output \g232761/u3_syn_4  ;
  output \g232768/u3_syn_4  ;
  output \g232777/u3_syn_4  ;
  output \g232785/u3_syn_4  ;
  output \g232793/u3_syn_4  ;
  output \g232801/u3_syn_4  ;
  output \g232809/u3_syn_4  ;
  output \g232815/u3_syn_4  ;
  output \g232823/u3_syn_4  ;
  output \g232833/u3_syn_4  ;
  output \g232841/u3_syn_4  ;
  output \g232846/u3_syn_4  ;
  output \g232851/u3_syn_4  ;
  output \g232865/u3_syn_4  ;
  output \g232873/u3_syn_4  ;
  output \g232881/u3_syn_4  ;
  output \g232882/u3_syn_4  ;
  output \g232895/u3_syn_4  ;
  output \g232904/u3_syn_4  ;
  output \g232913/u3_syn_4  ;
  output \g232921/u3_syn_4  ;
  output \g232928/u3_syn_4  ;
  output \g232934/u3_syn_4  ;
  output \g232945/u3_syn_4  ;
  output \g232953/u3_syn_4  ;
  output \g232954/u3_syn_4  ;
  output \g232969/u3_syn_4  ;
  output \g232977/u3_syn_4  ;
  output \g232981/u3_syn_4  ;
  output \g232993/u3_syn_4  ;
  output \g232995/u3_syn_4  ;
  output \g233009/u3_syn_4  ;
  output \g233017/u3_syn_4  ;
  output \g233025/u3_syn_4  ;
  output \g233033/u3_syn_4  ;
  output \g233041/u3_syn_4  ;
  output \g233047/u3_syn_4  ;
  output \g233057/u3_syn_4  ;
  output \g233065/u3_syn_4  ;
  output \g233073/u3_syn_4  ;
  output \g233081/u3_syn_4  ;
  output \g233087/u3_syn_4  ;
  output \g233097/u3_syn_4  ;
  output \g233105/u3_syn_4  ;
  output \g233113/u3_syn_4  ;
  output \g233121/u3_syn_4  ;
  output \g233128/u3_syn_4  ;
  output \g233134/u3_syn_4  ;
  output \g233144/u3_syn_4  ;
  output \g233153/u3_syn_4  ;
  output \g233161/u3_syn_4  ;
  output \g233169/u3_syn_4  ;
  output \g233177/u3_syn_4  ;
  output \g233185/u3_syn_4  ;
  output \g233193/u3_syn_4  ;
  output \g233201/u3_syn_4  ;
  output \g233209/u3_syn_4  ;
  output \g233217/u3_syn_4  ;
  output \g233219/u3_syn_4  ;
  output \g233229/u3_syn_4  ;
  output \g233241/u3_syn_4  ;
  output \g233249/u3_syn_4  ;
  output \g233257/u3_syn_4  ;
  output \g233265/u3_syn_4  ;
  output \g233273/u3_syn_4  ;
  output \g233281/u3_syn_4  ;
  output \g233289/u3_syn_4  ;
  output \g233297/u3_syn_4  ;
  output \g233305/u3_syn_4  ;
  output \g233313/u3_syn_4  ;
  output \g233321/u3_syn_4  ;
  output \g233329/u3_syn_4  ;
  output \g233337/u3_syn_4  ;
  output \g233345/u3_syn_4  ;
  output \g233353/u3_syn_4  ;
  output \g233361/u3_syn_4  ;
  output \g233369/u3_syn_4  ;
  output \g233377/u3_syn_4  ;
  output \g233382/u3_syn_4  ;
  output \g233392/u3_syn_4  ;
  output \g233394/u3_syn_4  ;
  output \g233409/u3_syn_4  ;
  output \g233417/u3_syn_4  ;
  output \g233425/u3_syn_4  ;
  output \g233433/u3_syn_4  ;
  output \g233441/u3_syn_4  ;
  output \g233449/u3_syn_4  ;
  output \g233453/u3_syn_4  ;
  output \g233465/u3_syn_4  ;
  output \g233473/u3_syn_4  ;
  output \g233481/u3_syn_4  ;
  output \g233489/u3_syn_4  ;
  output \g233497/u3_syn_4  ;
  output \g233505/u3_syn_4  ;
  output \g233513/u3_syn_4  ;
  output \g233516/u3_syn_4  ;
  output \g233529/u3_syn_4  ;
  output \g233531/u3_syn_4  ;
  output \g233546/u3_syn_4  ;
  output \g233554/u3_syn_4  ;
  output \g233562/u3_syn_4  ;
  output \g233570/u3_syn_4  ;
  output \g233578/u3_syn_4  ;
  output \g233586/u3_syn_4  ;
  output \g233594/u3_syn_4  ;
  output \g233602/u3_syn_4  ;
  output \g233603/u3_syn_4  ;
  output \g233618/u3_syn_4  ;
  output \g233626/u3_syn_4  ;
  output \g233634/u3_syn_4  ;
  output \g233642/u3_syn_4  ;
  output \g233650/u3_syn_4  ;
  output \g233658/u3_syn_4  ;
  output \g233666/u3_syn_4  ;
  output \g233674/u3_syn_4  ;
  output \g233682/u3_syn_4  ;
  output \g233690/u3_syn_4  ;
  output \g233698/u3_syn_4  ;
  output \g233706/u3_syn_4  ;
  output \g233714/u3_syn_4  ;
  output \g233722/u3_syn_4  ;
  output \g233730/u3_syn_4  ;
  output \g233738/u3_syn_4  ;
  output \g233746/u3_syn_4  ;
  output \g233754/u3_syn_4  ;
  output \g233762/u3_syn_4  ;
  output \g233770/u3_syn_4  ;
  output \g233778/u3_syn_4  ;
  output \g233783/u3_syn_4  ;
  output \g233794/u3_syn_4  ;
  output \g233802/u3_syn_4  ;
  output \g233806/u3_syn_4  ;
  output \g233818/u3_syn_4  ;
  output \g233826/u3_syn_4  ;
  output \g233828/u3_syn_4  ;
  output \g233838/u3_syn_4  ;
  output \g233850/u3_syn_4  ;
  output \g233858/u3_syn_4  ;
  output \g233860/u3_syn_4  ;
  output \g233870/u3_syn_4  ;
  output \g233881/u3_syn_4  ;
  output \g233890/u3_syn_4  ;
  output \g233899/u3_syn_4  ;
  output \g233908/u3_syn_4  ;
  output \g233917/u3_syn_4  ;
  output \g233919/u3_syn_4  ;
  output \g233927/u3_syn_4  ;
  output \g233935/u3_syn_4  ;
  output \g233943/u3_syn_4  ;
  output \g233945/u3_syn_4  ;
  output \g233953/u3_syn_4  ;
  output \g233961/u3_syn_4  ;
  output \g233969/u3_syn_4  ;
  output \g233977/u3_syn_4  ;
  output \g233985/u3_syn_4  ;
  output \g233993/u3_syn_4  ;
  output \g234001/u3_syn_4  ;
  output \g234008/u3_syn_4  ;
  output \g234009/u3_syn_4  ;
  output \g234024/u3_syn_4  ;
  output \g234032/u3_syn_4  ;
  output \g234038/u3_syn_4  ;
  output \g234056/u3_syn_4  ;
  output \g234063/u3_syn_4  ;
  output \g234071/u3_syn_4  ;
  output \g234079/u3_syn_4  ;
  output \g234098/u3_syn_4  ;
  output \g234106/u3_syn_4  ;
  output \g234114/u3_syn_4  ;
  output \g234122/u3_syn_4  ;
  output \g234130/u3_syn_4  ;
  output \g234138/u3_syn_4  ;
  output \g234145/u3_syn_4  ;
  output \g234156/u3_syn_4  ;
  output \g234162/u3_syn_4  ;
  output \g234171/u3_syn_4  ;
  output \g234183/u3_syn_4  ;
  output \g234248/u3_syn_4  ;
  output \g234265/u3_syn_4  ;
  output \g234273/u3_syn_4  ;
  output \g234281/u3_syn_4  ;
  output \g234289/u3_syn_4  ;
  output \g234297/u3_syn_4  ;
  output \g234306/u3_syn_4  ;
  output \g234314/u3_syn_4  ;
  output \g234322/u3_syn_4  ;
  output \g234331/u3_syn_4  ;
  output \g234339/u3_syn_4  ;
  output \g234347/u3_syn_4  ;
  output \g234355/u3_syn_4  ;
  output \g234363/u3_syn_4  ;
  output \g234371/u3_syn_4  ;
  output \g234379/u3_syn_4  ;
  output \g234387/u3_syn_4  ;
  output \g234395/u3_syn_4  ;
  output \g234403/u3_syn_4  ;
  output \g234411/u3_syn_4  ;
  output \g234419/u3_syn_4  ;
  output \g234427/u3_syn_4  ;
  output \g234435/u3_syn_4  ;
  output \g234443/u3_syn_4  ;
  output \g234451/u3_syn_4  ;
  output \g234459/u3_syn_4  ;
  output \g234467/u3_syn_4  ;
  output \g234475/u3_syn_4  ;
  output \g234483/u3_syn_4  ;
  output \g234491/u3_syn_4  ;
  output \g234499/u3_syn_4  ;
  output \g234507/u3_syn_4  ;
  output \g234515/u3_syn_4  ;
  output \g234523/u3_syn_4  ;
  output \g234531/u3_syn_4  ;
  output \g234539/u3_syn_4  ;
  output \g234547/u3_syn_4  ;
  output \g234555/u3_syn_4  ;
  output \g234563/u3_syn_4  ;
  output \g234571/u3_syn_4  ;
  output \g234579/u3_syn_4  ;
  output \g234587/u3_syn_4  ;
  output \g234595/u3_syn_4  ;
  output \g234604/u3_syn_4  ;
  output \g234612/u3_syn_4  ;
  output \g234620/u3_syn_4  ;
  output \g234628/u3_syn_4  ;
  output \g234636/u3_syn_4  ;
  output \g234644/u3_syn_4  ;
  output \g234652/u3_syn_4  ;
  output \g234660/u3_syn_4  ;
  output \g234668/u3_syn_4  ;
  output \g234676/u3_syn_4  ;
  output \g234684/u3_syn_4  ;
  output \g234692/u3_syn_4  ;
  output \g234700/u3_syn_4  ;
  output \g234708/u3_syn_4  ;
  output \g234716/u3_syn_4  ;
  output \g234725/u3_syn_4  ;
  output \g234733/u3_syn_4  ;
  output \g234741/u3_syn_4  ;
  output \g234749/u3_syn_4  ;
  output \g234757/u3_syn_4  ;
  output \g234765/u3_syn_4  ;
  output \g234773/u3_syn_4  ;
  output \g234781/u3_syn_4  ;
  output \g234789/u3_syn_4  ;
  output \g234798/u3_syn_4  ;
  output \g234806/u3_syn_4  ;
  output \g234814/u3_syn_4  ;
  output \g234822/u3_syn_4  ;
  output \g234830/u3_syn_4  ;
  output \g234838/u3_syn_4  ;
  output \g235911/u3_syn_4  ;
  output \g235912/u3_syn_4  ;
  output \g235920/u3_syn_4  ;
  output \g235928/u3_syn_4  ;
  output \g235936/u3_syn_4  ;
  output \g235944/u3_syn_4  ;
  output \g235952/u3_syn_4  ;
  output \g235960/u3_syn_4  ;
  output \g235968/u3_syn_4  ;
  output \g235976/u3_syn_4  ;
  output \g235984/u3_syn_4  ;
  output \g235992/u3_syn_4  ;
  output \g236000/u3_syn_4  ;
  output \g236008/u3_syn_4  ;
  output \g236016/u3_syn_4  ;
  output \g236021/u3_syn_4  ;
  output \g236025/u3_syn_4  ;
  output \g236033/u3_syn_4  ;
  output \g236041/u3_syn_4  ;
  output \g236049/u3_syn_4  ;
  output \g236057/u3_syn_4  ;
  output \g236065/u3_syn_4  ;
  output \g236073/u3_syn_4  ;
  output \g236081/u3_syn_4  ;
  output \g236089/u3_syn_4  ;
  output \g236097/u3_syn_4  ;
  output \g236105/u3_syn_4  ;
  output \g236113/u3_syn_4  ;
  output \g236121/u3_syn_4  ;
  output \g236129/u3_syn_4  ;
  output \g236137/u3_syn_4  ;
  output \g236145/u3_syn_4  ;
  output \g236153/u3_syn_4  ;
  output \g236161/u3_syn_4  ;
  output \g236169/u3_syn_4  ;
  output \g236177/u3_syn_4  ;
  output \g236185/u3_syn_4  ;
  output \g236193/u3_syn_4  ;
  output \g236196/u3_syn_4  ;
  output \g236198/u3_syn_4  ;
  output \g236203/u3_syn_4  ;
  output \g236211/u3_syn_4  ;
  output \g236219/u3_syn_4  ;
  output \g236220/u3_syn_4  ;
  output \g236229/u3_syn_4  ;
  output \g236232/u3_syn_4  ;
  output \g236238/u3_syn_4  ;
  output \g236246/u3_syn_4  ;
  output \g236255/u3_syn_4  ;
  output \g236263/u3_syn_4  ;
  output \g236271/u3_syn_4  ;
  output \g236275/u3_syn_4  ;
  output \g236280/u3_syn_4  ;
  output \g236288/u3_syn_4  ;
  output \g236296/u3_syn_4  ;
  output \g236304/u3_syn_4  ;
  output \g236305/u3_syn_4  ;
  output \g236306/u3_syn_4  ;
  output \g236315/u3_syn_4  ;
  output \g236323/u3_syn_4  ;
  output \g236331/u3_syn_4  ;
  output \g236334/u3_syn_4  ;
  output \g236340/u3_syn_4  ;
  output \g236348/u3_syn_4  ;
  output \g236357/u3_syn_4  ;
  output \g236359/u3_syn_4  ;
  output \g236367/u3_syn_4  ;
  output \g236374/u3_syn_4  ;
  output \g236376/u3_syn_4  ;
  output \g236377/u3_syn_4  ;
  output \g236385/u3_syn_4  ;
  output \g236393/u3_syn_4  ;
  output \g236402/u3_syn_4  ;
  output \g236410/u3_syn_4  ;
  output \g236419/u3_syn_4  ;
  output \g236427/u3_syn_4  ;
  output \g236433/u3_syn_4  ;
  output \g236436/u3_syn_4  ;
  output \g236444/u3_syn_4  ;
  output \g236452/u3_syn_4  ;
  output \g236460/u3_syn_4  ;
  output \g236468/u3_syn_4  ;
  output \g236476/u3_syn_4  ;
  output \g236484/u3_syn_4  ;
  output \g236492/u3_syn_4  ;
  output \g236500/u3_syn_4  ;
  output \g236508/u3_syn_4  ;
  output \g236516/u3_syn_4  ;
  output \g236518/u3_syn_4  ;
  output \g236525/u3_syn_4  ;
  output \g236533/u3_syn_4  ;
  output \g236542/u3_syn_4  ;
  output \g236550/u3_syn_4  ;
  output \g236559/u3_syn_4  ;
  output \g236567/u3_syn_4  ;
  output \g236575/u3_syn_4  ;
  output \g236583/u3_syn_4  ;
  output \g236591/u3_syn_4  ;
  output \g236599/u3_syn_4  ;
  output \g236607/u3_syn_4  ;
  output \g236608/u3_syn_4  ;
  output \g236616/u3_syn_4  ;
  output \g236624/u3_syn_4  ;
  output \g236632/u3_syn_4  ;
  output \g236640/u3_syn_4  ;
  output \g236647/u3_syn_4  ;
  output \g236649/u3_syn_4  ;
  output \g236659/u3_syn_4  ;
  output \g236671/u3_syn_4  ;
  output \g236677/u3_syn_4  ;
  output \g236688/u3_syn_4  ;
  output \g236696/u3_syn_4  ;
  output \g236705/u3_syn_4  ;
  output \g236712/u3_syn_4  ;
  output \g236718/u3_syn_4  ;
  output \g236729/u3_syn_4  ;
  output \g236732/u3_syn_4  ;
  output \g236745/u3_syn_4  ;
  output \g236753/u3_syn_4  ;
  output \g236761/u3_syn_4  ;
  output \g236769/u3_syn_4  ;
  output \g236777/u3_syn_4  ;
  output \g236779/u3_syn_4  ;
  output \g236788/u3_syn_4  ;
  output \g236800/u3_syn_4  ;
  output \g236802/u3_syn_4  ;
  output \g236805/u3_syn_4  ;
  output \g236813/u3_syn_4  ;
  output \g236825/u3_syn_4  ;
  output \g236829/u3_syn_4  ;
  output \g236837/u3_syn_4  ;
  output \g236849/u3_syn_4  ;
  output \g236854/u3_syn_4  ;
  output \g236860/u3_syn_4  ;
  output \g236872/u3_syn_4  ;
  output \g236878/u3_syn_4  ;
  output \g236884/u3_syn_4  ;
  output \g236896/u3_syn_4  ;
  output \g236903/u3_syn_4  ;
  output \g236908/u3_syn_4  ;
  output \g236920/u3_syn_4  ;
  output \g236930/u3_syn_4  ;
  output \g236939/u3_syn_4  ;
  output \g236947/u3_syn_4  ;
  output \g236949/u3_syn_4  ;
  output \g236956/u3_syn_4  ;
  output \g236962/u3_syn_4  ;
  output \g236965/u3_syn_4  ;
  output \g236980/u3_syn_4  ;
  output \g236988/u3_syn_4  ;
  output \g236989/u3_syn_4  ;
  output \g237004/u3_syn_4  ;
  output \g237005/u3_syn_4  ;
  output \g237020/u3_syn_4  ;
  output \g237021/u3_syn_4  ;
  output \g237033/u3_syn_4  ;
  output \g237044/u3_syn_4  ;
  output \g237045/u3_syn_4  ;
  output \g237056/u3_syn_4  ;
  output \g237068/u3_syn_4  ;
  output \g237076/u3_syn_4  ;
  output \g237084/u3_syn_4  ;
  output \g237092/u3_syn_4  ;
  output \g237095/u3_syn_4  ;
  output \g237107/u3_syn_4  ;
  output \g237110/u3_syn_4  ;
  output \g237119/u3_syn_4  ;
  output \g237131/u3_syn_4  ;
  output \g237135/u3_syn_4  ;
  output \g237148/u3_syn_4  ;
  output \g237152/u3_syn_4  ;
  output \g237165/u3_syn_4  ;
  output \g237168/u3_syn_4  ;
  output \g237180/u3_syn_4  ;
  output \g237185/u3_syn_4  ;
  output \g237192/u3_syn_4  ;
  output \g237204/u3_syn_4  ;
  output \g237209/u3_syn_4  ;
  output \g237215/u3_syn_4  ;
  output \g237229/u3_syn_4  ;
  output \g237231/u3_syn_4  ;
  output \g237245/u3_syn_4  ;
  output \g237251/u3_syn_4  ;
  output \g237260/u3_syn_4  ;
  output \g237262/u3_syn_4  ;
  output \g237277/u3_syn_4  ;
  output \g237281/u3_syn_4  ;
  output \g237293/u3_syn_4  ;
  output \g237294/u3_syn_4  ;
  output \g237310/u3_syn_4  ;
  output \g237311/u3_syn_4  ;
  output \g237323/u3_syn_4  ;
  output \g237334/u3_syn_4  ;
  output \g237342/u3_syn_4  ;
  output \g237350/u3_syn_4  ;
  output \g237353/u3_syn_4  ;
  output \g237359/u3_syn_4  ;
  output \g237367/u3_syn_4  ;
  output \g237368/u3_syn_4  ;
  output \g237378/u3_syn_4  ;
  output \g237391/u3_syn_4  ;
  output \g237392/u3_syn_4  ;
  output \g237403/u3_syn_4  ;
  output \g237415/u3_syn_4  ;
  output \g237417/u3_syn_4  ;
  output \g237431/u3_syn_4  ;
  output \g237439/u3_syn_4  ;
  output \g237440/u3_syn_4  ;
  output \g237454/u3_syn_4  ;
  output \g237457/u3_syn_4  ;
  output \g237472/u3_syn_4  ;
  output \g237480/u3_syn_4  ;
  output \g237488/u3_syn_4  ;
  output \g237496/u3_syn_4  ;
  output \g237499/u3_syn_4  ;
  output \g237512/u3_syn_4  ;
  output \g237515/u3_syn_4  ;
  output \g237525/u3_syn_4  ;
  output \g237529/u3_syn_4  ;
  output \g237535/u3_syn_4  ;
  output \g237541/u3_syn_4  ;
  output \g237553/u3_syn_4  ;
  output \g237561/u3_syn_4  ;
  output \g237569/u3_syn_4  ;
  output \g237575/u3_syn_4  ;
  output \g237578/u3_syn_4  ;
  output \g237581/u3_syn_4  ;
  output \g237591/u3_syn_4  ;
  output \g237602/u3_syn_4  ;
  output \g237610/u3_syn_4  ;
  output \g237617/u3_syn_4  ;
  output \g237623/u3_syn_4  ;
  output \g237633/u3_syn_4  ;
  output \g237635/u3_syn_4  ;
  output \g237648/u3_syn_4  ;
  output \g237658/u3_syn_4  ;
  output \g237659/u3_syn_4  ;
  output \g237660/u3_syn_4  ;
  output \g237668/u3_syn_4  ;
  output \g237675/u3_syn_4  ;
  output \g237684/u3_syn_4  ;
  output \g237692/u3_syn_4  ;
  output \g237693/u3_syn_4  ;
  output \g237705/u3_syn_4  ;
  output \g237716/u3_syn_4  ;
  output \g237717/u3_syn_4  ;
  output \g237729/u3_syn_4  ;
  output \g237740/u3_syn_4  ;
  output \g237741/u3_syn_4  ;
  output \g237756/u3_syn_4  ;
  output \g237764/u3_syn_4  ;
  output \g237768/u3_syn_4  ;
  output \g237780/u3_syn_4  ;
  output \g237782/u3_syn_4  ;
  output \g237792/u3_syn_4  ;
  output \g237804/u3_syn_4  ;
  output \g237812/u3_syn_4  ;
  output \g237820/u3_syn_4  ;
  output \g237828/u3_syn_4  ;
  output \g237836/u3_syn_4  ;
  output \g237844/u3_syn_4  ;
  output \g237852/u3_syn_4  ;
  output \g237860/u3_syn_4  ;
  output \g237868/u3_syn_4  ;
  output \g237876/u3_syn_4  ;
  output \g237884/u3_syn_4  ;
  output \g237888/u3_syn_4  ;
  output \g237895/u3_syn_4  ;
  output \g237907/u3_syn_4  ;
  output \g237916/u3_syn_4  ;
  output \g237924/u3_syn_4  ;
  output \g237931/u3_syn_4  ;
  output \g237940/u3_syn_4  ;
  output \g237949/u3_syn_4  ;
  output \g237950/u3_syn_4  ;
  output \g237955/u3_syn_4  ;
  output \g237961/u3_syn_4  ;
  output \g237965/u3_syn_4  ;
  output \g237975/u3_syn_4  ;
  output \g237983/u3_syn_4  ;
  output \g237989/u3_syn_4  ;
  output \g237999/u3_syn_4  ;
  output \g238007/u3_syn_4  ;
  output \g238015/u3_syn_4  ;
  output \g238017/u3_syn_4  ;
  output \g238033/u3_syn_4  ;
  output \g238035/u3_syn_4  ;
  output \g238049/u3_syn_4  ;
  output \g238057/u3_syn_4  ;
  output \g238065/u3_syn_4  ;
  output \g238072/u3_syn_4  ;
  output \g238081/u3_syn_4  ;
  output \g238082/u3_syn_4  ;
  output \g238097/u3_syn_4  ;
  output \g238105/u3_syn_4  ;
  output \g238113/u3_syn_4  ;
  output \g238114/u3_syn_4  ;
  output \g238129/u3_syn_4  ;
  output \g238137/u3_syn_4  ;
  output \g238145/u3_syn_4  ;
  output \g238153/u3_syn_4  ;
  output \g238161/u3_syn_4  ;
  output \g238163/u3_syn_4  ;
  output \g238177/u3_syn_4  ;
  output \g238179/u3_syn_4  ;
  output \g238194/u3_syn_4  ;
  output \g238197/u3_syn_4  ;
  output \g238209/u3_syn_4  ;
  output \g238213/u3_syn_4  ;
  output \g238225/u3_syn_4  ;
  output \g238229/u3_syn_4  ;
  output \g238237/u3_syn_4  ;
  output \g238250/u3_syn_4  ;
  output \g238257/u3_syn_4  ;
  output \g238263/u3_syn_4  ;
  output \g238269/u3_syn_4  ;
  output \g238282/u3_syn_4  ;
  output \g238285/u3_syn_4  ;
  output \g238298/u3_syn_4  ;
  output \g238301/u3_syn_4  ;
  output \g238314/u3_syn_4  ;
  output \g238316/u3_syn_4  ;
  output \g238329/u3_syn_4  ;
  output \g238338/u3_syn_4  ;
  output \g238346/u3_syn_4  ;
  output \g238351/u3_syn_4  ;
  output \g238356/u3_syn_4  ;
  output \g238368/u3_syn_4  ;
  output \g238378/u3_syn_4  ;
  output \g238386/u3_syn_4  ;
  output \g238394/u3_syn_4  ;
  output \g238402/u3_syn_4  ;
  output \g238409/u3_syn_4  ;
  output \g238412/u3_syn_4  ;
  output \g238427/u3_syn_4  ;
  output \g238429/u3_syn_4  ;
  output \g238443/u3_syn_4  ;
  output \g238448/u3_syn_4  ;
  output \g238457/u3_syn_4  ;
  output \g238460/u3_syn_4  ;
  output \g238472/u3_syn_4  ;
  output \g238484/u3_syn_4  ;
  output \g238492/u3_syn_4  ;
  output \g238500/u3_syn_4  ;
  output \g238505/u3_syn_4  ;
  output \g238516/u3_syn_4  ;
  output \g238524/u3_syn_4  ;
  output \g238532/u3_syn_4  ;
  output \g238534/u3_syn_4  ;
  output \g238544/u3_syn_4  ;
  output \g238549/u3_syn_4  ;
  output \g238550/u3_syn_4  ;
  output \g238565/u3_syn_4  ;
  output \g238566/u3_syn_4  ;
  output \g238582/u3_syn_4  ;
  output \g238583/u3_syn_4  ;
  output \g238594/u3_syn_4  ;
  output \g238606/u3_syn_4  ;
  output \g238614/u3_syn_4  ;
  output \g238615/u3_syn_4  ;
  output \g238619/u3_syn_4  ;
  output \g238631/u3_syn_4  ;
  output \g238639/u3_syn_4  ;
  output \g238647/u3_syn_4  ;
  output \g238649/u3_syn_4  ;
  output \g238659/u3_syn_4  ;
  output \g238670/u3_syn_4  ;
  output \g238671/u3_syn_4  ;
  output \g238680/u3_syn_4  ;
  output \g238688/u3_syn_4  ;
  output \g238691/u3_syn_4  ;
  output \g238696/u3_syn_4  ;
  output \g238705/u3_syn_4  ;
  output \g238708/u3_syn_4  ;
  output \g238721/u3_syn_4  ;
  output \g238724/u3_syn_4  ;
  output \g238736/u3_syn_4  ;
  output \g238745/u3_syn_4  ;
  output \g238753/u3_syn_4  ;
  output \g238757/u3_syn_4  ;
  output \g238764/u3_syn_4  ;
  output \g238776/u3_syn_4  ;
  output \g238781/u3_syn_4  ;
  output \g238787/u3_syn_4  ;
  output \g238799/u3_syn_4  ;
  output \g238807/u3_syn_4  ;
  output \g238811/u3_syn_4  ;
  output \g238824/u3_syn_4  ;
  output \g238830/u3_syn_4  ;
  output \g238841/u3_syn_4  ;
  output \g238843/u3_syn_4  ;
  output \g238855/u3_syn_4  ;
  output \g238859/u3_syn_4  ;
  output \g238863/u3_syn_4  ;
  output \g238868/u3_syn_4  ;
  output \g238880/u3_syn_4  ;
  output \g238888/u3_syn_4  ;
  output \g238892/u3_syn_4  ;
  output \g238903/u3_syn_4  ;
  output \g238911/u3_syn_4  ;
  output \g238915/u3_syn_4  ;
  output \g238927/u3_syn_4  ;
  output \g238937/u3_syn_4  ;
  output \g238945/u3_syn_4  ;
  output \g238953/u3_syn_4  ;
  output \g238961/u3_syn_4  ;
  output \g238970/u3_syn_4  ;
  output \g238971/u3_syn_4  ;
  output \g238983/u3_syn_4  ;
  output \g238994/u3_syn_4  ;
  output \g239002/u3_syn_4  ;
  output \g239009/u3_syn_4  ;
  output \g239015/u3_syn_4  ;
  output \g239025/u3_syn_4  ;
  output \g239030/u3_syn_4  ;
  output \g239041/u3_syn_4  ;
  output \g239048/u3_syn_4  ;
  output \g239053/u3_syn_4  ;
  output \g239065/u3_syn_4  ;
  output \g239073/u3_syn_4  ;
  output \g239081/u3_syn_4  ;
  output \g239082/u3_syn_4  ;
  output \g239093/u3_syn_4  ;
  output \g239105/u3_syn_4  ;
  output \g239108/u3_syn_4  ;
  output \g239117/u3_syn_4  ;
  output \g239129/u3_syn_4  ;
  output \g239137/u3_syn_4  ;
  output \g239139/u3_syn_4  ;
  output \g239148/u3_syn_4  ;
  output \g239160/u3_syn_4  ;
  output \g239162/u3_syn_4  ;
  output \g239172/u3_syn_4  ;
  output \g239184/u3_syn_4  ;
  output \g239187/u3_syn_4  ;
  output \g239189/u3_syn_4  ;
  output \g239201/u3_syn_4  ;
  output \g239208/u3_syn_4  ;
  output \g239217/u3_syn_4  ;
  output \g239219/u3_syn_4  ;
  output \g239226/u3_syn_4  ;
  output \g239234/u3_syn_4  ;
  output \g239242/u3_syn_4  ;
  output \g239246/u3_syn_4  ;
  output \g239257/u3_syn_4  ;
  output \g239258/u3_syn_4  ;
  output \g239263/u3_syn_4  ;
  output \g239275/u3_syn_4  ;
  output \g239277/u3_syn_4  ;
  output \g239291/u3_syn_4  ;
  output \g239296/u3_syn_4  ;
  output \g239308/u3_syn_4  ;
  output \g239311/u3_syn_4  ;
  output \g239322/u3_syn_4  ;
  output \g239329/u3_syn_4  ;
  output \g239338/u3_syn_4  ;
  output \g239339/u3_syn_4  ;
  output \g239346/u3_syn_4  ;
  output \g239351/u3_syn_4  ;
  output \g239363/u3_syn_4  ;
  output \g239370/u3_syn_4  ;
  output \g239375/u3_syn_4  ;
  output \g239387/u3_syn_4  ;
  output \g239395/u3_syn_4  ;
  output \g239418/u3_syn_4  ;
  output \g239439/u3_syn_4  ;
  output \g239442/u3_syn_4  ;
  output \g239454/u3_syn_4  ;
  output \g239464/u3_syn_4  ;
  output \g239470/u3_syn_4  ;
  output \g239481/u3_syn_4  ;
  output \g239487/u3_syn_4  ;
  output \g239497/u3_syn_4  ;
  output \g239520/u3_syn_4  ;
  output \g239532/u3_syn_4  ;
  output \g239543/u3_syn_4  ;
  output \g239551/u3_syn_4  ;
  output \g239552/u3_syn_4  ;
  output \g239567/u3_syn_4  ;
  output \g239575/u3_syn_4  ;
  output \g239579/u3_syn_4  ;
  output \g239592/u3_syn_4  ;
  output \g239594/u3_syn_4  ;
  output \g239608/u3_syn_4  ;
  output \g239626/u3_syn_4  ;
  output \g239634/u3_syn_4  ;
  output \g239646/u3_syn_4  ;
  output \g239649/u3_syn_4  ;
  output \g239657/u3_syn_4  ;
  output \g239670/u3_syn_4  ;
  output \g239673/u3_syn_4  ;
  output \g239686/u3_syn_4  ;
  output \g239694/u3_syn_4  ;
  output \g239695/u3_syn_4  ;
  output \g239701/u3_syn_4  ;
  output \g239705/u3_syn_4  ;
  output \g239709/u3_syn_4  ;
  output \g239715/u3_syn_4  ;
  output \g239717/u3_syn_4  ;
  output \g239726/u3_syn_4  ;
  output \g239734/u3_syn_4  ;
  output \g239735/u3_syn_4  ;
  output \g239743/u3_syn_4  ;
  output \g239760/u3_syn_4  ;
  output \g239768/u3_syn_4  ;
  output \g239776/u3_syn_4  ;
  output \g239784/u3_syn_4  ;
  output \g239793/u3_syn_4  ;
  output \g239801/u3_syn_4  ;
  output \g239817/u3_syn_4  ;
  output \g239818/u3_syn_4  ;
  output \g239848/u3_syn_4  ;
  output \g239856/u3_syn_4  ;
  output \g239872/u3_syn_4  ;
  output \g239880/u3_syn_4  ;
  output \g239888/u3_syn_4  ;
  output \g239896/u3_syn_4  ;
  output \g239904/u3_syn_4  ;
  output \g239912/u3_syn_4  ;
  output \g239920/u3_syn_4  ;
  output \g239928/u3_syn_4  ;
  output \g239936/u3_syn_4  ;
  output \g239951/u3_syn_4  ;
  output \g239963/u3_syn_4  ;
  output \g239979/u3_syn_4  ;
  output \g239986/u3_syn_4  ;
  output \g239999/u3_syn_4  ;
  output \g240000/u3_syn_4  ;
  output \g240008/u3_syn_4  ;
  output \g240012/u3_syn_4  ;
  output \g240018/u3_syn_4  ;
  output \g240026/u3_syn_4  ;
  output \g240034/u3_syn_4  ;
  output \g240042/u3_syn_4  ;
  output \g240050/u3_syn_4  ;
  output \g240074/u3_syn_4  ;
  output \g240091/u3_syn_4  ;
  output \g240122/u3_syn_4  ;
  output \g240147/u3_syn_4  ;
  output \g240209/u3_syn_4  ;
  output \g240219/u3_syn_4  ;
  output \g240259/u3_syn_4  ;
  output \g240334/u3_syn_4  ;
  output \g240406/u3_syn_4  ;
  output \g240416/u3_syn_4  ;
  output \g240424/u3_syn_4  ;
  output \g240432/u3_syn_4  ;
  output \g240440/u3_syn_4  ;
  output \g240448/u3_syn_4  ;
  output \g240456/u3_syn_4  ;
  output \g240464/u3_syn_4  ;
  output \g240472/u3_syn_4  ;
  output \g240480/u3_syn_4  ;
  output \g240488/u3_syn_4  ;
  output \g240496/u3_syn_4  ;
  output \g240504/u3_syn_4  ;
  output \g240512/u3_syn_4  ;
  output \g240520/u3_syn_4  ;
  output \g240530/u3_syn_4  ;
  output \g240538/u3_syn_4  ;
  output \g240547/u3_syn_4  ;
  output \g240555/u3_syn_4  ;
  output \g240563/u3_syn_4  ;
  output \g240571/u3_syn_4  ;
  output \g240579/u3_syn_4  ;
  output \g240587/u3_syn_4  ;
  output \g240595/u3_syn_4  ;
  output \g240603/u3_syn_4  ;
  output \g240611/u3_syn_4  ;
  output \g240619/u3_syn_4  ;
  output \g240627/u3_syn_4  ;
  output \g240635/u3_syn_4  ;
  output \g240643/u3_syn_4  ;
  output \g240651/u3_syn_4  ;
  output \g240659/u3_syn_4  ;
  output \g240667/u3_syn_4  ;
  output \g240675/u3_syn_4  ;
  output \g240683/u3_syn_4  ;
  output \g240691/u3_syn_4  ;
  output \g240699/u3_syn_4  ;
  output \g240707/u3_syn_4  ;
  output \g240715/u3_syn_4  ;
  output \g240723/u3_syn_4  ;
  output \g240731/u3_syn_4  ;
  output \g240739/u3_syn_4  ;
  output \g240747/u3_syn_4  ;
  output \g240755/u3_syn_4  ;
  output \g240763/u3_syn_4  ;
  output \g240771/u3_syn_4  ;
  output \g240779/u3_syn_4  ;
  output \g240787/u3_syn_4  ;
  output \g240795/u3_syn_4  ;
  output \g240803/u3_syn_4  ;
  output \g240811/u3_syn_4  ;
  output \g240819/u3_syn_4  ;
  output \g240827/u3_syn_4  ;
  output \g240835/u3_syn_4  ;
  output \g240843/u3_syn_4  ;
  output \g240851/u3_syn_4  ;
  output \g240859/u3_syn_4  ;
  output \g240867/u3_syn_4  ;
  output \g240875/u3_syn_4  ;
  output \g240883/u3_syn_4  ;
  output \g240891/u3_syn_4  ;
  output \g240899/u3_syn_4  ;
  output \g240907/u3_syn_4  ;
  output \g240915/u3_syn_4  ;
  output \g240923/u3_syn_4  ;
  output \g240931/u3_syn_4  ;
  output \g240939/u3_syn_4  ;
  output \g240947/u3_syn_4  ;
  output \g240955/u3_syn_4  ;
  output \g240963/u3_syn_4  ;
  output \g240971/u3_syn_4  ;
  output \g240979/u3_syn_4  ;
  output \g240987/u3_syn_4  ;
  output \g240995/u3_syn_4  ;
  output \g241003/u3_syn_4  ;
  output \g241011/u3_syn_4  ;
  output \g241019/u3_syn_4  ;
  output \g241027/u3_syn_4  ;
  output \g241036/u3_syn_4  ;
  output \g241044/u3_syn_4  ;
  output \g241052/u3_syn_4  ;
  output \g241060/u3_syn_4  ;
  output \g241068/u3_syn_4  ;
  output \g241076/u3_syn_4  ;
  output \g241084/u3_syn_4  ;
  output \g241092/u3_syn_4  ;
  output \g241100/u3_syn_4  ;
  output \g241108/u3_syn_4  ;
  output \g241116/u3_syn_4  ;
  output \g241124/u3_syn_4  ;
  output \g241132/u3_syn_4  ;
  output \g241140/u3_syn_4  ;
  output \g241148/u3_syn_4  ;
  output \g241156/u3_syn_4  ;
  output \g241164/u3_syn_4  ;
  output \g241172/u3_syn_4  ;
  output \g241180/u3_syn_4  ;
  output \g241188/u3_syn_4  ;
  output \g241196/u3_syn_4  ;
  output \g241205/u3_syn_4  ;
  output \g241213/u3_syn_4  ;
  output \g241221/u3_syn_4  ;
  output \g241229/u3_syn_4  ;
  output \g241237/u3_syn_4  ;
  output \g241245/u3_syn_4  ;
  output \g241253/u3_syn_4  ;
  output \g241261/u3_syn_4  ;
  output \g241269/u3_syn_4  ;
  output \g241277/u3_syn_4  ;
  output \g241285/u3_syn_4  ;
  output \g241293/u3_syn_4  ;
  output \g241301/u3_syn_4  ;
  output \g241309/u3_syn_4  ;
  output \g241317/u3_syn_4  ;
  output \g241325/u3_syn_4  ;
  output \g241333/u3_syn_4  ;
  output \g241341/u3_syn_4  ;
  output \g241349/u3_syn_4  ;
  output \g241358/u3_syn_4  ;
  output \g241366/u3_syn_4  ;
  output \g241374/u3_syn_4  ;
  output \g241382/u3_syn_4  ;
  output \g241390/u3_syn_4  ;
  output \g241398/u3_syn_4  ;
  output \g241406/u3_syn_4  ;
  output \g241415/u3_syn_4  ;
  output \g241424/u3_syn_4  ;
  output \g241433/u3_syn_4  ;
  output \g241441/u3_syn_4  ;
  output \g241449/u3_syn_4  ;
  output \g241459/u3_syn_4  ;
  output \g241470/u3_syn_4  ;
  output \g241480/u3_syn_4  ;
  output \g241489/u3_syn_4  ;
  output \g241497/u3_syn_4  ;
  output \g241505/u3_syn_4  ;
  output \g241513/u3_syn_4  ;
  output \g241545/_3_  ;
  output \g241580/_00_  ;
  output \g241737/_0_  ;
  output \g241752/_0_  ;
  output \g241755/_0_  ;
  output \g241767/_2__syn_2  ;
  output \g241781/_1__syn_2  ;
  output \g241782/_0_  ;
  output \g241803/_1__syn_2  ;
  output \g241805/_0_  ;
  output \g241812/_1__syn_2  ;
  output \g241814/_1__syn_2  ;
  output \g241816/_1__syn_2  ;
  output \g241819/_1__syn_2  ;
  output \g241822/_1__syn_2  ;
  output \g241823/_0_  ;
  output \g241833/_1__syn_2  ;
  output \g241843/_1__syn_2  ;
  output \g241844/_1__syn_2  ;
  output \g241848/_1__syn_2  ;
  output \g241855/_1__syn_2  ;
  output \g241868/_1__syn_2  ;
  output \g242013/_1__syn_2  ;
  output \g242015/_1__syn_2  ;
  output \g242017/_1__syn_2  ;
  output \g242021/_1__syn_2  ;
  output \g242039/_1__syn_2  ;
  output \g242081/_0_  ;
  output \g242086/_0_  ;
  output \g242101/_3_  ;
  output \g242116/_0_  ;
  output \g242135/_2_  ;
  output \g242147/_0_  ;
  output \g242158/_0_  ;
  output \g242196/_0_  ;
  output \g242202/_0_  ;
  output \g242203/_0_  ;
  output \g242204/_0_  ;
  output \g242212/_0_  ;
  output \g242226/_01_  ;
  output \g242281/_0_  ;
  output \g242407/_0_  ;
  output \g242410/_0_  ;
  output \g242426/_0_  ;
  output \g242438/_2_  ;
  output \g242466/_0_  ;
  output \g242530/_0_  ;
  output \g242532/_0_  ;
  output \g243397/_0_  ;
  output \g245925/_0_  ;
  output \g245932/_0_  ;
  output \g245933/_0_  ;
  output \g245986/_3_  ;
  output \g250157/_3_  ;
  output \g250202/_0_  ;
  output \g250246/_1_  ;
  output \g250248/_0_  ;
  output \g250250/_0_  ;
  output \g250305/_0_  ;
  output \g250323/_0_  ;
  output \g250373/_0_  ;
  output \g250377/_0_  ;
  output \g250412/_0_  ;
  output \g250413/_0_  ;
  output \g250418/_0_  ;
  output \g250419/_0_  ;
  output \g250421/_0_  ;
  output \g250433/_0_  ;
  output \g250448/_3_  ;
  output \g250567/_3_  ;
  output \g258965/_0_  ;
  output \g259006/_0_  ;
  output \g259471/_0_  ;
  output \g259473/_2_  ;
  output \g260557/_0_  ;
  output \g261035/_0_  ;
  output \g261095/_3_  ;
  output \g261207/_2__syn_2  ;
  output \g261754/_0_  ;
  output \g262017/_0_  ;
  output \g262045/_0_  ;
  output \g262046/_0_  ;
  output \g262100/_3_  ;
  output \g263539/_1_  ;
  output \g263574/_0_  ;
  output \g263858/_0_  ;
  output \g264104/_1_  ;
  output \g264107/_1_  ;
  output \g264117/_0_  ;
  output \g264282/_0_  ;
  output \g264511/_0_  ;
  output \g264541/_0_  ;
  output \g264562/_0_  ;
  output \g264618/_0_  ;
  output \g264660/_0_  ;
  output \g264681/_3_  ;
  output \g264727/_0_  ;
  output \g265013/_0_  ;
  output \g265084/_0_  ;
  output \g265378/_0_  ;
  output \g265413/_0_  ;
  output \g265446/_0_  ;
  output \g265486/_0_  ;
  output \g265524/_3_  ;
  output \g265528/_3_  ;
  output \g265548/_3_  ;
  output \g265579/_0_  ;
  output \g265768/_0_  ;
  output \g265801/_0_  ;
  output \g265819/_1_  ;
  output \g265853/_0_  ;
  output \g265933/_0_  ;
  output \g266022/_0_  ;
  output \g266183/_1_  ;
  output \g281909/_0_  ;
  output \g281965/_1_  ;
  output \g282284/_1_  ;
  output \g282639/_1_  ;
  output \g283047/_0_  ;
  output \g283157/_1_  ;
  output \g283184/_0_  ;
  output \g283334/_3_  ;
  output int_o_pad ;
  output \m_wb_adr_o[0]_pad  ;
  output \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2  ;
  output \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3  ;
  output \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3  ;
  output \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3  ;
  output \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3  ;
  output \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3  ;
  output \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3  ;
  output \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3  ;
  wire n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 ;
  assign n10512 = ~\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n10513 = ~\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n10514 = ~\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n10515 = n10513 & n10514 ;
  assign n10516 = ~\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n10517 = ~\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n10518 = n10516 & n10517 ;
  assign n10519 = n10515 & n10518 ;
  assign n10520 = ~\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n10521 = ~\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n10522 = n10520 & n10521 ;
  assign n10523 = ~\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n10524 = n10522 & n10523 ;
  assign n10525 = n10519 & n10524 ;
  assign n10526 = n10512 & n10525 ;
  assign n10527 = \rxethmac1_crcrx_Crc_reg[26]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[27]/NET0131  ;
  assign n10528 = ~\rxethmac1_crcrx_Crc_reg[28]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[2]/NET0131  ;
  assign n10529 = n10527 & n10528 ;
  assign n10530 = ~\rxethmac1_crcrx_Crc_reg[22]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[23]/NET0131  ;
  assign n10531 = \rxethmac1_crcrx_Crc_reg[24]/NET0131  & \rxethmac1_crcrx_Crc_reg[25]/NET0131  ;
  assign n10532 = n10530 & n10531 ;
  assign n10533 = n10529 & n10532 ;
  assign n10534 = \rxethmac1_crcrx_Crc_reg[6]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[7]/NET0131  ;
  assign n10535 = \rxethmac1_crcrx_Crc_reg[8]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[9]/NET0131  ;
  assign n10536 = n10534 & n10535 ;
  assign n10537 = \rxethmac1_crcrx_Crc_reg[30]/NET0131  & \rxethmac1_crcrx_Crc_reg[3]/NET0131  ;
  assign n10538 = \rxethmac1_crcrx_Crc_reg[4]/NET0131  & \rxethmac1_crcrx_Crc_reg[5]/NET0131  ;
  assign n10539 = n10537 & n10538 ;
  assign n10540 = n10536 & n10539 ;
  assign n10541 = n10533 & n10540 ;
  assign n10542 = \rxethmac1_crcrx_Crc_reg[11]/NET0131  & \rxethmac1_crcrx_Crc_reg[12]/NET0131  ;
  assign n10543 = ~\rxethmac1_crcrx_Crc_reg[13]/NET0131  & \rxethmac1_crcrx_Crc_reg[14]/NET0131  ;
  assign n10544 = n10542 & n10543 ;
  assign n10545 = ~\rxethmac1_crcrx_Crc_reg[29]/NET0131  & \rxethmac1_crcrx_Crc_reg[31]/NET0131  ;
  assign n10546 = \rxethmac1_crcrx_Crc_reg[0]/NET0131  & \rxethmac1_crcrx_Crc_reg[10]/NET0131  ;
  assign n10547 = n10545 & n10546 ;
  assign n10548 = n10544 & n10547 ;
  assign n10549 = ~\rxethmac1_crcrx_Crc_reg[19]/NET0131  & \rxethmac1_crcrx_Crc_reg[1]/NET0131  ;
  assign n10550 = ~\rxethmac1_crcrx_Crc_reg[20]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[21]/NET0131  ;
  assign n10551 = n10549 & n10550 ;
  assign n10552 = \rxethmac1_crcrx_Crc_reg[15]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[16]/NET0131  ;
  assign n10553 = ~\rxethmac1_crcrx_Crc_reg[17]/NET0131  & \rxethmac1_crcrx_Crc_reg[18]/NET0131  ;
  assign n10554 = n10552 & n10553 ;
  assign n10555 = n10551 & n10554 ;
  assign n10556 = n10548 & n10555 ;
  assign n10557 = n10541 & n10556 ;
  assign n10558 = ~n10526 & ~n10557 ;
  assign n10559 = \rxethmac1_rxstatem1_StateData0_reg/NET0131  & ~n10558 ;
  assign n10560 = ~\macstatus1_LatchedCrcError_reg/NET0131  & ~\rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n10561 = ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  & ~n10560 ;
  assign n10562 = ~n10559 & n10561 ;
  assign n10563 = \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  & n10522 ;
  assign n10564 = n10519 & n10563 ;
  assign n10565 = ~\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n10566 = ~\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n10567 = n10565 & n10566 ;
  assign n10568 = ~\rxethmac1_crcrx_Crc_reg[27]/NET0131  & n10567 ;
  assign n10569 = n10564 & n10568 ;
  assign n10570 = ~\rxethmac1_rxstatem1_StateIdle_reg/NET0131  & ~wb_rst_i_pad ;
  assign n10571 = \rxethmac1_CrcHash_reg[1]/P0001  & n10570 ;
  assign n10572 = n10567 & n10570 ;
  assign n10573 = n10564 & n10572 ;
  assign n10574 = ~n10571 & ~n10573 ;
  assign n10575 = ~n10569 & ~n10574 ;
  assign n10576 = ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  ;
  assign n10577 = ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  & n10576 ;
  assign n10578 = \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  & ~n10577 ;
  assign n10579 = ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  & ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  ;
  assign n10580 = n10576 & n10579 ;
  assign n10581 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & ~n10580 ;
  assign n10582 = ~n10578 & n10581 ;
  assign n10583 = ~\rxethmac1_crcrx_Crc_reg[27]/NET0131  & ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n10584 = ~n10582 & n10583 ;
  assign n10585 = ~\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n10586 = \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n10587 = \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n10588 = ~n10586 & ~n10587 ;
  assign n10589 = ~n10585 & n10588 ;
  assign n10590 = \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n10591 = ~\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n10592 = ~n10590 & ~n10591 ;
  assign n10593 = ~\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
  assign n10594 = ~\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n10595 = ~n10593 & ~n10594 ;
  assign n10596 = n10592 & n10595 ;
  assign n10597 = \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n10598 = \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n10599 = ~n10597 & ~n10598 ;
  assign n10600 = ~\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n10601 = ~\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n10602 = ~n10600 & ~n10601 ;
  assign n10603 = n10599 & n10602 ;
  assign n10604 = n10596 & n10603 ;
  assign n10605 = n10589 & n10604 ;
  assign n10606 = ~\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n10607 = ~\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n10608 = ~n10606 & ~n10607 ;
  assign n10609 = \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
  assign n10610 = ~\ethreg1_MODER_1_DataOut_reg[6]/NET0131  & ~n10609 ;
  assign n10611 = ~\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n10612 = \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n10613 = ~n10611 & ~n10612 ;
  assign n10614 = n10610 & n10613 ;
  assign n10615 = n10608 & n10614 ;
  assign n10616 = \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n10617 = \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n10618 = ~n10616 & ~n10617 ;
  assign n10619 = ~\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n10620 = \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n10621 = ~n10619 & ~n10620 ;
  assign n10622 = n10618 & n10621 ;
  assign n10623 = \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n10624 = ~\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n10625 = ~n10623 & ~n10624 ;
  assign n10626 = \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n10627 = \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n10628 = ~n10626 & ~n10627 ;
  assign n10629 = n10625 & n10628 ;
  assign n10630 = n10622 & n10629 ;
  assign n10631 = ~\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n10632 = ~\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n10633 = ~n10631 & ~n10632 ;
  assign n10634 = ~\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n10635 = \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n10636 = ~n10634 & ~n10635 ;
  assign n10637 = n10633 & n10636 ;
  assign n10638 = \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n10639 = ~\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n10640 = ~n10638 & ~n10639 ;
  assign n10641 = \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n10642 = ~\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n10643 = ~n10641 & ~n10642 ;
  assign n10644 = n10640 & n10643 ;
  assign n10645 = n10637 & n10644 ;
  assign n10646 = n10630 & n10645 ;
  assign n10647 = n10615 & n10646 ;
  assign n10648 = n10605 & n10647 ;
  assign n10649 = ~\rxethmac1_rxstatem1_StateData0_reg/NET0131  & ~\rxethmac1_rxstatem1_StateData1_reg/NET0131  ;
  assign n10650 = \ethreg1_MODER_0_DataOut_reg[7]/NET0131  & mtxen_pad_o_pad ;
  assign n10651 = \RxEnSync_reg/NET0131  & mrxdv_pad_i_pad ;
  assign n10652 = ~\ethreg1_MODER_0_DataOut_reg[7]/NET0131  & n10651 ;
  assign n10653 = ~n10650 & ~n10652 ;
  assign n10654 = ~n10649 & ~n10653 ;
  assign n10655 = \ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mtxd_pad_o[2]_pad  ;
  assign n10656 = ~\ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mrxd_pad_i[2]_pad  ;
  assign n10657 = ~n10655 & ~n10656 ;
  assign n10658 = \rxethmac1_crcrx_Crc_reg[29]/NET0131  & ~n10657 ;
  assign n10659 = ~\rxethmac1_crcrx_Crc_reg[29]/NET0131  & n10657 ;
  assign n10660 = ~n10658 & ~n10659 ;
  assign n10661 = n10654 & n10660 ;
  assign n10662 = ~n10648 & n10661 ;
  assign n10663 = ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  & ~n10582 ;
  assign n10664 = ~\rxethmac1_crcrx_Crc_reg[23]/NET0131  & n10663 ;
  assign n10665 = ~n10662 & n10664 ;
  assign n10666 = \rxethmac1_crcrx_Crc_reg[23]/NET0131  & n10663 ;
  assign n10667 = n10662 & n10666 ;
  assign n10668 = ~n10665 & ~n10667 ;
  assign n10669 = \ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mtxd_pad_o[1]_pad  ;
  assign n10670 = ~\ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mrxd_pad_i[1]_pad  ;
  assign n10671 = ~n10669 & ~n10670 ;
  assign n10672 = \rxethmac1_crcrx_Crc_reg[30]/NET0131  & ~n10671 ;
  assign n10673 = ~\rxethmac1_crcrx_Crc_reg[30]/NET0131  & n10671 ;
  assign n10674 = ~n10672 & ~n10673 ;
  assign n10675 = n10654 & n10674 ;
  assign n10676 = ~n10648 & n10675 ;
  assign n10677 = ~\rxethmac1_crcrx_Crc_reg[24]/NET0131  & n10663 ;
  assign n10678 = ~n10676 & n10677 ;
  assign n10679 = \rxethmac1_crcrx_Crc_reg[24]/NET0131  & n10663 ;
  assign n10680 = n10676 & n10679 ;
  assign n10681 = ~n10678 & ~n10680 ;
  assign n10682 = ~\rxethmac1_crcrx_Crc_reg[26]/NET0131  & n10567 ;
  assign n10683 = n10564 & n10682 ;
  assign n10684 = \rxethmac1_CrcHash_reg[0]/P0001  & n10570 ;
  assign n10685 = ~n10573 & ~n10684 ;
  assign n10686 = ~n10683 & ~n10685 ;
  assign n10687 = ~\ethreg1_MODER_1_DataOut_reg[7]/NET0131  & ~\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131  ;
  assign n10688 = ~\wishbone_TxStatus_reg[12]/NET0131  & n10687 ;
  assign n10689 = ~\ethreg1_MODER_1_DataOut_reg[5]/NET0131  & ~\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131  ;
  assign n10690 = ~\wishbone_TxStatus_reg[11]/NET0131  & n10689 ;
  assign n10691 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & \wishbone_TxEndFrm_reg/NET0131  ;
  assign n10692 = \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131  ;
  assign n10693 = ~n10691 & ~n10692 ;
  assign n10694 = \Collision_Tx2_reg/NET0131  & ~\ethreg1_MODER_1_DataOut_reg[2]/NET0131  ;
  assign n10695 = \txethmac1_txstatem1_StateData_reg[1]/NET0131  & ~n10694 ;
  assign n10696 = ~n10693 & n10695 ;
  assign n10697 = n10690 & n10696 ;
  assign n10698 = n10688 & n10697 ;
  assign n10699 = ~\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  & ~\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  ;
  assign n10700 = ~\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & ~\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  ;
  assign n10701 = n10699 & n10700 ;
  assign n10702 = ~\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & n10701 ;
  assign n10703 = \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & ~n10701 ;
  assign n10704 = ~n10702 & ~n10703 ;
  assign n10705 = ~\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  & ~\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  ;
  assign n10706 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & ~\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  ;
  assign n10707 = n10699 & n10706 ;
  assign n10708 = n10705 & n10707 ;
  assign n10709 = ~\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  & n10708 ;
  assign n10710 = n10704 & n10709 ;
  assign n10711 = ~\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & ~\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  ;
  assign n10712 = n10701 & n10711 ;
  assign n10713 = \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & ~n10712 ;
  assign n10714 = ~\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & n10711 ;
  assign n10715 = n10701 & n10714 ;
  assign n10716 = ~\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  & ~n10715 ;
  assign n10717 = ~n10713 & n10716 ;
  assign n10718 = n10710 & n10717 ;
  assign n10719 = ~\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & ~\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  ;
  assign n10720 = n10711 & n10719 ;
  assign n10721 = n10701 & n10720 ;
  assign n10722 = ~\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & ~\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  ;
  assign n10723 = ~n10721 & n10722 ;
  assign n10724 = \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & ~\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  ;
  assign n10725 = n10721 & n10724 ;
  assign n10726 = ~n10723 & ~n10725 ;
  assign n10727 = n10718 & ~n10726 ;
  assign n10728 = n10721 & n10722 ;
  assign n10729 = \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & ~n10728 ;
  assign n10730 = ~\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & n10722 ;
  assign n10731 = n10721 & n10730 ;
  assign n10732 = ~\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  & ~n10731 ;
  assign n10733 = ~n10729 & n10732 ;
  assign n10734 = n10727 & n10733 ;
  assign n10735 = ~\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & ~\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  ;
  assign n10736 = n10722 & n10735 ;
  assign n10737 = n10721 & n10736 ;
  assign n10738 = \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  & ~n10737 ;
  assign n10739 = ~\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  & n10737 ;
  assign n10740 = ~n10738 & ~n10739 ;
  assign n10741 = ~\txethmac1_txcounters1_NibCnt_reg[15]/NET0131  & ~n10740 ;
  assign n10742 = ~n10734 & n10741 ;
  assign n10743 = ~\txethmac1_txcounters1_NibCnt_reg[15]/NET0131  & n10740 ;
  assign n10744 = n10734 & n10743 ;
  assign n10745 = ~n10742 & ~n10744 ;
  assign n10746 = \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  & ~n10702 ;
  assign n10747 = ~\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & n10705 ;
  assign n10748 = n10707 & n10747 ;
  assign n10749 = ~n10712 & n10748 ;
  assign n10750 = ~n10746 & n10749 ;
  assign n10751 = ~\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & n10750 ;
  assign n10752 = \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  & ~n10715 ;
  assign n10753 = ~\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & ~n10721 ;
  assign n10754 = ~n10752 & n10753 ;
  assign n10755 = n10751 & n10754 ;
  assign n10756 = ~\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & n10721 ;
  assign n10757 = \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  & ~n10756 ;
  assign n10758 = ~\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & ~n10728 ;
  assign n10759 = ~n10757 & n10758 ;
  assign n10760 = n10755 & n10759 ;
  assign n10761 = \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  & ~n10731 ;
  assign n10762 = ~n10737 & ~n10761 ;
  assign n10763 = ~\txethmac1_txcounters1_NibCnt_reg[14]/NET0131  & ~n10762 ;
  assign n10764 = ~n10760 & n10763 ;
  assign n10765 = ~\txethmac1_txcounters1_NibCnt_reg[14]/NET0131  & n10762 ;
  assign n10766 = n10760 & n10765 ;
  assign n10767 = ~n10764 & ~n10766 ;
  assign n10768 = n10745 & n10767 ;
  assign n10769 = ~n10729 & ~n10731 ;
  assign n10770 = \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & ~n10769 ;
  assign n10771 = n10727 & n10770 ;
  assign n10772 = \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & n10769 ;
  assign n10773 = ~n10727 & n10772 ;
  assign n10774 = ~n10771 & ~n10773 ;
  assign n10775 = n10768 & ~n10774 ;
  assign n10776 = ~\txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & ~n10769 ;
  assign n10777 = ~n10727 & n10776 ;
  assign n10778 = ~\txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & n10769 ;
  assign n10779 = n10727 & n10778 ;
  assign n10780 = ~n10777 & ~n10779 ;
  assign n10781 = ~n10728 & ~n10757 ;
  assign n10782 = \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  & ~n10781 ;
  assign n10783 = n10755 & n10782 ;
  assign n10784 = \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  & n10781 ;
  assign n10785 = ~n10755 & n10784 ;
  assign n10786 = ~n10783 & ~n10785 ;
  assign n10787 = n10780 & ~n10786 ;
  assign n10788 = n10768 & n10787 ;
  assign n10789 = ~n10734 & ~n10740 ;
  assign n10790 = n10733 & n10740 ;
  assign n10791 = n10727 & n10790 ;
  assign n10792 = \txethmac1_txcounters1_NibCnt_reg[15]/NET0131  & ~n10791 ;
  assign n10793 = ~n10789 & n10792 ;
  assign n10794 = ~n10760 & ~n10762 ;
  assign n10795 = n10759 & n10762 ;
  assign n10796 = n10755 & n10795 ;
  assign n10797 = \txethmac1_txcounters1_NibCnt_reg[14]/NET0131  & ~n10796 ;
  assign n10798 = ~n10794 & n10797 ;
  assign n10799 = n10745 & n10798 ;
  assign n10800 = ~n10793 & ~n10799 ;
  assign n10801 = ~n10788 & n10800 ;
  assign n10802 = ~n10775 & n10801 ;
  assign n10803 = \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & ~n10721 ;
  assign n10804 = ~n10756 & ~n10803 ;
  assign n10805 = ~\txethmac1_txcounters1_NibCnt_reg[11]/NET0131  & ~n10804 ;
  assign n10806 = ~n10718 & n10805 ;
  assign n10807 = ~\txethmac1_txcounters1_NibCnt_reg[11]/NET0131  & n10804 ;
  assign n10808 = n10718 & n10807 ;
  assign n10809 = ~n10806 & ~n10808 ;
  assign n10810 = ~\txethmac1_txcounters1_NibCnt_reg[10]/NET0131  & n10718 ;
  assign n10811 = ~n10721 & ~n10752 ;
  assign n10812 = ~\txethmac1_txcounters1_NibCnt_reg[10]/NET0131  & ~n10811 ;
  assign n10813 = ~n10751 & n10812 ;
  assign n10814 = ~n10810 & ~n10813 ;
  assign n10815 = n10809 & n10814 ;
  assign n10816 = ~n10713 & ~n10715 ;
  assign n10817 = ~n10710 & ~n10816 ;
  assign n10818 = ~n10751 & ~n10817 ;
  assign n10819 = \txethmac1_txcounters1_NibCnt_reg[9]/NET0131  & n10818 ;
  assign n10820 = ~\txethmac1_txcounters1_NibCnt_reg[9]/NET0131  & ~n10818 ;
  assign n10821 = ~n10712 & ~n10746 ;
  assign n10822 = ~n10748 & ~n10821 ;
  assign n10823 = \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  & ~n10750 ;
  assign n10824 = ~n10822 & n10823 ;
  assign n10825 = ~n10820 & n10824 ;
  assign n10826 = ~n10819 & ~n10825 ;
  assign n10827 = n10815 & ~n10826 ;
  assign n10828 = \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  & ~n10804 ;
  assign n10829 = n10718 & n10828 ;
  assign n10830 = \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  & n10804 ;
  assign n10831 = ~n10718 & n10830 ;
  assign n10832 = ~n10829 & ~n10831 ;
  assign n10833 = ~n10751 & ~n10811 ;
  assign n10834 = \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  & ~n10718 ;
  assign n10835 = ~n10833 & n10834 ;
  assign n10836 = n10809 & n10835 ;
  assign n10837 = n10832 & ~n10836 ;
  assign n10838 = ~n10827 & n10837 ;
  assign n10839 = ~\txethmac1_txcounters1_NibCnt_reg[12]/NET0131  & ~n10781 ;
  assign n10840 = ~n10755 & n10839 ;
  assign n10841 = ~\txethmac1_txcounters1_NibCnt_reg[12]/NET0131  & n10781 ;
  assign n10842 = n10755 & n10841 ;
  assign n10843 = ~n10840 & ~n10842 ;
  assign n10844 = n10780 & n10843 ;
  assign n10845 = n10768 & n10844 ;
  assign n10846 = ~n10838 & n10845 ;
  assign n10847 = \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & ~n10708 ;
  assign n10848 = n10704 & n10847 ;
  assign n10849 = \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & n10708 ;
  assign n10850 = ~n10704 & n10849 ;
  assign n10851 = ~n10848 & ~n10850 ;
  assign n10852 = ~\txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & ~n10708 ;
  assign n10853 = ~n10704 & n10852 ;
  assign n10854 = ~\txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & n10708 ;
  assign n10855 = n10704 & n10854 ;
  assign n10856 = ~n10853 & ~n10855 ;
  assign n10857 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & ~n10705 ;
  assign n10858 = ~\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & ~\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  ;
  assign n10859 = ~n10857 & n10858 ;
  assign n10860 = ~\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & ~n10859 ;
  assign n10861 = ~\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  ;
  assign n10862 = ~\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  & n10861 ;
  assign n10863 = ~n10857 & n10862 ;
  assign n10864 = ~\txethmac1_txcounters1_NibCnt_reg[6]/NET0131  & ~n10863 ;
  assign n10865 = ~n10860 & n10864 ;
  assign n10866 = n10856 & ~n10865 ;
  assign n10867 = n10851 & ~n10866 ;
  assign n10868 = \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  & \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  ;
  assign n10869 = ~n10705 & ~n10868 ;
  assign n10870 = \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  & n10869 ;
  assign n10871 = \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
  assign n10872 = ~\txethmac1_txcounters1_NibCnt_reg[0]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
  assign n10873 = \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  & ~n10872 ;
  assign n10874 = ~n10871 & ~n10873 ;
  assign n10875 = ~n10870 & n10874 ;
  assign n10876 = ~\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n10877 = ~n10705 & n10876 ;
  assign n10878 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n10879 = n10705 & n10878 ;
  assign n10880 = ~n10877 & ~n10879 ;
  assign n10881 = ~\txethmac1_txcounters1_NibCnt_reg[2]/NET0131  & ~n10869 ;
  assign n10882 = n10880 & ~n10881 ;
  assign n10883 = ~n10875 & n10882 ;
  assign n10884 = ~\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & ~n10857 ;
  assign n10885 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  ;
  assign n10886 = ~n10705 & n10885 ;
  assign n10887 = \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  & ~n10886 ;
  assign n10888 = ~n10884 & n10887 ;
  assign n10889 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n10890 = ~n10705 & n10889 ;
  assign n10891 = ~\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n10892 = n10705 & n10891 ;
  assign n10893 = ~n10890 & ~n10892 ;
  assign n10894 = ~n10888 & n10893 ;
  assign n10895 = ~n10883 & n10894 ;
  assign n10896 = \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  ;
  assign n10897 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  ;
  assign n10898 = ~n10705 & n10897 ;
  assign n10899 = ~n10896 & ~n10898 ;
  assign n10900 = ~n10859 & n10899 ;
  assign n10901 = ~\txethmac1_txcounters1_NibCnt_reg[5]/NET0131  & ~n10900 ;
  assign n10902 = ~\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n10903 = ~n10857 & n10902 ;
  assign n10904 = \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n10905 = n10857 & n10904 ;
  assign n10906 = ~n10903 & ~n10905 ;
  assign n10907 = ~n10901 & n10906 ;
  assign n10908 = ~n10895 & n10907 ;
  assign n10909 = ~\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n10910 = ~n10859 & n10909 ;
  assign n10911 = \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n10912 = n10859 & n10911 ;
  assign n10913 = ~n10910 & ~n10912 ;
  assign n10914 = \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  & n10900 ;
  assign n10915 = n10913 & ~n10914 ;
  assign n10916 = n10851 & n10915 ;
  assign n10917 = ~n10908 & n10916 ;
  assign n10918 = ~n10867 & ~n10917 ;
  assign n10919 = ~\txethmac1_txcounters1_NibCnt_reg[8]/NET0131  & ~n10748 ;
  assign n10920 = ~n10821 & n10919 ;
  assign n10921 = ~\txethmac1_txcounters1_NibCnt_reg[8]/NET0131  & n10748 ;
  assign n10922 = n10821 & n10921 ;
  assign n10923 = ~n10920 & ~n10922 ;
  assign n10924 = ~n10820 & n10923 ;
  assign n10925 = n10815 & n10924 ;
  assign n10926 = n10918 & n10925 ;
  assign n10927 = n10845 & n10926 ;
  assign n10928 = ~n10846 & ~n10927 ;
  assign n10929 = n10802 & n10928 ;
  assign n10930 = ~n10739 & ~n10796 ;
  assign n10931 = ~\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  & ~n10738 ;
  assign n10932 = ~n10930 & n10931 ;
  assign n10933 = ~n10738 & ~n10930 ;
  assign n10934 = ~\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  & ~n10791 ;
  assign n10935 = ~n10933 & ~n10934 ;
  assign n10936 = ~n10932 & ~n10935 ;
  assign n10937 = n10697 & n10936 ;
  assign n10938 = ~n10929 & n10937 ;
  assign n10939 = ~n10698 & ~n10938 ;
  assign n10940 = \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  & n10871 ;
  assign n10941 = \txethmac1_txstatem1_StateFCS_reg/NET0131  & ~n10694 ;
  assign n10942 = n10940 & n10941 ;
  assign n10943 = \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n10944 = ~\ethreg1_MODER_1_DataOut_reg[6]/NET0131  & ~n10943 ;
  assign n10945 = ~\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n10946 = \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n10947 = ~n10945 & ~n10946 ;
  assign n10948 = \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n10949 = \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n10950 = ~n10948 & ~n10949 ;
  assign n10951 = n10947 & n10950 ;
  assign n10952 = n10944 & n10951 ;
  assign n10953 = ~\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n10954 = ~\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n10955 = ~n10953 & ~n10954 ;
  assign n10956 = \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n10957 = ~\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  ;
  assign n10958 = ~n10956 & ~n10957 ;
  assign n10959 = n10955 & n10958 ;
  assign n10960 = ~\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n10961 = \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n10962 = ~n10960 & ~n10961 ;
  assign n10963 = ~\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n10964 = \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n10965 = ~n10963 & ~n10964 ;
  assign n10966 = n10962 & n10965 ;
  assign n10967 = n10959 & n10966 ;
  assign n10968 = \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n10969 = ~\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n10970 = ~n10968 & ~n10969 ;
  assign n10971 = ~\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n10972 = \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n10973 = ~n10971 & ~n10972 ;
  assign n10974 = n10970 & n10973 ;
  assign n10975 = \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n10976 = \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n10977 = ~n10975 & ~n10976 ;
  assign n10978 = \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  ;
  assign n10979 = \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n10980 = ~n10978 & ~n10979 ;
  assign n10981 = n10977 & n10980 ;
  assign n10982 = n10974 & n10981 ;
  assign n10983 = n10967 & n10982 ;
  assign n10984 = n10952 & n10983 ;
  assign n10985 = \txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~\wishbone_TxUnderRun_reg/NET0131  ;
  assign n10986 = ~n10694 & n10985 ;
  assign n10987 = ~n10941 & ~n10986 ;
  assign n10988 = ~\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n10989 = ~\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n10990 = ~\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n10991 = ~n10989 & ~n10990 ;
  assign n10992 = ~n10988 & n10991 ;
  assign n10993 = \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n10994 = ~\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n10995 = ~n10993 & ~n10994 ;
  assign n10996 = ~\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n10997 = ~\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n10998 = ~n10996 & ~n10997 ;
  assign n10999 = n10995 & n10998 ;
  assign n11000 = \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n11001 = \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n11002 = ~n11000 & ~n11001 ;
  assign n11003 = ~\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n11004 = ~\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n11005 = ~n11003 & ~n11004 ;
  assign n11006 = n11002 & n11005 ;
  assign n11007 = n10999 & n11006 ;
  assign n11008 = n10992 & n11007 ;
  assign n11009 = ~n10987 & n11008 ;
  assign n11010 = n10984 & n11009 ;
  assign n11011 = ~n10942 & ~n11010 ;
  assign n11012 = \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11013 = \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n11014 = ~n11012 & ~n11013 ;
  assign n11015 = ~\ethreg1_IPGR1_0_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  assign n11016 = ~\ethreg1_IPGR1_0_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n11017 = ~n11015 & ~n11016 ;
  assign n11018 = ~n11014 & n11017 ;
  assign n11019 = ~\ethreg1_IPGR1_0_DataOut_reg[0]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  ;
  assign n11020 = \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  & n11019 ;
  assign n11021 = \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131  & ~n11020 ;
  assign n11022 = ~\txethmac1_txcounters1_NibCnt_reg[1]/NET0131  & ~n11019 ;
  assign n11023 = \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
  assign n11024 = ~n11022 & ~n11023 ;
  assign n11025 = ~n11021 & n11024 ;
  assign n11026 = ~\ethreg1_IPGR1_0_DataOut_reg[3]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11027 = ~\ethreg1_IPGR1_0_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
  assign n11028 = ~n11026 & ~n11027 ;
  assign n11029 = n11017 & n11028 ;
  assign n11030 = ~n11025 & n11029 ;
  assign n11031 = ~n11018 & ~n11030 ;
  assign n11032 = \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n11033 = \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  assign n11034 = ~n11032 & ~n11033 ;
  assign n11035 = n11031 & n11034 ;
  assign n11036 = ~\ethreg1_IPGR2_0_DataOut_reg[1]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
  assign n11037 = ~\ethreg1_IPGR2_0_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
  assign n11038 = ~n11036 & ~n11037 ;
  assign n11039 = \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  assign n11040 = \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n11041 = ~n11039 & ~n11040 ;
  assign n11042 = \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
  assign n11043 = \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11044 = ~n11042 & ~n11043 ;
  assign n11045 = n11041 & n11044 ;
  assign n11046 = n11038 & n11045 ;
  assign n11047 = ~\ethreg1_IPGR2_0_DataOut_reg[0]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  ;
  assign n11048 = ~\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n11049 = ~n11047 & ~n11048 ;
  assign n11050 = \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n11051 = ~\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11052 = ~n11050 & ~n11051 ;
  assign n11053 = n11049 & n11052 ;
  assign n11054 = ~\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n11055 = ~\ethreg1_IPGR2_0_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  assign n11056 = ~n11054 & ~n11055 ;
  assign n11057 = \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[0]/NET0131  ;
  assign n11058 = \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
  assign n11059 = ~n11057 & ~n11058 ;
  assign n11060 = n11056 & n11059 ;
  assign n11061 = n11053 & n11060 ;
  assign n11062 = n11046 & n11061 ;
  assign n11063 = \CarrierSense_Tx2_reg/NET0131  & ~\ethreg1_MODER_1_DataOut_reg[2]/NET0131  ;
  assign n11064 = ~\ethreg1_IPGR1_0_DataOut_reg[6]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n11065 = ~\txethmac1_txstatem1_Rule1_reg/NET0131  & \txethmac1_txstatem1_StateIPG_reg/NET0131  ;
  assign n11066 = ~n11064 & n11065 ;
  assign n11067 = n11063 & n11066 ;
  assign n11068 = ~n11062 & n11067 ;
  assign n11069 = ~n11035 & n11068 ;
  assign n11070 = \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  & \txethmac1_txstatem1_StateJam_reg/NET0131  ;
  assign n11071 = n10871 & n11070 ;
  assign n11072 = \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131  & ~\txethmac1_RetryCnt_reg[2]/NET0131  ;
  assign n11073 = ~\ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131  & \txethmac1_RetryCnt_reg[2]/NET0131  ;
  assign n11074 = ~n11072 & ~n11073 ;
  assign n11075 = \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131  & ~\txethmac1_RetryCnt_reg[3]/NET0131  ;
  assign n11076 = ~\ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131  & \txethmac1_RetryCnt_reg[3]/NET0131  ;
  assign n11077 = ~n11075 & ~n11076 ;
  assign n11078 = n11074 & n11077 ;
  assign n11079 = ~\ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131  & ~\txethmac1_RetryCnt_reg[1]/NET0131  ;
  assign n11080 = \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131  & \txethmac1_RetryCnt_reg[1]/NET0131  ;
  assign n11081 = ~n11079 & ~n11080 ;
  assign n11082 = ~\ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131  & ~\txethmac1_RetryCnt_reg[0]/NET0131  ;
  assign n11083 = \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131  & \txethmac1_RetryCnt_reg[0]/NET0131  ;
  assign n11084 = ~n11082 & ~n11083 ;
  assign n11085 = ~n11081 & ~n11084 ;
  assign n11086 = n11078 & n11085 ;
  assign n11087 = \txethmac1_ColWindow_reg/NET0131  & ~n11086 ;
  assign n11088 = ~\txethmac1_random1_RandomLatched_reg[6]/NET0131  & ~\txethmac1_random1_RandomLatched_reg[7]/NET0131  ;
  assign n11089 = ~\txethmac1_random1_RandomLatched_reg[8]/NET0131  & ~\txethmac1_random1_RandomLatched_reg[9]/NET0131  ;
  assign n11090 = n11088 & n11089 ;
  assign n11091 = ~\txethmac1_random1_RandomLatched_reg[0]/NET0131  & ~\txethmac1_random1_RandomLatched_reg[1]/NET0131  ;
  assign n11092 = ~\txethmac1_random1_RandomLatched_reg[2]/NET0131  & ~\txethmac1_random1_RandomLatched_reg[3]/NET0131  ;
  assign n11093 = ~\txethmac1_random1_RandomLatched_reg[4]/NET0131  & ~\txethmac1_random1_RandomLatched_reg[5]/NET0131  ;
  assign n11094 = n11092 & n11093 ;
  assign n11095 = n11091 & n11094 ;
  assign n11096 = n11090 & n11095 ;
  assign n11097 = ~\ethreg1_MODER_1_DataOut_reg[0]/NET0131  & ~n11096 ;
  assign n11098 = n11087 & n11097 ;
  assign n11099 = n11071 & ~n11098 ;
  assign n11100 = \txethmac1_random1_RandomLatched_reg[1]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n11101 = \txethmac1_random1_RandomLatched_reg[4]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n11102 = ~n11100 & ~n11101 ;
  assign n11103 = ~\txethmac1_random1_RandomLatched_reg[6]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n11104 = ~\txethmac1_random1_RandomLatched_reg[1]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n11105 = ~n11103 & ~n11104 ;
  assign n11106 = n11102 & n11105 ;
  assign n11107 = ~\txethmac1_random1_RandomLatched_reg[8]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11108 = \txethmac1_random1_RandomLatched_reg[9]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n11109 = ~n11107 & ~n11108 ;
  assign n11110 = ~\txethmac1_random1_RandomLatched_reg[3]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n11111 = \txethmac1_random1_RandomLatched_reg[8]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11112 = ~n11110 & ~n11111 ;
  assign n11113 = n11109 & n11112 ;
  assign n11114 = ~\txethmac1_random1_RandomLatched_reg[4]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n11115 = \txethmac1_random1_RandomLatched_reg[3]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n11116 = ~n11114 & ~n11115 ;
  assign n11117 = \txethmac1_random1_RandomLatched_reg[6]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n11118 = \txethmac1_random1_RandomLatched_reg[7]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n11119 = ~n11117 & ~n11118 ;
  assign n11120 = n11116 & n11119 ;
  assign n11121 = n11113 & n11120 ;
  assign n11122 = n11106 & n11121 ;
  assign n11123 = \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11124 = n10871 & n11123 ;
  assign n11125 = \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  assign n11126 = \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  & \txethmac1_txstatem1_StateBackOff_reg/NET0131  ;
  assign n11127 = n11125 & n11126 ;
  assign n11128 = n11124 & n11127 ;
  assign n11129 = \txethmac1_random1_RandomLatched_reg[2]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n11130 = \txethmac1_random1_RandomLatched_reg[0]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n11131 = ~n11129 & ~n11130 ;
  assign n11132 = ~\txethmac1_random1_RandomLatched_reg[2]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n11133 = ~\txethmac1_random1_RandomLatched_reg[9]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n11134 = ~n11132 & ~n11133 ;
  assign n11135 = n11131 & n11134 ;
  assign n11136 = ~\txethmac1_random1_RandomLatched_reg[5]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11137 = \txethmac1_random1_RandomLatched_reg[5]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11138 = ~n11136 & ~n11137 ;
  assign n11139 = ~\txethmac1_random1_RandomLatched_reg[0]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n11140 = ~\txethmac1_random1_RandomLatched_reg[7]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n11141 = ~n11139 & ~n11140 ;
  assign n11142 = ~n11138 & n11141 ;
  assign n11143 = n11135 & n11142 ;
  assign n11144 = n11128 & n11143 ;
  assign n11145 = n11122 & n11144 ;
  assign n11146 = \txethmac1_txstatem1_StateIdle_reg/NET0131  & n11063 ;
  assign n11147 = \txethmac1_txstatem1_StateBackOff_reg/NET0131  & \wishbone_TxUnderRun_reg/NET0131  ;
  assign n11148 = ~n11146 & ~n11147 ;
  assign n11149 = ~n11145 & n11148 ;
  assign n11150 = ~n11099 & n11149 ;
  assign n11151 = ~n11069 & n11150 ;
  assign n11152 = n11011 & n11151 ;
  assign n11153 = n10939 & n11152 ;
  assign n11154 = ~n10690 & n10696 ;
  assign n11155 = n10688 & n11154 ;
  assign n11156 = n10936 & n11154 ;
  assign n11157 = ~n10929 & n11156 ;
  assign n11158 = ~n11155 & ~n11157 ;
  assign n11159 = \txethmac1_txstatem1_StatePAD_reg/NET0131  & ~n10694 ;
  assign n11160 = ~n10690 & n11159 ;
  assign n11161 = n10936 & n11160 ;
  assign n11162 = ~n10929 & n11161 ;
  assign n11163 = \txethmac1_txstatem1_StateData_reg[0]/NET0131  & \wishbone_TxUnderRun_reg/NET0131  ;
  assign n11164 = ~n10694 & n11163 ;
  assign n11165 = ~n10694 & ~n11164 ;
  assign n11166 = \txethmac1_txstatem1_StatePreamble_reg/NET0131  & n11124 ;
  assign n11167 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & ~\txethmac1_txstatem1_StatePAD_reg/NET0131  ;
  assign n11168 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~\txethmac1_txstatem1_StateData_reg[1]/NET0131  ;
  assign n11169 = n11167 & n11168 ;
  assign n11170 = ~n11166 & n11169 ;
  assign n11171 = ~n11165 & ~n11170 ;
  assign n11172 = ~\txethmac1_txcounters1_NibCnt_reg[11]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  ;
  assign n11173 = ~\txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11174 = n11172 & n11173 ;
  assign n11175 = ~\ethreg1_MODER_1_DataOut_reg[1]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  ;
  assign n11176 = n11125 & n11175 ;
  assign n11177 = n11174 & n11176 ;
  assign n11178 = ~\txethmac1_txcounters1_NibCnt_reg[6]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  ;
  assign n11179 = \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[9]/NET0131  ;
  assign n11180 = n11178 & n11179 ;
  assign n11181 = n10940 & n11180 ;
  assign n11182 = n11177 & n11181 ;
  assign n11183 = \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  ;
  assign n11184 = ~\maccontrol1_receivecontrol1_Pause_reg/NET0131  & ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11185 = \wishbone_TxStartFrm_reg/NET0131  & n11184 ;
  assign n11186 = ~n11183 & ~n11185 ;
  assign n11187 = \txethmac1_txstatem1_StateDefer_reg/NET0131  & n11186 ;
  assign n11188 = n11182 & n11187 ;
  assign n11189 = \txethmac1_txstatem1_StateDefer_reg/NET0131  & ~n11063 ;
  assign n11190 = ~n11182 & n11189 ;
  assign n11191 = ~\txethmac1_txstatem1_StateIdle_reg/NET0131  & ~n11071 ;
  assign n11192 = ~n11166 & n11191 ;
  assign n11193 = ~n11190 & n11192 ;
  assign n11194 = ~n11188 & n11193 ;
  assign n11195 = ~n11171 & n11194 ;
  assign n11196 = ~n11162 & n11195 ;
  assign n11197 = n11158 & n11196 ;
  assign n11198 = n11153 & n11197 ;
  assign n11199 = \txethmac1_txstatem1_StateDefer_reg/NET0131  & ~n11186 ;
  assign n11200 = ~n11182 & n11199 ;
  assign n11201 = ~\txethmac1_txstatem1_StatePreamble_reg/NET0131  & n11168 ;
  assign n11202 = ~\txethmac1_txstatem1_StateJam_reg/NET0131  & n11167 ;
  assign n11203 = n11201 & n11202 ;
  assign n11204 = ~\txethmac1_txstatem1_StateBackOff_reg/NET0131  & ~\txethmac1_txstatem1_StateIPG_reg/NET0131  ;
  assign n11205 = n11203 & n11204 ;
  assign n11206 = ~n11200 & n11205 ;
  assign n11207 = \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  & ~n11206 ;
  assign n11208 = ~\txethmac1_txcounters1_NibCnt_reg[0]/NET0131  & n11205 ;
  assign n11209 = ~n11200 & n11208 ;
  assign n11210 = ~n11207 & ~n11209 ;
  assign n11211 = n11198 & n11210 ;
  assign n11212 = \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  & n11125 ;
  assign n11213 = n11124 & n11212 ;
  assign n11214 = ~n11206 & n11213 ;
  assign n11215 = \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[9]/NET0131  ;
  assign n11216 = \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  & n11215 ;
  assign n11217 = n11214 & n11216 ;
  assign n11218 = \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  & n11217 ;
  assign n11219 = ~\txethmac1_txcounters1_NibCnt_reg[11]/NET0131  & ~n11218 ;
  assign n11220 = \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  ;
  assign n11221 = n11217 & n11220 ;
  assign n11222 = ~n11219 & ~n11221 ;
  assign n11223 = n11198 & n11222 ;
  assign n11224 = ~\txethmac1_txcounters1_NibCnt_reg[12]/NET0131  & ~n11221 ;
  assign n11225 = \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  ;
  assign n11226 = \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  & n11225 ;
  assign n11227 = n11217 & n11226 ;
  assign n11228 = ~n11224 & ~n11227 ;
  assign n11229 = n11198 & n11228 ;
  assign n11230 = ~\txethmac1_txcounters1_NibCnt_reg[10]/NET0131  & ~n11217 ;
  assign n11231 = ~n11218 & ~n11230 ;
  assign n11232 = n11198 & n11231 ;
  assign n11233 = ~\txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & ~n11227 ;
  assign n11234 = \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & n11227 ;
  assign n11235 = ~n11233 & ~n11234 ;
  assign n11236 = n11198 & n11235 ;
  assign n11237 = ~\txethmac1_txcounters1_NibCnt_reg[14]/NET0131  & ~n11234 ;
  assign n11238 = \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[14]/NET0131  ;
  assign n11239 = n11227 & n11238 ;
  assign n11240 = ~n11237 & ~n11239 ;
  assign n11241 = n11198 & n11240 ;
  assign n11242 = ~\txethmac1_txcounters1_NibCnt_reg[15]/NET0131  & ~n11239 ;
  assign n11243 = \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[15]/NET0131  ;
  assign n11244 = \txethmac1_txcounters1_NibCnt_reg[14]/NET0131  & n11243 ;
  assign n11245 = n11227 & n11244 ;
  assign n11246 = ~n11242 & ~n11245 ;
  assign n11247 = n11198 & n11246 ;
  assign n11248 = ~\txethmac1_txcounters1_NibCnt_reg[1]/NET0131  & n11205 ;
  assign n11249 = ~n11200 & n11248 ;
  assign n11250 = ~n10872 & ~n11249 ;
  assign n11251 = n10871 & ~n11206 ;
  assign n11252 = n11250 & ~n11251 ;
  assign n11253 = n11198 & n11252 ;
  assign n11254 = ~\txethmac1_txcounters1_NibCnt_reg[2]/NET0131  & ~n10871 ;
  assign n11255 = ~\txethmac1_txcounters1_NibCnt_reg[2]/NET0131  & n11205 ;
  assign n11256 = ~n11200 & n11255 ;
  assign n11257 = ~n11254 & ~n11256 ;
  assign n11258 = n10940 & ~n11206 ;
  assign n11259 = n11257 & ~n11258 ;
  assign n11260 = n11198 & n11259 ;
  assign n11261 = n11124 & ~n11206 ;
  assign n11262 = ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  & ~n10940 ;
  assign n11263 = ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  & n11205 ;
  assign n11264 = ~n11200 & n11263 ;
  assign n11265 = ~n11262 & ~n11264 ;
  assign n11266 = ~n11261 & n11265 ;
  assign n11267 = n11198 & n11266 ;
  assign n11268 = \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  & n11124 ;
  assign n11269 = ~n11206 & n11268 ;
  assign n11270 = ~\txethmac1_txcounters1_NibCnt_reg[4]/NET0131  & ~n11124 ;
  assign n11271 = ~\txethmac1_txcounters1_NibCnt_reg[4]/NET0131  & n11205 ;
  assign n11272 = ~n11200 & n11271 ;
  assign n11273 = ~n11270 & ~n11272 ;
  assign n11274 = ~n11269 & n11273 ;
  assign n11275 = n11198 & n11274 ;
  assign n11276 = n11124 & n11125 ;
  assign n11277 = ~n11206 & n11276 ;
  assign n11278 = ~\txethmac1_txcounters1_NibCnt_reg[5]/NET0131  & ~n11269 ;
  assign n11279 = ~n11277 & ~n11278 ;
  assign n11280 = n11198 & n11279 ;
  assign n11281 = ~\txethmac1_txcounters1_NibCnt_reg[6]/NET0131  & ~n11277 ;
  assign n11282 = ~n11214 & ~n11281 ;
  assign n11283 = n11198 & n11282 ;
  assign n11284 = \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & n11214 ;
  assign n11285 = ~\txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & ~n11214 ;
  assign n11286 = ~n11284 & ~n11285 ;
  assign n11287 = n11198 & n11286 ;
  assign n11288 = \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  ;
  assign n11289 = n11214 & n11288 ;
  assign n11290 = ~\txethmac1_txcounters1_NibCnt_reg[8]/NET0131  & ~n11284 ;
  assign n11291 = ~n11289 & ~n11290 ;
  assign n11292 = n11198 & n11291 ;
  assign n11293 = ~\txethmac1_txcounters1_NibCnt_reg[9]/NET0131  & ~n11289 ;
  assign n11294 = ~n11217 & ~n11293 ;
  assign n11295 = n11198 & n11294 ;
  assign n11296 = ~\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  & ~\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131  ;
  assign n11297 = ~\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  & n11296 ;
  assign n11298 = ~\txethmac1_txstatem1_StateIdle_reg/NET0131  & ~\txethmac1_txstatem1_StatePreamble_reg/NET0131  ;
  assign n11299 = ~\txethmac1_txcrc_Crc_reg[26]/NET0131  & n11298 ;
  assign n11300 = n11297 & n11299 ;
  assign n11301 = ~\txethmac1_txcrc_Crc_reg[27]/NET0131  & n11298 ;
  assign n11302 = n11297 & n11301 ;
  assign n11303 = ~\txethmac1_txstatem1_Rule1_reg/NET0131  & ~n11048 ;
  assign n11304 = ~n11041 & n11303 ;
  assign n11305 = ~n11050 & n11051 ;
  assign n11306 = n11038 & ~n11059 ;
  assign n11307 = n11044 & ~n11050 ;
  assign n11308 = ~n11306 & n11307 ;
  assign n11309 = ~n11305 & ~n11308 ;
  assign n11310 = n11056 & n11303 ;
  assign n11311 = n11309 & n11310 ;
  assign n11312 = ~n11304 & ~n11311 ;
  assign n11313 = ~\ethreg1_IPGT_0_DataOut_reg[6]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n11314 = \txethmac1_txstatem1_Rule1_reg/NET0131  & ~n11313 ;
  assign n11315 = \txethmac1_txstatem1_StateIPG_reg/NET0131  & ~n11314 ;
  assign n11316 = \ethreg1_IPGT_0_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11317 = \ethreg1_IPGT_0_DataOut_reg[4]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n11318 = ~n11316 & ~n11317 ;
  assign n11319 = ~\ethreg1_IPGT_0_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  assign n11320 = ~\ethreg1_IPGT_0_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
  assign n11321 = ~n11319 & ~n11320 ;
  assign n11322 = ~n11318 & n11321 ;
  assign n11323 = ~\ethreg1_IPGT_0_DataOut_reg[1]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
  assign n11324 = \ethreg1_IPGT_0_DataOut_reg[0]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[0]/NET0131  ;
  assign n11325 = ~n11323 & n11324 ;
  assign n11326 = \ethreg1_IPGT_0_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
  assign n11327 = \ethreg1_IPGT_0_DataOut_reg[1]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
  assign n11328 = ~n11326 & ~n11327 ;
  assign n11329 = ~n11325 & n11328 ;
  assign n11330 = ~\ethreg1_IPGT_0_DataOut_reg[3]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
  assign n11331 = ~\ethreg1_IPGT_0_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
  assign n11332 = ~n11330 & ~n11331 ;
  assign n11333 = n11321 & n11332 ;
  assign n11334 = ~n11329 & n11333 ;
  assign n11335 = ~n11322 & ~n11334 ;
  assign n11336 = \ethreg1_IPGT_0_DataOut_reg[6]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
  assign n11337 = \ethreg1_IPGT_0_DataOut_reg[5]/NET0131  & ~\txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
  assign n11338 = ~n11336 & ~n11337 ;
  assign n11339 = \txethmac1_txstatem1_StateIPG_reg/NET0131  & n11338 ;
  assign n11340 = n11335 & n11339 ;
  assign n11341 = ~n11315 & ~n11340 ;
  assign n11342 = n11312 & ~n11341 ;
  assign n11343 = ~\txethmac1_txstatem1_StateIdle_reg/NET0131  & ~n11342 ;
  assign n11344 = \txethmac1_txstatem1_StateIdle_reg/NET0131  & n11183 ;
  assign n11345 = \txethmac1_txstatem1_StateIdle_reg/NET0131  & \wishbone_TxStartFrm_reg/NET0131  ;
  assign n11346 = n11184 & n11345 ;
  assign n11347 = ~n11344 & ~n11346 ;
  assign n11348 = ~n11063 & ~n11347 ;
  assign n11349 = ~n11343 & ~n11348 ;
  assign n11350 = n11153 & n11349 ;
  assign n11351 = ~\txethmac1_txstatem1_StateDefer_reg/NET0131  & n11153 ;
  assign n11352 = ~n11190 & ~n11351 ;
  assign n11353 = ~n10648 & n10654 ;
  assign n11354 = \ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mtxd_pad_o[3]_pad  ;
  assign n11355 = ~\ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mrxd_pad_i[3]_pad  ;
  assign n11356 = ~n11354 & ~n11355 ;
  assign n11357 = \rxethmac1_crcrx_Crc_reg[28]/NET0131  & ~n11356 ;
  assign n11358 = ~\rxethmac1_crcrx_Crc_reg[28]/NET0131  & n11356 ;
  assign n11359 = ~n11357 & ~n11358 ;
  assign n11360 = ~n10660 & ~n11359 ;
  assign n11361 = n10660 & n11359 ;
  assign n11362 = ~n11360 & ~n11361 ;
  assign n11363 = ~\rxethmac1_crcrx_Crc_reg[19]/NET0131  & n11362 ;
  assign n11364 = n11353 & n11363 ;
  assign n11365 = ~\rxethmac1_crcrx_Crc_reg[19]/NET0131  & n10663 ;
  assign n11366 = n10663 & n11362 ;
  assign n11367 = n11353 & n11366 ;
  assign n11368 = ~n11365 & ~n11367 ;
  assign n11369 = ~n11364 & ~n11368 ;
  assign n11370 = ~n10660 & n10674 ;
  assign n11371 = n10660 & ~n10674 ;
  assign n11372 = ~n11370 & ~n11371 ;
  assign n11373 = ~\rxethmac1_crcrx_Crc_reg[20]/NET0131  & ~n11372 ;
  assign n11374 = n11353 & n11373 ;
  assign n11375 = ~\rxethmac1_crcrx_Crc_reg[20]/NET0131  & n10663 ;
  assign n11376 = n10663 & ~n11372 ;
  assign n11377 = n11353 & n11376 ;
  assign n11378 = ~n11375 & ~n11377 ;
  assign n11379 = ~n11374 & ~n11378 ;
  assign n11380 = ~\rxethmac1_crcrx_Crc_reg[26]/NET0131  & ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n11381 = ~n10582 & n11380 ;
  assign n11382 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & ~n11162 ;
  assign n11383 = n11158 & n11382 ;
  assign n11384 = ~n11171 & ~n11383 ;
  assign n11385 = n11153 & n11384 ;
  assign n11386 = ~\txethmac1_txstatem1_StateJam_reg/NET0131  & n11165 ;
  assign n11387 = ~\txethmac1_txstatem1_StateJam_reg/NET0131  & n11169 ;
  assign n11388 = ~n11166 & n11387 ;
  assign n11389 = ~n11386 & ~n11388 ;
  assign n11390 = \txethmac1_ColWindow_reg/NET0131  & n11071 ;
  assign n11391 = ~n11086 & n11390 ;
  assign n11392 = n11097 & n11391 ;
  assign n11393 = n11389 & ~n11392 ;
  assign n11394 = n11153 & n11393 ;
  assign n11395 = ~n11162 & ~n11171 ;
  assign n11396 = n11158 & n11395 ;
  assign n11397 = ~n10929 & n10936 ;
  assign n11398 = ~n10688 & n10696 ;
  assign n11399 = ~n11397 & n11398 ;
  assign n11400 = ~\txethmac1_txstatem1_StatePAD_reg/NET0131  & ~n11399 ;
  assign n11401 = n11396 & ~n11400 ;
  assign n11402 = ~\txethmac1_StopExcessiveDeferOccured_reg/NET0131  & \txethmac1_txstatem1_StateDefer_reg/NET0131  ;
  assign n11403 = ~n11186 & n11402 ;
  assign n11404 = n11182 & n11403 ;
  assign n11405 = ~\wishbone_TxUnderRun_reg/NET0131  & ~n11071 ;
  assign n11406 = \txethmac1_ColWindow_reg/NET0131  & ~\wishbone_TxUnderRun_reg/NET0131  ;
  assign n11407 = ~n11086 & n11406 ;
  assign n11408 = ~n11405 & ~n11407 ;
  assign n11409 = ~n11404 & ~n11408 ;
  assign n11410 = n11011 & n11409 ;
  assign n11411 = n10939 & n11410 ;
  assign n11412 = ~n11097 & n11390 ;
  assign n11413 = ~n11145 & ~n11412 ;
  assign n11414 = \txethmac1_RetryCnt_reg[0]/NET0131  & ~n11413 ;
  assign n11415 = ~\txethmac1_RetryCnt_reg[0]/NET0131  & n11413 ;
  assign n11416 = ~n11414 & ~n11415 ;
  assign n11417 = n11411 & n11416 ;
  assign n11418 = \txethmac1_RetryCnt_reg[0]/NET0131  & \txethmac1_RetryCnt_reg[1]/NET0131  ;
  assign n11419 = ~n11413 & n11418 ;
  assign n11420 = ~\txethmac1_RetryCnt_reg[2]/NET0131  & ~n11419 ;
  assign n11421 = \txethmac1_RetryCnt_reg[2]/NET0131  & n11418 ;
  assign n11422 = ~n11413 & n11421 ;
  assign n11423 = ~n11420 & ~n11422 ;
  assign n11424 = n11411 & n11423 ;
  assign n11425 = ~\txethmac1_RetryCnt_reg[3]/NET0131  & ~n11422 ;
  assign n11426 = \txethmac1_RetryCnt_reg[2]/NET0131  & \txethmac1_RetryCnt_reg[3]/NET0131  ;
  assign n11427 = n11418 & n11426 ;
  assign n11428 = ~n11413 & n11427 ;
  assign n11429 = ~n11425 & ~n11428 ;
  assign n11430 = n11411 & n11429 ;
  assign n11431 = ~\txethmac1_RetryCnt_reg[1]/NET0131  & ~n11414 ;
  assign n11432 = ~n11419 & ~n11431 ;
  assign n11433 = n11411 & n11432 ;
  assign n11434 = ~\maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11435 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & \txethmac1_txstatem1_StateData_reg[1]/NET0131  ;
  assign n11436 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[7]/NET0131  ;
  assign n11437 = n11435 & ~n11436 ;
  assign n11438 = ~n11434 & n11437 ;
  assign n11439 = ~\maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11440 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[3]/NET0131  ;
  assign n11441 = \txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n11440 ;
  assign n11442 = ~n11439 & n11441 ;
  assign n11443 = ~n11438 & ~n11442 ;
  assign n11444 = ~\txethmac1_txcrc_Crc_reg[28]/NET0131  & ~n11443 ;
  assign n11445 = \txethmac1_txcrc_Crc_reg[28]/NET0131  & n11443 ;
  assign n11446 = ~n11444 & ~n11445 ;
  assign n11447 = ~\maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11448 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[4]/NET0131  ;
  assign n11449 = n11435 & ~n11448 ;
  assign n11450 = ~n11447 & n11449 ;
  assign n11451 = ~\maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11452 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[0]/NET0131  ;
  assign n11453 = \txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n11452 ;
  assign n11454 = ~n11451 & n11453 ;
  assign n11455 = ~n11450 & ~n11454 ;
  assign n11456 = \txethmac1_txcrc_Crc_reg[31]/NET0131  & ~n11455 ;
  assign n11457 = ~\txethmac1_txcrc_Crc_reg[31]/NET0131  & n11455 ;
  assign n11458 = ~n11456 & ~n11457 ;
  assign n11459 = n11446 & ~n11458 ;
  assign n11460 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & ~n11459 ;
  assign n11461 = ~n11446 & n11458 ;
  assign n11462 = ~\txethmac1_txcrc_Crc_reg[22]/NET0131  & ~n11461 ;
  assign n11463 = n11460 & n11462 ;
  assign n11464 = n11297 & n11298 ;
  assign n11465 = ~\txethmac1_txcrc_Crc_reg[22]/NET0131  & n11464 ;
  assign n11466 = ~n11461 & n11464 ;
  assign n11467 = n11460 & n11466 ;
  assign n11468 = ~n11465 & ~n11467 ;
  assign n11469 = ~n11463 & ~n11468 ;
  assign n11470 = ~\maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11471 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[2]/NET0131  ;
  assign n11472 = \txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n11471 ;
  assign n11473 = ~n11470 & n11472 ;
  assign n11474 = ~\maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11475 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[6]/NET0131  ;
  assign n11476 = n11435 & ~n11475 ;
  assign n11477 = ~n11474 & n11476 ;
  assign n11478 = ~n11473 & ~n11477 ;
  assign n11479 = ~\txethmac1_txcrc_Crc_reg[29]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11480 = ~n11478 & n11479 ;
  assign n11481 = \txethmac1_txcrc_Crc_reg[29]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11482 = n11478 & n11481 ;
  assign n11483 = ~n11480 & ~n11482 ;
  assign n11484 = \txethmac1_txcrc_Crc_reg[23]/NET0131  & n11483 ;
  assign n11485 = ~\txethmac1_txcrc_Crc_reg[23]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11486 = ~\txethmac1_txcrc_Crc_reg[29]/NET0131  & n11485 ;
  assign n11487 = ~n11478 & n11486 ;
  assign n11488 = \txethmac1_txcrc_Crc_reg[29]/NET0131  & n11485 ;
  assign n11489 = n11478 & n11488 ;
  assign n11490 = ~n11487 & ~n11489 ;
  assign n11491 = n11464 & n11490 ;
  assign n11492 = ~n11484 & n11491 ;
  assign n11493 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[5]/NET0131  ;
  assign n11494 = \txethmac1_txstatem1_StateData_reg[1]/NET0131  & ~n11493 ;
  assign n11495 = ~\maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11496 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n11495 ;
  assign n11497 = n11494 & n11496 ;
  assign n11498 = ~\maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n11499 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\wishbone_TxData_reg[1]/NET0131  ;
  assign n11500 = \txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n11499 ;
  assign n11501 = ~n11498 & n11500 ;
  assign n11502 = ~n11497 & ~n11501 ;
  assign n11503 = ~\txethmac1_txcrc_Crc_reg[30]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11504 = ~n11502 & n11503 ;
  assign n11505 = \txethmac1_txcrc_Crc_reg[30]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11506 = n11502 & n11505 ;
  assign n11507 = ~n11504 & ~n11506 ;
  assign n11508 = \txethmac1_txcrc_Crc_reg[24]/NET0131  & n11507 ;
  assign n11509 = ~\txethmac1_txcrc_Crc_reg[24]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11510 = ~\txethmac1_txcrc_Crc_reg[30]/NET0131  & n11509 ;
  assign n11511 = ~n11502 & n11510 ;
  assign n11512 = \txethmac1_txcrc_Crc_reg[30]/NET0131  & n11509 ;
  assign n11513 = n11502 & n11512 ;
  assign n11514 = ~n11511 & ~n11513 ;
  assign n11515 = n11464 & n11514 ;
  assign n11516 = ~n11508 & n11515 ;
  assign n11517 = ~\txethmac1_txstatem1_StateIPG_reg/NET0131  & ~n11190 ;
  assign n11518 = ~n11342 & ~n11517 ;
  assign n11519 = n11153 & n11518 ;
  assign n11520 = ~\txethmac1_txstatem1_StateBackOff_reg/NET0131  & ~n11392 ;
  assign n11521 = n11153 & ~n11520 ;
  assign n11522 = \ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mtxd_pad_o[0]_pad  ;
  assign n11523 = ~\ethreg1_MODER_0_DataOut_reg[7]/NET0131  & \mrxd_pad_i[0]_pad  ;
  assign n11524 = ~n11522 & ~n11523 ;
  assign n11525 = \rxethmac1_crcrx_Crc_reg[31]/NET0131  & ~n11524 ;
  assign n11526 = ~\rxethmac1_crcrx_Crc_reg[31]/NET0131  & n11524 ;
  assign n11527 = ~n11525 & ~n11526 ;
  assign n11528 = ~n11359 & n11527 ;
  assign n11529 = n11359 & ~n11527 ;
  assign n11530 = ~n11528 & ~n11529 ;
  assign n11531 = n11353 & ~n11530 ;
  assign n11532 = ~\rxethmac1_crcrx_Crc_reg[22]/NET0131  & n10663 ;
  assign n11533 = ~n11531 & n11532 ;
  assign n11534 = \rxethmac1_crcrx_Crc_reg[22]/NET0131  & n10663 ;
  assign n11535 = n11531 & n11534 ;
  assign n11536 = ~n11533 & ~n11535 ;
  assign n11537 = \txethmac1_txcrc_Crc_reg[31]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11538 = n11455 & n11537 ;
  assign n11539 = ~\txethmac1_txcrc_Crc_reg[31]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11540 = ~n11455 & n11539 ;
  assign n11541 = ~n11538 & ~n11540 ;
  assign n11542 = \txethmac1_txcrc_Crc_reg[25]/NET0131  & n11541 ;
  assign n11543 = ~\txethmac1_txcrc_Crc_reg[25]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11544 = ~\txethmac1_txcrc_Crc_reg[31]/NET0131  & n11543 ;
  assign n11545 = ~n11455 & n11544 ;
  assign n11546 = \txethmac1_txcrc_Crc_reg[31]/NET0131  & n11543 ;
  assign n11547 = n11455 & n11546 ;
  assign n11548 = ~n11545 & ~n11547 ;
  assign n11549 = n11464 & n11548 ;
  assign n11550 = ~n11542 & n11549 ;
  assign n11551 = ~n11010 & ~n11164 ;
  assign n11552 = \txethmac1_ColWindow_reg/NET0131  & n11086 ;
  assign n11553 = n11171 & n11552 ;
  assign n11554 = ~\txethmac1_ColWindow_reg/NET0131  & ~n11164 ;
  assign n11555 = ~n11165 & n11554 ;
  assign n11556 = ~n11170 & n11555 ;
  assign n11557 = ~n11404 & ~n11556 ;
  assign n11558 = ~n11553 & n11557 ;
  assign n11559 = n11551 & n11558 ;
  assign n11560 = ~n10942 & n11559 ;
  assign n11561 = n10939 & n11560 ;
  assign n11562 = ~\txethmac1_TxDone_reg/NET0131  & ~n10942 ;
  assign n11563 = n10939 & n11562 ;
  assign n11564 = ~\txethmac1_StatusLatch_reg/NET0131  & n11183 ;
  assign n11565 = ~\txethmac1_StatusLatch_reg/NET0131  & \wishbone_TxStartFrm_reg/NET0131  ;
  assign n11566 = n11184 & n11565 ;
  assign n11567 = ~n11564 & ~n11566 ;
  assign n11568 = ~n11563 & n11567 ;
  assign n11569 = ~\ethreg1_ResetTxCIrq_sync2_reg/NET0131  & \ethreg1_SetTxCIrq_txclk_reg/NET0131  ;
  assign n11570 = \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  & \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131  ;
  assign n11571 = ~n11569 & ~n11570 ;
  assign n11572 = ~n10942 & ~n11569 ;
  assign n11573 = n10939 & n11572 ;
  assign n11574 = ~n11571 & ~n11573 ;
  assign n11575 = n10654 & n11527 ;
  assign n11576 = ~n10648 & n11575 ;
  assign n11577 = ~\rxethmac1_crcrx_Crc_reg[15]/NET0131  & n10663 ;
  assign n11578 = ~n11576 & n11577 ;
  assign n11579 = \rxethmac1_crcrx_Crc_reg[15]/NET0131  & n10663 ;
  assign n11580 = n11576 & n11579 ;
  assign n11581 = ~n11578 & ~n11580 ;
  assign n11582 = ~\rxethmac1_crcrx_Crc_reg[16]/NET0131  & ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n11583 = ~n10582 & n11582 ;
  assign n11584 = ~\txethmac1_txcrc_Crc_reg[28]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11585 = ~n11443 & n11584 ;
  assign n11586 = \txethmac1_txcrc_Crc_reg[28]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11587 = n11443 & n11586 ;
  assign n11588 = ~n11585 & ~n11587 ;
  assign n11589 = \txethmac1_txcrc_Crc_reg[18]/NET0131  & n11588 ;
  assign n11590 = ~\txethmac1_txcrc_Crc_reg[18]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11591 = ~\txethmac1_txcrc_Crc_reg[28]/NET0131  & n11590 ;
  assign n11592 = ~n11443 & n11591 ;
  assign n11593 = \txethmac1_txcrc_Crc_reg[28]/NET0131  & n11590 ;
  assign n11594 = n11443 & n11593 ;
  assign n11595 = ~n11592 & ~n11594 ;
  assign n11596 = n11464 & n11595 ;
  assign n11597 = ~n11589 & n11596 ;
  assign n11598 = ~n11443 & ~n11478 ;
  assign n11599 = n11443 & n11478 ;
  assign n11600 = ~n11598 & ~n11599 ;
  assign n11601 = \txethmac1_txcrc_Crc_reg[28]/NET0131  & ~\txethmac1_txcrc_Crc_reg[29]/NET0131  ;
  assign n11602 = ~\txethmac1_txcrc_Crc_reg[28]/NET0131  & \txethmac1_txcrc_Crc_reg[29]/NET0131  ;
  assign n11603 = ~n11601 & ~n11602 ;
  assign n11604 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & ~n11603 ;
  assign n11605 = ~n11600 & n11604 ;
  assign n11606 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n11603 ;
  assign n11607 = n11600 & n11606 ;
  assign n11608 = ~n11605 & ~n11607 ;
  assign n11609 = \txethmac1_txcrc_Crc_reg[19]/NET0131  & n11608 ;
  assign n11610 = ~\txethmac1_txcrc_Crc_reg[19]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11611 = ~n11603 & n11610 ;
  assign n11612 = ~n11600 & n11611 ;
  assign n11613 = n11603 & n11610 ;
  assign n11614 = n11600 & n11613 ;
  assign n11615 = ~n11612 & ~n11614 ;
  assign n11616 = n11464 & n11615 ;
  assign n11617 = ~n11609 & n11616 ;
  assign n11618 = \txethmac1_txcrc_Crc_reg[29]/NET0131  & ~n11478 ;
  assign n11619 = ~\txethmac1_txcrc_Crc_reg[29]/NET0131  & n11478 ;
  assign n11620 = ~n11618 & ~n11619 ;
  assign n11621 = \txethmac1_txcrc_Crc_reg[30]/NET0131  & ~n11502 ;
  assign n11622 = ~\txethmac1_txcrc_Crc_reg[30]/NET0131  & n11502 ;
  assign n11623 = ~n11621 & ~n11622 ;
  assign n11624 = n11620 & n11623 ;
  assign n11625 = ~n11620 & ~n11623 ;
  assign n11626 = ~n11624 & ~n11625 ;
  assign n11627 = ~\txethmac1_txcrc_Crc_reg[20]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n11628 = n11626 & n11627 ;
  assign n11629 = ~\txethmac1_txcrc_Crc_reg[20]/NET0131  & n11464 ;
  assign n11630 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n11464 ;
  assign n11631 = n11626 & n11630 ;
  assign n11632 = ~n11629 & ~n11631 ;
  assign n11633 = ~n11628 & ~n11632 ;
  assign n11634 = n10654 & n11359 ;
  assign n11635 = ~n10648 & n11634 ;
  assign n11636 = ~\rxethmac1_crcrx_Crc_reg[12]/NET0131  & n10663 ;
  assign n11637 = ~n11635 & n11636 ;
  assign n11638 = \rxethmac1_crcrx_Crc_reg[12]/NET0131  & n10663 ;
  assign n11639 = n11635 & n11638 ;
  assign n11640 = ~n11637 & ~n11639 ;
  assign n11641 = ~\rxethmac1_crcrx_Crc_reg[18]/NET0131  & n10663 ;
  assign n11642 = ~n11635 & n11641 ;
  assign n11643 = \rxethmac1_crcrx_Crc_reg[18]/NET0131  & n10663 ;
  assign n11644 = n11635 & n11643 ;
  assign n11645 = ~n11642 & ~n11644 ;
  assign n11646 = n11458 & n11623 ;
  assign n11647 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & ~n11646 ;
  assign n11648 = ~n11458 & ~n11623 ;
  assign n11649 = ~\txethmac1_txcrc_Crc_reg[21]/NET0131  & ~n11648 ;
  assign n11650 = n11647 & n11649 ;
  assign n11651 = ~\txethmac1_txcrc_Crc_reg[21]/NET0131  & n11464 ;
  assign n11652 = n11464 & ~n11648 ;
  assign n11653 = n11647 & n11652 ;
  assign n11654 = ~n11651 & ~n11653 ;
  assign n11655 = ~n11650 & ~n11654 ;
  assign n11656 = ~\rxethmac1_crcrx_Crc_reg[11]/NET0131  & n10663 ;
  assign n11657 = ~n11576 & n11656 ;
  assign n11658 = \rxethmac1_crcrx_Crc_reg[11]/NET0131  & n10663 ;
  assign n11659 = n11576 & n11658 ;
  assign n11660 = ~n11657 & ~n11659 ;
  assign n11661 = \ethreg1_ResetRxCIrq_sync2_reg/NET0131  & ~\ethreg1_ResetRxCIrq_sync3_reg/NET0131  ;
  assign n11662 = \ethreg1_SetRxCIrq_rxclk_reg/NET0131  & ~n11661 ;
  assign n11663 = \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n11664 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n11665 = n11663 & n11664 ;
  assign n11666 = \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n11667 = \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  & n11666 ;
  assign n11668 = n11665 & n11667 ;
  assign n11669 = \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n11670 = \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  & n11669 ;
  assign n11671 = n11668 & n11670 ;
  assign n11672 = \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n11673 = \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  & n11672 ;
  assign n11674 = n11671 & n11673 ;
  assign n11675 = \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  & n11674 ;
  assign n11676 = n10638 & ~n11675 ;
  assign n11677 = \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n11678 = n11675 & n11677 ;
  assign n11679 = ~n11676 & ~n11678 ;
  assign n11680 = ~\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  & ~n11675 ;
  assign n11681 = \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n11682 = n11674 & n11681 ;
  assign n11683 = ~\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  & ~n11682 ;
  assign n11684 = ~n11680 & n11683 ;
  assign n11685 = n10598 & ~n11674 ;
  assign n11686 = \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n11687 = n11674 & n11686 ;
  assign n11688 = ~n11685 & ~n11687 ;
  assign n11689 = ~n11684 & ~n11688 ;
  assign n11690 = \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  & n11671 ;
  assign n11691 = ~\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  & ~n11690 ;
  assign n11692 = \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n11693 = n11671 & n11692 ;
  assign n11694 = ~\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  & ~n11693 ;
  assign n11695 = ~n11691 & n11694 ;
  assign n11696 = n10624 & ~n11671 ;
  assign n11697 = ~\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n11698 = n11671 & n11697 ;
  assign n11699 = ~n11696 & ~n11698 ;
  assign n11700 = ~n11695 & n11699 ;
  assign n11701 = n10617 & ~n11693 ;
  assign n11702 = \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n11703 = n11693 & n11702 ;
  assign n11704 = ~n11701 & ~n11703 ;
  assign n11705 = n10641 & ~n11690 ;
  assign n11706 = \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n11707 = n11690 & n11706 ;
  assign n11708 = ~n11705 & ~n11707 ;
  assign n11709 = n11704 & n11708 ;
  assign n11710 = ~n11700 & n11709 ;
  assign n11711 = n10597 & ~n11668 ;
  assign n11712 = \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11713 = n11668 & n11712 ;
  assign n11714 = ~n11711 & ~n11713 ;
  assign n11715 = \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  & n11668 ;
  assign n11716 = n10620 & ~n11715 ;
  assign n11717 = \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n11718 = n11715 & n11717 ;
  assign n11719 = ~n11716 & ~n11718 ;
  assign n11720 = n11714 & n11719 ;
  assign n11721 = \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n11722 = n11668 & n11721 ;
  assign n11723 = ~\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  & ~n11722 ;
  assign n11724 = ~\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  & ~n11671 ;
  assign n11725 = ~n11723 & n11724 ;
  assign n11726 = ~\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  & ~n11715 ;
  assign n11727 = ~\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  & ~n11722 ;
  assign n11728 = ~n11726 & n11727 ;
  assign n11729 = ~n11725 & ~n11728 ;
  assign n11730 = ~n11720 & n11729 ;
  assign n11731 = \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  & n11665 ;
  assign n11732 = ~\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  & ~n11731 ;
  assign n11733 = \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n11734 = n11665 & n11733 ;
  assign n11735 = ~\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  & ~n11734 ;
  assign n11736 = ~n11732 & n11735 ;
  assign n11737 = n10611 & ~n11665 ;
  assign n11738 = ~\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11739 = n11665 & n11738 ;
  assign n11740 = ~n11737 & ~n11739 ;
  assign n11741 = ~n11736 & n11740 ;
  assign n11742 = n10586 & ~n11734 ;
  assign n11743 = \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n11744 = n11734 & n11743 ;
  assign n11745 = ~n11742 & ~n11744 ;
  assign n11746 = n10587 & ~n11731 ;
  assign n11747 = \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n11748 = n11731 & n11747 ;
  assign n11749 = ~n11746 & ~n11748 ;
  assign n11750 = n11745 & n11749 ;
  assign n11751 = ~n11741 & n11750 ;
  assign n11752 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n11753 = ~\ethreg1_MODER_1_DataOut_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n11754 = ~n11752 & ~n11753 ;
  assign n11755 = ~\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  & ~n10612 ;
  assign n11756 = ~n10608 & n11755 ;
  assign n11757 = ~n11754 & ~n11756 ;
  assign n11758 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & n11663 ;
  assign n11759 = ~\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  & ~n11752 ;
  assign n11760 = ~n11758 & ~n11759 ;
  assign n11761 = \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  & ~n11760 ;
  assign n11762 = ~n10608 & ~n10612 ;
  assign n11763 = \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  & ~n11762 ;
  assign n11764 = ~n11761 & ~n11763 ;
  assign n11765 = ~n11757 & n11764 ;
  assign n11766 = ~\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  & ~n11758 ;
  assign n11767 = ~\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  & ~n11665 ;
  assign n11768 = ~n11766 & n11767 ;
  assign n11769 = ~\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  & n11760 ;
  assign n11770 = ~n11768 & ~n11769 ;
  assign n11771 = ~n11765 & n11770 ;
  assign n11772 = n10626 & ~n11665 ;
  assign n11773 = \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11774 = n11665 & n11773 ;
  assign n11775 = ~n11772 & ~n11774 ;
  assign n11776 = n10616 & ~n11758 ;
  assign n11777 = \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n11778 = n11758 & n11777 ;
  assign n11779 = ~n11776 & ~n11778 ;
  assign n11780 = n11775 & n11779 ;
  assign n11781 = n11750 & n11780 ;
  assign n11782 = ~n11771 & n11781 ;
  assign n11783 = ~n11751 & ~n11782 ;
  assign n11784 = ~\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  & ~n11734 ;
  assign n11785 = ~\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  & ~n11668 ;
  assign n11786 = ~n11784 & n11785 ;
  assign n11787 = n10600 & ~n11668 ;
  assign n11788 = ~\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11789 = n11668 & n11788 ;
  assign n11790 = ~n11787 & ~n11789 ;
  assign n11791 = ~n11786 & n11790 ;
  assign n11792 = n11729 & n11791 ;
  assign n11793 = n11783 & n11792 ;
  assign n11794 = ~n11730 & ~n11793 ;
  assign n11795 = n10609 & ~n11722 ;
  assign n11796 = \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
  assign n11797 = n11722 & n11796 ;
  assign n11798 = ~n11795 & ~n11797 ;
  assign n11799 = n10627 & ~n11671 ;
  assign n11800 = \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n11801 = n11671 & n11800 ;
  assign n11802 = ~n11799 & ~n11801 ;
  assign n11803 = n11798 & n11802 ;
  assign n11804 = n11709 & n11803 ;
  assign n11805 = n11794 & n11804 ;
  assign n11806 = ~n11710 & ~n11805 ;
  assign n11807 = ~\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  & ~n11693 ;
  assign n11808 = ~\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  & ~n11674 ;
  assign n11809 = ~n11807 & n11808 ;
  assign n11810 = n10594 & ~n11674 ;
  assign n11811 = ~\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n11812 = n11674 & n11811 ;
  assign n11813 = ~n11810 & ~n11812 ;
  assign n11814 = ~n11809 & n11813 ;
  assign n11815 = ~n11684 & n11814 ;
  assign n11816 = n11806 & n11815 ;
  assign n11817 = ~n11689 & ~n11816 ;
  assign n11818 = n11679 & n11817 ;
  assign n11819 = \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n11820 = ~n11675 & n11819 ;
  assign n11821 = \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n11822 = n11675 & n11821 ;
  assign n11823 = ~n11820 & ~n11822 ;
  assign n11824 = \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n11825 = ~n11674 & n11824 ;
  assign n11826 = \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n11827 = n11674 & n11826 ;
  assign n11828 = ~n11825 & ~n11827 ;
  assign n11829 = \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n11830 = ~n11693 & n11829 ;
  assign n11831 = \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n11832 = n11693 & n11831 ;
  assign n11833 = ~n11830 & ~n11832 ;
  assign n11834 = n11828 & n11833 ;
  assign n11835 = n11823 & n11834 ;
  assign n11836 = ~\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  & ~n11682 ;
  assign n11837 = ~n11680 & n11836 ;
  assign n11838 = ~\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n11839 = ~n11674 & n11838 ;
  assign n11840 = ~\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n11841 = n11674 & n11840 ;
  assign n11842 = ~n11839 & ~n11841 ;
  assign n11843 = n11823 & ~n11842 ;
  assign n11844 = ~n11837 & ~n11843 ;
  assign n11845 = ~n11835 & n11844 ;
  assign n11846 = ~\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n11847 = ~n11671 & n11846 ;
  assign n11848 = ~\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n11849 = n11671 & n11848 ;
  assign n11850 = ~n11847 & ~n11849 ;
  assign n11851 = ~\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & ~n11671 ;
  assign n11852 = ~n11723 & n11851 ;
  assign n11853 = n11850 & ~n11852 ;
  assign n11854 = \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n11855 = ~n11671 & n11854 ;
  assign n11856 = \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n11857 = n11671 & n11856 ;
  assign n11858 = ~n11855 & ~n11857 ;
  assign n11859 = \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n11860 = ~n11690 & n11859 ;
  assign n11861 = \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n11862 = n11690 & n11861 ;
  assign n11863 = ~n11860 & ~n11862 ;
  assign n11864 = n11858 & n11863 ;
  assign n11865 = ~n11853 & n11864 ;
  assign n11866 = \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11867 = ~n11668 & n11866 ;
  assign n11868 = \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11869 = n11668 & n11868 ;
  assign n11870 = ~n11867 & ~n11869 ;
  assign n11871 = ~\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11872 = ~n11668 & n11871 ;
  assign n11873 = ~\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n11874 = n11668 & n11873 ;
  assign n11875 = ~n11872 & ~n11874 ;
  assign n11876 = ~\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  & ~n11722 ;
  assign n11877 = ~n11726 & n11876 ;
  assign n11878 = n11875 & ~n11877 ;
  assign n11879 = ~n11870 & n11878 ;
  assign n11880 = ~\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11881 = ~n11665 & n11880 ;
  assign n11882 = ~\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11883 = n11665 & n11882 ;
  assign n11884 = ~n11881 & ~n11883 ;
  assign n11885 = ~\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & ~n11734 ;
  assign n11886 = ~n11732 & n11885 ;
  assign n11887 = n11884 & ~n11886 ;
  assign n11888 = \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n11889 = ~n11734 & n11888 ;
  assign n11890 = \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n11891 = n11734 & n11890 ;
  assign n11892 = ~n11889 & ~n11891 ;
  assign n11893 = \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n11894 = ~n11731 & n11893 ;
  assign n11895 = \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
  assign n11896 = n11731 & n11895 ;
  assign n11897 = ~n11894 & ~n11896 ;
  assign n11898 = n11892 & n11897 ;
  assign n11899 = ~n11887 & n11898 ;
  assign n11900 = ~\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & n11754 ;
  assign n11901 = ~\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n11902 = \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n11903 = \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n11904 = ~n11902 & ~n11903 ;
  assign n11905 = ~n11901 & ~n11904 ;
  assign n11906 = ~n11900 & n11905 ;
  assign n11907 = \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & ~n11760 ;
  assign n11908 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & ~n11754 ;
  assign n11909 = ~n11907 & ~n11908 ;
  assign n11910 = ~n11906 & n11909 ;
  assign n11911 = ~\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  & ~n11665 ;
  assign n11912 = ~n11766 & n11911 ;
  assign n11913 = ~\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & n11760 ;
  assign n11914 = ~n11912 & ~n11913 ;
  assign n11915 = ~n11910 & n11914 ;
  assign n11916 = \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11917 = ~n11665 & n11916 ;
  assign n11918 = \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n11919 = n11665 & n11918 ;
  assign n11920 = ~n11917 & ~n11919 ;
  assign n11921 = \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n11922 = ~n11758 & n11921 ;
  assign n11923 = \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n11924 = n11758 & n11923 ;
  assign n11925 = ~n11922 & ~n11924 ;
  assign n11926 = n11920 & n11925 ;
  assign n11927 = n11898 & n11926 ;
  assign n11928 = ~n11915 & n11927 ;
  assign n11929 = ~n11899 & ~n11928 ;
  assign n11930 = ~\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  & ~n11668 ;
  assign n11931 = ~n11784 & n11930 ;
  assign n11932 = n11878 & ~n11931 ;
  assign n11933 = n11929 & n11932 ;
  assign n11934 = ~n11879 & ~n11933 ;
  assign n11935 = \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
  assign n11936 = ~n11722 & n11935 ;
  assign n11937 = \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
  assign n11938 = n11722 & n11937 ;
  assign n11939 = ~n11936 & ~n11938 ;
  assign n11940 = \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n11941 = ~n11715 & n11940 ;
  assign n11942 = \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n11943 = n11715 & n11942 ;
  assign n11944 = ~n11941 & ~n11943 ;
  assign n11945 = n11939 & n11944 ;
  assign n11946 = n11864 & n11945 ;
  assign n11947 = n11934 & n11946 ;
  assign n11948 = ~n11865 & ~n11947 ;
  assign n11949 = ~\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  & ~n11674 ;
  assign n11950 = ~n11807 & n11949 ;
  assign n11951 = ~\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & ~n11693 ;
  assign n11952 = ~n11691 & n11951 ;
  assign n11953 = ~n11950 & ~n11952 ;
  assign n11954 = n11844 & n11953 ;
  assign n11955 = n11948 & n11954 ;
  assign n11956 = ~n11845 & ~n11955 ;
  assign n11957 = \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n11958 = ~\macstatus1_LatchedCrcError_reg/NET0131  & \macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n11959 = n11957 & n11958 ;
  assign n11960 = n11956 & n11959 ;
  assign n11961 = ~n11818 & n11960 ;
  assign n11962 = ~n11662 & ~n11961 ;
  assign n11963 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131  ;
  assign n11964 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  ;
  assign n11965 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  ;
  assign n11966 = n11964 & n11965 ;
  assign n11967 = n11963 & n11966 ;
  assign n11968 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  ;
  assign n11969 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131  ;
  assign n11970 = n11968 & n11969 ;
  assign n11971 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131  ;
  assign n11972 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131  ;
  assign n11973 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  ;
  assign n11974 = n11972 & n11973 ;
  assign n11975 = n11971 & n11974 ;
  assign n11976 = n11970 & n11975 ;
  assign n11977 = n11967 & n11976 ;
  assign n11978 = \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  & \maccontrol1_receivecontrol1_Divider2_reg/NET0131  ;
  assign n11979 = \maccontrol1_receivecontrol1_Pause_reg/NET0131  & \maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131  ;
  assign n11980 = n11978 & n11979 ;
  assign n11981 = \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  & \maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131  ;
  assign n11982 = \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131  & n11981 ;
  assign n11983 = n11980 & n11982 ;
  assign n11984 = \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  & \maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131  ;
  assign n11985 = n11983 & n11984 ;
  assign n11986 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131  ;
  assign n11987 = n11985 & n11986 ;
  assign n11988 = ~n11977 & n11987 ;
  assign n11989 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  & n11988 ;
  assign n11990 = \maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  & ~n11989 ;
  assign n11991 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  ;
  assign n11992 = n11988 & n11991 ;
  assign n11993 = ~n11990 & ~n11992 ;
  assign n11994 = ~n11961 & n11993 ;
  assign n11995 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131  & n11959 ;
  assign n11996 = n11956 & n11995 ;
  assign n11997 = ~n11818 & n11996 ;
  assign n11998 = ~n11994 & ~n11997 ;
  assign n11999 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  & n11985 ;
  assign n12000 = ~n11977 & n11999 ;
  assign n12001 = \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  & ~n11985 ;
  assign n12002 = \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  & n11967 ;
  assign n12003 = n11976 & n12002 ;
  assign n12004 = ~n12001 & ~n12003 ;
  assign n12005 = ~n12000 & n12004 ;
  assign n12006 = ~n11961 & n12005 ;
  assign n12007 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131  & n11959 ;
  assign n12008 = n11956 & n12007 ;
  assign n12009 = ~n11818 & n12008 ;
  assign n12010 = ~n12006 & ~n12009 ;
  assign n12011 = n11971 & n11991 ;
  assign n12012 = n11988 & n12011 ;
  assign n12013 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131  ;
  assign n12014 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  & n12013 ;
  assign n12015 = n12012 & n12014 ;
  assign n12016 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  & n12015 ;
  assign n12017 = \maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131  & ~n12016 ;
  assign n12018 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  ;
  assign n12019 = n12015 & n12018 ;
  assign n12020 = ~n12017 & ~n12019 ;
  assign n12021 = ~n11961 & n12020 ;
  assign n12022 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131  & n11959 ;
  assign n12023 = n11956 & n12022 ;
  assign n12024 = ~n11818 & n12023 ;
  assign n12025 = ~n12021 & ~n12024 ;
  assign n12026 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  ;
  assign n12027 = n11963 & n12026 ;
  assign n12028 = n12015 & n12027 ;
  assign n12029 = \maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  & ~n12028 ;
  assign n12030 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  & n12028 ;
  assign n12031 = ~n12029 & ~n12030 ;
  assign n12032 = ~n11961 & n12031 ;
  assign n12033 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131  & n11959 ;
  assign n12034 = n11956 & n12033 ;
  assign n12035 = ~n11818 & n12034 ;
  assign n12036 = ~n12032 & ~n12035 ;
  assign n12037 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  & n11963 ;
  assign n12038 = n12015 & n12037 ;
  assign n12039 = \maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131  & ~n12019 ;
  assign n12040 = ~n12038 & ~n12039 ;
  assign n12041 = ~n11961 & n12040 ;
  assign n12042 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131  & n11959 ;
  assign n12043 = n11956 & n12042 ;
  assign n12044 = ~n11818 & n12043 ;
  assign n12045 = ~n12041 & ~n12044 ;
  assign n12046 = \maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131  & ~n12000 ;
  assign n12047 = ~n11988 & ~n12046 ;
  assign n12048 = ~n11961 & n12047 ;
  assign n12049 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131  & n11959 ;
  assign n12050 = n11956 & n12049 ;
  assign n12051 = ~n11818 & n12050 ;
  assign n12052 = ~n12048 & ~n12051 ;
  assign n12053 = n11967 & n12015 ;
  assign n12054 = \maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131  & ~n12053 ;
  assign n12055 = ~n11961 & n12054 ;
  assign n12056 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131  & n11959 ;
  assign n12057 = n11956 & n12056 ;
  assign n12058 = ~n11818 & n12057 ;
  assign n12059 = ~n12055 & ~n12058 ;
  assign n12060 = \maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  & ~n11988 ;
  assign n12061 = ~n11989 & ~n12060 ;
  assign n12062 = ~n11961 & n12061 ;
  assign n12063 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131  & n11959 ;
  assign n12064 = n11956 & n12063 ;
  assign n12065 = ~n11818 & n12064 ;
  assign n12066 = ~n12062 & ~n12065 ;
  assign n12067 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  ;
  assign n12068 = n12012 & n12067 ;
  assign n12069 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  & n12012 ;
  assign n12070 = \maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  & ~n12069 ;
  assign n12071 = ~n12068 & ~n12070 ;
  assign n12072 = ~n11961 & n12071 ;
  assign n12073 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131  & n11959 ;
  assign n12074 = n11956 & n12073 ;
  assign n12075 = ~n11818 & n12074 ;
  assign n12076 = ~n12072 & ~n12075 ;
  assign n12077 = \maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  & ~n12015 ;
  assign n12078 = ~n12016 & ~n12077 ;
  assign n12079 = ~n11961 & n12078 ;
  assign n12080 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131  & n11959 ;
  assign n12081 = n11956 & n12080 ;
  assign n12082 = ~n11818 & n12081 ;
  assign n12083 = ~n12079 & ~n12082 ;
  assign n12084 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131  ;
  assign n12085 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  & n12084 ;
  assign n12086 = n11988 & n12085 ;
  assign n12087 = \maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131  & ~n11992 ;
  assign n12088 = ~n12086 & ~n12087 ;
  assign n12089 = ~n11961 & n12088 ;
  assign n12090 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131  & n11959 ;
  assign n12091 = n11956 & n12090 ;
  assign n12092 = ~n11818 & n12091 ;
  assign n12093 = ~n12089 & ~n12092 ;
  assign n12094 = \maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131  & ~n12086 ;
  assign n12095 = ~n12012 & ~n12094 ;
  assign n12096 = ~n11961 & n12095 ;
  assign n12097 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131  & n11959 ;
  assign n12098 = n11956 & n12097 ;
  assign n12099 = ~n11818 & n12098 ;
  assign n12100 = ~n12096 & ~n12099 ;
  assign n12101 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131  & ~n12030 ;
  assign n12102 = ~\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  & \maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131  ;
  assign n12103 = n12028 & n12102 ;
  assign n12104 = ~n12101 & ~n12103 ;
  assign n12105 = ~n11961 & ~n12104 ;
  assign n12106 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131  & n11959 ;
  assign n12107 = n11956 & n12106 ;
  assign n12108 = ~n11818 & n12107 ;
  assign n12109 = ~n12105 & ~n12108 ;
  assign n12110 = \maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131  & ~n12068 ;
  assign n12111 = ~n12015 & ~n12110 ;
  assign n12112 = ~n11961 & n12111 ;
  assign n12113 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131  & n11959 ;
  assign n12114 = n11956 & n12113 ;
  assign n12115 = ~n11818 & n12114 ;
  assign n12116 = ~n12112 & ~n12115 ;
  assign n12117 = \maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131  & ~n12038 ;
  assign n12118 = ~n12028 & ~n12117 ;
  assign n12119 = ~n11961 & n12118 ;
  assign n12120 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131  & n11959 ;
  assign n12121 = n11956 & n12120 ;
  assign n12122 = ~n11818 & n12121 ;
  assign n12123 = ~n12119 & ~n12122 ;
  assign n12124 = \maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  & ~n12012 ;
  assign n12125 = ~n12069 & ~n12124 ;
  assign n12126 = ~n11961 & n12125 ;
  assign n12127 = ~\maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131  & n11959 ;
  assign n12128 = n11956 & n12127 ;
  assign n12129 = ~n11818 & n12128 ;
  assign n12130 = ~n12126 & ~n12129 ;
  assign n12131 = n10674 & n11527 ;
  assign n12132 = ~n10674 & ~n11527 ;
  assign n12133 = ~n12131 & ~n12132 ;
  assign n12134 = n10660 & n12133 ;
  assign n12135 = ~n10660 & ~n12133 ;
  assign n12136 = ~n12134 & ~n12135 ;
  assign n12137 = n11353 & n12136 ;
  assign n12138 = ~\rxethmac1_crcrx_Crc_reg[9]/NET0131  & n10663 ;
  assign n12139 = ~n12137 & n12138 ;
  assign n12140 = \rxethmac1_crcrx_Crc_reg[9]/NET0131  & n10663 ;
  assign n12141 = n12137 & n12140 ;
  assign n12142 = ~n12139 & ~n12141 ;
  assign n12143 = \txethmac1_txcrc_Crc_reg[14]/NET0131  & n11507 ;
  assign n12144 = ~\txethmac1_txcrc_Crc_reg[14]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n12145 = ~\txethmac1_txcrc_Crc_reg[30]/NET0131  & n12144 ;
  assign n12146 = ~n11502 & n12145 ;
  assign n12147 = \txethmac1_txcrc_Crc_reg[30]/NET0131  & n12144 ;
  assign n12148 = n11502 & n12147 ;
  assign n12149 = ~n12146 & ~n12148 ;
  assign n12150 = n11464 & n12149 ;
  assign n12151 = ~n12143 & n12150 ;
  assign n12152 = \txethmac1_txcrc_Crc_reg[15]/NET0131  & n11541 ;
  assign n12153 = ~\txethmac1_txcrc_Crc_reg[15]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n12154 = ~\txethmac1_txcrc_Crc_reg[31]/NET0131  & n12153 ;
  assign n12155 = ~n11455 & n12154 ;
  assign n12156 = \txethmac1_txcrc_Crc_reg[31]/NET0131  & n12153 ;
  assign n12157 = n11455 & n12156 ;
  assign n12158 = ~n12155 & ~n12157 ;
  assign n12159 = n11464 & n12158 ;
  assign n12160 = ~n12152 & n12159 ;
  assign n12161 = ~\txethmac1_txcrc_Crc_reg[16]/NET0131  & n11298 ;
  assign n12162 = n11297 & n12161 ;
  assign n12163 = \rxethmac1_rxstatem1_StateData1_reg/NET0131  & ~n10650 ;
  assign n12164 = ~n10652 & n12163 ;
  assign n12165 = \rxethmac1_rxstatem1_StateData0_reg/NET0131  & n10653 ;
  assign n12166 = \rxethmac1_rxstatem1_StateData0_reg/NET0131  & n10605 ;
  assign n12167 = n10647 & n12166 ;
  assign n12168 = ~n12165 & ~n12167 ;
  assign n12169 = ~n12164 & n12168 ;
  assign n12170 = n11956 & ~n12169 ;
  assign n12171 = ~\macstatus1_ShortFrame_reg/NET0131  & ~n12164 ;
  assign n12172 = n12168 & n12171 ;
  assign n12173 = ~\macstatus1_LoadRxStatus_reg/NET0131  & ~n12172 ;
  assign n12174 = ~n12170 & n12173 ;
  assign n12175 = ~n11359 & n11372 ;
  assign n12176 = n11359 & ~n11372 ;
  assign n12177 = ~n12175 & ~n12176 ;
  assign n12178 = n11353 & n12177 ;
  assign n12179 = ~\rxethmac1_crcrx_Crc_reg[8]/NET0131  & n10663 ;
  assign n12180 = ~n12178 & n12179 ;
  assign n12181 = \rxethmac1_crcrx_Crc_reg[8]/NET0131  & n10663 ;
  assign n12182 = n12178 & n12181 ;
  assign n12183 = ~n12180 & ~n12182 ;
  assign n12184 = ~\rxethmac1_crcrx_Crc_reg[14]/NET0131  & n10663 ;
  assign n12185 = ~n10676 & n12184 ;
  assign n12186 = \rxethmac1_crcrx_Crc_reg[14]/NET0131  & n10663 ;
  assign n12187 = n10676 & n12186 ;
  assign n12188 = ~n12185 & ~n12187 ;
  assign n12189 = ~\txethmac1_txcrc_Crc_reg[17]/NET0131  & n11298 ;
  assign n12190 = n11297 & n12189 ;
  assign n12191 = \macstatus1_ReceivedPacketTooBig_reg/NET0131  & ~n12164 ;
  assign n12192 = n12168 & n12191 ;
  assign n12193 = ~\ethreg1_MODER_1_DataOut_reg[6]/NET0131  & ~n12169 ;
  assign n12194 = n11679 & n12193 ;
  assign n12195 = n11817 & n12194 ;
  assign n12196 = ~n12192 & ~n12195 ;
  assign n12197 = ~\macstatus1_LoadRxStatus_reg/NET0131  & ~n12196 ;
  assign n12198 = \txethmac1_txcrc_Crc_reg[12]/NET0131  & n11588 ;
  assign n12199 = ~\txethmac1_txcrc_Crc_reg[12]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n12200 = ~\txethmac1_txcrc_Crc_reg[28]/NET0131  & n12199 ;
  assign n12201 = ~n11443 & n12200 ;
  assign n12202 = \txethmac1_txcrc_Crc_reg[28]/NET0131  & n12199 ;
  assign n12203 = n11443 & n12202 ;
  assign n12204 = ~n12201 & ~n12203 ;
  assign n12205 = n11464 & n12204 ;
  assign n12206 = ~n12198 & n12205 ;
  assign n12207 = ~n10657 & n11524 ;
  assign n12208 = n10657 & ~n11524 ;
  assign n12209 = ~n12207 & ~n12208 ;
  assign n12210 = \rxethmac1_crcrx_Crc_reg[29]/NET0131  & ~\rxethmac1_crcrx_Crc_reg[31]/NET0131  ;
  assign n12211 = ~n10545 & ~n12210 ;
  assign n12212 = n11359 & ~n12211 ;
  assign n12213 = ~n11359 & n12211 ;
  assign n12214 = ~n12212 & ~n12213 ;
  assign n12215 = n12209 & ~n12214 ;
  assign n12216 = ~n12209 & n12214 ;
  assign n12217 = ~n12215 & ~n12216 ;
  assign n12218 = n11353 & n12217 ;
  assign n12219 = ~\rxethmac1_crcrx_Crc_reg[7]/NET0131  & n10663 ;
  assign n12220 = ~n12218 & n12219 ;
  assign n12221 = \rxethmac1_crcrx_Crc_reg[7]/NET0131  & n10663 ;
  assign n12222 = n12218 & n12221 ;
  assign n12223 = ~n12220 & ~n12222 ;
  assign n12224 = \txethmac1_txcrc_Crc_reg[13]/NET0131  & n11483 ;
  assign n12225 = ~\txethmac1_txcrc_Crc_reg[13]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n12226 = ~\txethmac1_txcrc_Crc_reg[29]/NET0131  & n12225 ;
  assign n12227 = ~n11478 & n12226 ;
  assign n12228 = \txethmac1_txcrc_Crc_reg[29]/NET0131  & n12225 ;
  assign n12229 = n11478 & n12228 ;
  assign n12230 = ~n12227 & ~n12229 ;
  assign n12231 = n11464 & n12230 ;
  assign n12232 = ~n12224 & n12231 ;
  assign n12233 = ~\rxethmac1_crcrx_Crc_reg[5]/NET0131  & ~n11372 ;
  assign n12234 = n11353 & n12233 ;
  assign n12235 = ~\rxethmac1_crcrx_Crc_reg[5]/NET0131  & n10663 ;
  assign n12236 = ~n11377 & ~n12235 ;
  assign n12237 = ~n12234 & ~n12236 ;
  assign n12238 = ~\txethmac1_txcrc_Crc_reg[10]/NET0131  & ~n11648 ;
  assign n12239 = n11647 & n12238 ;
  assign n12240 = ~\txethmac1_txcrc_Crc_reg[10]/NET0131  & n11464 ;
  assign n12241 = n11647 & n11652 ;
  assign n12242 = ~n12240 & ~n12241 ;
  assign n12243 = ~n12239 & ~n12242 ;
  assign n12244 = \txethmac1_txcrc_Crc_reg[11]/NET0131  & n11541 ;
  assign n12245 = ~\txethmac1_txcrc_Crc_reg[11]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n12246 = ~\txethmac1_txcrc_Crc_reg[31]/NET0131  & n12245 ;
  assign n12247 = ~n11455 & n12246 ;
  assign n12248 = \txethmac1_txcrc_Crc_reg[31]/NET0131  & n12245 ;
  assign n12249 = n11455 & n12248 ;
  assign n12250 = ~n12247 & ~n12249 ;
  assign n12251 = n11464 & n12250 ;
  assign n12252 = ~n12244 & n12251 ;
  assign n12253 = ~\rxethmac1_crcrx_Crc_reg[10]/NET0131  & n12133 ;
  assign n12254 = n11353 & n12253 ;
  assign n12255 = ~\rxethmac1_crcrx_Crc_reg[10]/NET0131  & n10663 ;
  assign n12256 = n10663 & n12133 ;
  assign n12257 = n11353 & n12256 ;
  assign n12258 = ~n12255 & ~n12257 ;
  assign n12259 = ~n12254 & ~n12258 ;
  assign n12260 = ~\rxethmac1_crcrx_Crc_reg[4]/NET0131  & n10663 ;
  assign n12261 = ~n12218 & n12260 ;
  assign n12262 = \rxethmac1_crcrx_Crc_reg[4]/NET0131  & n10663 ;
  assign n12263 = n12218 & n12262 ;
  assign n12264 = ~n12261 & ~n12263 ;
  assign n12265 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  & ~\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n12266 = \maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131  & \rxethmac1_RxValid_reg/NET0131  ;
  assign n12267 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  & n12266 ;
  assign n12268 = n12265 & n12267 ;
  assign n12269 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & ~\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  ;
  assign n12270 = ~\rxethmac1_RxData_reg[4]/NET0131  & ~\rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12271 = ~\rxethmac1_RxData_reg[6]/NET0131  & n12270 ;
  assign n12272 = ~\rxethmac1_RxData_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12273 = ~\rxethmac1_RxData_reg[7]/NET0131  & n12272 ;
  assign n12274 = n12271 & n12273 ;
  assign n12275 = \rxethmac1_RxData_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12276 = n12274 & n12275 ;
  assign n12277 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  & \rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12278 = \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12279 = ~n12277 & ~n12278 ;
  assign n12280 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  & \rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12281 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  & \rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12282 = ~n12280 & ~n12281 ;
  assign n12283 = n12279 & n12282 ;
  assign n12284 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12285 = \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  & \rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12286 = ~n12284 & ~n12285 ;
  assign n12287 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  & ~\rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12288 = \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12289 = ~n12287 & ~n12288 ;
  assign n12290 = ~n12286 & ~n12289 ;
  assign n12291 = n12283 & n12290 ;
  assign n12292 = \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  & ~\rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12293 = \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  & ~\rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12294 = ~n12292 & ~n12293 ;
  assign n12295 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  & \rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12296 = \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12297 = ~n12295 & ~n12296 ;
  assign n12298 = n12294 & n12297 ;
  assign n12299 = \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  & ~\rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12300 = \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12301 = ~n12299 & ~n12300 ;
  assign n12302 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  & \rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12303 = ~\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  & \rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12304 = ~n12302 & ~n12303 ;
  assign n12305 = n12301 & n12304 ;
  assign n12306 = n12298 & n12305 ;
  assign n12307 = n12291 & n12306 ;
  assign n12308 = ~n12276 & ~n12307 ;
  assign n12309 = n12269 & ~n12308 ;
  assign n12310 = ~\rxethmac1_RxData_reg[6]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12311 = n12270 & n12310 ;
  assign n12312 = ~\rxethmac1_RxData_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12313 = n12272 & n12312 ;
  assign n12314 = n12311 & n12313 ;
  assign n12315 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  & \rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12316 = \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  & ~\rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12317 = ~n12315 & ~n12316 ;
  assign n12318 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  & \rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12319 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  & \rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12320 = ~n12318 & ~n12319 ;
  assign n12321 = n12317 & n12320 ;
  assign n12322 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12323 = \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  & \rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12324 = ~n12322 & ~n12323 ;
  assign n12325 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12326 = \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  & \rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12327 = ~n12325 & ~n12326 ;
  assign n12328 = ~n12324 & ~n12327 ;
  assign n12329 = n12321 & n12328 ;
  assign n12330 = \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12331 = \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12332 = ~n12330 & ~n12331 ;
  assign n12333 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  & \rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12334 = \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  & ~\rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12335 = ~n12333 & ~n12334 ;
  assign n12336 = n12332 & n12335 ;
  assign n12337 = \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  & ~\rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12338 = \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  & ~\rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12339 = ~n12337 & ~n12338 ;
  assign n12340 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12341 = ~\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  & \rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12342 = ~n12340 & ~n12341 ;
  assign n12343 = n12339 & n12342 ;
  assign n12344 = n12336 & n12343 ;
  assign n12345 = n12329 & n12344 ;
  assign n12346 = ~n12314 & ~n12345 ;
  assign n12347 = \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & ~\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  ;
  assign n12348 = \maccontrol1_receivecontrol1_AddressOK_reg/NET0131  & n12347 ;
  assign n12349 = ~n12346 & n12348 ;
  assign n12350 = ~n12309 & ~n12349 ;
  assign n12351 = n12268 & ~n12350 ;
  assign n12352 = ~\maccontrol1_receivecontrol1_AddressOK_reg/NET0131  & ~n12351 ;
  assign n12353 = \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  & ~\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  ;
  assign n12354 = n12266 & n12353 ;
  assign n12355 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  & ~\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n12356 = n12354 & n12355 ;
  assign n12357 = ~\macstatus1_ReceiveEnd_reg/NET0131  & ~n12356 ;
  assign n12358 = ~n12268 & n12357 ;
  assign n12359 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  & \rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12360 = \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12361 = ~n12359 & ~n12360 ;
  assign n12362 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  & \rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12363 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  & \rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12364 = ~n12362 & ~n12363 ;
  assign n12365 = n12361 & n12364 ;
  assign n12366 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  & ~\rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12367 = \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  & \rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12368 = ~n12366 & ~n12367 ;
  assign n12369 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  & ~\rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12370 = \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12371 = ~n12369 & ~n12370 ;
  assign n12372 = ~n12368 & ~n12371 ;
  assign n12373 = n12365 & n12372 ;
  assign n12374 = \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12375 = \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  & ~\rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12376 = ~n12374 & ~n12375 ;
  assign n12377 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  & \rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12378 = \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12379 = ~n12377 & ~n12378 ;
  assign n12380 = n12376 & n12379 ;
  assign n12381 = \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  & ~\rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12382 = \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12383 = ~n12381 & ~n12382 ;
  assign n12384 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  & \rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12385 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  & \rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12386 = ~n12384 & ~n12385 ;
  assign n12387 = n12383 & n12386 ;
  assign n12388 = n12380 & n12387 ;
  assign n12389 = n12373 & n12388 ;
  assign n12390 = ~n12276 & ~n12389 ;
  assign n12391 = n12347 & ~n12390 ;
  assign n12392 = n12274 & n12312 ;
  assign n12393 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  & \rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12394 = \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12395 = ~n12393 & ~n12394 ;
  assign n12396 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  & \rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12397 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  & \rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12398 = ~n12396 & ~n12397 ;
  assign n12399 = n12395 & n12398 ;
  assign n12400 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12401 = \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  & \rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12402 = ~n12400 & ~n12401 ;
  assign n12403 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  & ~\rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12404 = \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  & \rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12405 = ~n12403 & ~n12404 ;
  assign n12406 = ~n12402 & ~n12405 ;
  assign n12407 = n12399 & n12406 ;
  assign n12408 = \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  & ~\rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12409 = \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  & ~\rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12410 = ~n12408 & ~n12409 ;
  assign n12411 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  & \rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12412 = \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12413 = ~n12411 & ~n12412 ;
  assign n12414 = n12410 & n12413 ;
  assign n12415 = \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12416 = \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  & ~\rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12417 = ~n12415 & ~n12416 ;
  assign n12418 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  & \rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12419 = ~\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12420 = ~n12418 & ~n12419 ;
  assign n12421 = n12417 & n12420 ;
  assign n12422 = n12414 & n12421 ;
  assign n12423 = n12407 & n12422 ;
  assign n12424 = ~n12392 & ~n12423 ;
  assign n12425 = n12269 & ~n12424 ;
  assign n12426 = ~n12391 & ~n12425 ;
  assign n12427 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  & n12354 ;
  assign n12428 = ~n12268 & n12427 ;
  assign n12429 = ~n12426 & n12428 ;
  assign n12430 = ~n12358 & ~n12429 ;
  assign n12431 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  & \rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12432 = \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12433 = ~n12431 & ~n12432 ;
  assign n12434 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  & \rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12435 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  & \rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12436 = ~n12434 & ~n12435 ;
  assign n12437 = n12433 & n12436 ;
  assign n12438 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  & ~\rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12439 = \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  & \rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12440 = ~n12438 & ~n12439 ;
  assign n12441 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12442 = \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  & \rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12443 = ~n12441 & ~n12442 ;
  assign n12444 = ~n12440 & ~n12443 ;
  assign n12445 = n12437 & n12444 ;
  assign n12446 = \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  & ~\rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12447 = \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12448 = ~n12446 & ~n12447 ;
  assign n12449 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  & \rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12450 = \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  & ~\rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12451 = ~n12449 & ~n12450 ;
  assign n12452 = n12448 & n12451 ;
  assign n12453 = \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12454 = \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  & ~\rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12455 = ~n12453 & ~n12454 ;
  assign n12456 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12457 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  & \rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12458 = ~n12456 & ~n12457 ;
  assign n12459 = n12455 & n12458 ;
  assign n12460 = n12452 & n12459 ;
  assign n12461 = n12445 & n12460 ;
  assign n12462 = \rxethmac1_RxData_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12463 = \rxethmac1_RxData_reg[6]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12464 = n12462 & n12463 ;
  assign n12465 = n12270 & n12312 ;
  assign n12466 = n12464 & n12465 ;
  assign n12467 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & ~n12466 ;
  assign n12468 = ~n12461 & n12467 ;
  assign n12469 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  & \rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12470 = \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  & ~\rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12471 = ~n12469 & ~n12470 ;
  assign n12472 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  & \rxethmac1_RxData_reg[7]/NET0131  ;
  assign n12473 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  & \rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12474 = ~n12472 & ~n12473 ;
  assign n12475 = n12471 & n12474 ;
  assign n12476 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  & ~\rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12477 = \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  & \rxethmac1_RxData_reg[1]/NET0131  ;
  assign n12478 = ~n12476 & ~n12477 ;
  assign n12479 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  & ~\rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12480 = \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  & \rxethmac1_RxData_reg[4]/NET0131  ;
  assign n12481 = ~n12479 & ~n12480 ;
  assign n12482 = ~n12478 & ~n12481 ;
  assign n12483 = n12475 & n12482 ;
  assign n12484 = \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  & ~\rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12485 = \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  & ~\rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12486 = ~n12484 & ~n12485 ;
  assign n12487 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  & \rxethmac1_RxData_reg[5]/NET0131  ;
  assign n12488 = \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  & ~\rxethmac1_RxData_reg[0]/NET0131  ;
  assign n12489 = ~n12487 & ~n12488 ;
  assign n12490 = n12486 & n12489 ;
  assign n12491 = \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  & ~\rxethmac1_RxData_reg[2]/NET0131  ;
  assign n12492 = \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  & ~\rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12493 = ~n12491 & ~n12492 ;
  assign n12494 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  & \rxethmac1_RxData_reg[6]/NET0131  ;
  assign n12495 = ~\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  & \rxethmac1_RxData_reg[3]/NET0131  ;
  assign n12496 = ~n12494 & ~n12495 ;
  assign n12497 = n12493 & n12496 ;
  assign n12498 = n12490 & n12497 ;
  assign n12499 = n12483 & n12498 ;
  assign n12500 = \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & ~n12392 ;
  assign n12501 = ~n12499 & n12500 ;
  assign n12502 = \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  & n12265 ;
  assign n12503 = n12267 & n12502 ;
  assign n12504 = ~n12501 & n12503 ;
  assign n12505 = ~n12468 & n12504 ;
  assign n12506 = ~n12351 & ~n12505 ;
  assign n12507 = n12430 & n12506 ;
  assign n12508 = ~n12352 & ~n12507 ;
  assign n12509 = ~\rxethmac1_crcrx_Crc_reg[25]/NET0131  & n10663 ;
  assign n12510 = ~n11576 & n12509 ;
  assign n12511 = \rxethmac1_crcrx_Crc_reg[25]/NET0131  & n10663 ;
  assign n12512 = n11576 & n12511 ;
  assign n12513 = ~n12510 & ~n12512 ;
  assign n12514 = \WillTransmit_q2_reg/P0001  & ~\ethreg1_MODER_1_DataOut_reg[2]/NET0131  ;
  assign n12515 = \rxethmac1_rxstatem1_StateIdle_reg/NET0131  & n12514 ;
  assign n12516 = ~n10657 & n10671 ;
  assign n12517 = ~n11524 & n12516 ;
  assign n12518 = \rxethmac1_rxstatem1_StateSFD_reg/NET0131  & ~n11356 ;
  assign n12519 = n12517 & n12518 ;
  assign n12520 = ~\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  ;
  assign n12521 = ~\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  & \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131  ;
  assign n12522 = \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131  & n12521 ;
  assign n12523 = n12520 & n12522 ;
  assign n12524 = ~\ethreg1_MODER_0_DataOut_reg[6]/NET0131  & ~n12523 ;
  assign n12525 = n12519 & n12524 ;
  assign n12526 = ~n12515 & ~n12525 ;
  assign n12527 = ~n12167 & n12526 ;
  assign n12528 = ~n10653 & ~n12527 ;
  assign n12529 = \rxethmac1_rxstatem1_StateData1_reg/NET0131  & ~n10653 ;
  assign n12530 = ~n10653 & ~n12524 ;
  assign n12531 = n12519 & n12530 ;
  assign n12532 = ~n12529 & ~n12531 ;
  assign n12533 = ~\rxethmac1_rxstatem1_StateDrop_reg/NET0131  & ~\rxethmac1_rxstatem1_StatePreamble_reg/NET0131  ;
  assign n12534 = ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  & n12533 ;
  assign n12535 = n10649 & n12534 ;
  assign n12536 = n10653 & ~n12535 ;
  assign n12537 = n12532 & ~n12536 ;
  assign n12538 = n11356 & ~n11524 ;
  assign n12539 = n12516 & n12538 ;
  assign n12540 = \rxethmac1_rxstatem1_StateIdle_reg/NET0131  & ~n12514 ;
  assign n12541 = ~n10653 & n12540 ;
  assign n12542 = ~n12539 & n12541 ;
  assign n12543 = ~\rxethmac1_rxstatem1_StatePreamble_reg/NET0131  & ~n12540 ;
  assign n12544 = ~n10653 & ~n12543 ;
  assign n12545 = n12539 & n12544 ;
  assign n12546 = ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  & ~n12545 ;
  assign n12547 = ~n12542 & ~n12546 ;
  assign n12548 = n12537 & n12547 ;
  assign n12549 = ~n12528 & n12548 ;
  assign n12550 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & ~n11446 ;
  assign n12551 = ~n11626 & n12550 ;
  assign n12552 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n11446 ;
  assign n12553 = n11626 & n12552 ;
  assign n12554 = ~n12551 & ~n12553 ;
  assign n12555 = \txethmac1_txcrc_Crc_reg[8]/NET0131  & n12554 ;
  assign n12556 = ~\txethmac1_txcrc_Crc_reg[8]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n12557 = ~n11446 & n12556 ;
  assign n12558 = ~n11626 & n12557 ;
  assign n12559 = n11446 & n12556 ;
  assign n12560 = n11626 & n12559 ;
  assign n12561 = ~n12558 & ~n12560 ;
  assign n12562 = n11464 & n12561 ;
  assign n12563 = ~n12555 & n12562 ;
  assign n12564 = ~n11359 & ~n12133 ;
  assign n12565 = n11359 & n12133 ;
  assign n12566 = ~n12564 & ~n12565 ;
  assign n12567 = n11353 & n12566 ;
  assign n12568 = ~\rxethmac1_crcrx_Crc_reg[3]/NET0131  & n10663 ;
  assign n12569 = ~n12567 & n12568 ;
  assign n12570 = \rxethmac1_crcrx_Crc_reg[3]/NET0131  & n10663 ;
  assign n12571 = n12567 & n12570 ;
  assign n12572 = ~n12569 & ~n12571 ;
  assign n12573 = ~\rxethmac1_rxstatem1_StatePreamble_reg/NET0131  & ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n12574 = ~n12540 & n12573 ;
  assign n12575 = \rxethmac1_rxstatem1_StateData1_reg/NET0131  & ~n10581 ;
  assign n12576 = n12574 & ~n12575 ;
  assign n12577 = \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  & n11663 ;
  assign n12578 = \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  & n11733 ;
  assign n12579 = n12577 & n12578 ;
  assign n12580 = \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n12581 = \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  & n12580 ;
  assign n12582 = n12579 & n12581 ;
  assign n12583 = \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  & n11692 ;
  assign n12584 = \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n12585 = \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n12586 = n12584 & n12585 ;
  assign n12587 = n12583 & n12586 ;
  assign n12588 = n12574 & n12587 ;
  assign n12589 = n12582 & n12588 ;
  assign n12590 = ~n12576 & ~n12589 ;
  assign n12591 = ~n10653 & ~n12519 ;
  assign n12592 = n12590 & n12591 ;
  assign n12593 = ~n12167 & n12592 ;
  assign n12594 = \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  & n12593 ;
  assign n12595 = ~n12167 & ~n12519 ;
  assign n12596 = ~n10653 & ~n12595 ;
  assign n12597 = ~\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  & ~n12593 ;
  assign n12598 = ~n12596 & ~n12597 ;
  assign n12599 = ~n12594 & n12598 ;
  assign n12600 = \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  & n12580 ;
  assign n12601 = n12579 & n12600 ;
  assign n12602 = n12593 & n12601 ;
  assign n12603 = \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  & n12602 ;
  assign n12604 = ~\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  & ~n12603 ;
  assign n12605 = \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  & n12584 ;
  assign n12606 = n12580 & n12605 ;
  assign n12607 = n12579 & n12606 ;
  assign n12608 = n12593 & n12607 ;
  assign n12609 = ~n12596 & ~n12608 ;
  assign n12610 = ~n12604 & n12609 ;
  assign n12611 = \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  & n12608 ;
  assign n12612 = ~\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  & ~n12608 ;
  assign n12613 = ~n12596 & ~n12612 ;
  assign n12614 = ~n12611 & n12613 ;
  assign n12615 = n11692 & n12608 ;
  assign n12616 = ~\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  & ~n12615 ;
  assign n12617 = n12583 & n12608 ;
  assign n12618 = ~n12596 & ~n12617 ;
  assign n12619 = ~n12616 & n12618 ;
  assign n12620 = ~\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  & ~n12611 ;
  assign n12621 = ~n12596 & ~n12615 ;
  assign n12622 = ~n12620 & n12621 ;
  assign n12623 = ~\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  & ~n12617 ;
  assign n12624 = n12579 & n12580 ;
  assign n12625 = n12587 & n12624 ;
  assign n12626 = n12593 & n12625 ;
  assign n12627 = ~n12596 & ~n12626 ;
  assign n12628 = ~n12623 & n12627 ;
  assign n12629 = \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  & n12626 ;
  assign n12630 = ~\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  & ~n12626 ;
  assign n12631 = ~n12596 & ~n12630 ;
  assign n12632 = ~n12629 & n12631 ;
  assign n12633 = ~\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  & ~n12594 ;
  assign n12634 = n12580 & n12593 ;
  assign n12635 = ~n12596 & ~n12634 ;
  assign n12636 = ~n12633 & n12635 ;
  assign n12637 = ~\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  & ~n12634 ;
  assign n12638 = \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  & n12580 ;
  assign n12639 = n12593 & n12638 ;
  assign n12640 = ~n12596 & ~n12639 ;
  assign n12641 = ~n12637 & n12640 ;
  assign n12642 = ~\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  & ~n12639 ;
  assign n12643 = \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  & n12638 ;
  assign n12644 = n12593 & n12643 ;
  assign n12645 = ~n12596 & ~n12644 ;
  assign n12646 = ~n12642 & n12645 ;
  assign n12647 = ~\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  & ~n12644 ;
  assign n12648 = n12577 & n12580 ;
  assign n12649 = n12593 & n12648 ;
  assign n12650 = ~n12596 & ~n12649 ;
  assign n12651 = ~n12647 & n12650 ;
  assign n12652 = ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  & ~n12649 ;
  assign n12653 = \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  & n12580 ;
  assign n12654 = n12577 & n12653 ;
  assign n12655 = n12593 & n12654 ;
  assign n12656 = ~n12596 & ~n12655 ;
  assign n12657 = ~n12652 & n12656 ;
  assign n12658 = \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  & n12655 ;
  assign n12659 = ~\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  & ~n12655 ;
  assign n12660 = ~n12596 & ~n12659 ;
  assign n12661 = ~n12658 & n12660 ;
  assign n12662 = ~\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  & ~n12658 ;
  assign n12663 = n12593 & n12624 ;
  assign n12664 = ~n12596 & ~n12663 ;
  assign n12665 = ~n12662 & n12664 ;
  assign n12666 = ~\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  & ~n12663 ;
  assign n12667 = ~n12596 & ~n12602 ;
  assign n12668 = ~n12666 & n12667 ;
  assign n12669 = ~\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  & ~n12602 ;
  assign n12670 = ~n12596 & ~n12603 ;
  assign n12671 = ~n12669 & n12670 ;
  assign n12672 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n11458 ;
  assign n12673 = ~n11626 & n12672 ;
  assign n12674 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & ~n11458 ;
  assign n12675 = n11626 & n12674 ;
  assign n12676 = ~n12673 & ~n12675 ;
  assign n12677 = \txethmac1_txcrc_Crc_reg[9]/NET0131  & n12676 ;
  assign n12678 = ~\txethmac1_txcrc_Crc_reg[9]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n12679 = n11458 & n12678 ;
  assign n12680 = ~n11626 & n12679 ;
  assign n12681 = ~n11458 & n12678 ;
  assign n12682 = n11626 & n12681 ;
  assign n12683 = ~n12680 & ~n12682 ;
  assign n12684 = n11464 & n12683 ;
  assign n12685 = ~n12677 & n12684 ;
  assign n12686 = ~n12528 & n12537 ;
  assign n12687 = \rxethmac1_rxstatem1_StateData0_reg/NET0131  & ~n10653 ;
  assign n12688 = ~n10648 & n12687 ;
  assign n12689 = ~\rxethmac1_rxstatem1_StateData1_reg/NET0131  & ~n12688 ;
  assign n12690 = n12686 & ~n12689 ;
  assign n12691 = ~n10653 & n12518 ;
  assign n12692 = n12517 & n12691 ;
  assign n12693 = ~\rxethmac1_rxstatem1_StateIdle_reg/NET0131  & ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n12694 = n12533 & n12693 ;
  assign n12695 = ~\ethreg1_MODER_0_DataOut_reg[6]/NET0131  & ~n12694 ;
  assign n12696 = ~n12523 & n12695 ;
  assign n12697 = \rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131  & ~\rxethmac1_rxstatem1_StateDrop_reg/NET0131  ;
  assign n12698 = n12696 & n12697 ;
  assign n12699 = ~n12692 & n12698 ;
  assign n12700 = \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  & \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131  ;
  assign n12701 = \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  & n12700 ;
  assign n12702 = n12699 & n12701 ;
  assign n12703 = ~\rxethmac1_rxstatem1_StateDrop_reg/NET0131  & ~n12692 ;
  assign n12704 = \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131  & n12703 ;
  assign n12705 = ~n12702 & n12704 ;
  assign n12706 = ~\rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131  & n12703 ;
  assign n12707 = n12702 & n12706 ;
  assign n12708 = ~n12705 & ~n12707 ;
  assign n12709 = \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  & n12699 ;
  assign n12710 = ~\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  & ~n12709 ;
  assign n12711 = \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  & \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  ;
  assign n12712 = n12699 & n12711 ;
  assign n12713 = n12703 & ~n12712 ;
  assign n12714 = ~n12710 & n12713 ;
  assign n12715 = ~\rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131  & ~n12712 ;
  assign n12716 = ~n12702 & n12703 ;
  assign n12717 = ~n12715 & n12716 ;
  assign n12718 = ~n12696 & n12697 ;
  assign n12719 = ~n12692 & n12718 ;
  assign n12720 = ~\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131  & ~\rxethmac1_rxstatem1_StateDrop_reg/NET0131  ;
  assign n12721 = n12696 & n12720 ;
  assign n12722 = ~n12692 & n12721 ;
  assign n12723 = ~n12719 & ~n12722 ;
  assign n12724 = \wishbone_TxPointerLSB_reg[0]/NET0131  & \wishbone_TxPointerLSB_reg[1]/NET0131  ;
  assign n12725 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & \txethmac1_TxUsedData_reg/NET0131  ;
  assign n12726 = \wishbone_TxStartFrm_reg/NET0131  & n12725 ;
  assign n12727 = n12724 & n12726 ;
  assign n12728 = \wishbone_Flop_reg/NET0131  & n12725 ;
  assign n12729 = \wishbone_TxData_reg[1]/NET0131  & ~n12728 ;
  assign n12730 = ~n12727 & n12729 ;
  assign n12731 = \wishbone_TxByteCnt_reg[0]/NET0131  & \wishbone_TxByteCnt_reg[1]/NET0131  ;
  assign n12732 = \wishbone_TxDataLatched_reg[1]/NET0131  & n12731 ;
  assign n12733 = \wishbone_TxByteCnt_reg[0]/NET0131  & ~\wishbone_TxByteCnt_reg[1]/NET0131  ;
  assign n12734 = \wishbone_TxDataLatched_reg[17]/NET0131  & n12733 ;
  assign n12735 = ~n12732 & ~n12734 ;
  assign n12736 = ~\wishbone_TxByteCnt_reg[0]/NET0131  & \wishbone_TxByteCnt_reg[1]/NET0131  ;
  assign n12737 = \wishbone_TxDataLatched_reg[9]/NET0131  & n12736 ;
  assign n12738 = ~\wishbone_TxByteCnt_reg[0]/NET0131  & ~\wishbone_TxByteCnt_reg[1]/NET0131  ;
  assign n12739 = \wishbone_TxDataLatched_reg[25]/NET0131  & n12738 ;
  assign n12740 = ~n12737 & ~n12739 ;
  assign n12741 = n12735 & n12740 ;
  assign n12742 = ~n12727 & n12728 ;
  assign n12743 = ~n12741 & n12742 ;
  assign n12744 = ~n12730 & ~n12743 ;
  assign n12745 = \wishbone_tx_fifo_data_out_reg[25]/P0001  & n12724 ;
  assign n12746 = n12726 & n12745 ;
  assign n12747 = ~\wishbone_TxStartFrm_reg/NET0131  & \wishbone_TxStartFrm_sync2_reg/NET0131  ;
  assign n12748 = ~n12746 & ~n12747 ;
  assign n12749 = n12744 & n12748 ;
  assign n12750 = ~\wishbone_TxPointerLSB_reg[0]/NET0131  & ~\wishbone_TxPointerLSB_reg[1]/NET0131  ;
  assign n12751 = \wishbone_tx_fifo_data_out_reg[25]/P0001  & n12750 ;
  assign n12752 = n12747 & ~n12751 ;
  assign n12753 = ~\wishbone_TxPointerLSB_reg[0]/NET0131  & \wishbone_TxPointerLSB_reg[1]/NET0131  ;
  assign n12754 = \wishbone_tx_fifo_data_out_reg[9]/P0001  & n12753 ;
  assign n12755 = \wishbone_tx_fifo_data_out_reg[1]/P0001  & n12724 ;
  assign n12756 = \wishbone_TxPointerLSB_reg[0]/NET0131  & ~\wishbone_TxPointerLSB_reg[1]/NET0131  ;
  assign n12757 = \wishbone_tx_fifo_data_out_reg[17]/P0001  & n12756 ;
  assign n12758 = ~n12755 & ~n12757 ;
  assign n12759 = ~n12754 & n12758 ;
  assign n12760 = n12752 & n12759 ;
  assign n12761 = ~n12749 & ~n12760 ;
  assign n12762 = \wishbone_TxData_reg[2]/NET0131  & ~n12728 ;
  assign n12763 = ~n12727 & n12762 ;
  assign n12764 = \wishbone_TxDataLatched_reg[10]/NET0131  & n12736 ;
  assign n12765 = \wishbone_TxDataLatched_reg[26]/NET0131  & n12738 ;
  assign n12766 = ~n12764 & ~n12765 ;
  assign n12767 = \wishbone_TxDataLatched_reg[2]/NET0131  & n12731 ;
  assign n12768 = \wishbone_TxDataLatched_reg[18]/NET0131  & n12733 ;
  assign n12769 = ~n12767 & ~n12768 ;
  assign n12770 = n12766 & n12769 ;
  assign n12771 = n12742 & ~n12770 ;
  assign n12772 = ~n12763 & ~n12771 ;
  assign n12773 = \wishbone_tx_fifo_data_out_reg[26]/P0001  & n12724 ;
  assign n12774 = n12726 & n12773 ;
  assign n12775 = ~n12747 & ~n12774 ;
  assign n12776 = n12772 & n12775 ;
  assign n12777 = \wishbone_tx_fifo_data_out_reg[26]/P0001  & n12750 ;
  assign n12778 = n12747 & ~n12777 ;
  assign n12779 = \wishbone_tx_fifo_data_out_reg[10]/P0001  & n12753 ;
  assign n12780 = \wishbone_tx_fifo_data_out_reg[2]/P0001  & n12724 ;
  assign n12781 = \wishbone_tx_fifo_data_out_reg[18]/P0001  & n12756 ;
  assign n12782 = ~n12780 & ~n12781 ;
  assign n12783 = ~n12779 & n12782 ;
  assign n12784 = n12778 & n12783 ;
  assign n12785 = ~n12776 & ~n12784 ;
  assign n12786 = \wishbone_TxData_reg[3]/NET0131  & ~n12728 ;
  assign n12787 = ~n12727 & n12786 ;
  assign n12788 = \wishbone_TxDataLatched_reg[3]/NET0131  & n12731 ;
  assign n12789 = \wishbone_TxDataLatched_reg[19]/NET0131  & n12733 ;
  assign n12790 = ~n12788 & ~n12789 ;
  assign n12791 = \wishbone_TxDataLatched_reg[11]/NET0131  & n12736 ;
  assign n12792 = \wishbone_TxDataLatched_reg[27]/NET0131  & n12738 ;
  assign n12793 = ~n12791 & ~n12792 ;
  assign n12794 = n12790 & n12793 ;
  assign n12795 = n12742 & ~n12794 ;
  assign n12796 = ~n12787 & ~n12795 ;
  assign n12797 = \wishbone_tx_fifo_data_out_reg[27]/P0001  & n12724 ;
  assign n12798 = n12726 & n12797 ;
  assign n12799 = ~n12747 & ~n12798 ;
  assign n12800 = n12796 & n12799 ;
  assign n12801 = \wishbone_tx_fifo_data_out_reg[27]/P0001  & n12750 ;
  assign n12802 = n12747 & ~n12801 ;
  assign n12803 = \wishbone_tx_fifo_data_out_reg[11]/P0001  & n12753 ;
  assign n12804 = \wishbone_tx_fifo_data_out_reg[3]/P0001  & n12724 ;
  assign n12805 = \wishbone_tx_fifo_data_out_reg[19]/P0001  & n12756 ;
  assign n12806 = ~n12804 & ~n12805 ;
  assign n12807 = ~n12803 & n12806 ;
  assign n12808 = n12802 & n12807 ;
  assign n12809 = ~n12800 & ~n12808 ;
  assign n12810 = \wishbone_TxData_reg[4]/NET0131  & ~n12728 ;
  assign n12811 = ~n12727 & n12810 ;
  assign n12812 = \wishbone_TxDataLatched_reg[4]/NET0131  & n12731 ;
  assign n12813 = \wishbone_TxDataLatched_reg[20]/NET0131  & n12733 ;
  assign n12814 = ~n12812 & ~n12813 ;
  assign n12815 = \wishbone_TxDataLatched_reg[12]/NET0131  & n12736 ;
  assign n12816 = \wishbone_TxDataLatched_reg[28]/NET0131  & n12738 ;
  assign n12817 = ~n12815 & ~n12816 ;
  assign n12818 = n12814 & n12817 ;
  assign n12819 = n12742 & ~n12818 ;
  assign n12820 = ~n12811 & ~n12819 ;
  assign n12821 = \wishbone_tx_fifo_data_out_reg[28]/P0001  & n12724 ;
  assign n12822 = n12726 & n12821 ;
  assign n12823 = ~n12747 & ~n12822 ;
  assign n12824 = n12820 & n12823 ;
  assign n12825 = \wishbone_tx_fifo_data_out_reg[28]/P0001  & n12750 ;
  assign n12826 = n12747 & ~n12825 ;
  assign n12827 = \wishbone_tx_fifo_data_out_reg[12]/P0001  & n12753 ;
  assign n12828 = \wishbone_tx_fifo_data_out_reg[4]/P0001  & n12724 ;
  assign n12829 = \wishbone_tx_fifo_data_out_reg[20]/P0001  & n12756 ;
  assign n12830 = ~n12828 & ~n12829 ;
  assign n12831 = ~n12827 & n12830 ;
  assign n12832 = n12826 & n12831 ;
  assign n12833 = ~n12824 & ~n12832 ;
  assign n12834 = \wishbone_TxData_reg[0]/NET0131  & ~n12728 ;
  assign n12835 = ~n12727 & n12834 ;
  assign n12836 = \wishbone_TxDataLatched_reg[8]/NET0131  & n12736 ;
  assign n12837 = \wishbone_TxDataLatched_reg[24]/NET0131  & n12738 ;
  assign n12838 = ~n12836 & ~n12837 ;
  assign n12839 = \wishbone_TxDataLatched_reg[0]/NET0131  & n12731 ;
  assign n12840 = \wishbone_TxDataLatched_reg[16]/NET0131  & n12733 ;
  assign n12841 = ~n12839 & ~n12840 ;
  assign n12842 = n12838 & n12841 ;
  assign n12843 = n12742 & ~n12842 ;
  assign n12844 = ~n12835 & ~n12843 ;
  assign n12845 = \wishbone_tx_fifo_data_out_reg[24]/P0001  & n12724 ;
  assign n12846 = n12726 & n12845 ;
  assign n12847 = ~n12747 & ~n12846 ;
  assign n12848 = n12844 & n12847 ;
  assign n12849 = \wishbone_tx_fifo_data_out_reg[24]/P0001  & n12750 ;
  assign n12850 = n12747 & ~n12849 ;
  assign n12851 = \wishbone_tx_fifo_data_out_reg[8]/P0001  & n12753 ;
  assign n12852 = \wishbone_tx_fifo_data_out_reg[0]/P0001  & n12724 ;
  assign n12853 = \wishbone_tx_fifo_data_out_reg[16]/P0001  & n12756 ;
  assign n12854 = ~n12852 & ~n12853 ;
  assign n12855 = ~n12851 & n12854 ;
  assign n12856 = n12850 & n12855 ;
  assign n12857 = ~n12848 & ~n12856 ;
  assign n12858 = \wishbone_TxData_reg[6]/NET0131  & ~n12728 ;
  assign n12859 = ~n12727 & n12858 ;
  assign n12860 = \wishbone_TxDataLatched_reg[6]/NET0131  & n12731 ;
  assign n12861 = \wishbone_TxDataLatched_reg[22]/NET0131  & n12733 ;
  assign n12862 = ~n12860 & ~n12861 ;
  assign n12863 = \wishbone_TxDataLatched_reg[14]/NET0131  & n12736 ;
  assign n12864 = \wishbone_TxDataLatched_reg[30]/NET0131  & n12738 ;
  assign n12865 = ~n12863 & ~n12864 ;
  assign n12866 = n12862 & n12865 ;
  assign n12867 = n12742 & ~n12866 ;
  assign n12868 = ~n12859 & ~n12867 ;
  assign n12869 = \wishbone_tx_fifo_data_out_reg[30]/P0001  & n12724 ;
  assign n12870 = n12726 & n12869 ;
  assign n12871 = ~n12747 & ~n12870 ;
  assign n12872 = n12868 & n12871 ;
  assign n12873 = \wishbone_tx_fifo_data_out_reg[30]/P0001  & n12750 ;
  assign n12874 = n12747 & ~n12873 ;
  assign n12875 = \wishbone_tx_fifo_data_out_reg[14]/P0001  & n12753 ;
  assign n12876 = \wishbone_tx_fifo_data_out_reg[6]/P0001  & n12724 ;
  assign n12877 = \wishbone_tx_fifo_data_out_reg[22]/P0001  & n12756 ;
  assign n12878 = ~n12876 & ~n12877 ;
  assign n12879 = ~n12875 & n12878 ;
  assign n12880 = n12874 & n12879 ;
  assign n12881 = ~n12872 & ~n12880 ;
  assign n12882 = \wishbone_TxData_reg[5]/NET0131  & ~n12728 ;
  assign n12883 = ~n12727 & n12882 ;
  assign n12884 = \wishbone_TxDataLatched_reg[5]/NET0131  & n12731 ;
  assign n12885 = \wishbone_TxDataLatched_reg[21]/NET0131  & n12733 ;
  assign n12886 = ~n12884 & ~n12885 ;
  assign n12887 = \wishbone_TxDataLatched_reg[13]/NET0131  & n12736 ;
  assign n12888 = \wishbone_TxDataLatched_reg[29]/NET0131  & n12738 ;
  assign n12889 = ~n12887 & ~n12888 ;
  assign n12890 = n12886 & n12889 ;
  assign n12891 = n12742 & ~n12890 ;
  assign n12892 = ~n12883 & ~n12891 ;
  assign n12893 = \wishbone_tx_fifo_data_out_reg[29]/P0001  & n12724 ;
  assign n12894 = n12726 & n12893 ;
  assign n12895 = ~n12747 & ~n12894 ;
  assign n12896 = n12892 & n12895 ;
  assign n12897 = \wishbone_tx_fifo_data_out_reg[29]/P0001  & n12750 ;
  assign n12898 = n12747 & ~n12897 ;
  assign n12899 = \wishbone_tx_fifo_data_out_reg[13]/P0001  & n12753 ;
  assign n12900 = \wishbone_tx_fifo_data_out_reg[5]/P0001  & n12724 ;
  assign n12901 = \wishbone_tx_fifo_data_out_reg[21]/P0001  & n12756 ;
  assign n12902 = ~n12900 & ~n12901 ;
  assign n12903 = ~n12899 & n12902 ;
  assign n12904 = n12898 & n12903 ;
  assign n12905 = ~n12896 & ~n12904 ;
  assign n12906 = \wishbone_TxData_reg[7]/NET0131  & ~n12728 ;
  assign n12907 = ~n12727 & n12906 ;
  assign n12908 = \wishbone_TxDataLatched_reg[7]/NET0131  & n12731 ;
  assign n12909 = \wishbone_TxDataLatched_reg[23]/NET0131  & n12733 ;
  assign n12910 = ~n12908 & ~n12909 ;
  assign n12911 = \wishbone_TxDataLatched_reg[15]/NET0131  & n12736 ;
  assign n12912 = \wishbone_TxDataLatched_reg[31]/NET0131  & n12738 ;
  assign n12913 = ~n12911 & ~n12912 ;
  assign n12914 = n12910 & n12913 ;
  assign n12915 = n12742 & ~n12914 ;
  assign n12916 = ~n12907 & ~n12915 ;
  assign n12917 = \wishbone_tx_fifo_data_out_reg[31]/P0001  & n12724 ;
  assign n12918 = n12726 & n12917 ;
  assign n12919 = ~n12747 & ~n12918 ;
  assign n12920 = n12916 & n12919 ;
  assign n12921 = \wishbone_tx_fifo_data_out_reg[31]/P0001  & n12750 ;
  assign n12922 = n12747 & ~n12921 ;
  assign n12923 = \wishbone_tx_fifo_data_out_reg[15]/P0001  & n12753 ;
  assign n12924 = \wishbone_tx_fifo_data_out_reg[7]/P0001  & n12724 ;
  assign n12925 = \wishbone_tx_fifo_data_out_reg[23]/P0001  & n12756 ;
  assign n12926 = ~n12924 & ~n12925 ;
  assign n12927 = ~n12923 & n12926 ;
  assign n12928 = n12922 & n12927 ;
  assign n12929 = ~n12920 & ~n12928 ;
  assign n12930 = ~\rxethmac1_crcrx_Crc_reg[1]/NET0131  & n10663 ;
  assign n12931 = ~n12218 & n12930 ;
  assign n12932 = \rxethmac1_crcrx_Crc_reg[1]/NET0131  & n10663 ;
  assign n12933 = n12218 & n12932 ;
  assign n12934 = ~n12931 & ~n12933 ;
  assign n12935 = \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  & ~\rxethmac1_rxstatem1_StateDrop_reg/NET0131  ;
  assign n12936 = ~n12692 & n12935 ;
  assign n12937 = ~n12699 & n12936 ;
  assign n12938 = ~\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  & ~\rxethmac1_rxstatem1_StateDrop_reg/NET0131  ;
  assign n12939 = ~n12692 & n12938 ;
  assign n12940 = n12699 & n12939 ;
  assign n12941 = ~n12937 & ~n12940 ;
  assign n12942 = ~\rxethmac1_rxstatem1_StateIdle_reg/NET0131  & n10649 ;
  assign n12943 = n12534 & n12942 ;
  assign n12944 = n10653 & ~n12943 ;
  assign n12945 = \txethmac1_txcrc_Crc_reg[30]/NET0131  & ~\txethmac1_txcrc_Crc_reg[31]/NET0131  ;
  assign n12946 = ~\txethmac1_txcrc_Crc_reg[30]/NET0131  & \txethmac1_txcrc_Crc_reg[31]/NET0131  ;
  assign n12947 = ~n12945 & ~n12946 ;
  assign n12948 = ~n11502 & ~n12947 ;
  assign n12949 = ~n11455 & n12948 ;
  assign n12950 = ~n11446 & n12949 ;
  assign n12951 = n11502 & ~n12947 ;
  assign n12952 = ~n11455 & n12951 ;
  assign n12953 = n11446 & n12952 ;
  assign n12954 = ~n12950 & ~n12953 ;
  assign n12955 = n11455 & n12948 ;
  assign n12956 = n11446 & n12955 ;
  assign n12957 = n11455 & n12951 ;
  assign n12958 = ~n11446 & n12957 ;
  assign n12959 = ~n12956 & ~n12958 ;
  assign n12960 = n12954 & n12959 ;
  assign n12961 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n12960 ;
  assign n12962 = ~n11502 & n12947 ;
  assign n12963 = ~n11455 & n12962 ;
  assign n12964 = n11446 & n12963 ;
  assign n12965 = n11502 & n12947 ;
  assign n12966 = ~n11455 & n12965 ;
  assign n12967 = ~n11446 & n12966 ;
  assign n12968 = ~n12964 & ~n12967 ;
  assign n12969 = n11455 & n12962 ;
  assign n12970 = ~n11446 & n12969 ;
  assign n12971 = n11455 & n12965 ;
  assign n12972 = n11446 & n12971 ;
  assign n12973 = ~n12970 & ~n12972 ;
  assign n12974 = n12968 & n12973 ;
  assign n12975 = ~\txethmac1_txcrc_Crc_reg[6]/NET0131  & n12974 ;
  assign n12976 = n12961 & n12975 ;
  assign n12977 = ~\txethmac1_txcrc_Crc_reg[6]/NET0131  & n11464 ;
  assign n12978 = n11464 & n12974 ;
  assign n12979 = n12961 & n12978 ;
  assign n12980 = ~n12977 & ~n12979 ;
  assign n12981 = ~n12976 & ~n12980 ;
  assign n12982 = \txethmac1_txcrc_Crc_reg[29]/NET0131  & ~\txethmac1_txcrc_Crc_reg[31]/NET0131  ;
  assign n12983 = ~\txethmac1_txcrc_Crc_reg[29]/NET0131  & \txethmac1_txcrc_Crc_reg[31]/NET0131  ;
  assign n12984 = ~n12982 & ~n12983 ;
  assign n12985 = ~n11478 & ~n12984 ;
  assign n12986 = ~n11455 & n12985 ;
  assign n12987 = ~n11446 & n12986 ;
  assign n12988 = n11478 & ~n12984 ;
  assign n12989 = ~n11455 & n12988 ;
  assign n12990 = n11446 & n12989 ;
  assign n12991 = ~n12987 & ~n12990 ;
  assign n12992 = n11455 & n12985 ;
  assign n12993 = n11446 & n12992 ;
  assign n12994 = n11455 & n12988 ;
  assign n12995 = ~n11446 & n12994 ;
  assign n12996 = ~n12993 & ~n12995 ;
  assign n12997 = n12991 & n12996 ;
  assign n12998 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n12997 ;
  assign n12999 = ~n11478 & n12984 ;
  assign n13000 = ~n11455 & n12999 ;
  assign n13001 = n11446 & n13000 ;
  assign n13002 = n11478 & n12984 ;
  assign n13003 = ~n11455 & n13002 ;
  assign n13004 = ~n11446 & n13003 ;
  assign n13005 = ~n13001 & ~n13004 ;
  assign n13006 = n11455 & n12999 ;
  assign n13007 = ~n11446 & n13006 ;
  assign n13008 = n11455 & n13002 ;
  assign n13009 = n11446 & n13008 ;
  assign n13010 = ~n13007 & ~n13009 ;
  assign n13011 = n13005 & n13010 ;
  assign n13012 = ~\txethmac1_txcrc_Crc_reg[7]/NET0131  & n13011 ;
  assign n13013 = n12998 & n13012 ;
  assign n13014 = ~\txethmac1_txcrc_Crc_reg[7]/NET0131  & n11464 ;
  assign n13015 = n11464 & n13011 ;
  assign n13016 = n12998 & n13015 ;
  assign n13017 = ~n13014 & ~n13016 ;
  assign n13018 = ~n13013 & ~n13017 ;
  assign n13019 = ~\rxethmac1_RxEndFrm_reg/NET0131  & ~\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131  ;
  assign n13020 = \rxethmac1_Broadcast_reg/NET0131  & n13019 ;
  assign n13021 = ~\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  & n10522 ;
  assign n13022 = n10519 & n13021 ;
  assign n13023 = \rxethmac1_LatchedByte_reg[4]/NET0131  & \rxethmac1_LatchedByte_reg[5]/NET0131  ;
  assign n13024 = \rxethmac1_LatchedByte_reg[6]/NET0131  & \rxethmac1_LatchedByte_reg[7]/NET0131  ;
  assign n13025 = n13023 & n13024 ;
  assign n13026 = \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n13027 = n10565 & n13026 ;
  assign n13028 = n13025 & n13027 ;
  assign n13029 = n13022 & n13028 ;
  assign n13030 = ~n13020 & ~n13029 ;
  assign n13031 = n10519 & n10522 ;
  assign n13032 = \rxethmac1_LatchedByte_reg[0]/NET0131  & \rxethmac1_LatchedByte_reg[1]/NET0131  ;
  assign n13033 = \rxethmac1_LatchedByte_reg[2]/NET0131  & \rxethmac1_LatchedByte_reg[3]/NET0131  ;
  assign n13034 = n13032 & n13033 ;
  assign n13035 = n13025 & n13034 ;
  assign n13036 = n10565 & ~n12638 ;
  assign n13037 = ~n13035 & n13036 ;
  assign n13038 = n13031 & n13037 ;
  assign n13039 = ~n13030 & ~n13038 ;
  assign n13040 = ~n12528 & ~n12536 ;
  assign n13041 = ~\rxethmac1_rxstatem1_StateData0_reg/NET0131  & n12532 ;
  assign n13042 = ~n12688 & ~n13041 ;
  assign n13043 = n13040 & n13042 ;
  assign n13044 = ~n10653 & n12539 ;
  assign n13045 = ~\rxethmac1_rxstatem1_StatePreamble_reg/NET0131  & ~n12542 ;
  assign n13046 = ~n13044 & ~n13045 ;
  assign n13047 = ~n12536 & n13046 ;
  assign n13048 = ~n12528 & n13047 ;
  assign n13049 = n10566 & ~n10649 ;
  assign n13050 = n10525 & n13049 ;
  assign n13051 = ~\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  & ~n10649 ;
  assign n13052 = n10512 & n13051 ;
  assign n13053 = n10564 & n13052 ;
  assign n13054 = ~n10649 & n12580 ;
  assign n13055 = n10525 & n13054 ;
  assign n13056 = n12461 & n13053 ;
  assign n13057 = ~n13055 & ~n13056 ;
  assign n13058 = n13053 & n13057 ;
  assign n13059 = n13026 & n13051 ;
  assign n13060 = n10564 & n13059 ;
  assign n13061 = n10566 & n13051 ;
  assign n13062 = n10564 & n13061 ;
  assign n13063 = n12423 & n13062 ;
  assign n13064 = ~n13060 & n13063 ;
  assign n13065 = n12580 & n13051 ;
  assign n13066 = n10564 & n13065 ;
  assign n13067 = ~n13019 & ~n13066 ;
  assign n13068 = ~n13062 & ~n13067 ;
  assign n13069 = ~n12389 & n13066 ;
  assign n13070 = ~n13060 & ~n13069 ;
  assign n13071 = n13068 & n13070 ;
  assign n13072 = ~n13064 & ~n13071 ;
  assign n13073 = n12499 & n13060 ;
  assign n13074 = n13057 & ~n13073 ;
  assign n13075 = n13072 & n13074 ;
  assign n13076 = ~n13058 & ~n13075 ;
  assign n13077 = ~n12345 & n13055 ;
  assign n13078 = \rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131  & ~n13077 ;
  assign n13079 = n13076 & n13078 ;
  assign n13080 = ~n13050 & ~n13079 ;
  assign n13081 = ~n12307 & n13050 ;
  assign n13082 = ~n13080 & ~n13081 ;
  assign n13083 = ~\rxethmac1_rxstatem1_StateDrop_reg/NET0131  & ~n12515 ;
  assign n13084 = ~n12525 & n13083 ;
  assign n13085 = ~n12167 & n13084 ;
  assign n13086 = ~n10653 & ~n13085 ;
  assign n13087 = ~\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131  ;
  assign n13088 = ~\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131  & ~n13087 ;
  assign n13089 = ~\macstatus1_InvalidSymbol_reg/NET0131  & \macstatus1_LatchedMRxErr_reg/NET0131  ;
  assign n13090 = ~\ethreg1_MODER_2_DataOut_reg[0]/NET0131  & \macstatus1_ShortFrame_reg/NET0131  ;
  assign n13091 = ~\RxAbortRst_reg/NET0131  & \RxAbort_latch_reg/NET0131  ;
  assign n13092 = ~n13090 & ~n13091 ;
  assign n13093 = ~n13089 & n13092 ;
  assign n13094 = n13088 & n13093 ;
  assign n13095 = \m_wb_adr_o[2]_pad  & \m_wb_adr_o[3]_pad  ;
  assign n13096 = \m_wb_adr_o[4]_pad  & \m_wb_adr_o[5]_pad  ;
  assign n13097 = n13095 & n13096 ;
  assign n13098 = \m_wb_adr_o[6]_pad  & \m_wb_adr_o[8]_pad  ;
  assign n13099 = \m_wb_adr_o[7]_pad  & n13098 ;
  assign n13100 = n13097 & n13099 ;
  assign n13101 = \m_wb_adr_o[10]_pad  & \m_wb_adr_o[9]_pad  ;
  assign n13102 = \m_wb_adr_o[11]_pad  & n13101 ;
  assign n13103 = n13100 & n13102 ;
  assign n13104 = \m_wb_adr_o[13]_pad  & \m_wb_adr_o[14]_pad  ;
  assign n13105 = \m_wb_adr_o[12]_pad  & \m_wb_adr_o[15]_pad  ;
  assign n13106 = n13104 & n13105 ;
  assign n13107 = n13103 & n13106 ;
  assign n13108 = \m_wb_adr_o[17]_pad  & \m_wb_adr_o[18]_pad  ;
  assign n13109 = \m_wb_adr_o[16]_pad  & \m_wb_adr_o[19]_pad  ;
  assign n13110 = n13108 & n13109 ;
  assign n13111 = n13107 & n13110 ;
  assign n13112 = \m_wb_adr_o[20]_pad  & \m_wb_adr_o[21]_pad  ;
  assign n13113 = \m_wb_adr_o[22]_pad  & \m_wb_adr_o[23]_pad  ;
  assign n13114 = \m_wb_adr_o[24]_pad  & n13113 ;
  assign n13115 = \m_wb_adr_o[25]_pad  & \m_wb_adr_o[26]_pad  ;
  assign n13116 = n13114 & n13115 ;
  assign n13117 = n13112 & n13116 ;
  assign n13118 = n13111 & n13117 ;
  assign n13119 = \m_wb_adr_o[27]_pad  & \m_wb_adr_o[28]_pad  ;
  assign n13120 = \m_wb_adr_o[29]_pad  & n13119 ;
  assign n13121 = n13118 & n13120 ;
  assign n13122 = ~\m_wb_adr_o[30]_pad  & ~n13121 ;
  assign n13123 = \m_wb_adr_o[29]_pad  & \m_wb_adr_o[30]_pad  ;
  assign n13124 = n13119 & n13123 ;
  assign n13125 = n13118 & n13124 ;
  assign n13126 = ~\wishbone_rx_fifo_cnt_reg[0]/NET0131  & ~\wishbone_rx_fifo_cnt_reg[1]/NET0131  ;
  assign n13127 = ~\wishbone_rx_fifo_cnt_reg[2]/NET0131  & n13126 ;
  assign n13128 = ~\wishbone_rx_fifo_cnt_reg[3]/NET0131  & ~\wishbone_rx_fifo_cnt_reg[4]/NET0131  ;
  assign n13129 = n13127 & n13128 ;
  assign n13130 = \wishbone_rx_burst_en_reg/NET0131  & ~n13129 ;
  assign n13131 = ~m_wb_ack_i_pad & ~m_wb_err_i_pad ;
  assign n13132 = \wishbone_MasterWbRX_reg/NET0131  & \wishbone_cyc_cleared_reg/NET0131  ;
  assign n13133 = ~n13131 & n13132 ;
  assign n13134 = \wishbone_MasterWbRX_reg/NET0131  & ~\wishbone_cyc_cleared_reg/NET0131  ;
  assign n13135 = n13131 & n13134 ;
  assign n13136 = ~n13133 & ~n13135 ;
  assign n13137 = n13130 & n13136 ;
  assign n13138 = ~\wishbone_MasterWbRX_reg/NET0131  & \wishbone_cyc_cleared_reg/NET0131  ;
  assign n13139 = \wishbone_MasterWbTX_reg/NET0131  & ~n13138 ;
  assign n13140 = ~\wishbone_MasterWbTX_reg/NET0131  & n13138 ;
  assign n13141 = ~\wishbone_MasterWbRX_reg/NET0131  & ~n13131 ;
  assign n13142 = ~n13140 & ~n13141 ;
  assign n13143 = ~n13139 & n13142 ;
  assign n13144 = ~\wishbone_rx_burst_cnt_reg[0]/NET0131  & ~\wishbone_rx_burst_cnt_reg[1]/NET0131  ;
  assign n13145 = ~\wishbone_RxPointerMSB_reg[30]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n13146 = n13144 & n13145 ;
  assign n13147 = ~\wishbone_BlockReadTxDataFromMemory_reg/NET0131  & \wishbone_ReadTxDataFromMemory_reg/NET0131  ;
  assign n13148 = \wishbone_MasterWbRX_reg/NET0131  & n13147 ;
  assign n13149 = n13131 & n13148 ;
  assign n13150 = ~n13146 & ~n13149 ;
  assign n13151 = n13143 & n13150 ;
  assign n13152 = n13137 & n13151 ;
  assign n13153 = n13131 & ~n13138 ;
  assign n13154 = ~n13134 & n13153 ;
  assign n13155 = \wishbone_tx_burst_en_reg/NET0131  & n13147 ;
  assign n13156 = ~\wishbone_MasterWbTX_reg/NET0131  & n13155 ;
  assign n13157 = n13154 & n13156 ;
  assign n13158 = ~\wishbone_MasterWbRX_reg/NET0131  & ~\wishbone_cyc_cleared_reg/NET0131  ;
  assign n13159 = ~n13131 & n13158 ;
  assign n13160 = n13131 & n13138 ;
  assign n13161 = ~n13159 & ~n13160 ;
  assign n13162 = \wishbone_MasterWbTX_reg/NET0131  & n13155 ;
  assign n13163 = ~n13161 & n13162 ;
  assign n13164 = ~n13157 & ~n13163 ;
  assign n13165 = ~\wishbone_MasterWbRX_reg/NET0131  & n13131 ;
  assign n13166 = ~n13129 & n13165 ;
  assign n13167 = ~\wishbone_tx_burst_cnt_reg[0]/NET0131  & ~\wishbone_tx_burst_cnt_reg[1]/NET0131  ;
  assign n13168 = ~\wishbone_tx_burst_cnt_reg[2]/NET0131  & n13167 ;
  assign n13169 = ~n13166 & ~n13168 ;
  assign n13170 = ~n13164 & n13169 ;
  assign n13171 = ~n13152 & ~n13170 ;
  assign n13172 = ~n13125 & ~n13171 ;
  assign n13173 = ~n13122 & n13172 ;
  assign n13174 = ~n13164 & ~n13166 ;
  assign n13175 = ~\wishbone_tx_burst_en_reg/NET0131  & n13147 ;
  assign n13176 = ~\wishbone_MasterWbRX_reg/NET0131  & ~\wishbone_MasterWbTX_reg/NET0131  ;
  assign n13177 = ~\wishbone_cyc_cleared_reg/NET0131  & n13131 ;
  assign n13178 = n13176 & n13177 ;
  assign n13179 = n13129 & n13178 ;
  assign n13180 = n13175 & n13179 ;
  assign n13181 = ~\wishbone_MasterWbRX_reg/NET0131  & ~n13129 ;
  assign n13182 = \wishbone_cyc_cleared_reg/NET0131  & n13131 ;
  assign n13183 = \wishbone_MasterWbRX_reg/NET0131  & \wishbone_MasterWbTX_reg/NET0131  ;
  assign n13184 = ~n13176 & ~n13183 ;
  assign n13185 = n13182 & n13184 ;
  assign n13186 = n13175 & n13185 ;
  assign n13187 = ~n13181 & n13186 ;
  assign n13188 = ~n13180 & ~n13187 ;
  assign n13189 = ~n13174 & n13188 ;
  assign n13190 = n13143 & ~n13149 ;
  assign n13191 = n13137 & n13190 ;
  assign n13192 = ~\wishbone_rx_burst_en_reg/NET0131  & ~n13129 ;
  assign n13193 = ~n13148 & n13185 ;
  assign n13194 = ~n13178 & ~n13193 ;
  assign n13195 = n13192 & ~n13194 ;
  assign n13196 = ~n13191 & ~n13195 ;
  assign n13197 = n13189 & n13196 ;
  assign n13198 = \m_wb_adr_o[30]_pad  & n13197 ;
  assign n13199 = ~n13166 & n13168 ;
  assign n13200 = ~n13164 & n13199 ;
  assign n13201 = n13188 & ~n13200 ;
  assign n13202 = \wishbone_TxPointerMSB_reg[30]/NET0131  & ~n13201 ;
  assign n13203 = ~\wishbone_rx_burst_cnt_reg[2]/NET0131  & n13144 ;
  assign n13204 = ~n13192 & ~n13203 ;
  assign n13205 = ~n13178 & ~n13203 ;
  assign n13206 = ~n13193 & n13205 ;
  assign n13207 = ~n13204 & ~n13206 ;
  assign n13208 = \wishbone_RxPointerMSB_reg[30]/NET0131  & n13207 ;
  assign n13209 = ~n13196 & n13208 ;
  assign n13210 = ~n13202 & ~n13209 ;
  assign n13211 = ~n13198 & n13210 ;
  assign n13212 = ~n13173 & n13211 ;
  assign n13213 = \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & n12275 ;
  assign n13214 = n12274 & n13213 ;
  assign n13215 = ~n12347 & ~n13214 ;
  assign n13216 = \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  & \rxethmac1_RxValid_reg/NET0131  ;
  assign n13217 = n12265 & n13216 ;
  assign n13218 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  & n13217 ;
  assign n13219 = \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  & \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n13220 = n12354 & n13219 ;
  assign n13221 = ~n13218 & ~n13220 ;
  assign n13222 = n13215 & ~n13221 ;
  assign n13223 = \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131  & ~n13222 ;
  assign n13224 = \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  & n12354 ;
  assign n13225 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  ;
  assign n13226 = n12312 & n13225 ;
  assign n13227 = n12274 & n13226 ;
  assign n13228 = n13224 & n13227 ;
  assign n13229 = ~n13223 & ~n13228 ;
  assign n13230 = ~\wishbone_bd_ram_raddr_reg[0]/P0001  & ~\wishbone_bd_ram_raddr_reg[1]/NET0131  ;
  assign n13231 = \wishbone_bd_ram_raddr_reg[2]/NET0131  & ~\wishbone_bd_ram_raddr_reg[3]/P0001  ;
  assign n13232 = n13230 & n13231 ;
  assign n13233 = ~\wishbone_bd_ram_raddr_reg[4]/NET0131  & \wishbone_bd_ram_raddr_reg[5]/NET0131  ;
  assign n13234 = ~\wishbone_bd_ram_raddr_reg[6]/NET0131  & \wishbone_bd_ram_raddr_reg[7]/NET0131  ;
  assign n13235 = n13233 & n13234 ;
  assign n13236 = n13232 & n13235 ;
  assign n13237 = \wishbone_bd_ram_mem3_reg[164][28]/P0001  & n13236 ;
  assign n13238 = ~\wishbone_bd_ram_raddr_reg[6]/NET0131  & ~\wishbone_bd_ram_raddr_reg[7]/NET0131  ;
  assign n13239 = ~\wishbone_bd_ram_raddr_reg[4]/NET0131  & ~\wishbone_bd_ram_raddr_reg[5]/NET0131  ;
  assign n13240 = n13238 & n13239 ;
  assign n13241 = \wishbone_bd_ram_raddr_reg[0]/P0001  & ~\wishbone_bd_ram_raddr_reg[1]/NET0131  ;
  assign n13242 = n13231 & n13241 ;
  assign n13243 = n13240 & n13242 ;
  assign n13244 = \wishbone_bd_ram_mem3_reg[5][28]/P0001  & n13243 ;
  assign n13245 = ~n13237 & ~n13244 ;
  assign n13246 = \wishbone_bd_ram_raddr_reg[4]/NET0131  & ~\wishbone_bd_ram_raddr_reg[5]/NET0131  ;
  assign n13247 = n13238 & n13246 ;
  assign n13248 = \wishbone_bd_ram_raddr_reg[0]/P0001  & \wishbone_bd_ram_raddr_reg[1]/NET0131  ;
  assign n13249 = ~\wishbone_bd_ram_raddr_reg[2]/NET0131  & \wishbone_bd_ram_raddr_reg[3]/P0001  ;
  assign n13250 = n13248 & n13249 ;
  assign n13251 = n13247 & n13250 ;
  assign n13252 = \wishbone_bd_ram_mem3_reg[27][28]/P0001  & n13251 ;
  assign n13253 = ~\wishbone_bd_ram_raddr_reg[2]/NET0131  & ~\wishbone_bd_ram_raddr_reg[3]/P0001  ;
  assign n13254 = n13248 & n13253 ;
  assign n13255 = n13235 & n13254 ;
  assign n13256 = \wishbone_bd_ram_mem3_reg[163][28]/P0001  & n13255 ;
  assign n13257 = ~n13252 & ~n13256 ;
  assign n13258 = n13245 & n13257 ;
  assign n13259 = n13230 & n13253 ;
  assign n13260 = \wishbone_bd_ram_raddr_reg[4]/NET0131  & \wishbone_bd_ram_raddr_reg[5]/NET0131  ;
  assign n13261 = n13234 & n13260 ;
  assign n13262 = n13259 & n13261 ;
  assign n13263 = \wishbone_bd_ram_mem3_reg[176][28]/P0001  & n13262 ;
  assign n13264 = ~\wishbone_bd_ram_raddr_reg[0]/P0001  & \wishbone_bd_ram_raddr_reg[1]/NET0131  ;
  assign n13265 = n13249 & n13264 ;
  assign n13266 = \wishbone_bd_ram_raddr_reg[6]/NET0131  & \wishbone_bd_ram_raddr_reg[7]/NET0131  ;
  assign n13267 = n13239 & n13266 ;
  assign n13268 = n13265 & n13267 ;
  assign n13269 = \wishbone_bd_ram_mem3_reg[202][28]/P0001  & n13268 ;
  assign n13270 = ~n13263 & ~n13269 ;
  assign n13271 = n13235 & n13259 ;
  assign n13272 = \wishbone_bd_ram_mem3_reg[160][28]/P0001  & n13271 ;
  assign n13273 = \wishbone_bd_ram_raddr_reg[2]/NET0131  & \wishbone_bd_ram_raddr_reg[3]/P0001  ;
  assign n13274 = n13264 & n13273 ;
  assign n13275 = \wishbone_bd_ram_raddr_reg[6]/NET0131  & ~\wishbone_bd_ram_raddr_reg[7]/NET0131  ;
  assign n13276 = n13239 & n13275 ;
  assign n13277 = n13274 & n13276 ;
  assign n13278 = \wishbone_bd_ram_mem3_reg[78][28]/P0001  & n13277 ;
  assign n13279 = ~n13272 & ~n13278 ;
  assign n13280 = n13270 & n13279 ;
  assign n13281 = n13258 & n13280 ;
  assign n13282 = n13260 & n13266 ;
  assign n13283 = n13274 & n13282 ;
  assign n13284 = \wishbone_bd_ram_mem3_reg[254][28]/P0001  & n13283 ;
  assign n13285 = n13230 & n13273 ;
  assign n13286 = n13234 & n13239 ;
  assign n13287 = n13285 & n13286 ;
  assign n13288 = \wishbone_bd_ram_mem3_reg[140][28]/P0001  & n13287 ;
  assign n13289 = ~n13284 & ~n13288 ;
  assign n13290 = n13233 & n13238 ;
  assign n13291 = n13285 & n13290 ;
  assign n13292 = \wishbone_bd_ram_mem3_reg[44][28]/P0001  & n13291 ;
  assign n13293 = n13234 & n13246 ;
  assign n13294 = n13274 & n13293 ;
  assign n13295 = \wishbone_bd_ram_mem3_reg[158][28]/P0001  & n13294 ;
  assign n13296 = ~n13292 & ~n13295 ;
  assign n13297 = n13289 & n13296 ;
  assign n13298 = n13274 & n13290 ;
  assign n13299 = \wishbone_bd_ram_mem3_reg[46][28]/P0001  & n13298 ;
  assign n13300 = n13253 & n13264 ;
  assign n13301 = n13261 & n13300 ;
  assign n13302 = \wishbone_bd_ram_mem3_reg[178][28]/P0001  & n13301 ;
  assign n13303 = ~n13299 & ~n13302 ;
  assign n13304 = n13233 & n13275 ;
  assign n13305 = n13241 & n13273 ;
  assign n13306 = n13304 & n13305 ;
  assign n13307 = \wishbone_bd_ram_mem3_reg[109][28]/P0001  & n13306 ;
  assign n13308 = n13241 & n13249 ;
  assign n13309 = n13293 & n13308 ;
  assign n13310 = \wishbone_bd_ram_mem3_reg[153][28]/P0001  & n13309 ;
  assign n13311 = ~n13307 & ~n13310 ;
  assign n13312 = n13303 & n13311 ;
  assign n13313 = n13297 & n13312 ;
  assign n13314 = n13281 & n13313 ;
  assign n13315 = n13246 & n13275 ;
  assign n13316 = n13248 & n13273 ;
  assign n13317 = n13315 & n13316 ;
  assign n13318 = \wishbone_bd_ram_mem3_reg[95][28]/P0001  & n13317 ;
  assign n13319 = n13231 & n13248 ;
  assign n13320 = n13304 & n13319 ;
  assign n13321 = \wishbone_bd_ram_mem3_reg[103][28]/P0001  & n13320 ;
  assign n13322 = ~n13318 & ~n13321 ;
  assign n13323 = n13241 & n13253 ;
  assign n13324 = n13247 & n13323 ;
  assign n13325 = \wishbone_bd_ram_mem3_reg[17][28]/P0001  & n13324 ;
  assign n13326 = n13238 & n13260 ;
  assign n13327 = n13316 & n13326 ;
  assign n13328 = \wishbone_bd_ram_mem3_reg[63][28]/P0001  & n13327 ;
  assign n13329 = ~n13325 & ~n13328 ;
  assign n13330 = n13322 & n13329 ;
  assign n13331 = n13233 & n13266 ;
  assign n13332 = n13308 & n13331 ;
  assign n13333 = \wishbone_bd_ram_mem3_reg[233][28]/P0001  & n13332 ;
  assign n13334 = n13246 & n13266 ;
  assign n13335 = n13316 & n13334 ;
  assign n13336 = \wishbone_bd_ram_mem3_reg[223][28]/P0001  & n13335 ;
  assign n13337 = ~n13333 & ~n13336 ;
  assign n13338 = n13231 & n13264 ;
  assign n13339 = n13276 & n13338 ;
  assign n13340 = \wishbone_bd_ram_mem3_reg[70][28]/P0001  & n13339 ;
  assign n13341 = n13265 & n13290 ;
  assign n13342 = \wishbone_bd_ram_mem3_reg[42][28]/P0001  & n13341 ;
  assign n13343 = ~n13340 & ~n13342 ;
  assign n13344 = n13337 & n13343 ;
  assign n13345 = n13330 & n13344 ;
  assign n13346 = n13230 & n13249 ;
  assign n13347 = n13315 & n13346 ;
  assign n13348 = \wishbone_bd_ram_mem3_reg[88][28]/P0001  & n13347 ;
  assign n13349 = n13316 & n13331 ;
  assign n13350 = \wishbone_bd_ram_mem3_reg[239][28]/P0001  & n13349 ;
  assign n13351 = ~n13348 & ~n13350 ;
  assign n13352 = n13259 & n13282 ;
  assign n13353 = \wishbone_bd_ram_mem3_reg[240][28]/P0001  & n13352 ;
  assign n13354 = n13240 & n13254 ;
  assign n13355 = \wishbone_bd_ram_mem3_reg[3][28]/P0001  & n13354 ;
  assign n13356 = ~n13353 & ~n13355 ;
  assign n13357 = n13351 & n13356 ;
  assign n13358 = n13254 & n13286 ;
  assign n13359 = \wishbone_bd_ram_mem3_reg[131][28]/P0001  & n13358 ;
  assign n13360 = n13235 & n13305 ;
  assign n13361 = \wishbone_bd_ram_mem3_reg[173][28]/P0001  & n13360 ;
  assign n13362 = ~n13359 & ~n13361 ;
  assign n13363 = n13319 & n13331 ;
  assign n13364 = \wishbone_bd_ram_mem3_reg[231][28]/P0001  & n13363 ;
  assign n13365 = n13261 & n13274 ;
  assign n13366 = \wishbone_bd_ram_mem3_reg[190][28]/P0001  & n13365 ;
  assign n13367 = ~n13364 & ~n13366 ;
  assign n13368 = n13362 & n13367 ;
  assign n13369 = n13357 & n13368 ;
  assign n13370 = n13345 & n13369 ;
  assign n13371 = n13314 & n13370 ;
  assign n13372 = n13261 & n13308 ;
  assign n13373 = \wishbone_bd_ram_mem3_reg[185][28]/P0001  & n13372 ;
  assign n13374 = n13300 & n13315 ;
  assign n13375 = \wishbone_bd_ram_mem3_reg[82][28]/P0001  & n13374 ;
  assign n13376 = ~n13373 & ~n13375 ;
  assign n13377 = n13235 & n13285 ;
  assign n13378 = \wishbone_bd_ram_mem3_reg[172][28]/P0001  & n13377 ;
  assign n13379 = n13232 & n13276 ;
  assign n13380 = \wishbone_bd_ram_mem3_reg[68][28]/P0001  & n13379 ;
  assign n13381 = ~n13378 & ~n13380 ;
  assign n13382 = n13376 & n13381 ;
  assign n13383 = n13282 & n13300 ;
  assign n13384 = \wishbone_bd_ram_mem3_reg[242][28]/P0001  & n13383 ;
  assign n13385 = n13232 & n13315 ;
  assign n13386 = \wishbone_bd_ram_mem3_reg[84][28]/P0001  & n13385 ;
  assign n13387 = ~n13384 & ~n13386 ;
  assign n13388 = n13254 & n13331 ;
  assign n13389 = \wishbone_bd_ram_mem3_reg[227][28]/P0001  & n13388 ;
  assign n13390 = n13259 & n13267 ;
  assign n13391 = \wishbone_bd_ram_mem3_reg[192][28]/P0001  & n13390 ;
  assign n13392 = ~n13389 & ~n13391 ;
  assign n13393 = n13387 & n13392 ;
  assign n13394 = n13382 & n13393 ;
  assign n13395 = n13260 & n13275 ;
  assign n13396 = n13305 & n13395 ;
  assign n13397 = \wishbone_bd_ram_mem3_reg[125][28]/P0001  & n13396 ;
  assign n13398 = n13265 & n13286 ;
  assign n13399 = \wishbone_bd_ram_mem3_reg[138][28]/P0001  & n13398 ;
  assign n13400 = ~n13397 & ~n13399 ;
  assign n13401 = n13232 & n13304 ;
  assign n13402 = \wishbone_bd_ram_mem3_reg[100][28]/P0001  & n13401 ;
  assign n13403 = n13265 & n13293 ;
  assign n13404 = \wishbone_bd_ram_mem3_reg[154][28]/P0001  & n13403 ;
  assign n13405 = ~n13402 & ~n13404 ;
  assign n13406 = n13400 & n13405 ;
  assign n13407 = n13261 & n13285 ;
  assign n13408 = \wishbone_bd_ram_mem3_reg[188][28]/P0001  & n13407 ;
  assign n13409 = n13315 & n13323 ;
  assign n13410 = \wishbone_bd_ram_mem3_reg[81][28]/P0001  & n13409 ;
  assign n13411 = ~n13408 & ~n13410 ;
  assign n13412 = n13247 & n13305 ;
  assign n13413 = \wishbone_bd_ram_mem3_reg[29][28]/P0001  & n13412 ;
  assign n13414 = n13267 & n13274 ;
  assign n13415 = \wishbone_bd_ram_mem3_reg[206][28]/P0001  & n13414 ;
  assign n13416 = ~n13413 & ~n13415 ;
  assign n13417 = n13411 & n13416 ;
  assign n13418 = n13406 & n13417 ;
  assign n13419 = n13394 & n13418 ;
  assign n13420 = n13290 & n13305 ;
  assign n13421 = \wishbone_bd_ram_mem3_reg[45][28]/P0001  & n13420 ;
  assign n13422 = n13235 & n13250 ;
  assign n13423 = \wishbone_bd_ram_mem3_reg[171][28]/P0001  & n13422 ;
  assign n13424 = ~n13421 & ~n13423 ;
  assign n13425 = n13259 & n13304 ;
  assign n13426 = \wishbone_bd_ram_mem3_reg[96][28]/P0001  & n13425 ;
  assign n13427 = n13286 & n13300 ;
  assign n13428 = \wishbone_bd_ram_mem3_reg[130][28]/P0001  & n13427 ;
  assign n13429 = ~n13426 & ~n13428 ;
  assign n13430 = n13424 & n13429 ;
  assign n13431 = n13282 & n13308 ;
  assign n13432 = \wishbone_bd_ram_mem3_reg[249][28]/P0001  & n13431 ;
  assign n13433 = n13259 & n13331 ;
  assign n13434 = \wishbone_bd_ram_mem3_reg[224][28]/P0001  & n13433 ;
  assign n13435 = ~n13432 & ~n13434 ;
  assign n13436 = n13290 & n13316 ;
  assign n13437 = \wishbone_bd_ram_mem3_reg[47][28]/P0001  & n13436 ;
  assign n13438 = n13242 & n13247 ;
  assign n13439 = \wishbone_bd_ram_mem3_reg[21][28]/P0001  & n13438 ;
  assign n13440 = ~n13437 & ~n13439 ;
  assign n13441 = n13435 & n13440 ;
  assign n13442 = n13430 & n13441 ;
  assign n13443 = n13300 & n13334 ;
  assign n13444 = \wishbone_bd_ram_mem3_reg[210][28]/P0001  & n13443 ;
  assign n13445 = n13293 & n13305 ;
  assign n13446 = \wishbone_bd_ram_mem3_reg[157][28]/P0001  & n13445 ;
  assign n13447 = ~n13444 & ~n13446 ;
  assign n13448 = n13274 & n13286 ;
  assign n13449 = \wishbone_bd_ram_mem3_reg[142][28]/P0001  & n13448 ;
  assign n13450 = n13290 & n13300 ;
  assign n13451 = \wishbone_bd_ram_mem3_reg[34][28]/P0001  & n13450 ;
  assign n13452 = ~n13449 & ~n13451 ;
  assign n13453 = n13447 & n13452 ;
  assign n13454 = n13254 & n13315 ;
  assign n13455 = \wishbone_bd_ram_mem3_reg[83][28]/P0001  & n13454 ;
  assign n13456 = n13276 & n13308 ;
  assign n13457 = \wishbone_bd_ram_mem3_reg[73][28]/P0001  & n13456 ;
  assign n13458 = ~n13455 & ~n13457 ;
  assign n13459 = n13240 & n13346 ;
  assign n13460 = \wishbone_bd_ram_mem3_reg[8][28]/P0001  & n13459 ;
  assign n13461 = n13286 & n13316 ;
  assign n13462 = \wishbone_bd_ram_mem3_reg[143][28]/P0001  & n13461 ;
  assign n13463 = ~n13460 & ~n13462 ;
  assign n13464 = n13458 & n13463 ;
  assign n13465 = n13453 & n13464 ;
  assign n13466 = n13442 & n13465 ;
  assign n13467 = n13419 & n13466 ;
  assign n13468 = n13371 & n13467 ;
  assign n13469 = n13242 & n13293 ;
  assign n13470 = \wishbone_bd_ram_mem3_reg[149][28]/P0001  & n13469 ;
  assign n13471 = n13304 & n13316 ;
  assign n13472 = \wishbone_bd_ram_mem3_reg[111][28]/P0001  & n13471 ;
  assign n13473 = ~n13470 & ~n13472 ;
  assign n13474 = n13232 & n13282 ;
  assign n13475 = \wishbone_bd_ram_mem3_reg[244][28]/P0001  & n13474 ;
  assign n13476 = n13250 & n13304 ;
  assign n13477 = \wishbone_bd_ram_mem3_reg[107][28]/P0001  & n13476 ;
  assign n13478 = ~n13475 & ~n13477 ;
  assign n13479 = n13473 & n13478 ;
  assign n13480 = n13285 & n13331 ;
  assign n13481 = \wishbone_bd_ram_mem3_reg[236][28]/P0001  & n13480 ;
  assign n13482 = n13259 & n13395 ;
  assign n13483 = \wishbone_bd_ram_mem3_reg[112][28]/P0001  & n13482 ;
  assign n13484 = ~n13481 & ~n13483 ;
  assign n13485 = n13315 & n13338 ;
  assign n13486 = \wishbone_bd_ram_mem3_reg[86][28]/P0001  & n13485 ;
  assign n13487 = n13242 & n13276 ;
  assign n13488 = \wishbone_bd_ram_mem3_reg[69][28]/P0001  & n13487 ;
  assign n13489 = ~n13486 & ~n13488 ;
  assign n13490 = n13484 & n13489 ;
  assign n13491 = n13479 & n13490 ;
  assign n13492 = n13242 & n13286 ;
  assign n13493 = \wishbone_bd_ram_mem3_reg[133][28]/P0001  & n13492 ;
  assign n13494 = n13286 & n13338 ;
  assign n13495 = \wishbone_bd_ram_mem3_reg[134][28]/P0001  & n13494 ;
  assign n13496 = ~n13493 & ~n13495 ;
  assign n13497 = n13232 & n13331 ;
  assign n13498 = \wishbone_bd_ram_mem3_reg[228][28]/P0001  & n13497 ;
  assign n13499 = n13267 & n13319 ;
  assign n13500 = \wishbone_bd_ram_mem3_reg[199][28]/P0001  & n13499 ;
  assign n13501 = ~n13498 & ~n13500 ;
  assign n13502 = n13496 & n13501 ;
  assign n13503 = n13304 & n13308 ;
  assign n13504 = \wishbone_bd_ram_mem3_reg[105][28]/P0001  & n13503 ;
  assign n13505 = n13235 & n13323 ;
  assign n13506 = \wishbone_bd_ram_mem3_reg[161][28]/P0001  & n13505 ;
  assign n13507 = ~n13504 & ~n13506 ;
  assign n13508 = n13259 & n13293 ;
  assign n13509 = \wishbone_bd_ram_mem3_reg[144][28]/P0001  & n13508 ;
  assign n13510 = n13331 & n13346 ;
  assign n13511 = \wishbone_bd_ram_mem3_reg[232][28]/P0001  & n13510 ;
  assign n13512 = ~n13509 & ~n13511 ;
  assign n13513 = n13507 & n13512 ;
  assign n13514 = n13502 & n13513 ;
  assign n13515 = n13491 & n13514 ;
  assign n13516 = n13259 & n13315 ;
  assign n13517 = \wishbone_bd_ram_mem3_reg[80][28]/P0001  & n13516 ;
  assign n13518 = n13250 & n13331 ;
  assign n13519 = \wishbone_bd_ram_mem3_reg[235][28]/P0001  & n13518 ;
  assign n13520 = ~n13517 & ~n13519 ;
  assign n13521 = n13247 & n13265 ;
  assign n13522 = \wishbone_bd_ram_mem3_reg[26][28]/P0001  & n13521 ;
  assign n13523 = n13254 & n13290 ;
  assign n13524 = \wishbone_bd_ram_mem3_reg[35][28]/P0001  & n13523 ;
  assign n13525 = ~n13522 & ~n13524 ;
  assign n13526 = n13520 & n13525 ;
  assign n13527 = n13232 & n13240 ;
  assign n13528 = \wishbone_bd_ram_mem3_reg[4][28]/P0001  & n13527 ;
  assign n13529 = n13274 & n13326 ;
  assign n13530 = \wishbone_bd_ram_mem3_reg[62][28]/P0001  & n13529 ;
  assign n13531 = ~n13528 & ~n13530 ;
  assign n13532 = n13247 & n13300 ;
  assign n13533 = \wishbone_bd_ram_mem3_reg[18][28]/P0001  & n13532 ;
  assign n13534 = n13304 & n13338 ;
  assign n13535 = \wishbone_bd_ram_mem3_reg[102][28]/P0001  & n13534 ;
  assign n13536 = ~n13533 & ~n13535 ;
  assign n13537 = n13531 & n13536 ;
  assign n13538 = n13526 & n13537 ;
  assign n13539 = n13240 & n13259 ;
  assign n13540 = \wishbone_bd_ram_mem3_reg[0][28]/P0001  & n13539 ;
  assign n13541 = n13235 & n13308 ;
  assign n13542 = \wishbone_bd_ram_mem3_reg[169][28]/P0001  & n13541 ;
  assign n13543 = ~n13540 & ~n13542 ;
  assign n13544 = n13305 & n13326 ;
  assign n13545 = \wishbone_bd_ram_mem3_reg[61][28]/P0001  & n13544 ;
  assign n13546 = n13240 & n13319 ;
  assign n13547 = \wishbone_bd_ram_mem3_reg[7][28]/P0001  & n13546 ;
  assign n13548 = ~n13545 & ~n13547 ;
  assign n13549 = n13543 & n13548 ;
  assign n13550 = n13346 & n13395 ;
  assign n13551 = \wishbone_bd_ram_mem3_reg[120][28]/P0001  & n13550 ;
  assign n13552 = n13242 & n13331 ;
  assign n13553 = \wishbone_bd_ram_mem3_reg[229][28]/P0001  & n13552 ;
  assign n13554 = ~n13551 & ~n13553 ;
  assign n13555 = n13265 & n13304 ;
  assign n13556 = \wishbone_bd_ram_mem3_reg[106][28]/P0001  & n13555 ;
  assign n13557 = n13242 & n13395 ;
  assign n13558 = \wishbone_bd_ram_mem3_reg[117][28]/P0001  & n13557 ;
  assign n13559 = ~n13556 & ~n13558 ;
  assign n13560 = n13554 & n13559 ;
  assign n13561 = n13549 & n13560 ;
  assign n13562 = n13538 & n13561 ;
  assign n13563 = n13515 & n13562 ;
  assign n13564 = n13265 & n13276 ;
  assign n13565 = \wishbone_bd_ram_mem3_reg[74][28]/P0001  & n13564 ;
  assign n13566 = n13250 & n13286 ;
  assign n13567 = \wishbone_bd_ram_mem3_reg[139][28]/P0001  & n13566 ;
  assign n13568 = ~n13565 & ~n13567 ;
  assign n13569 = n13300 & n13304 ;
  assign n13570 = \wishbone_bd_ram_mem3_reg[98][28]/P0001  & n13569 ;
  assign n13571 = n13282 & n13319 ;
  assign n13572 = \wishbone_bd_ram_mem3_reg[247][28]/P0001  & n13571 ;
  assign n13573 = ~n13570 & ~n13572 ;
  assign n13574 = n13568 & n13573 ;
  assign n13575 = n13254 & n13282 ;
  assign n13576 = \wishbone_bd_ram_mem3_reg[243][28]/P0001  & n13575 ;
  assign n13577 = n13250 & n13334 ;
  assign n13578 = \wishbone_bd_ram_mem3_reg[219][28]/P0001  & n13577 ;
  assign n13579 = ~n13576 & ~n13578 ;
  assign n13580 = n13240 & n13308 ;
  assign n13581 = \wishbone_bd_ram_mem3_reg[9][28]/P0001  & n13580 ;
  assign n13582 = n13276 & n13346 ;
  assign n13583 = \wishbone_bd_ram_mem3_reg[72][28]/P0001  & n13582 ;
  assign n13584 = ~n13581 & ~n13583 ;
  assign n13585 = n13579 & n13584 ;
  assign n13586 = n13574 & n13585 ;
  assign n13587 = n13242 & n13261 ;
  assign n13588 = \wishbone_bd_ram_mem3_reg[181][28]/P0001  & n13587 ;
  assign n13589 = n13338 & n13395 ;
  assign n13590 = \wishbone_bd_ram_mem3_reg[118][28]/P0001  & n13589 ;
  assign n13591 = ~n13588 & ~n13590 ;
  assign n13592 = n13267 & n13338 ;
  assign n13593 = \wishbone_bd_ram_mem3_reg[198][28]/P0001  & n13592 ;
  assign n13594 = n13242 & n13267 ;
  assign n13595 = \wishbone_bd_ram_mem3_reg[197][28]/P0001  & n13594 ;
  assign n13596 = ~n13593 & ~n13595 ;
  assign n13597 = n13591 & n13596 ;
  assign n13598 = n13261 & n13338 ;
  assign n13599 = \wishbone_bd_ram_mem3_reg[182][28]/P0001  & n13598 ;
  assign n13600 = n13267 & n13308 ;
  assign n13601 = \wishbone_bd_ram_mem3_reg[201][28]/P0001  & n13600 ;
  assign n13602 = ~n13599 & ~n13601 ;
  assign n13603 = n13276 & n13300 ;
  assign n13604 = \wishbone_bd_ram_mem3_reg[66][28]/P0001  & n13603 ;
  assign n13605 = n13250 & n13276 ;
  assign n13606 = \wishbone_bd_ram_mem3_reg[75][28]/P0001  & n13605 ;
  assign n13607 = ~n13604 & ~n13606 ;
  assign n13608 = n13602 & n13607 ;
  assign n13609 = n13597 & n13608 ;
  assign n13610 = n13586 & n13609 ;
  assign n13611 = n13326 & n13346 ;
  assign n13612 = \wishbone_bd_ram_mem3_reg[56][28]/P0001  & n13611 ;
  assign n13613 = n13250 & n13326 ;
  assign n13614 = \wishbone_bd_ram_mem3_reg[59][28]/P0001  & n13613 ;
  assign n13615 = ~n13612 & ~n13614 ;
  assign n13616 = n13261 & n13265 ;
  assign n13617 = \wishbone_bd_ram_mem3_reg[186][28]/P0001  & n13616 ;
  assign n13618 = n13319 & n13326 ;
  assign n13619 = \wishbone_bd_ram_mem3_reg[55][28]/P0001  & n13618 ;
  assign n13620 = ~n13617 & ~n13619 ;
  assign n13621 = n13615 & n13620 ;
  assign n13622 = n13326 & n13338 ;
  assign n13623 = \wishbone_bd_ram_mem3_reg[54][28]/P0001  & n13622 ;
  assign n13624 = n13267 & n13300 ;
  assign n13625 = \wishbone_bd_ram_mem3_reg[194][28]/P0001  & n13624 ;
  assign n13626 = ~n13623 & ~n13625 ;
  assign n13627 = n13293 & n13316 ;
  assign n13628 = \wishbone_bd_ram_mem3_reg[159][28]/P0001  & n13627 ;
  assign n13629 = n13286 & n13323 ;
  assign n13630 = \wishbone_bd_ram_mem3_reg[129][28]/P0001  & n13629 ;
  assign n13631 = ~n13628 & ~n13630 ;
  assign n13632 = n13626 & n13631 ;
  assign n13633 = n13621 & n13632 ;
  assign n13634 = n13232 & n13334 ;
  assign n13635 = \wishbone_bd_ram_mem3_reg[212][28]/P0001  & n13634 ;
  assign n13636 = n13276 & n13319 ;
  assign n13637 = \wishbone_bd_ram_mem3_reg[71][28]/P0001  & n13636 ;
  assign n13638 = ~n13635 & ~n13637 ;
  assign n13639 = n13232 & n13290 ;
  assign n13640 = \wishbone_bd_ram_mem3_reg[36][28]/P0001  & n13639 ;
  assign n13641 = n13305 & n13334 ;
  assign n13642 = \wishbone_bd_ram_mem3_reg[221][28]/P0001  & n13641 ;
  assign n13643 = ~n13640 & ~n13642 ;
  assign n13644 = n13638 & n13643 ;
  assign n13645 = n13261 & n13319 ;
  assign n13646 = \wishbone_bd_ram_mem3_reg[183][28]/P0001  & n13645 ;
  assign n13647 = n13282 & n13346 ;
  assign n13648 = \wishbone_bd_ram_mem3_reg[248][28]/P0001  & n13647 ;
  assign n13649 = ~n13646 & ~n13648 ;
  assign n13650 = n13232 & n13261 ;
  assign n13651 = \wishbone_bd_ram_mem3_reg[180][28]/P0001  & n13650 ;
  assign n13652 = n13259 & n13286 ;
  assign n13653 = \wishbone_bd_ram_mem3_reg[128][28]/P0001  & n13652 ;
  assign n13654 = ~n13651 & ~n13653 ;
  assign n13655 = n13649 & n13654 ;
  assign n13656 = n13644 & n13655 ;
  assign n13657 = n13633 & n13656 ;
  assign n13658 = n13610 & n13657 ;
  assign n13659 = n13563 & n13658 ;
  assign n13660 = n13468 & n13659 ;
  assign n13661 = n13290 & n13346 ;
  assign n13662 = \wishbone_bd_ram_mem3_reg[40][28]/P0001  & n13661 ;
  assign n13663 = n13254 & n13276 ;
  assign n13664 = \wishbone_bd_ram_mem3_reg[67][28]/P0001  & n13663 ;
  assign n13665 = ~n13662 & ~n13664 ;
  assign n13666 = n13293 & n13338 ;
  assign n13667 = \wishbone_bd_ram_mem3_reg[150][28]/P0001  & n13666 ;
  assign n13668 = n13300 & n13331 ;
  assign n13669 = \wishbone_bd_ram_mem3_reg[226][28]/P0001  & n13668 ;
  assign n13670 = ~n13667 & ~n13669 ;
  assign n13671 = n13665 & n13670 ;
  assign n13672 = n13286 & n13319 ;
  assign n13673 = \wishbone_bd_ram_mem3_reg[135][28]/P0001  & n13672 ;
  assign n13674 = n13235 & n13316 ;
  assign n13675 = \wishbone_bd_ram_mem3_reg[175][28]/P0001  & n13674 ;
  assign n13676 = ~n13673 & ~n13675 ;
  assign n13677 = n13265 & n13282 ;
  assign n13678 = \wishbone_bd_ram_mem3_reg[250][28]/P0001  & n13677 ;
  assign n13679 = n13265 & n13395 ;
  assign n13680 = \wishbone_bd_ram_mem3_reg[122][28]/P0001  & n13679 ;
  assign n13681 = ~n13678 & ~n13680 ;
  assign n13682 = n13676 & n13681 ;
  assign n13683 = n13671 & n13682 ;
  assign n13684 = n13304 & n13346 ;
  assign n13685 = \wishbone_bd_ram_mem3_reg[104][28]/P0001  & n13684 ;
  assign n13686 = n13300 & n13326 ;
  assign n13687 = \wishbone_bd_ram_mem3_reg[50][28]/P0001  & n13686 ;
  assign n13688 = ~n13685 & ~n13687 ;
  assign n13689 = n13323 & n13334 ;
  assign n13690 = \wishbone_bd_ram_mem3_reg[209][28]/P0001  & n13689 ;
  assign n13691 = n13315 & n13319 ;
  assign n13692 = \wishbone_bd_ram_mem3_reg[87][28]/P0001  & n13691 ;
  assign n13693 = ~n13690 & ~n13692 ;
  assign n13694 = n13688 & n13693 ;
  assign n13695 = n13247 & n13259 ;
  assign n13696 = \wishbone_bd_ram_mem3_reg[16][28]/P0001  & n13695 ;
  assign n13697 = n13293 & n13319 ;
  assign n13698 = \wishbone_bd_ram_mem3_reg[151][28]/P0001  & n13697 ;
  assign n13699 = ~n13696 & ~n13698 ;
  assign n13700 = n13254 & n13267 ;
  assign n13701 = \wishbone_bd_ram_mem3_reg[195][28]/P0001  & n13700 ;
  assign n13702 = n13254 & n13293 ;
  assign n13703 = \wishbone_bd_ram_mem3_reg[147][28]/P0001  & n13702 ;
  assign n13704 = ~n13701 & ~n13703 ;
  assign n13705 = n13699 & n13704 ;
  assign n13706 = n13694 & n13705 ;
  assign n13707 = n13683 & n13706 ;
  assign n13708 = n13282 & n13305 ;
  assign n13709 = \wishbone_bd_ram_mem3_reg[253][28]/P0001  & n13708 ;
  assign n13710 = n13242 & n13290 ;
  assign n13711 = \wishbone_bd_ram_mem3_reg[37][28]/P0001  & n13710 ;
  assign n13712 = ~n13709 & ~n13711 ;
  assign n13713 = n13247 & n13274 ;
  assign n13714 = \wishbone_bd_ram_mem3_reg[30][28]/P0001  & n13713 ;
  assign n13715 = n13293 & n13323 ;
  assign n13716 = \wishbone_bd_ram_mem3_reg[145][28]/P0001  & n13715 ;
  assign n13717 = ~n13714 & ~n13716 ;
  assign n13718 = n13712 & n13717 ;
  assign n13719 = n13323 & n13331 ;
  assign n13720 = \wishbone_bd_ram_mem3_reg[225][28]/P0001  & n13719 ;
  assign n13721 = n13274 & n13334 ;
  assign n13722 = \wishbone_bd_ram_mem3_reg[222][28]/P0001  & n13721 ;
  assign n13723 = ~n13720 & ~n13722 ;
  assign n13724 = n13304 & n13323 ;
  assign n13725 = \wishbone_bd_ram_mem3_reg[97][28]/P0001  & n13724 ;
  assign n13726 = n13235 & n13300 ;
  assign n13727 = \wishbone_bd_ram_mem3_reg[162][28]/P0001  & n13726 ;
  assign n13728 = ~n13725 & ~n13727 ;
  assign n13729 = n13723 & n13728 ;
  assign n13730 = n13718 & n13729 ;
  assign n13731 = n13308 & n13326 ;
  assign n13732 = \wishbone_bd_ram_mem3_reg[57][28]/P0001  & n13731 ;
  assign n13733 = n13240 & n13285 ;
  assign n13734 = \wishbone_bd_ram_mem3_reg[12][28]/P0001  & n13733 ;
  assign n13735 = ~n13732 & ~n13734 ;
  assign n13736 = n13259 & n13290 ;
  assign n13737 = \wishbone_bd_ram_mem3_reg[32][28]/P0001  & n13736 ;
  assign n13738 = n13250 & n13293 ;
  assign n13739 = \wishbone_bd_ram_mem3_reg[155][28]/P0001  & n13738 ;
  assign n13740 = ~n13737 & ~n13739 ;
  assign n13741 = n13735 & n13740 ;
  assign n13742 = n13247 & n13308 ;
  assign n13743 = \wishbone_bd_ram_mem3_reg[25][28]/P0001  & n13742 ;
  assign n13744 = n13247 & n13338 ;
  assign n13745 = \wishbone_bd_ram_mem3_reg[22][28]/P0001  & n13744 ;
  assign n13746 = ~n13743 & ~n13745 ;
  assign n13747 = n13254 & n13395 ;
  assign n13748 = \wishbone_bd_ram_mem3_reg[115][28]/P0001  & n13747 ;
  assign n13749 = n13250 & n13395 ;
  assign n13750 = \wishbone_bd_ram_mem3_reg[123][28]/P0001  & n13749 ;
  assign n13751 = ~n13748 & ~n13750 ;
  assign n13752 = n13746 & n13751 ;
  assign n13753 = n13741 & n13752 ;
  assign n13754 = n13730 & n13753 ;
  assign n13755 = n13707 & n13754 ;
  assign n13756 = n13250 & n13261 ;
  assign n13757 = \wishbone_bd_ram_mem3_reg[187][28]/P0001  & n13756 ;
  assign n13758 = n13247 & n13316 ;
  assign n13759 = \wishbone_bd_ram_mem3_reg[31][28]/P0001  & n13758 ;
  assign n13760 = ~n13757 & ~n13759 ;
  assign n13761 = n13250 & n13290 ;
  assign n13762 = \wishbone_bd_ram_mem3_reg[43][28]/P0001  & n13761 ;
  assign n13763 = n13300 & n13395 ;
  assign n13764 = \wishbone_bd_ram_mem3_reg[114][28]/P0001  & n13763 ;
  assign n13765 = ~n13762 & ~n13764 ;
  assign n13766 = n13760 & n13765 ;
  assign n13767 = n13308 & n13334 ;
  assign n13768 = \wishbone_bd_ram_mem3_reg[217][28]/P0001  & n13767 ;
  assign n13769 = n13285 & n13293 ;
  assign n13770 = \wishbone_bd_ram_mem3_reg[156][28]/P0001  & n13769 ;
  assign n13771 = ~n13768 & ~n13770 ;
  assign n13772 = n13242 & n13304 ;
  assign n13773 = \wishbone_bd_ram_mem3_reg[101][28]/P0001  & n13772 ;
  assign n13774 = n13240 & n13250 ;
  assign n13775 = \wishbone_bd_ram_mem3_reg[11][28]/P0001  & n13774 ;
  assign n13776 = ~n13773 & ~n13775 ;
  assign n13777 = n13771 & n13776 ;
  assign n13778 = n13766 & n13777 ;
  assign n13779 = n13276 & n13316 ;
  assign n13780 = \wishbone_bd_ram_mem3_reg[79][28]/P0001  & n13779 ;
  assign n13781 = n13265 & n13331 ;
  assign n13782 = \wishbone_bd_ram_mem3_reg[234][28]/P0001  & n13781 ;
  assign n13783 = ~n13780 & ~n13782 ;
  assign n13784 = n13242 & n13315 ;
  assign n13785 = \wishbone_bd_ram_mem3_reg[85][28]/P0001  & n13784 ;
  assign n13786 = n13274 & n13395 ;
  assign n13787 = \wishbone_bd_ram_mem3_reg[126][28]/P0001  & n13786 ;
  assign n13788 = ~n13785 & ~n13787 ;
  assign n13789 = n13783 & n13788 ;
  assign n13790 = n13285 & n13326 ;
  assign n13791 = \wishbone_bd_ram_mem3_reg[60][28]/P0001  & n13790 ;
  assign n13792 = n13265 & n13334 ;
  assign n13793 = \wishbone_bd_ram_mem3_reg[218][28]/P0001  & n13792 ;
  assign n13794 = ~n13791 & ~n13793 ;
  assign n13795 = n13235 & n13346 ;
  assign n13796 = \wishbone_bd_ram_mem3_reg[168][28]/P0001  & n13795 ;
  assign n13797 = n13240 & n13316 ;
  assign n13798 = \wishbone_bd_ram_mem3_reg[15][28]/P0001  & n13797 ;
  assign n13799 = ~n13796 & ~n13798 ;
  assign n13800 = n13794 & n13799 ;
  assign n13801 = n13789 & n13800 ;
  assign n13802 = n13778 & n13801 ;
  assign n13803 = n13316 & n13395 ;
  assign n13804 = \wishbone_bd_ram_mem3_reg[127][28]/P0001  & n13803 ;
  assign n13805 = n13254 & n13334 ;
  assign n13806 = \wishbone_bd_ram_mem3_reg[211][28]/P0001  & n13805 ;
  assign n13807 = ~n13804 & ~n13806 ;
  assign n13808 = n13286 & n13308 ;
  assign n13809 = \wishbone_bd_ram_mem3_reg[137][28]/P0001  & n13808 ;
  assign n13810 = n13247 & n13285 ;
  assign n13811 = \wishbone_bd_ram_mem3_reg[28][28]/P0001  & n13810 ;
  assign n13812 = ~n13809 & ~n13811 ;
  assign n13813 = n13807 & n13812 ;
  assign n13814 = n13285 & n13304 ;
  assign n13815 = \wishbone_bd_ram_mem3_reg[108][28]/P0001  & n13814 ;
  assign n13816 = n13250 & n13267 ;
  assign n13817 = \wishbone_bd_ram_mem3_reg[203][28]/P0001  & n13816 ;
  assign n13818 = ~n13815 & ~n13817 ;
  assign n13819 = n13274 & n13331 ;
  assign n13820 = \wishbone_bd_ram_mem3_reg[238][28]/P0001  & n13819 ;
  assign n13821 = n13267 & n13285 ;
  assign n13822 = \wishbone_bd_ram_mem3_reg[204][28]/P0001  & n13821 ;
  assign n13823 = ~n13820 & ~n13822 ;
  assign n13824 = n13818 & n13823 ;
  assign n13825 = n13813 & n13824 ;
  assign n13826 = n13267 & n13316 ;
  assign n13827 = \wishbone_bd_ram_mem3_reg[207][28]/P0001  & n13826 ;
  assign n13828 = n13290 & n13338 ;
  assign n13829 = \wishbone_bd_ram_mem3_reg[38][28]/P0001  & n13828 ;
  assign n13830 = ~n13827 & ~n13829 ;
  assign n13831 = n13276 & n13285 ;
  assign n13832 = \wishbone_bd_ram_mem3_reg[76][28]/P0001  & n13831 ;
  assign n13833 = n13274 & n13315 ;
  assign n13834 = \wishbone_bd_ram_mem3_reg[94][28]/P0001  & n13833 ;
  assign n13835 = ~n13832 & ~n13834 ;
  assign n13836 = n13830 & n13835 ;
  assign n13837 = n13240 & n13265 ;
  assign n13838 = \wishbone_bd_ram_mem3_reg[10][28]/P0001  & n13837 ;
  assign n13839 = n13232 & n13247 ;
  assign n13840 = \wishbone_bd_ram_mem3_reg[20][28]/P0001  & n13839 ;
  assign n13841 = ~n13838 & ~n13840 ;
  assign n13842 = n13276 & n13323 ;
  assign n13843 = \wishbone_bd_ram_mem3_reg[65][28]/P0001  & n13842 ;
  assign n13844 = n13240 & n13305 ;
  assign n13845 = \wishbone_bd_ram_mem3_reg[13][28]/P0001  & n13844 ;
  assign n13846 = ~n13843 & ~n13845 ;
  assign n13847 = n13841 & n13846 ;
  assign n13848 = n13836 & n13847 ;
  assign n13849 = n13825 & n13848 ;
  assign n13850 = n13802 & n13849 ;
  assign n13851 = n13755 & n13850 ;
  assign n13852 = n13286 & n13305 ;
  assign n13853 = \wishbone_bd_ram_mem3_reg[141][28]/P0001  & n13852 ;
  assign n13854 = n13282 & n13323 ;
  assign n13855 = \wishbone_bd_ram_mem3_reg[241][28]/P0001  & n13854 ;
  assign n13856 = ~n13853 & ~n13855 ;
  assign n13857 = n13247 & n13319 ;
  assign n13858 = \wishbone_bd_ram_mem3_reg[23][28]/P0001  & n13857 ;
  assign n13859 = n13285 & n13315 ;
  assign n13860 = \wishbone_bd_ram_mem3_reg[92][28]/P0001  & n13859 ;
  assign n13861 = ~n13858 & ~n13860 ;
  assign n13862 = n13856 & n13861 ;
  assign n13863 = n13261 & n13323 ;
  assign n13864 = \wishbone_bd_ram_mem3_reg[177][28]/P0001  & n13863 ;
  assign n13865 = n13232 & n13395 ;
  assign n13866 = \wishbone_bd_ram_mem3_reg[116][28]/P0001  & n13865 ;
  assign n13867 = ~n13864 & ~n13866 ;
  assign n13868 = n13232 & n13293 ;
  assign n13869 = \wishbone_bd_ram_mem3_reg[148][28]/P0001  & n13868 ;
  assign n13870 = n13242 & n13334 ;
  assign n13871 = \wishbone_bd_ram_mem3_reg[213][28]/P0001  & n13870 ;
  assign n13872 = ~n13869 & ~n13871 ;
  assign n13873 = n13867 & n13872 ;
  assign n13874 = n13862 & n13873 ;
  assign n13875 = n13242 & n13326 ;
  assign n13876 = \wishbone_bd_ram_mem3_reg[53][28]/P0001  & n13875 ;
  assign n13877 = n13242 & n13282 ;
  assign n13878 = \wishbone_bd_ram_mem3_reg[245][28]/P0001  & n13877 ;
  assign n13879 = ~n13876 & ~n13878 ;
  assign n13880 = n13254 & n13326 ;
  assign n13881 = \wishbone_bd_ram_mem3_reg[51][28]/P0001  & n13880 ;
  assign n13882 = n13323 & n13395 ;
  assign n13883 = \wishbone_bd_ram_mem3_reg[113][28]/P0001  & n13882 ;
  assign n13884 = ~n13881 & ~n13883 ;
  assign n13885 = n13879 & n13884 ;
  assign n13886 = n13247 & n13254 ;
  assign n13887 = \wishbone_bd_ram_mem3_reg[19][28]/P0001  & n13886 ;
  assign n13888 = n13240 & n13323 ;
  assign n13889 = \wishbone_bd_ram_mem3_reg[1][28]/P0001  & n13888 ;
  assign n13890 = ~n13887 & ~n13889 ;
  assign n13891 = n13305 & n13315 ;
  assign n13892 = \wishbone_bd_ram_mem3_reg[93][28]/P0001  & n13891 ;
  assign n13893 = n13290 & n13319 ;
  assign n13894 = \wishbone_bd_ram_mem3_reg[39][28]/P0001  & n13893 ;
  assign n13895 = ~n13892 & ~n13894 ;
  assign n13896 = n13890 & n13895 ;
  assign n13897 = n13885 & n13896 ;
  assign n13898 = n13874 & n13897 ;
  assign n13899 = n13235 & n13274 ;
  assign n13900 = \wishbone_bd_ram_mem3_reg[174][28]/P0001  & n13899 ;
  assign n13901 = n13319 & n13334 ;
  assign n13902 = \wishbone_bd_ram_mem3_reg[215][28]/P0001  & n13901 ;
  assign n13903 = ~n13900 & ~n13902 ;
  assign n13904 = n13259 & n13276 ;
  assign n13905 = \wishbone_bd_ram_mem3_reg[64][28]/P0001  & n13904 ;
  assign n13906 = n13265 & n13315 ;
  assign n13907 = \wishbone_bd_ram_mem3_reg[90][28]/P0001  & n13906 ;
  assign n13908 = ~n13905 & ~n13907 ;
  assign n13909 = n13903 & n13908 ;
  assign n13910 = n13308 & n13315 ;
  assign n13911 = \wishbone_bd_ram_mem3_reg[89][28]/P0001  & n13910 ;
  assign n13912 = n13293 & n13346 ;
  assign n13913 = \wishbone_bd_ram_mem3_reg[152][28]/P0001  & n13912 ;
  assign n13914 = ~n13911 & ~n13913 ;
  assign n13915 = n13240 & n13338 ;
  assign n13916 = \wishbone_bd_ram_mem3_reg[6][28]/P0001  & n13915 ;
  assign n13917 = n13259 & n13326 ;
  assign n13918 = \wishbone_bd_ram_mem3_reg[48][28]/P0001  & n13917 ;
  assign n13919 = ~n13916 & ~n13918 ;
  assign n13920 = n13914 & n13919 ;
  assign n13921 = n13909 & n13920 ;
  assign n13922 = n13267 & n13346 ;
  assign n13923 = \wishbone_bd_ram_mem3_reg[200][28]/P0001  & n13922 ;
  assign n13924 = n13305 & n13331 ;
  assign n13925 = \wishbone_bd_ram_mem3_reg[237][28]/P0001  & n13924 ;
  assign n13926 = ~n13923 & ~n13925 ;
  assign n13927 = n13232 & n13286 ;
  assign n13928 = \wishbone_bd_ram_mem3_reg[132][28]/P0001  & n13927 ;
  assign n13929 = n13323 & n13326 ;
  assign n13930 = \wishbone_bd_ram_mem3_reg[49][28]/P0001  & n13929 ;
  assign n13931 = ~n13928 & ~n13930 ;
  assign n13932 = n13926 & n13931 ;
  assign n13933 = n13290 & n13323 ;
  assign n13934 = \wishbone_bd_ram_mem3_reg[33][28]/P0001  & n13933 ;
  assign n13935 = n13276 & n13305 ;
  assign n13936 = \wishbone_bd_ram_mem3_reg[77][28]/P0001  & n13935 ;
  assign n13937 = ~n13934 & ~n13936 ;
  assign n13938 = n13334 & n13338 ;
  assign n13939 = \wishbone_bd_ram_mem3_reg[214][28]/P0001  & n13938 ;
  assign n13940 = n13235 & n13319 ;
  assign n13941 = \wishbone_bd_ram_mem3_reg[167][28]/P0001  & n13940 ;
  assign n13942 = ~n13939 & ~n13941 ;
  assign n13943 = n13937 & n13942 ;
  assign n13944 = n13932 & n13943 ;
  assign n13945 = n13921 & n13944 ;
  assign n13946 = n13898 & n13945 ;
  assign n13947 = n13267 & n13305 ;
  assign n13948 = \wishbone_bd_ram_mem3_reg[205][28]/P0001  & n13947 ;
  assign n13949 = n13265 & n13326 ;
  assign n13950 = \wishbone_bd_ram_mem3_reg[58][28]/P0001  & n13949 ;
  assign n13951 = ~n13948 & ~n13950 ;
  assign n13952 = n13282 & n13316 ;
  assign n13953 = \wishbone_bd_ram_mem3_reg[255][28]/P0001  & n13952 ;
  assign n13954 = n13250 & n13315 ;
  assign n13955 = \wishbone_bd_ram_mem3_reg[91][28]/P0001  & n13954 ;
  assign n13956 = ~n13953 & ~n13955 ;
  assign n13957 = n13951 & n13956 ;
  assign n13958 = n13293 & n13300 ;
  assign n13959 = \wishbone_bd_ram_mem3_reg[146][28]/P0001  & n13958 ;
  assign n13960 = n13261 & n13346 ;
  assign n13961 = \wishbone_bd_ram_mem3_reg[184][28]/P0001  & n13960 ;
  assign n13962 = ~n13959 & ~n13961 ;
  assign n13963 = n13286 & n13346 ;
  assign n13964 = \wishbone_bd_ram_mem3_reg[136][28]/P0001  & n13963 ;
  assign n13965 = n13285 & n13334 ;
  assign n13966 = \wishbone_bd_ram_mem3_reg[220][28]/P0001  & n13965 ;
  assign n13967 = ~n13964 & ~n13966 ;
  assign n13968 = n13962 & n13967 ;
  assign n13969 = n13957 & n13968 ;
  assign n13970 = n13247 & n13346 ;
  assign n13971 = \wishbone_bd_ram_mem3_reg[24][28]/P0001  & n13970 ;
  assign n13972 = n13240 & n13274 ;
  assign n13973 = \wishbone_bd_ram_mem3_reg[14][28]/P0001  & n13972 ;
  assign n13974 = ~n13971 & ~n13973 ;
  assign n13975 = n13240 & n13300 ;
  assign n13976 = \wishbone_bd_ram_mem3_reg[2][28]/P0001  & n13975 ;
  assign n13977 = n13232 & n13267 ;
  assign n13978 = \wishbone_bd_ram_mem3_reg[196][28]/P0001  & n13977 ;
  assign n13979 = ~n13976 & ~n13978 ;
  assign n13980 = n13974 & n13979 ;
  assign n13981 = n13282 & n13338 ;
  assign n13982 = \wishbone_bd_ram_mem3_reg[246][28]/P0001  & n13981 ;
  assign n13983 = n13308 & n13395 ;
  assign n13984 = \wishbone_bd_ram_mem3_reg[121][28]/P0001  & n13983 ;
  assign n13985 = ~n13982 & ~n13984 ;
  assign n13986 = n13282 & n13285 ;
  assign n13987 = \wishbone_bd_ram_mem3_reg[252][28]/P0001  & n13986 ;
  assign n13988 = n13232 & n13326 ;
  assign n13989 = \wishbone_bd_ram_mem3_reg[52][28]/P0001  & n13988 ;
  assign n13990 = ~n13987 & ~n13989 ;
  assign n13991 = n13985 & n13990 ;
  assign n13992 = n13980 & n13991 ;
  assign n13993 = n13969 & n13992 ;
  assign n13994 = n13331 & n13338 ;
  assign n13995 = \wishbone_bd_ram_mem3_reg[230][28]/P0001  & n13994 ;
  assign n13996 = n13254 & n13304 ;
  assign n13997 = \wishbone_bd_ram_mem3_reg[99][28]/P0001  & n13996 ;
  assign n13998 = ~n13995 & ~n13997 ;
  assign n13999 = n13235 & n13338 ;
  assign n14000 = \wishbone_bd_ram_mem3_reg[166][28]/P0001  & n13999 ;
  assign n14001 = n13261 & n13305 ;
  assign n14002 = \wishbone_bd_ram_mem3_reg[189][28]/P0001  & n14001 ;
  assign n14003 = ~n14000 & ~n14002 ;
  assign n14004 = n13998 & n14003 ;
  assign n14005 = n13334 & n13346 ;
  assign n14006 = \wishbone_bd_ram_mem3_reg[216][28]/P0001  & n14005 ;
  assign n14007 = n13235 & n13265 ;
  assign n14008 = \wishbone_bd_ram_mem3_reg[170][28]/P0001  & n14007 ;
  assign n14009 = ~n14006 & ~n14008 ;
  assign n14010 = n13259 & n13334 ;
  assign n14011 = \wishbone_bd_ram_mem3_reg[208][28]/P0001  & n14010 ;
  assign n14012 = n13261 & n13316 ;
  assign n14013 = \wishbone_bd_ram_mem3_reg[191][28]/P0001  & n14012 ;
  assign n14014 = ~n14011 & ~n14013 ;
  assign n14015 = n14009 & n14014 ;
  assign n14016 = n14004 & n14015 ;
  assign n14017 = n13290 & n13308 ;
  assign n14018 = \wishbone_bd_ram_mem3_reg[41][28]/P0001  & n14017 ;
  assign n14019 = n13250 & n13282 ;
  assign n14020 = \wishbone_bd_ram_mem3_reg[251][28]/P0001  & n14019 ;
  assign n14021 = ~n14018 & ~n14020 ;
  assign n14022 = n13267 & n13323 ;
  assign n14023 = \wishbone_bd_ram_mem3_reg[193][28]/P0001  & n14022 ;
  assign n14024 = n13285 & n13395 ;
  assign n14025 = \wishbone_bd_ram_mem3_reg[124][28]/P0001  & n14024 ;
  assign n14026 = ~n14023 & ~n14025 ;
  assign n14027 = n14021 & n14026 ;
  assign n14028 = n13235 & n13242 ;
  assign n14029 = \wishbone_bd_ram_mem3_reg[165][28]/P0001  & n14028 ;
  assign n14030 = n13274 & n13304 ;
  assign n14031 = \wishbone_bd_ram_mem3_reg[110][28]/P0001  & n14030 ;
  assign n14032 = ~n14029 & ~n14031 ;
  assign n14033 = n13319 & n13395 ;
  assign n14034 = \wishbone_bd_ram_mem3_reg[119][28]/P0001  & n14033 ;
  assign n14035 = n13254 & n13261 ;
  assign n14036 = \wishbone_bd_ram_mem3_reg[179][28]/P0001  & n14035 ;
  assign n14037 = ~n14034 & ~n14036 ;
  assign n14038 = n14032 & n14037 ;
  assign n14039 = n14027 & n14038 ;
  assign n14040 = n14016 & n14039 ;
  assign n14041 = n13993 & n14040 ;
  assign n14042 = n13946 & n14041 ;
  assign n14043 = n13851 & n14042 ;
  assign n14044 = n13660 & n14043 ;
  assign n14045 = \wishbone_TxEn_q_reg/NET0131  & \wishbone_TxEn_reg/NET0131  ;
  assign n14046 = \wishbone_TxBDRead_reg/NET0131  & n14045 ;
  assign n14047 = ~wb_rst_i_pad & n14046 ;
  assign n14048 = ~n14044 & n14047 ;
  assign n14049 = m_wb_ack_i_pad & \wishbone_MasterWbTX_reg/NET0131  ;
  assign n14050 = \wishbone_TxLength_reg[12]/NET0131  & ~n14049 ;
  assign n14051 = ~n14046 & n14050 ;
  assign n14052 = ~\wishbone_TxLength_reg[7]/NET0131  & ~\wishbone_TxLength_reg[8]/NET0131  ;
  assign n14053 = ~\wishbone_TxLength_reg[9]/NET0131  & n14052 ;
  assign n14054 = ~\wishbone_TxLength_reg[2]/NET0131  & ~\wishbone_TxLength_reg[3]/NET0131  ;
  assign n14055 = ~\wishbone_TxLength_reg[4]/NET0131  & n14054 ;
  assign n14056 = ~\wishbone_TxLength_reg[5]/NET0131  & ~\wishbone_TxLength_reg[6]/NET0131  ;
  assign n14057 = n14055 & n14056 ;
  assign n14058 = n14053 & n14057 ;
  assign n14059 = ~\wishbone_TxLength_reg[10]/NET0131  & ~\wishbone_TxLength_reg[11]/NET0131  ;
  assign n14060 = ~\wishbone_TxLength_reg[14]/NET0131  & n14059 ;
  assign n14061 = ~\wishbone_TxLength_reg[12]/NET0131  & ~\wishbone_TxLength_reg[13]/NET0131  ;
  assign n14062 = ~\wishbone_TxLength_reg[15]/NET0131  & n14061 ;
  assign n14063 = n14060 & n14062 ;
  assign n14064 = n14058 & n14063 ;
  assign n14065 = ~n14046 & n14049 ;
  assign n14066 = ~n14064 & n14065 ;
  assign n14067 = ~n14051 & ~n14066 ;
  assign n14068 = \wishbone_TxLength_reg[0]/NET0131  & \wishbone_TxPointerLSB_rst_reg[0]/NET0131  ;
  assign n14069 = ~\wishbone_TxLength_reg[1]/NET0131  & ~n14068 ;
  assign n14070 = \wishbone_TxLength_reg[1]/NET0131  & n14068 ;
  assign n14071 = ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  & ~n14070 ;
  assign n14072 = ~n14069 & ~n14071 ;
  assign n14073 = n14053 & n14059 ;
  assign n14074 = n14057 & n14073 ;
  assign n14075 = ~n14072 & n14074 ;
  assign n14076 = ~\wishbone_TxLength_reg[12]/NET0131  & ~n14051 ;
  assign n14077 = ~n14075 & n14076 ;
  assign n14078 = \wishbone_TxLength_reg[12]/NET0131  & ~n14051 ;
  assign n14079 = n14075 & n14078 ;
  assign n14080 = ~n14077 & ~n14079 ;
  assign n14081 = ~n14067 & n14080 ;
  assign n14082 = ~n14048 & ~n14081 ;
  assign n14083 = \wishbone_bd_ram_mem3_reg[77][29]/P0001  & n13935 ;
  assign n14084 = \wishbone_bd_ram_mem3_reg[42][29]/P0001  & n13341 ;
  assign n14085 = ~n14083 & ~n14084 ;
  assign n14086 = \wishbone_bd_ram_mem3_reg[65][29]/P0001  & n13842 ;
  assign n14087 = \wishbone_bd_ram_mem3_reg[70][29]/P0001  & n13339 ;
  assign n14088 = ~n14086 & ~n14087 ;
  assign n14089 = n14085 & n14088 ;
  assign n14090 = \wishbone_bd_ram_mem3_reg[202][29]/P0001  & n13268 ;
  assign n14091 = \wishbone_bd_ram_mem3_reg[111][29]/P0001  & n13471 ;
  assign n14092 = ~n14090 & ~n14091 ;
  assign n14093 = \wishbone_bd_ram_mem3_reg[160][29]/P0001  & n13271 ;
  assign n14094 = \wishbone_bd_ram_mem3_reg[127][29]/P0001  & n13803 ;
  assign n14095 = ~n14093 & ~n14094 ;
  assign n14096 = n14092 & n14095 ;
  assign n14097 = n14089 & n14096 ;
  assign n14098 = \wishbone_bd_ram_mem3_reg[71][29]/P0001  & n13636 ;
  assign n14099 = \wishbone_bd_ram_mem3_reg[113][29]/P0001  & n13882 ;
  assign n14100 = ~n14098 & ~n14099 ;
  assign n14101 = \wishbone_bd_ram_mem3_reg[86][29]/P0001  & n13485 ;
  assign n14102 = \wishbone_bd_ram_mem3_reg[158][29]/P0001  & n13294 ;
  assign n14103 = ~n14101 & ~n14102 ;
  assign n14104 = n14100 & n14103 ;
  assign n14105 = \wishbone_bd_ram_mem3_reg[46][29]/P0001  & n13298 ;
  assign n14106 = \wishbone_bd_ram_mem3_reg[112][29]/P0001  & n13482 ;
  assign n14107 = ~n14105 & ~n14106 ;
  assign n14108 = \wishbone_bd_ram_mem3_reg[36][29]/P0001  & n13639 ;
  assign n14109 = \wishbone_bd_ram_mem3_reg[90][29]/P0001  & n13906 ;
  assign n14110 = ~n14108 & ~n14109 ;
  assign n14111 = n14107 & n14110 ;
  assign n14112 = n14104 & n14111 ;
  assign n14113 = n14097 & n14112 ;
  assign n14114 = \wishbone_bd_ram_mem3_reg[125][29]/P0001  & n13396 ;
  assign n14115 = \wishbone_bd_ram_mem3_reg[121][29]/P0001  & n13983 ;
  assign n14116 = ~n14114 & ~n14115 ;
  assign n14117 = \wishbone_bd_ram_mem3_reg[4][29]/P0001  & n13527 ;
  assign n14118 = \wishbone_bd_ram_mem3_reg[81][29]/P0001  & n13409 ;
  assign n14119 = ~n14117 & ~n14118 ;
  assign n14120 = n14116 & n14119 ;
  assign n14121 = \wishbone_bd_ram_mem3_reg[233][29]/P0001  & n13332 ;
  assign n14122 = \wishbone_bd_ram_mem3_reg[191][29]/P0001  & n14012 ;
  assign n14123 = ~n14121 & ~n14122 ;
  assign n14124 = \wishbone_bd_ram_mem3_reg[83][29]/P0001  & n13454 ;
  assign n14125 = \wishbone_bd_ram_mem3_reg[27][29]/P0001  & n13251 ;
  assign n14126 = ~n14124 & ~n14125 ;
  assign n14127 = n14123 & n14126 ;
  assign n14128 = n14120 & n14127 ;
  assign n14129 = \wishbone_bd_ram_mem3_reg[104][29]/P0001  & n13684 ;
  assign n14130 = \wishbone_bd_ram_mem3_reg[201][29]/P0001  & n13600 ;
  assign n14131 = ~n14129 & ~n14130 ;
  assign n14132 = \wishbone_bd_ram_mem3_reg[75][29]/P0001  & n13605 ;
  assign n14133 = \wishbone_bd_ram_mem3_reg[2][29]/P0001  & n13975 ;
  assign n14134 = ~n14132 & ~n14133 ;
  assign n14135 = n14131 & n14134 ;
  assign n14136 = \wishbone_bd_ram_mem3_reg[67][29]/P0001  & n13663 ;
  assign n14137 = \wishbone_bd_ram_mem3_reg[106][29]/P0001  & n13555 ;
  assign n14138 = ~n14136 & ~n14137 ;
  assign n14139 = \wishbone_bd_ram_mem3_reg[174][29]/P0001  & n13899 ;
  assign n14140 = \wishbone_bd_ram_mem3_reg[181][29]/P0001  & n13587 ;
  assign n14141 = ~n14139 & ~n14140 ;
  assign n14142 = n14138 & n14141 ;
  assign n14143 = n14135 & n14142 ;
  assign n14144 = n14128 & n14143 ;
  assign n14145 = n14113 & n14144 ;
  assign n14146 = \wishbone_bd_ram_mem3_reg[224][29]/P0001  & n13433 ;
  assign n14147 = \wishbone_bd_ram_mem3_reg[188][29]/P0001  & n13407 ;
  assign n14148 = ~n14146 & ~n14147 ;
  assign n14149 = \wishbone_bd_ram_mem3_reg[105][29]/P0001  & n13503 ;
  assign n14150 = \wishbone_bd_ram_mem3_reg[58][29]/P0001  & n13949 ;
  assign n14151 = ~n14149 & ~n14150 ;
  assign n14152 = n14148 & n14151 ;
  assign n14153 = \wishbone_bd_ram_mem3_reg[199][29]/P0001  & n13499 ;
  assign n14154 = \wishbone_bd_ram_mem3_reg[49][29]/P0001  & n13929 ;
  assign n14155 = ~n14153 & ~n14154 ;
  assign n14156 = \wishbone_bd_ram_mem3_reg[250][29]/P0001  & n13677 ;
  assign n14157 = \wishbone_bd_ram_mem3_reg[126][29]/P0001  & n13786 ;
  assign n14158 = ~n14156 & ~n14157 ;
  assign n14159 = n14155 & n14158 ;
  assign n14160 = n14152 & n14159 ;
  assign n14161 = \wishbone_bd_ram_mem3_reg[143][29]/P0001  & n13461 ;
  assign n14162 = \wishbone_bd_ram_mem3_reg[147][29]/P0001  & n13702 ;
  assign n14163 = ~n14161 & ~n14162 ;
  assign n14164 = \wishbone_bd_ram_mem3_reg[100][29]/P0001  & n13401 ;
  assign n14165 = \wishbone_bd_ram_mem3_reg[94][29]/P0001  & n13833 ;
  assign n14166 = ~n14164 & ~n14165 ;
  assign n14167 = n14163 & n14166 ;
  assign n14168 = \wishbone_bd_ram_mem3_reg[193][29]/P0001  & n14022 ;
  assign n14169 = \wishbone_bd_ram_mem3_reg[178][29]/P0001  & n13301 ;
  assign n14170 = ~n14168 & ~n14169 ;
  assign n14171 = \wishbone_bd_ram_mem3_reg[47][29]/P0001  & n13436 ;
  assign n14172 = \wishbone_bd_ram_mem3_reg[225][29]/P0001  & n13719 ;
  assign n14173 = ~n14171 & ~n14172 ;
  assign n14174 = n14170 & n14173 ;
  assign n14175 = n14167 & n14174 ;
  assign n14176 = n14160 & n14175 ;
  assign n14177 = \wishbone_bd_ram_mem3_reg[123][29]/P0001  & n13749 ;
  assign n14178 = \wishbone_bd_ram_mem3_reg[192][29]/P0001  & n13390 ;
  assign n14179 = ~n14177 & ~n14178 ;
  assign n14180 = \wishbone_bd_ram_mem3_reg[173][29]/P0001  & n13360 ;
  assign n14181 = \wishbone_bd_ram_mem3_reg[120][29]/P0001  & n13550 ;
  assign n14182 = ~n14180 & ~n14181 ;
  assign n14183 = n14179 & n14182 ;
  assign n14184 = \wishbone_bd_ram_mem3_reg[253][29]/P0001  & n13708 ;
  assign n14185 = \wishbone_bd_ram_mem3_reg[243][29]/P0001  & n13575 ;
  assign n14186 = ~n14184 & ~n14185 ;
  assign n14187 = \wishbone_bd_ram_mem3_reg[57][29]/P0001  & n13731 ;
  assign n14188 = \wishbone_bd_ram_mem3_reg[44][29]/P0001  & n13291 ;
  assign n14189 = ~n14187 & ~n14188 ;
  assign n14190 = n14186 & n14189 ;
  assign n14191 = n14183 & n14190 ;
  assign n14192 = \wishbone_bd_ram_mem3_reg[210][29]/P0001  & n13443 ;
  assign n14193 = \wishbone_bd_ram_mem3_reg[85][29]/P0001  & n13784 ;
  assign n14194 = ~n14192 & ~n14193 ;
  assign n14195 = \wishbone_bd_ram_mem3_reg[134][29]/P0001  & n13494 ;
  assign n14196 = \wishbone_bd_ram_mem3_reg[95][29]/P0001  & n13317 ;
  assign n14197 = ~n14195 & ~n14196 ;
  assign n14198 = n14194 & n14197 ;
  assign n14199 = \wishbone_bd_ram_mem3_reg[48][29]/P0001  & n13917 ;
  assign n14200 = \wishbone_bd_ram_mem3_reg[35][29]/P0001  & n13523 ;
  assign n14201 = ~n14199 & ~n14200 ;
  assign n14202 = \wishbone_bd_ram_mem3_reg[24][29]/P0001  & n13970 ;
  assign n14203 = \wishbone_bd_ram_mem3_reg[231][29]/P0001  & n13363 ;
  assign n14204 = ~n14202 & ~n14203 ;
  assign n14205 = n14201 & n14204 ;
  assign n14206 = n14198 & n14205 ;
  assign n14207 = n14191 & n14206 ;
  assign n14208 = n14176 & n14207 ;
  assign n14209 = n14145 & n14208 ;
  assign n14210 = \wishbone_bd_ram_mem3_reg[80][29]/P0001  & n13516 ;
  assign n14211 = \wishbone_bd_ram_mem3_reg[91][29]/P0001  & n13954 ;
  assign n14212 = ~n14210 & ~n14211 ;
  assign n14213 = \wishbone_bd_ram_mem3_reg[212][29]/P0001  & n13634 ;
  assign n14214 = \wishbone_bd_ram_mem3_reg[107][29]/P0001  & n13476 ;
  assign n14215 = ~n14213 & ~n14214 ;
  assign n14216 = n14212 & n14215 ;
  assign n14217 = \wishbone_bd_ram_mem3_reg[247][29]/P0001  & n13571 ;
  assign n14218 = \wishbone_bd_ram_mem3_reg[222][29]/P0001  & n13721 ;
  assign n14219 = ~n14217 & ~n14218 ;
  assign n14220 = \wishbone_bd_ram_mem3_reg[34][29]/P0001  & n13450 ;
  assign n14221 = \wishbone_bd_ram_mem3_reg[17][29]/P0001  & n13324 ;
  assign n14222 = ~n14220 & ~n14221 ;
  assign n14223 = n14219 & n14222 ;
  assign n14224 = n14216 & n14223 ;
  assign n14225 = \wishbone_bd_ram_mem3_reg[139][29]/P0001  & n13566 ;
  assign n14226 = \wishbone_bd_ram_mem3_reg[142][29]/P0001  & n13448 ;
  assign n14227 = ~n14225 & ~n14226 ;
  assign n14228 = \wishbone_bd_ram_mem3_reg[198][29]/P0001  & n13592 ;
  assign n14229 = \wishbone_bd_ram_mem3_reg[244][29]/P0001  & n13474 ;
  assign n14230 = ~n14228 & ~n14229 ;
  assign n14231 = n14227 & n14230 ;
  assign n14232 = \wishbone_bd_ram_mem3_reg[169][29]/P0001  & n13541 ;
  assign n14233 = \wishbone_bd_ram_mem3_reg[149][29]/P0001  & n13469 ;
  assign n14234 = ~n14232 & ~n14233 ;
  assign n14235 = \wishbone_bd_ram_mem3_reg[182][29]/P0001  & n13598 ;
  assign n14236 = \wishbone_bd_ram_mem3_reg[154][29]/P0001  & n13403 ;
  assign n14237 = ~n14235 & ~n14236 ;
  assign n14238 = n14234 & n14237 ;
  assign n14239 = n14231 & n14238 ;
  assign n14240 = n14224 & n14239 ;
  assign n14241 = \wishbone_bd_ram_mem3_reg[144][29]/P0001  & n13508 ;
  assign n14242 = \wishbone_bd_ram_mem3_reg[61][29]/P0001  & n13544 ;
  assign n14243 = ~n14241 & ~n14242 ;
  assign n14244 = \wishbone_bd_ram_mem3_reg[135][29]/P0001  & n13672 ;
  assign n14245 = \wishbone_bd_ram_mem3_reg[66][29]/P0001  & n13603 ;
  assign n14246 = ~n14244 & ~n14245 ;
  assign n14247 = n14243 & n14246 ;
  assign n14248 = \wishbone_bd_ram_mem3_reg[175][29]/P0001  & n13674 ;
  assign n14249 = \wishbone_bd_ram_mem3_reg[141][29]/P0001  & n13852 ;
  assign n14250 = ~n14248 & ~n14249 ;
  assign n14251 = \wishbone_bd_ram_mem3_reg[189][29]/P0001  & n14001 ;
  assign n14252 = \wishbone_bd_ram_mem3_reg[185][29]/P0001  & n13372 ;
  assign n14253 = ~n14251 & ~n14252 ;
  assign n14254 = n14250 & n14253 ;
  assign n14255 = n14247 & n14254 ;
  assign n14256 = \wishbone_bd_ram_mem3_reg[13][29]/P0001  & n13844 ;
  assign n14257 = \wishbone_bd_ram_mem3_reg[162][29]/P0001  & n13726 ;
  assign n14258 = ~n14256 & ~n14257 ;
  assign n14259 = \wishbone_bd_ram_mem3_reg[131][29]/P0001  & n13358 ;
  assign n14260 = \wishbone_bd_ram_mem3_reg[22][29]/P0001  & n13744 ;
  assign n14261 = ~n14259 & ~n14260 ;
  assign n14262 = n14258 & n14261 ;
  assign n14263 = \wishbone_bd_ram_mem3_reg[103][29]/P0001  & n13320 ;
  assign n14264 = \wishbone_bd_ram_mem3_reg[240][29]/P0001  & n13352 ;
  assign n14265 = ~n14263 & ~n14264 ;
  assign n14266 = \wishbone_bd_ram_mem3_reg[170][29]/P0001  & n14007 ;
  assign n14267 = \wishbone_bd_ram_mem3_reg[136][29]/P0001  & n13963 ;
  assign n14268 = ~n14266 & ~n14267 ;
  assign n14269 = n14265 & n14268 ;
  assign n14270 = n14262 & n14269 ;
  assign n14271 = n14255 & n14270 ;
  assign n14272 = n14240 & n14271 ;
  assign n14273 = \wishbone_bd_ram_mem3_reg[6][29]/P0001  & n13915 ;
  assign n14274 = \wishbone_bd_ram_mem3_reg[110][29]/P0001  & n14030 ;
  assign n14275 = ~n14273 & ~n14274 ;
  assign n14276 = \wishbone_bd_ram_mem3_reg[89][29]/P0001  & n13910 ;
  assign n14277 = \wishbone_bd_ram_mem3_reg[64][29]/P0001  & n13904 ;
  assign n14278 = ~n14276 & ~n14277 ;
  assign n14279 = n14275 & n14278 ;
  assign n14280 = \wishbone_bd_ram_mem3_reg[220][29]/P0001  & n13965 ;
  assign n14281 = \wishbone_bd_ram_mem3_reg[216][29]/P0001  & n14005 ;
  assign n14282 = ~n14280 & ~n14281 ;
  assign n14283 = \wishbone_bd_ram_mem3_reg[12][29]/P0001  & n13733 ;
  assign n14284 = \wishbone_bd_ram_mem3_reg[56][29]/P0001  & n13611 ;
  assign n14285 = ~n14283 & ~n14284 ;
  assign n14286 = n14282 & n14285 ;
  assign n14287 = n14279 & n14286 ;
  assign n14288 = \wishbone_bd_ram_mem3_reg[194][29]/P0001  & n13624 ;
  assign n14289 = \wishbone_bd_ram_mem3_reg[39][29]/P0001  & n13893 ;
  assign n14290 = ~n14288 & ~n14289 ;
  assign n14291 = \wishbone_bd_ram_mem3_reg[237][29]/P0001  & n13924 ;
  assign n14292 = \wishbone_bd_ram_mem3_reg[204][29]/P0001  & n13821 ;
  assign n14293 = ~n14291 & ~n14292 ;
  assign n14294 = n14290 & n14293 ;
  assign n14295 = \wishbone_bd_ram_mem3_reg[171][29]/P0001  & n13422 ;
  assign n14296 = \wishbone_bd_ram_mem3_reg[239][29]/P0001  & n13349 ;
  assign n14297 = ~n14295 & ~n14296 ;
  assign n14298 = \wishbone_bd_ram_mem3_reg[93][29]/P0001  & n13891 ;
  assign n14299 = \wishbone_bd_ram_mem3_reg[59][29]/P0001  & n13613 ;
  assign n14300 = ~n14298 & ~n14299 ;
  assign n14301 = n14297 & n14300 ;
  assign n14302 = n14294 & n14301 ;
  assign n14303 = n14287 & n14302 ;
  assign n14304 = \wishbone_bd_ram_mem3_reg[38][29]/P0001  & n13828 ;
  assign n14305 = \wishbone_bd_ram_mem3_reg[45][29]/P0001  & n13420 ;
  assign n14306 = ~n14304 & ~n14305 ;
  assign n14307 = \wishbone_bd_ram_mem3_reg[195][29]/P0001  & n13700 ;
  assign n14308 = \wishbone_bd_ram_mem3_reg[196][29]/P0001  & n13977 ;
  assign n14309 = ~n14307 & ~n14308 ;
  assign n14310 = n14306 & n14309 ;
  assign n14311 = \wishbone_bd_ram_mem3_reg[101][29]/P0001  & n13772 ;
  assign n14312 = \wishbone_bd_ram_mem3_reg[226][29]/P0001  & n13668 ;
  assign n14313 = ~n14311 & ~n14312 ;
  assign n14314 = \wishbone_bd_ram_mem3_reg[159][29]/P0001  & n13627 ;
  assign n14315 = \wishbone_bd_ram_mem3_reg[116][29]/P0001  & n13865 ;
  assign n14316 = ~n14314 & ~n14315 ;
  assign n14317 = n14313 & n14316 ;
  assign n14318 = n14310 & n14317 ;
  assign n14319 = \wishbone_bd_ram_mem3_reg[203][29]/P0001  & n13816 ;
  assign n14320 = \wishbone_bd_ram_mem3_reg[117][29]/P0001  & n13557 ;
  assign n14321 = ~n14319 & ~n14320 ;
  assign n14322 = \wishbone_bd_ram_mem3_reg[73][29]/P0001  & n13456 ;
  assign n14323 = \wishbone_bd_ram_mem3_reg[251][29]/P0001  & n14019 ;
  assign n14324 = ~n14322 & ~n14323 ;
  assign n14325 = n14321 & n14324 ;
  assign n14326 = \wishbone_bd_ram_mem3_reg[183][29]/P0001  & n13645 ;
  assign n14327 = \wishbone_bd_ram_mem3_reg[252][29]/P0001  & n13986 ;
  assign n14328 = ~n14326 & ~n14327 ;
  assign n14329 = \wishbone_bd_ram_mem3_reg[180][29]/P0001  & n13650 ;
  assign n14330 = \wishbone_bd_ram_mem3_reg[29][29]/P0001  & n13412 ;
  assign n14331 = ~n14329 & ~n14330 ;
  assign n14332 = n14328 & n14331 ;
  assign n14333 = n14325 & n14332 ;
  assign n14334 = n14318 & n14333 ;
  assign n14335 = n14303 & n14334 ;
  assign n14336 = n14272 & n14335 ;
  assign n14337 = n14209 & n14336 ;
  assign n14338 = \wishbone_bd_ram_mem3_reg[40][29]/P0001  & n13661 ;
  assign n14339 = \wishbone_bd_ram_mem3_reg[1][29]/P0001  & n13888 ;
  assign n14340 = ~n14338 & ~n14339 ;
  assign n14341 = \wishbone_bd_ram_mem3_reg[82][29]/P0001  & n13374 ;
  assign n14342 = \wishbone_bd_ram_mem3_reg[206][29]/P0001  & n13414 ;
  assign n14343 = ~n14341 & ~n14342 ;
  assign n14344 = n14340 & n14343 ;
  assign n14345 = \wishbone_bd_ram_mem3_reg[157][29]/P0001  & n13445 ;
  assign n14346 = \wishbone_bd_ram_mem3_reg[8][29]/P0001  & n13459 ;
  assign n14347 = ~n14345 & ~n14346 ;
  assign n14348 = \wishbone_bd_ram_mem3_reg[213][29]/P0001  & n13870 ;
  assign n14349 = \wishbone_bd_ram_mem3_reg[63][29]/P0001  & n13327 ;
  assign n14350 = ~n14348 & ~n14349 ;
  assign n14351 = n14347 & n14350 ;
  assign n14352 = n14344 & n14351 ;
  assign n14353 = \wishbone_bd_ram_mem3_reg[166][29]/P0001  & n13999 ;
  assign n14354 = \wishbone_bd_ram_mem3_reg[69][29]/P0001  & n13487 ;
  assign n14355 = ~n14353 & ~n14354 ;
  assign n14356 = \wishbone_bd_ram_mem3_reg[84][29]/P0001  & n13385 ;
  assign n14357 = \wishbone_bd_ram_mem3_reg[53][29]/P0001  & n13875 ;
  assign n14358 = ~n14356 & ~n14357 ;
  assign n14359 = n14355 & n14358 ;
  assign n14360 = \wishbone_bd_ram_mem3_reg[148][29]/P0001  & n13868 ;
  assign n14361 = \wishbone_bd_ram_mem3_reg[98][29]/P0001  & n13569 ;
  assign n14362 = ~n14360 & ~n14361 ;
  assign n14363 = \wishbone_bd_ram_mem3_reg[186][29]/P0001  & n13616 ;
  assign n14364 = \wishbone_bd_ram_mem3_reg[7][29]/P0001  & n13546 ;
  assign n14365 = ~n14363 & ~n14364 ;
  assign n14366 = n14362 & n14365 ;
  assign n14367 = n14359 & n14366 ;
  assign n14368 = n14352 & n14367 ;
  assign n14369 = \wishbone_bd_ram_mem3_reg[221][29]/P0001  & n13641 ;
  assign n14370 = \wishbone_bd_ram_mem3_reg[0][29]/P0001  & n13539 ;
  assign n14371 = ~n14369 & ~n14370 ;
  assign n14372 = \wishbone_bd_ram_mem3_reg[50][29]/P0001  & n13686 ;
  assign n14373 = \wishbone_bd_ram_mem3_reg[230][29]/P0001  & n13994 ;
  assign n14374 = ~n14372 & ~n14373 ;
  assign n14375 = n14371 & n14374 ;
  assign n14376 = \wishbone_bd_ram_mem3_reg[190][29]/P0001  & n13365 ;
  assign n14377 = \wishbone_bd_ram_mem3_reg[232][29]/P0001  & n13510 ;
  assign n14378 = ~n14376 & ~n14377 ;
  assign n14379 = \wishbone_bd_ram_mem3_reg[228][29]/P0001  & n13497 ;
  assign n14380 = \wishbone_bd_ram_mem3_reg[214][29]/P0001  & n13938 ;
  assign n14381 = ~n14379 & ~n14380 ;
  assign n14382 = n14378 & n14381 ;
  assign n14383 = n14375 & n14382 ;
  assign n14384 = \wishbone_bd_ram_mem3_reg[119][29]/P0001  & n14033 ;
  assign n14385 = \wishbone_bd_ram_mem3_reg[9][29]/P0001  & n13580 ;
  assign n14386 = ~n14384 & ~n14385 ;
  assign n14387 = \wishbone_bd_ram_mem3_reg[215][29]/P0001  & n13901 ;
  assign n14388 = \wishbone_bd_ram_mem3_reg[74][29]/P0001  & n13564 ;
  assign n14389 = ~n14387 & ~n14388 ;
  assign n14390 = n14386 & n14389 ;
  assign n14391 = \wishbone_bd_ram_mem3_reg[32][29]/P0001  & n13736 ;
  assign n14392 = \wishbone_bd_ram_mem3_reg[41][29]/P0001  & n14017 ;
  assign n14393 = ~n14391 & ~n14392 ;
  assign n14394 = \wishbone_bd_ram_mem3_reg[51][29]/P0001  & n13880 ;
  assign n14395 = \wishbone_bd_ram_mem3_reg[208][29]/P0001  & n14010 ;
  assign n14396 = ~n14394 & ~n14395 ;
  assign n14397 = n14393 & n14396 ;
  assign n14398 = n14390 & n14397 ;
  assign n14399 = n14383 & n14398 ;
  assign n14400 = n14368 & n14399 ;
  assign n14401 = \wishbone_bd_ram_mem3_reg[249][29]/P0001  & n13431 ;
  assign n14402 = \wishbone_bd_ram_mem3_reg[15][29]/P0001  & n13797 ;
  assign n14403 = ~n14401 & ~n14402 ;
  assign n14404 = \wishbone_bd_ram_mem3_reg[68][29]/P0001  & n13379 ;
  assign n14405 = \wishbone_bd_ram_mem3_reg[72][29]/P0001  & n13582 ;
  assign n14406 = ~n14404 & ~n14405 ;
  assign n14407 = n14403 & n14406 ;
  assign n14408 = \wishbone_bd_ram_mem3_reg[87][29]/P0001  & n13691 ;
  assign n14409 = \wishbone_bd_ram_mem3_reg[130][29]/P0001  & n13427 ;
  assign n14410 = ~n14408 & ~n14409 ;
  assign n14411 = \wishbone_bd_ram_mem3_reg[138][29]/P0001  & n13398 ;
  assign n14412 = \wishbone_bd_ram_mem3_reg[115][29]/P0001  & n13747 ;
  assign n14413 = ~n14411 & ~n14412 ;
  assign n14414 = n14410 & n14413 ;
  assign n14415 = n14407 & n14414 ;
  assign n14416 = \wishbone_bd_ram_mem3_reg[43][29]/P0001  & n13761 ;
  assign n14417 = \wishbone_bd_ram_mem3_reg[241][29]/P0001  & n13854 ;
  assign n14418 = ~n14416 & ~n14417 ;
  assign n14419 = \wishbone_bd_ram_mem3_reg[118][29]/P0001  & n13589 ;
  assign n14420 = \wishbone_bd_ram_mem3_reg[242][29]/P0001  & n13383 ;
  assign n14421 = ~n14419 & ~n14420 ;
  assign n14422 = n14418 & n14421 ;
  assign n14423 = \wishbone_bd_ram_mem3_reg[60][29]/P0001  & n13790 ;
  assign n14424 = \wishbone_bd_ram_mem3_reg[168][29]/P0001  & n13795 ;
  assign n14425 = ~n14423 & ~n14424 ;
  assign n14426 = \wishbone_bd_ram_mem3_reg[122][29]/P0001  & n13679 ;
  assign n14427 = \wishbone_bd_ram_mem3_reg[109][29]/P0001  & n13306 ;
  assign n14428 = ~n14426 & ~n14427 ;
  assign n14429 = n14425 & n14428 ;
  assign n14430 = n14422 & n14429 ;
  assign n14431 = n14415 & n14430 ;
  assign n14432 = \wishbone_bd_ram_mem3_reg[108][29]/P0001  & n13814 ;
  assign n14433 = \wishbone_bd_ram_mem3_reg[211][29]/P0001  & n13805 ;
  assign n14434 = ~n14432 & ~n14433 ;
  assign n14435 = \wishbone_bd_ram_mem3_reg[97][29]/P0001  & n13724 ;
  assign n14436 = \wishbone_bd_ram_mem3_reg[19][29]/P0001  & n13886 ;
  assign n14437 = ~n14435 & ~n14436 ;
  assign n14438 = n14434 & n14437 ;
  assign n14439 = \wishbone_bd_ram_mem3_reg[145][29]/P0001  & n13715 ;
  assign n14440 = \wishbone_bd_ram_mem3_reg[114][29]/P0001  & n13763 ;
  assign n14441 = ~n14439 & ~n14440 ;
  assign n14442 = \wishbone_bd_ram_mem3_reg[246][29]/P0001  & n13981 ;
  assign n14443 = \wishbone_bd_ram_mem3_reg[255][29]/P0001  & n13952 ;
  assign n14444 = ~n14442 & ~n14443 ;
  assign n14445 = n14441 & n14444 ;
  assign n14446 = n14438 & n14445 ;
  assign n14447 = \wishbone_bd_ram_mem3_reg[207][29]/P0001  & n13826 ;
  assign n14448 = \wishbone_bd_ram_mem3_reg[20][29]/P0001  & n13839 ;
  assign n14449 = ~n14447 & ~n14448 ;
  assign n14450 = \wishbone_bd_ram_mem3_reg[25][29]/P0001  & n13742 ;
  assign n14451 = \wishbone_bd_ram_mem3_reg[238][29]/P0001  & n13819 ;
  assign n14452 = ~n14450 & ~n14451 ;
  assign n14453 = n14449 & n14452 ;
  assign n14454 = \wishbone_bd_ram_mem3_reg[11][29]/P0001  & n13774 ;
  assign n14455 = \wishbone_bd_ram_mem3_reg[161][29]/P0001  & n13505 ;
  assign n14456 = ~n14454 & ~n14455 ;
  assign n14457 = \wishbone_bd_ram_mem3_reg[21][29]/P0001  & n13438 ;
  assign n14458 = \wishbone_bd_ram_mem3_reg[33][29]/P0001  & n13933 ;
  assign n14459 = ~n14457 & ~n14458 ;
  assign n14460 = n14456 & n14459 ;
  assign n14461 = n14453 & n14460 ;
  assign n14462 = n14446 & n14461 ;
  assign n14463 = n14431 & n14462 ;
  assign n14464 = n14400 & n14463 ;
  assign n14465 = \wishbone_bd_ram_mem3_reg[62][29]/P0001  & n13529 ;
  assign n14466 = \wishbone_bd_ram_mem3_reg[248][29]/P0001  & n13647 ;
  assign n14467 = ~n14465 & ~n14466 ;
  assign n14468 = \wishbone_bd_ram_mem3_reg[152][29]/P0001  & n13912 ;
  assign n14469 = \wishbone_bd_ram_mem3_reg[172][29]/P0001  & n13377 ;
  assign n14470 = ~n14468 & ~n14469 ;
  assign n14471 = n14467 & n14470 ;
  assign n14472 = \wishbone_bd_ram_mem3_reg[146][29]/P0001  & n13958 ;
  assign n14473 = \wishbone_bd_ram_mem3_reg[54][29]/P0001  & n13622 ;
  assign n14474 = ~n14472 & ~n14473 ;
  assign n14475 = \wishbone_bd_ram_mem3_reg[128][29]/P0001  & n13652 ;
  assign n14476 = \wishbone_bd_ram_mem3_reg[229][29]/P0001  & n13552 ;
  assign n14477 = ~n14475 & ~n14476 ;
  assign n14478 = n14474 & n14477 ;
  assign n14479 = n14471 & n14478 ;
  assign n14480 = \wishbone_bd_ram_mem3_reg[165][29]/P0001  & n14028 ;
  assign n14481 = \wishbone_bd_ram_mem3_reg[254][29]/P0001  & n13283 ;
  assign n14482 = ~n14480 & ~n14481 ;
  assign n14483 = \wishbone_bd_ram_mem3_reg[76][29]/P0001  & n13831 ;
  assign n14484 = \wishbone_bd_ram_mem3_reg[179][29]/P0001  & n14035 ;
  assign n14485 = ~n14483 & ~n14484 ;
  assign n14486 = n14482 & n14485 ;
  assign n14487 = \wishbone_bd_ram_mem3_reg[28][29]/P0001  & n13810 ;
  assign n14488 = \wishbone_bd_ram_mem3_reg[3][29]/P0001  & n13354 ;
  assign n14489 = ~n14487 & ~n14488 ;
  assign n14490 = \wishbone_bd_ram_mem3_reg[137][29]/P0001  & n13808 ;
  assign n14491 = \wishbone_bd_ram_mem3_reg[78][29]/P0001  & n13277 ;
  assign n14492 = ~n14490 & ~n14491 ;
  assign n14493 = n14489 & n14492 ;
  assign n14494 = n14486 & n14493 ;
  assign n14495 = n14479 & n14494 ;
  assign n14496 = \wishbone_bd_ram_mem3_reg[151][29]/P0001  & n13697 ;
  assign n14497 = \wishbone_bd_ram_mem3_reg[14][29]/P0001  & n13972 ;
  assign n14498 = ~n14496 & ~n14497 ;
  assign n14499 = \wishbone_bd_ram_mem3_reg[26][29]/P0001  & n13521 ;
  assign n14500 = \wishbone_bd_ram_mem3_reg[200][29]/P0001  & n13922 ;
  assign n14501 = ~n14499 & ~n14500 ;
  assign n14502 = n14498 & n14501 ;
  assign n14503 = \wishbone_bd_ram_mem3_reg[102][29]/P0001  & n13534 ;
  assign n14504 = \wishbone_bd_ram_mem3_reg[129][29]/P0001  & n13629 ;
  assign n14505 = ~n14503 & ~n14504 ;
  assign n14506 = \wishbone_bd_ram_mem3_reg[10][29]/P0001  & n13837 ;
  assign n14507 = \wishbone_bd_ram_mem3_reg[163][29]/P0001  & n13255 ;
  assign n14508 = ~n14506 & ~n14507 ;
  assign n14509 = n14505 & n14508 ;
  assign n14510 = n14502 & n14509 ;
  assign n14511 = \wishbone_bd_ram_mem3_reg[205][29]/P0001  & n13947 ;
  assign n14512 = \wishbone_bd_ram_mem3_reg[176][29]/P0001  & n13262 ;
  assign n14513 = ~n14511 & ~n14512 ;
  assign n14514 = \wishbone_bd_ram_mem3_reg[23][29]/P0001  & n13857 ;
  assign n14515 = \wishbone_bd_ram_mem3_reg[164][29]/P0001  & n13236 ;
  assign n14516 = ~n14514 & ~n14515 ;
  assign n14517 = n14513 & n14516 ;
  assign n14518 = \wishbone_bd_ram_mem3_reg[18][29]/P0001  & n13532 ;
  assign n14519 = \wishbone_bd_ram_mem3_reg[88][29]/P0001  & n13347 ;
  assign n14520 = ~n14518 & ~n14519 ;
  assign n14521 = \wishbone_bd_ram_mem3_reg[219][29]/P0001  & n13577 ;
  assign n14522 = \wishbone_bd_ram_mem3_reg[167][29]/P0001  & n13940 ;
  assign n14523 = ~n14521 & ~n14522 ;
  assign n14524 = n14520 & n14523 ;
  assign n14525 = n14517 & n14524 ;
  assign n14526 = n14510 & n14525 ;
  assign n14527 = n14495 & n14526 ;
  assign n14528 = \wishbone_bd_ram_mem3_reg[236][29]/P0001  & n13480 ;
  assign n14529 = \wishbone_bd_ram_mem3_reg[79][29]/P0001  & n13779 ;
  assign n14530 = ~n14528 & ~n14529 ;
  assign n14531 = \wishbone_bd_ram_mem3_reg[140][29]/P0001  & n13287 ;
  assign n14532 = \wishbone_bd_ram_mem3_reg[124][29]/P0001  & n14024 ;
  assign n14533 = ~n14531 & ~n14532 ;
  assign n14534 = n14530 & n14533 ;
  assign n14535 = \wishbone_bd_ram_mem3_reg[177][29]/P0001  & n13863 ;
  assign n14536 = \wishbone_bd_ram_mem3_reg[133][29]/P0001  & n13492 ;
  assign n14537 = ~n14535 & ~n14536 ;
  assign n14538 = \wishbone_bd_ram_mem3_reg[218][29]/P0001  & n13792 ;
  assign n14539 = \wishbone_bd_ram_mem3_reg[235][29]/P0001  & n13518 ;
  assign n14540 = ~n14538 & ~n14539 ;
  assign n14541 = n14537 & n14540 ;
  assign n14542 = n14534 & n14541 ;
  assign n14543 = \wishbone_bd_ram_mem3_reg[5][29]/P0001  & n13243 ;
  assign n14544 = \wishbone_bd_ram_mem3_reg[31][29]/P0001  & n13758 ;
  assign n14545 = ~n14543 & ~n14544 ;
  assign n14546 = \wishbone_bd_ram_mem3_reg[30][29]/P0001  & n13713 ;
  assign n14547 = \wishbone_bd_ram_mem3_reg[184][29]/P0001  & n13960 ;
  assign n14548 = ~n14546 & ~n14547 ;
  assign n14549 = n14545 & n14548 ;
  assign n14550 = \wishbone_bd_ram_mem3_reg[245][29]/P0001  & n13877 ;
  assign n14551 = \wishbone_bd_ram_mem3_reg[16][29]/P0001  & n13695 ;
  assign n14552 = ~n14550 & ~n14551 ;
  assign n14553 = \wishbone_bd_ram_mem3_reg[227][29]/P0001  & n13388 ;
  assign n14554 = \wishbone_bd_ram_mem3_reg[52][29]/P0001  & n13988 ;
  assign n14555 = ~n14553 & ~n14554 ;
  assign n14556 = n14552 & n14555 ;
  assign n14557 = n14549 & n14556 ;
  assign n14558 = n14542 & n14557 ;
  assign n14559 = \wishbone_bd_ram_mem3_reg[153][29]/P0001  & n13309 ;
  assign n14560 = \wishbone_bd_ram_mem3_reg[155][29]/P0001  & n13738 ;
  assign n14561 = ~n14559 & ~n14560 ;
  assign n14562 = \wishbone_bd_ram_mem3_reg[96][29]/P0001  & n13425 ;
  assign n14563 = \wishbone_bd_ram_mem3_reg[156][29]/P0001  & n13769 ;
  assign n14564 = ~n14562 & ~n14563 ;
  assign n14565 = n14561 & n14564 ;
  assign n14566 = \wishbone_bd_ram_mem3_reg[217][29]/P0001  & n13767 ;
  assign n14567 = \wishbone_bd_ram_mem3_reg[209][29]/P0001  & n13689 ;
  assign n14568 = ~n14566 & ~n14567 ;
  assign n14569 = \wishbone_bd_ram_mem3_reg[150][29]/P0001  & n13666 ;
  assign n14570 = \wishbone_bd_ram_mem3_reg[223][29]/P0001  & n13335 ;
  assign n14571 = ~n14569 & ~n14570 ;
  assign n14572 = n14568 & n14571 ;
  assign n14573 = n14565 & n14572 ;
  assign n14574 = \wishbone_bd_ram_mem3_reg[55][29]/P0001  & n13618 ;
  assign n14575 = \wishbone_bd_ram_mem3_reg[99][29]/P0001  & n13996 ;
  assign n14576 = ~n14574 & ~n14575 ;
  assign n14577 = \wishbone_bd_ram_mem3_reg[234][29]/P0001  & n13781 ;
  assign n14578 = \wishbone_bd_ram_mem3_reg[187][29]/P0001  & n13756 ;
  assign n14579 = ~n14577 & ~n14578 ;
  assign n14580 = n14576 & n14579 ;
  assign n14581 = \wishbone_bd_ram_mem3_reg[92][29]/P0001  & n13859 ;
  assign n14582 = \wishbone_bd_ram_mem3_reg[132][29]/P0001  & n13927 ;
  assign n14583 = ~n14581 & ~n14582 ;
  assign n14584 = \wishbone_bd_ram_mem3_reg[37][29]/P0001  & n13710 ;
  assign n14585 = \wishbone_bd_ram_mem3_reg[197][29]/P0001  & n13594 ;
  assign n14586 = ~n14584 & ~n14585 ;
  assign n14587 = n14583 & n14586 ;
  assign n14588 = n14580 & n14587 ;
  assign n14589 = n14573 & n14588 ;
  assign n14590 = n14558 & n14589 ;
  assign n14591 = n14527 & n14590 ;
  assign n14592 = n14464 & n14591 ;
  assign n14593 = n14337 & n14592 ;
  assign n14594 = n14047 & ~n14593 ;
  assign n14595 = ~n14046 & ~n14049 ;
  assign n14596 = ~\wishbone_TxLength_reg[12]/NET0131  & n14075 ;
  assign n14597 = n14066 & ~n14596 ;
  assign n14598 = ~n14595 & ~n14597 ;
  assign n14599 = \wishbone_TxLength_reg[13]/NET0131  & ~n14598 ;
  assign n14600 = n14061 & n14075 ;
  assign n14601 = n14066 & n14600 ;
  assign n14602 = ~n14599 & ~n14601 ;
  assign n14603 = ~n14594 & n14602 ;
  assign n14604 = \wishbone_bd_ram_mem3_reg[64][30]/P0001  & n13904 ;
  assign n14605 = \wishbone_bd_ram_mem3_reg[211][30]/P0001  & n13805 ;
  assign n14606 = ~n14604 & ~n14605 ;
  assign n14607 = \wishbone_bd_ram_mem3_reg[1][30]/P0001  & n13888 ;
  assign n14608 = \wishbone_bd_ram_mem3_reg[10][30]/P0001  & n13837 ;
  assign n14609 = ~n14607 & ~n14608 ;
  assign n14610 = n14606 & n14609 ;
  assign n14611 = \wishbone_bd_ram_mem3_reg[132][30]/P0001  & n13927 ;
  assign n14612 = \wishbone_bd_ram_mem3_reg[237][30]/P0001  & n13924 ;
  assign n14613 = ~n14611 & ~n14612 ;
  assign n14614 = \wishbone_bd_ram_mem3_reg[119][30]/P0001  & n14033 ;
  assign n14615 = \wishbone_bd_ram_mem3_reg[242][30]/P0001  & n13383 ;
  assign n14616 = ~n14614 & ~n14615 ;
  assign n14617 = n14613 & n14616 ;
  assign n14618 = n14610 & n14617 ;
  assign n14619 = \wishbone_bd_ram_mem3_reg[206][30]/P0001  & n13414 ;
  assign n14620 = \wishbone_bd_ram_mem3_reg[175][30]/P0001  & n13674 ;
  assign n14621 = ~n14619 & ~n14620 ;
  assign n14622 = \wishbone_bd_ram_mem3_reg[77][30]/P0001  & n13935 ;
  assign n14623 = \wishbone_bd_ram_mem3_reg[232][30]/P0001  & n13510 ;
  assign n14624 = ~n14622 & ~n14623 ;
  assign n14625 = n14621 & n14624 ;
  assign n14626 = \wishbone_bd_ram_mem3_reg[109][30]/P0001  & n13306 ;
  assign n14627 = \wishbone_bd_ram_mem3_reg[181][30]/P0001  & n13587 ;
  assign n14628 = ~n14626 & ~n14627 ;
  assign n14629 = \wishbone_bd_ram_mem3_reg[74][30]/P0001  & n13564 ;
  assign n14630 = \wishbone_bd_ram_mem3_reg[192][30]/P0001  & n13390 ;
  assign n14631 = ~n14629 & ~n14630 ;
  assign n14632 = n14628 & n14631 ;
  assign n14633 = n14625 & n14632 ;
  assign n14634 = n14618 & n14633 ;
  assign n14635 = \wishbone_bd_ram_mem3_reg[104][30]/P0001  & n13684 ;
  assign n14636 = \wishbone_bd_ram_mem3_reg[102][30]/P0001  & n13534 ;
  assign n14637 = ~n14635 & ~n14636 ;
  assign n14638 = \wishbone_bd_ram_mem3_reg[50][30]/P0001  & n13686 ;
  assign n14639 = \wishbone_bd_ram_mem3_reg[163][30]/P0001  & n13255 ;
  assign n14640 = ~n14638 & ~n14639 ;
  assign n14641 = n14637 & n14640 ;
  assign n14642 = \wishbone_bd_ram_mem3_reg[226][30]/P0001  & n13668 ;
  assign n14643 = \wishbone_bd_ram_mem3_reg[199][30]/P0001  & n13499 ;
  assign n14644 = ~n14642 & ~n14643 ;
  assign n14645 = \wishbone_bd_ram_mem3_reg[32][30]/P0001  & n13736 ;
  assign n14646 = \wishbone_bd_ram_mem3_reg[67][30]/P0001  & n13663 ;
  assign n14647 = ~n14645 & ~n14646 ;
  assign n14648 = n14644 & n14647 ;
  assign n14649 = n14641 & n14648 ;
  assign n14650 = \wishbone_bd_ram_mem3_reg[182][30]/P0001  & n13598 ;
  assign n14651 = \wishbone_bd_ram_mem3_reg[227][30]/P0001  & n13388 ;
  assign n14652 = ~n14650 & ~n14651 ;
  assign n14653 = \wishbone_bd_ram_mem3_reg[216][30]/P0001  & n14005 ;
  assign n14654 = \wishbone_bd_ram_mem3_reg[43][30]/P0001  & n13761 ;
  assign n14655 = ~n14653 & ~n14654 ;
  assign n14656 = n14652 & n14655 ;
  assign n14657 = \wishbone_bd_ram_mem3_reg[58][30]/P0001  & n13949 ;
  assign n14658 = \wishbone_bd_ram_mem3_reg[205][30]/P0001  & n13947 ;
  assign n14659 = ~n14657 & ~n14658 ;
  assign n14660 = \wishbone_bd_ram_mem3_reg[144][30]/P0001  & n13508 ;
  assign n14661 = \wishbone_bd_ram_mem3_reg[215][30]/P0001  & n13901 ;
  assign n14662 = ~n14660 & ~n14661 ;
  assign n14663 = n14659 & n14662 ;
  assign n14664 = n14656 & n14663 ;
  assign n14665 = n14649 & n14664 ;
  assign n14666 = n14634 & n14665 ;
  assign n14667 = \wishbone_bd_ram_mem3_reg[173][30]/P0001  & n13360 ;
  assign n14668 = \wishbone_bd_ram_mem3_reg[123][30]/P0001  & n13749 ;
  assign n14669 = ~n14667 & ~n14668 ;
  assign n14670 = \wishbone_bd_ram_mem3_reg[193][30]/P0001  & n14022 ;
  assign n14671 = \wishbone_bd_ram_mem3_reg[3][30]/P0001  & n13354 ;
  assign n14672 = ~n14670 & ~n14671 ;
  assign n14673 = n14669 & n14672 ;
  assign n14674 = \wishbone_bd_ram_mem3_reg[183][30]/P0001  & n13645 ;
  assign n14675 = \wishbone_bd_ram_mem3_reg[131][30]/P0001  & n13358 ;
  assign n14676 = ~n14674 & ~n14675 ;
  assign n14677 = \wishbone_bd_ram_mem3_reg[213][30]/P0001  & n13870 ;
  assign n14678 = \wishbone_bd_ram_mem3_reg[156][30]/P0001  & n13769 ;
  assign n14679 = ~n14677 & ~n14678 ;
  assign n14680 = n14676 & n14679 ;
  assign n14681 = n14673 & n14680 ;
  assign n14682 = \wishbone_bd_ram_mem3_reg[107][30]/P0001  & n13476 ;
  assign n14683 = \wishbone_bd_ram_mem3_reg[73][30]/P0001  & n13456 ;
  assign n14684 = ~n14682 & ~n14683 ;
  assign n14685 = \wishbone_bd_ram_mem3_reg[208][30]/P0001  & n14010 ;
  assign n14686 = \wishbone_bd_ram_mem3_reg[241][30]/P0001  & n13854 ;
  assign n14687 = ~n14685 & ~n14686 ;
  assign n14688 = n14684 & n14687 ;
  assign n14689 = \wishbone_bd_ram_mem3_reg[154][30]/P0001  & n13403 ;
  assign n14690 = \wishbone_bd_ram_mem3_reg[252][30]/P0001  & n13986 ;
  assign n14691 = ~n14689 & ~n14690 ;
  assign n14692 = \wishbone_bd_ram_mem3_reg[72][30]/P0001  & n13582 ;
  assign n14693 = \wishbone_bd_ram_mem3_reg[229][30]/P0001  & n13552 ;
  assign n14694 = ~n14692 & ~n14693 ;
  assign n14695 = n14691 & n14694 ;
  assign n14696 = n14688 & n14695 ;
  assign n14697 = n14681 & n14696 ;
  assign n14698 = \wishbone_bd_ram_mem3_reg[83][30]/P0001  & n13454 ;
  assign n14699 = \wishbone_bd_ram_mem3_reg[130][30]/P0001  & n13427 ;
  assign n14700 = ~n14698 & ~n14699 ;
  assign n14701 = \wishbone_bd_ram_mem3_reg[98][30]/P0001  & n13569 ;
  assign n14702 = \wishbone_bd_ram_mem3_reg[146][30]/P0001  & n13958 ;
  assign n14703 = ~n14701 & ~n14702 ;
  assign n14704 = n14700 & n14703 ;
  assign n14705 = \wishbone_bd_ram_mem3_reg[210][30]/P0001  & n13443 ;
  assign n14706 = \wishbone_bd_ram_mem3_reg[180][30]/P0001  & n13650 ;
  assign n14707 = ~n14705 & ~n14706 ;
  assign n14708 = \wishbone_bd_ram_mem3_reg[56][30]/P0001  & n13611 ;
  assign n14709 = \wishbone_bd_ram_mem3_reg[27][30]/P0001  & n13251 ;
  assign n14710 = ~n14708 & ~n14709 ;
  assign n14711 = n14707 & n14710 ;
  assign n14712 = n14704 & n14711 ;
  assign n14713 = \wishbone_bd_ram_mem3_reg[196][30]/P0001  & n13977 ;
  assign n14714 = \wishbone_bd_ram_mem3_reg[61][30]/P0001  & n13544 ;
  assign n14715 = ~n14713 & ~n14714 ;
  assign n14716 = \wishbone_bd_ram_mem3_reg[116][30]/P0001  & n13865 ;
  assign n14717 = \wishbone_bd_ram_mem3_reg[148][30]/P0001  & n13868 ;
  assign n14718 = ~n14716 & ~n14717 ;
  assign n14719 = n14715 & n14718 ;
  assign n14720 = \wishbone_bd_ram_mem3_reg[66][30]/P0001  & n13603 ;
  assign n14721 = \wishbone_bd_ram_mem3_reg[15][30]/P0001  & n13797 ;
  assign n14722 = ~n14720 & ~n14721 ;
  assign n14723 = \wishbone_bd_ram_mem3_reg[33][30]/P0001  & n13933 ;
  assign n14724 = \wishbone_bd_ram_mem3_reg[174][30]/P0001  & n13899 ;
  assign n14725 = ~n14723 & ~n14724 ;
  assign n14726 = n14722 & n14725 ;
  assign n14727 = n14719 & n14726 ;
  assign n14728 = n14712 & n14727 ;
  assign n14729 = n14697 & n14728 ;
  assign n14730 = n14666 & n14729 ;
  assign n14731 = \wishbone_bd_ram_mem3_reg[34][30]/P0001  & n13450 ;
  assign n14732 = \wishbone_bd_ram_mem3_reg[169][30]/P0001  & n13541 ;
  assign n14733 = ~n14731 & ~n14732 ;
  assign n14734 = \wishbone_bd_ram_mem3_reg[200][30]/P0001  & n13922 ;
  assign n14735 = \wishbone_bd_ram_mem3_reg[230][30]/P0001  & n13994 ;
  assign n14736 = ~n14734 & ~n14735 ;
  assign n14737 = n14733 & n14736 ;
  assign n14738 = \wishbone_bd_ram_mem3_reg[255][30]/P0001  & n13952 ;
  assign n14739 = \wishbone_bd_ram_mem3_reg[87][30]/P0001  & n13691 ;
  assign n14740 = ~n14738 & ~n14739 ;
  assign n14741 = \wishbone_bd_ram_mem3_reg[0][30]/P0001  & n13539 ;
  assign n14742 = \wishbone_bd_ram_mem3_reg[18][30]/P0001  & n13532 ;
  assign n14743 = ~n14741 & ~n14742 ;
  assign n14744 = n14740 & n14743 ;
  assign n14745 = n14737 & n14744 ;
  assign n14746 = \wishbone_bd_ram_mem3_reg[186][30]/P0001  & n13616 ;
  assign n14747 = \wishbone_bd_ram_mem3_reg[136][30]/P0001  & n13963 ;
  assign n14748 = ~n14746 & ~n14747 ;
  assign n14749 = \wishbone_bd_ram_mem3_reg[158][30]/P0001  & n13294 ;
  assign n14750 = \wishbone_bd_ram_mem3_reg[212][30]/P0001  & n13634 ;
  assign n14751 = ~n14749 & ~n14750 ;
  assign n14752 = n14748 & n14751 ;
  assign n14753 = \wishbone_bd_ram_mem3_reg[112][30]/P0001  & n13482 ;
  assign n14754 = \wishbone_bd_ram_mem3_reg[86][30]/P0001  & n13485 ;
  assign n14755 = ~n14753 & ~n14754 ;
  assign n14756 = \wishbone_bd_ram_mem3_reg[153][30]/P0001  & n13309 ;
  assign n14757 = \wishbone_bd_ram_mem3_reg[234][30]/P0001  & n13781 ;
  assign n14758 = ~n14756 & ~n14757 ;
  assign n14759 = n14755 & n14758 ;
  assign n14760 = n14752 & n14759 ;
  assign n14761 = n14745 & n14760 ;
  assign n14762 = \wishbone_bd_ram_mem3_reg[20][30]/P0001  & n13839 ;
  assign n14763 = \wishbone_bd_ram_mem3_reg[224][30]/P0001  & n13433 ;
  assign n14764 = ~n14762 & ~n14763 ;
  assign n14765 = \wishbone_bd_ram_mem3_reg[60][30]/P0001  & n13790 ;
  assign n14766 = \wishbone_bd_ram_mem3_reg[36][30]/P0001  & n13639 ;
  assign n14767 = ~n14765 & ~n14766 ;
  assign n14768 = n14764 & n14767 ;
  assign n14769 = \wishbone_bd_ram_mem3_reg[164][30]/P0001  & n13236 ;
  assign n14770 = \wishbone_bd_ram_mem3_reg[135][30]/P0001  & n13672 ;
  assign n14771 = ~n14769 & ~n14770 ;
  assign n14772 = \wishbone_bd_ram_mem3_reg[19][30]/P0001  & n13886 ;
  assign n14773 = \wishbone_bd_ram_mem3_reg[103][30]/P0001  & n13320 ;
  assign n14774 = ~n14772 & ~n14773 ;
  assign n14775 = n14771 & n14774 ;
  assign n14776 = n14768 & n14775 ;
  assign n14777 = \wishbone_bd_ram_mem3_reg[9][30]/P0001  & n13580 ;
  assign n14778 = \wishbone_bd_ram_mem3_reg[97][30]/P0001  & n13724 ;
  assign n14779 = ~n14777 & ~n14778 ;
  assign n14780 = \wishbone_bd_ram_mem3_reg[149][30]/P0001  & n13469 ;
  assign n14781 = \wishbone_bd_ram_mem3_reg[28][30]/P0001  & n13810 ;
  assign n14782 = ~n14780 & ~n14781 ;
  assign n14783 = n14779 & n14782 ;
  assign n14784 = \wishbone_bd_ram_mem3_reg[89][30]/P0001  & n13910 ;
  assign n14785 = \wishbone_bd_ram_mem3_reg[250][30]/P0001  & n13677 ;
  assign n14786 = ~n14784 & ~n14785 ;
  assign n14787 = \wishbone_bd_ram_mem3_reg[185][30]/P0001  & n13372 ;
  assign n14788 = \wishbone_bd_ram_mem3_reg[100][30]/P0001  & n13401 ;
  assign n14789 = ~n14787 & ~n14788 ;
  assign n14790 = n14786 & n14789 ;
  assign n14791 = n14783 & n14790 ;
  assign n14792 = n14776 & n14791 ;
  assign n14793 = n14761 & n14792 ;
  assign n14794 = \wishbone_bd_ram_mem3_reg[129][30]/P0001  & n13629 ;
  assign n14795 = \wishbone_bd_ram_mem3_reg[91][30]/P0001  & n13954 ;
  assign n14796 = ~n14794 & ~n14795 ;
  assign n14797 = \wishbone_bd_ram_mem3_reg[166][30]/P0001  & n13999 ;
  assign n14798 = \wishbone_bd_ram_mem3_reg[204][30]/P0001  & n13821 ;
  assign n14799 = ~n14797 & ~n14798 ;
  assign n14800 = n14796 & n14799 ;
  assign n14801 = \wishbone_bd_ram_mem3_reg[236][30]/P0001  & n13480 ;
  assign n14802 = \wishbone_bd_ram_mem3_reg[187][30]/P0001  & n13756 ;
  assign n14803 = ~n14801 & ~n14802 ;
  assign n14804 = \wishbone_bd_ram_mem3_reg[13][30]/P0001  & n13844 ;
  assign n14805 = \wishbone_bd_ram_mem3_reg[26][30]/P0001  & n13521 ;
  assign n14806 = ~n14804 & ~n14805 ;
  assign n14807 = n14803 & n14806 ;
  assign n14808 = n14800 & n14807 ;
  assign n14809 = \wishbone_bd_ram_mem3_reg[178][30]/P0001  & n13301 ;
  assign n14810 = \wishbone_bd_ram_mem3_reg[157][30]/P0001  & n13445 ;
  assign n14811 = ~n14809 & ~n14810 ;
  assign n14812 = \wishbone_bd_ram_mem3_reg[176][30]/P0001  & n13262 ;
  assign n14813 = \wishbone_bd_ram_mem3_reg[235][30]/P0001  & n13518 ;
  assign n14814 = ~n14812 & ~n14813 ;
  assign n14815 = n14811 & n14814 ;
  assign n14816 = \wishbone_bd_ram_mem3_reg[96][30]/P0001  & n13425 ;
  assign n14817 = \wishbone_bd_ram_mem3_reg[190][30]/P0001  & n13365 ;
  assign n14818 = ~n14816 & ~n14817 ;
  assign n14819 = \wishbone_bd_ram_mem3_reg[92][30]/P0001  & n13859 ;
  assign n14820 = \wishbone_bd_ram_mem3_reg[117][30]/P0001  & n13557 ;
  assign n14821 = ~n14819 & ~n14820 ;
  assign n14822 = n14818 & n14821 ;
  assign n14823 = n14815 & n14822 ;
  assign n14824 = n14808 & n14823 ;
  assign n14825 = \wishbone_bd_ram_mem3_reg[47][30]/P0001  & n13436 ;
  assign n14826 = \wishbone_bd_ram_mem3_reg[54][30]/P0001  & n13622 ;
  assign n14827 = ~n14825 & ~n14826 ;
  assign n14828 = \wishbone_bd_ram_mem3_reg[139][30]/P0001  & n13566 ;
  assign n14829 = \wishbone_bd_ram_mem3_reg[239][30]/P0001  & n13349 ;
  assign n14830 = ~n14828 & ~n14829 ;
  assign n14831 = n14827 & n14830 ;
  assign n14832 = \wishbone_bd_ram_mem3_reg[59][30]/P0001  & n13613 ;
  assign n14833 = \wishbone_bd_ram_mem3_reg[134][30]/P0001  & n13494 ;
  assign n14834 = ~n14832 & ~n14833 ;
  assign n14835 = \wishbone_bd_ram_mem3_reg[23][30]/P0001  & n13857 ;
  assign n14836 = \wishbone_bd_ram_mem3_reg[142][30]/P0001  & n13448 ;
  assign n14837 = ~n14835 & ~n14836 ;
  assign n14838 = n14834 & n14837 ;
  assign n14839 = n14831 & n14838 ;
  assign n14840 = \wishbone_bd_ram_mem3_reg[179][30]/P0001  & n14035 ;
  assign n14841 = \wishbone_bd_ram_mem3_reg[53][30]/P0001  & n13875 ;
  assign n14842 = ~n14840 & ~n14841 ;
  assign n14843 = \wishbone_bd_ram_mem3_reg[6][30]/P0001  & n13915 ;
  assign n14844 = \wishbone_bd_ram_mem3_reg[254][30]/P0001  & n13283 ;
  assign n14845 = ~n14843 & ~n14844 ;
  assign n14846 = n14842 & n14845 ;
  assign n14847 = \wishbone_bd_ram_mem3_reg[243][30]/P0001  & n13575 ;
  assign n14848 = \wishbone_bd_ram_mem3_reg[219][30]/P0001  & n13577 ;
  assign n14849 = ~n14847 & ~n14848 ;
  assign n14850 = \wishbone_bd_ram_mem3_reg[189][30]/P0001  & n14001 ;
  assign n14851 = \wishbone_bd_ram_mem3_reg[141][30]/P0001  & n13852 ;
  assign n14852 = ~n14850 & ~n14851 ;
  assign n14853 = n14849 & n14852 ;
  assign n14854 = n14846 & n14853 ;
  assign n14855 = n14839 & n14854 ;
  assign n14856 = n14824 & n14855 ;
  assign n14857 = n14793 & n14856 ;
  assign n14858 = n14730 & n14857 ;
  assign n14859 = \wishbone_bd_ram_mem3_reg[42][30]/P0001  & n13341 ;
  assign n14860 = \wishbone_bd_ram_mem3_reg[128][30]/P0001  & n13652 ;
  assign n14861 = ~n14859 & ~n14860 ;
  assign n14862 = \wishbone_bd_ram_mem3_reg[137][30]/P0001  & n13808 ;
  assign n14863 = \wishbone_bd_ram_mem3_reg[251][30]/P0001  & n14019 ;
  assign n14864 = ~n14862 & ~n14863 ;
  assign n14865 = n14861 & n14864 ;
  assign n14866 = \wishbone_bd_ram_mem3_reg[85][30]/P0001  & n13784 ;
  assign n14867 = \wishbone_bd_ram_mem3_reg[2][30]/P0001  & n13975 ;
  assign n14868 = ~n14866 & ~n14867 ;
  assign n14869 = \wishbone_bd_ram_mem3_reg[238][30]/P0001  & n13819 ;
  assign n14870 = \wishbone_bd_ram_mem3_reg[218][30]/P0001  & n13792 ;
  assign n14871 = ~n14869 & ~n14870 ;
  assign n14872 = n14868 & n14871 ;
  assign n14873 = n14865 & n14872 ;
  assign n14874 = \wishbone_bd_ram_mem3_reg[108][30]/P0001  & n13814 ;
  assign n14875 = \wishbone_bd_ram_mem3_reg[21][30]/P0001  & n13438 ;
  assign n14876 = ~n14874 & ~n14875 ;
  assign n14877 = \wishbone_bd_ram_mem3_reg[114][30]/P0001  & n13763 ;
  assign n14878 = \wishbone_bd_ram_mem3_reg[155][30]/P0001  & n13738 ;
  assign n14879 = ~n14877 & ~n14878 ;
  assign n14880 = n14876 & n14879 ;
  assign n14881 = \wishbone_bd_ram_mem3_reg[80][30]/P0001  & n13516 ;
  assign n14882 = \wishbone_bd_ram_mem3_reg[231][30]/P0001  & n13363 ;
  assign n14883 = ~n14881 & ~n14882 ;
  assign n14884 = \wishbone_bd_ram_mem3_reg[198][30]/P0001  & n13592 ;
  assign n14885 = \wishbone_bd_ram_mem3_reg[25][30]/P0001  & n13742 ;
  assign n14886 = ~n14884 & ~n14885 ;
  assign n14887 = n14883 & n14886 ;
  assign n14888 = n14880 & n14887 ;
  assign n14889 = n14873 & n14888 ;
  assign n14890 = \wishbone_bd_ram_mem3_reg[245][30]/P0001  & n13877 ;
  assign n14891 = \wishbone_bd_ram_mem3_reg[17][30]/P0001  & n13324 ;
  assign n14892 = ~n14890 & ~n14891 ;
  assign n14893 = \wishbone_bd_ram_mem3_reg[69][30]/P0001  & n13487 ;
  assign n14894 = \wishbone_bd_ram_mem3_reg[160][30]/P0001  & n13271 ;
  assign n14895 = ~n14893 & ~n14894 ;
  assign n14896 = n14892 & n14895 ;
  assign n14897 = \wishbone_bd_ram_mem3_reg[201][30]/P0001  & n13600 ;
  assign n14898 = \wishbone_bd_ram_mem3_reg[167][30]/P0001  & n13940 ;
  assign n14899 = ~n14897 & ~n14898 ;
  assign n14900 = \wishbone_bd_ram_mem3_reg[105][30]/P0001  & n13503 ;
  assign n14901 = \wishbone_bd_ram_mem3_reg[111][30]/P0001  & n13471 ;
  assign n14902 = ~n14900 & ~n14901 ;
  assign n14903 = n14899 & n14902 ;
  assign n14904 = n14896 & n14903 ;
  assign n14905 = \wishbone_bd_ram_mem3_reg[223][30]/P0001  & n13335 ;
  assign n14906 = \wishbone_bd_ram_mem3_reg[30][30]/P0001  & n13713 ;
  assign n14907 = ~n14905 & ~n14906 ;
  assign n14908 = \wishbone_bd_ram_mem3_reg[165][30]/P0001  & n14028 ;
  assign n14909 = \wishbone_bd_ram_mem3_reg[70][30]/P0001  & n13339 ;
  assign n14910 = ~n14908 & ~n14909 ;
  assign n14911 = n14907 & n14910 ;
  assign n14912 = \wishbone_bd_ram_mem3_reg[51][30]/P0001  & n13880 ;
  assign n14913 = \wishbone_bd_ram_mem3_reg[81][30]/P0001  & n13409 ;
  assign n14914 = ~n14912 & ~n14913 ;
  assign n14915 = \wishbone_bd_ram_mem3_reg[76][30]/P0001  & n13831 ;
  assign n14916 = \wishbone_bd_ram_mem3_reg[159][30]/P0001  & n13627 ;
  assign n14917 = ~n14915 & ~n14916 ;
  assign n14918 = n14914 & n14917 ;
  assign n14919 = n14911 & n14918 ;
  assign n14920 = n14904 & n14919 ;
  assign n14921 = n14889 & n14920 ;
  assign n14922 = \wishbone_bd_ram_mem3_reg[214][30]/P0001  & n13938 ;
  assign n14923 = \wishbone_bd_ram_mem3_reg[172][30]/P0001  & n13377 ;
  assign n14924 = ~n14922 & ~n14923 ;
  assign n14925 = \wishbone_bd_ram_mem3_reg[24][30]/P0001  & n13970 ;
  assign n14926 = \wishbone_bd_ram_mem3_reg[170][30]/P0001  & n14007 ;
  assign n14927 = ~n14925 & ~n14926 ;
  assign n14928 = n14924 & n14927 ;
  assign n14929 = \wishbone_bd_ram_mem3_reg[240][30]/P0001  & n13352 ;
  assign n14930 = \wishbone_bd_ram_mem3_reg[151][30]/P0001  & n13697 ;
  assign n14931 = ~n14929 & ~n14930 ;
  assign n14932 = \wishbone_bd_ram_mem3_reg[195][30]/P0001  & n13700 ;
  assign n14933 = \wishbone_bd_ram_mem3_reg[46][30]/P0001  & n13298 ;
  assign n14934 = ~n14932 & ~n14933 ;
  assign n14935 = n14931 & n14934 ;
  assign n14936 = n14928 & n14935 ;
  assign n14937 = \wishbone_bd_ram_mem3_reg[44][30]/P0001  & n13291 ;
  assign n14938 = \wishbone_bd_ram_mem3_reg[133][30]/P0001  & n13492 ;
  assign n14939 = ~n14937 & ~n14938 ;
  assign n14940 = \wishbone_bd_ram_mem3_reg[57][30]/P0001  & n13731 ;
  assign n14941 = \wishbone_bd_ram_mem3_reg[106][30]/P0001  & n13555 ;
  assign n14942 = ~n14940 & ~n14941 ;
  assign n14943 = n14939 & n14942 ;
  assign n14944 = \wishbone_bd_ram_mem3_reg[161][30]/P0001  & n13505 ;
  assign n14945 = \wishbone_bd_ram_mem3_reg[99][30]/P0001  & n13996 ;
  assign n14946 = ~n14944 & ~n14945 ;
  assign n14947 = \wishbone_bd_ram_mem3_reg[101][30]/P0001  & n13772 ;
  assign n14948 = \wishbone_bd_ram_mem3_reg[233][30]/P0001  & n13332 ;
  assign n14949 = ~n14947 & ~n14948 ;
  assign n14950 = n14946 & n14949 ;
  assign n14951 = n14943 & n14950 ;
  assign n14952 = n14936 & n14951 ;
  assign n14953 = \wishbone_bd_ram_mem3_reg[113][30]/P0001  & n13882 ;
  assign n14954 = \wishbone_bd_ram_mem3_reg[197][30]/P0001  & n13594 ;
  assign n14955 = ~n14953 & ~n14954 ;
  assign n14956 = \wishbone_bd_ram_mem3_reg[152][30]/P0001  & n13912 ;
  assign n14957 = \wishbone_bd_ram_mem3_reg[22][30]/P0001  & n13744 ;
  assign n14958 = ~n14956 & ~n14957 ;
  assign n14959 = n14955 & n14958 ;
  assign n14960 = \wishbone_bd_ram_mem3_reg[84][30]/P0001  & n13385 ;
  assign n14961 = \wishbone_bd_ram_mem3_reg[244][30]/P0001  & n13474 ;
  assign n14962 = ~n14960 & ~n14961 ;
  assign n14963 = \wishbone_bd_ram_mem3_reg[221][30]/P0001  & n13641 ;
  assign n14964 = \wishbone_bd_ram_mem3_reg[203][30]/P0001  & n13816 ;
  assign n14965 = ~n14963 & ~n14964 ;
  assign n14966 = n14962 & n14965 ;
  assign n14967 = n14959 & n14966 ;
  assign n14968 = \wishbone_bd_ram_mem3_reg[253][30]/P0001  & n13708 ;
  assign n14969 = \wishbone_bd_ram_mem3_reg[79][30]/P0001  & n13779 ;
  assign n14970 = ~n14968 & ~n14969 ;
  assign n14971 = \wishbone_bd_ram_mem3_reg[55][30]/P0001  & n13618 ;
  assign n14972 = \wishbone_bd_ram_mem3_reg[222][30]/P0001  & n13721 ;
  assign n14973 = ~n14971 & ~n14972 ;
  assign n14974 = n14970 & n14973 ;
  assign n14975 = \wishbone_bd_ram_mem3_reg[48][30]/P0001  & n13917 ;
  assign n14976 = \wishbone_bd_ram_mem3_reg[52][30]/P0001  & n13988 ;
  assign n14977 = ~n14975 & ~n14976 ;
  assign n14978 = \wishbone_bd_ram_mem3_reg[5][30]/P0001  & n13243 ;
  assign n14979 = \wishbone_bd_ram_mem3_reg[78][30]/P0001  & n13277 ;
  assign n14980 = ~n14978 & ~n14979 ;
  assign n14981 = n14977 & n14980 ;
  assign n14982 = n14974 & n14981 ;
  assign n14983 = n14967 & n14982 ;
  assign n14984 = n14952 & n14983 ;
  assign n14985 = n14921 & n14984 ;
  assign n14986 = \wishbone_bd_ram_mem3_reg[29][30]/P0001  & n13412 ;
  assign n14987 = \wishbone_bd_ram_mem3_reg[184][30]/P0001  & n13960 ;
  assign n14988 = ~n14986 & ~n14987 ;
  assign n14989 = \wishbone_bd_ram_mem3_reg[82][30]/P0001  & n13374 ;
  assign n14990 = \wishbone_bd_ram_mem3_reg[63][30]/P0001  & n13327 ;
  assign n14991 = ~n14989 & ~n14990 ;
  assign n14992 = n14988 & n14991 ;
  assign n14993 = \wishbone_bd_ram_mem3_reg[143][30]/P0001  & n13461 ;
  assign n14994 = \wishbone_bd_ram_mem3_reg[75][30]/P0001  & n13605 ;
  assign n14995 = ~n14993 & ~n14994 ;
  assign n14996 = \wishbone_bd_ram_mem3_reg[118][30]/P0001  & n13589 ;
  assign n14997 = \wishbone_bd_ram_mem3_reg[194][30]/P0001  & n13624 ;
  assign n14998 = ~n14996 & ~n14997 ;
  assign n14999 = n14995 & n14998 ;
  assign n15000 = n14992 & n14999 ;
  assign n15001 = \wishbone_bd_ram_mem3_reg[45][30]/P0001  & n13420 ;
  assign n15002 = \wishbone_bd_ram_mem3_reg[225][30]/P0001  & n13719 ;
  assign n15003 = ~n15001 & ~n15002 ;
  assign n15004 = \wishbone_bd_ram_mem3_reg[35][30]/P0001  & n13523 ;
  assign n15005 = \wishbone_bd_ram_mem3_reg[127][30]/P0001  & n13803 ;
  assign n15006 = ~n15004 & ~n15005 ;
  assign n15007 = n15003 & n15006 ;
  assign n15008 = \wishbone_bd_ram_mem3_reg[115][30]/P0001  & n13747 ;
  assign n15009 = \wishbone_bd_ram_mem3_reg[37][30]/P0001  & n13710 ;
  assign n15010 = ~n15008 & ~n15009 ;
  assign n15011 = \wishbone_bd_ram_mem3_reg[7][30]/P0001  & n13546 ;
  assign n15012 = \wishbone_bd_ram_mem3_reg[68][30]/P0001  & n13379 ;
  assign n15013 = ~n15011 & ~n15012 ;
  assign n15014 = n15010 & n15013 ;
  assign n15015 = n15007 & n15014 ;
  assign n15016 = n15000 & n15015 ;
  assign n15017 = \wishbone_bd_ram_mem3_reg[121][30]/P0001  & n13983 ;
  assign n15018 = \wishbone_bd_ram_mem3_reg[11][30]/P0001  & n13774 ;
  assign n15019 = ~n15017 & ~n15018 ;
  assign n15020 = \wishbone_bd_ram_mem3_reg[49][30]/P0001  & n13929 ;
  assign n15021 = \wishbone_bd_ram_mem3_reg[145][30]/P0001  & n13715 ;
  assign n15022 = ~n15020 & ~n15021 ;
  assign n15023 = n15019 & n15022 ;
  assign n15024 = \wishbone_bd_ram_mem3_reg[125][30]/P0001  & n13396 ;
  assign n15025 = \wishbone_bd_ram_mem3_reg[122][30]/P0001  & n13679 ;
  assign n15026 = ~n15024 & ~n15025 ;
  assign n15027 = \wishbone_bd_ram_mem3_reg[147][30]/P0001  & n13702 ;
  assign n15028 = \wishbone_bd_ram_mem3_reg[31][30]/P0001  & n13758 ;
  assign n15029 = ~n15027 & ~n15028 ;
  assign n15030 = n15026 & n15029 ;
  assign n15031 = n15023 & n15030 ;
  assign n15032 = \wishbone_bd_ram_mem3_reg[220][30]/P0001  & n13965 ;
  assign n15033 = \wishbone_bd_ram_mem3_reg[188][30]/P0001  & n13407 ;
  assign n15034 = ~n15032 & ~n15033 ;
  assign n15035 = \wishbone_bd_ram_mem3_reg[12][30]/P0001  & n13733 ;
  assign n15036 = \wishbone_bd_ram_mem3_reg[38][30]/P0001  & n13828 ;
  assign n15037 = ~n15035 & ~n15036 ;
  assign n15038 = n15034 & n15037 ;
  assign n15039 = \wishbone_bd_ram_mem3_reg[8][30]/P0001  & n13459 ;
  assign n15040 = \wishbone_bd_ram_mem3_reg[39][30]/P0001  & n13893 ;
  assign n15041 = ~n15039 & ~n15040 ;
  assign n15042 = \wishbone_bd_ram_mem3_reg[246][30]/P0001  & n13981 ;
  assign n15043 = \wishbone_bd_ram_mem3_reg[138][30]/P0001  & n13398 ;
  assign n15044 = ~n15042 & ~n15043 ;
  assign n15045 = n15041 & n15044 ;
  assign n15046 = n15038 & n15045 ;
  assign n15047 = n15031 & n15046 ;
  assign n15048 = n15016 & n15047 ;
  assign n15049 = \wishbone_bd_ram_mem3_reg[209][30]/P0001  & n13689 ;
  assign n15050 = \wishbone_bd_ram_mem3_reg[4][30]/P0001  & n13527 ;
  assign n15051 = ~n15049 & ~n15050 ;
  assign n15052 = \wishbone_bd_ram_mem3_reg[191][30]/P0001  & n14012 ;
  assign n15053 = \wishbone_bd_ram_mem3_reg[228][30]/P0001  & n13497 ;
  assign n15054 = ~n15052 & ~n15053 ;
  assign n15055 = n15051 & n15054 ;
  assign n15056 = \wishbone_bd_ram_mem3_reg[120][30]/P0001  & n13550 ;
  assign n15057 = \wishbone_bd_ram_mem3_reg[202][30]/P0001  & n13268 ;
  assign n15058 = ~n15056 & ~n15057 ;
  assign n15059 = \wishbone_bd_ram_mem3_reg[168][30]/P0001  & n13795 ;
  assign n15060 = \wishbone_bd_ram_mem3_reg[247][30]/P0001  & n13571 ;
  assign n15061 = ~n15059 & ~n15060 ;
  assign n15062 = n15058 & n15061 ;
  assign n15063 = n15055 & n15062 ;
  assign n15064 = \wishbone_bd_ram_mem3_reg[88][30]/P0001  & n13347 ;
  assign n15065 = \wishbone_bd_ram_mem3_reg[41][30]/P0001  & n14017 ;
  assign n15066 = ~n15064 & ~n15065 ;
  assign n15067 = \wishbone_bd_ram_mem3_reg[40][30]/P0001  & n13661 ;
  assign n15068 = \wishbone_bd_ram_mem3_reg[94][30]/P0001  & n13833 ;
  assign n15069 = ~n15067 & ~n15068 ;
  assign n15070 = n15066 & n15069 ;
  assign n15071 = \wishbone_bd_ram_mem3_reg[217][30]/P0001  & n13767 ;
  assign n15072 = \wishbone_bd_ram_mem3_reg[62][30]/P0001  & n13529 ;
  assign n15073 = ~n15071 & ~n15072 ;
  assign n15074 = \wishbone_bd_ram_mem3_reg[207][30]/P0001  & n13826 ;
  assign n15075 = \wishbone_bd_ram_mem3_reg[16][30]/P0001  & n13695 ;
  assign n15076 = ~n15074 & ~n15075 ;
  assign n15077 = n15073 & n15076 ;
  assign n15078 = n15070 & n15077 ;
  assign n15079 = n15063 & n15078 ;
  assign n15080 = \wishbone_bd_ram_mem3_reg[171][30]/P0001  & n13422 ;
  assign n15081 = \wishbone_bd_ram_mem3_reg[150][30]/P0001  & n13666 ;
  assign n15082 = ~n15080 & ~n15081 ;
  assign n15083 = \wishbone_bd_ram_mem3_reg[95][30]/P0001  & n13317 ;
  assign n15084 = \wishbone_bd_ram_mem3_reg[90][30]/P0001  & n13906 ;
  assign n15085 = ~n15083 & ~n15084 ;
  assign n15086 = n15082 & n15085 ;
  assign n15087 = \wishbone_bd_ram_mem3_reg[248][30]/P0001  & n13647 ;
  assign n15088 = \wishbone_bd_ram_mem3_reg[126][30]/P0001  & n13786 ;
  assign n15089 = ~n15087 & ~n15088 ;
  assign n15090 = \wishbone_bd_ram_mem3_reg[93][30]/P0001  & n13891 ;
  assign n15091 = \wishbone_bd_ram_mem3_reg[140][30]/P0001  & n13287 ;
  assign n15092 = ~n15090 & ~n15091 ;
  assign n15093 = n15089 & n15092 ;
  assign n15094 = n15086 & n15093 ;
  assign n15095 = \wishbone_bd_ram_mem3_reg[14][30]/P0001  & n13972 ;
  assign n15096 = \wishbone_bd_ram_mem3_reg[249][30]/P0001  & n13431 ;
  assign n15097 = ~n15095 & ~n15096 ;
  assign n15098 = \wishbone_bd_ram_mem3_reg[162][30]/P0001  & n13726 ;
  assign n15099 = \wishbone_bd_ram_mem3_reg[110][30]/P0001  & n14030 ;
  assign n15100 = ~n15098 & ~n15099 ;
  assign n15101 = n15097 & n15100 ;
  assign n15102 = \wishbone_bd_ram_mem3_reg[71][30]/P0001  & n13636 ;
  assign n15103 = \wishbone_bd_ram_mem3_reg[124][30]/P0001  & n14024 ;
  assign n15104 = ~n15102 & ~n15103 ;
  assign n15105 = \wishbone_bd_ram_mem3_reg[65][30]/P0001  & n13842 ;
  assign n15106 = \wishbone_bd_ram_mem3_reg[177][30]/P0001  & n13863 ;
  assign n15107 = ~n15105 & ~n15106 ;
  assign n15108 = n15104 & n15107 ;
  assign n15109 = n15101 & n15108 ;
  assign n15110 = n15094 & n15109 ;
  assign n15111 = n15079 & n15110 ;
  assign n15112 = n15048 & n15111 ;
  assign n15113 = n14985 & n15112 ;
  assign n15114 = n14858 & n15113 ;
  assign n15115 = n14047 & ~n15114 ;
  assign n15116 = ~\wishbone_TxLength_reg[14]/NET0131  & ~n14601 ;
  assign n15117 = n14066 & ~n14600 ;
  assign n15118 = \wishbone_TxLength_reg[14]/NET0131  & ~n14595 ;
  assign n15119 = ~n15117 & n15118 ;
  assign n15120 = ~n15116 & ~n15119 ;
  assign n15121 = ~n15115 & ~n15120 ;
  assign n15122 = ~\rxethmac1_crcrx_Crc_reg[6]/NET0131  & n10663 ;
  assign n15123 = ~n12567 & n15122 ;
  assign n15124 = \rxethmac1_crcrx_Crc_reg[6]/NET0131  & n10663 ;
  assign n15125 = n12567 & n15124 ;
  assign n15126 = ~n15123 & ~n15125 ;
  assign n15127 = ~\rxethmac1_crcrx_Crc_reg[0]/NET0131  & n10663 ;
  assign n15128 = ~n12567 & n15127 ;
  assign n15129 = \rxethmac1_crcrx_Crc_reg[0]/NET0131  & n10663 ;
  assign n15130 = n12567 & n15129 ;
  assign n15131 = ~n15128 & ~n15130 ;
  assign n15132 = \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  & ~n11167 ;
  assign n15133 = ~\txethmac1_txstatem1_StateData_reg[1]/NET0131  & ~n15132 ;
  assign n15134 = ~n11128 & n15133 ;
  assign n15135 = \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n15136 = \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n15137 = \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  & n15136 ;
  assign n15138 = n15135 & n15137 ;
  assign n15139 = \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n15140 = \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n15141 = n15139 & n15140 ;
  assign n15142 = \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n15143 = \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  & n15142 ;
  assign n15144 = n15141 & n15143 ;
  assign n15145 = n15138 & n15144 ;
  assign n15146 = \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n15147 = \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  ;
  assign n15148 = n15146 & n15147 ;
  assign n15149 = ~n11128 & n15148 ;
  assign n15150 = n15145 & n15149 ;
  assign n15151 = ~n15134 & ~n15150 ;
  assign n15152 = \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n15153 = \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  & n15152 ;
  assign n15154 = n15151 & n15153 ;
  assign n15155 = \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
  assign n15156 = n15138 & n15155 ;
  assign n15157 = n15154 & n15156 ;
  assign n15158 = \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  & n15146 ;
  assign n15159 = n15142 & n15158 ;
  assign n15160 = n15157 & n15159 ;
  assign n15161 = ~\txethmac1_PacketFinished_q_reg/NET0131  & n11347 ;
  assign n15162 = ~n11392 & n15161 ;
  assign n15163 = \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  & n15162 ;
  assign n15164 = ~n15160 & n15163 ;
  assign n15165 = ~\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  & n15162 ;
  assign n15166 = n15160 & n15165 ;
  assign n15167 = ~n15164 & ~n15166 ;
  assign n15168 = \wishbone_TxPointerMSB_reg[2]/NET0131  & ~n13201 ;
  assign n15169 = \m_wb_adr_o[2]_pad  & ~n13203 ;
  assign n15170 = ~n13195 & n15169 ;
  assign n15171 = ~n13196 & ~n15170 ;
  assign n15172 = \wishbone_RxPointerMSB_reg[2]/NET0131  & n15171 ;
  assign n15173 = ~n15168 & ~n15172 ;
  assign n15174 = ~n13149 & ~n13203 ;
  assign n15175 = n13143 & n15174 ;
  assign n15176 = n13137 & n15175 ;
  assign n15177 = ~n13170 & ~n15176 ;
  assign n15178 = \wishbone_TxPointerMSB_reg[2]/NET0131  & ~n13166 ;
  assign n15179 = ~n13164 & n15178 ;
  assign n15180 = n15177 & ~n15179 ;
  assign n15181 = ~\m_wb_adr_o[2]_pad  & ~n15180 ;
  assign n15182 = \m_wb_adr_o[2]_pad  & n13197 ;
  assign n15183 = ~n15181 & ~n15182 ;
  assign n15184 = n15173 & n15183 ;
  assign n15185 = \wishbone_bd_ram_mem3_reg[143][24]/P0001  & n13461 ;
  assign n15186 = \wishbone_bd_ram_mem3_reg[8][24]/P0001  & n13459 ;
  assign n15187 = ~n15185 & ~n15186 ;
  assign n15188 = \wishbone_bd_ram_mem3_reg[142][24]/P0001  & n13448 ;
  assign n15189 = \wishbone_bd_ram_mem3_reg[115][24]/P0001  & n13747 ;
  assign n15190 = ~n15188 & ~n15189 ;
  assign n15191 = n15187 & n15190 ;
  assign n15192 = \wishbone_bd_ram_mem3_reg[111][24]/P0001  & n13471 ;
  assign n15193 = \wishbone_bd_ram_mem3_reg[228][24]/P0001  & n13497 ;
  assign n15194 = ~n15192 & ~n15193 ;
  assign n15195 = \wishbone_bd_ram_mem3_reg[47][24]/P0001  & n13436 ;
  assign n15196 = \wishbone_bd_ram_mem3_reg[185][24]/P0001  & n13372 ;
  assign n15197 = ~n15195 & ~n15196 ;
  assign n15198 = n15194 & n15197 ;
  assign n15199 = n15191 & n15198 ;
  assign n15200 = \wishbone_bd_ram_mem3_reg[249][24]/P0001  & n13431 ;
  assign n15201 = \wishbone_bd_ram_mem3_reg[106][24]/P0001  & n13555 ;
  assign n15202 = ~n15200 & ~n15201 ;
  assign n15203 = \wishbone_bd_ram_mem3_reg[65][24]/P0001  & n13842 ;
  assign n15204 = \wishbone_bd_ram_mem3_reg[150][24]/P0001  & n13666 ;
  assign n15205 = ~n15203 & ~n15204 ;
  assign n15206 = n15202 & n15205 ;
  assign n15207 = \wishbone_bd_ram_mem3_reg[154][24]/P0001  & n13403 ;
  assign n15208 = \wishbone_bd_ram_mem3_reg[129][24]/P0001  & n13629 ;
  assign n15209 = ~n15207 & ~n15208 ;
  assign n15210 = \wishbone_bd_ram_mem3_reg[172][24]/P0001  & n13377 ;
  assign n15211 = \wishbone_bd_ram_mem3_reg[28][24]/P0001  & n13810 ;
  assign n15212 = ~n15210 & ~n15211 ;
  assign n15213 = n15209 & n15212 ;
  assign n15214 = n15206 & n15213 ;
  assign n15215 = n15199 & n15214 ;
  assign n15216 = \wishbone_bd_ram_mem3_reg[171][24]/P0001  & n13422 ;
  assign n15217 = \wishbone_bd_ram_mem3_reg[40][24]/P0001  & n13661 ;
  assign n15218 = ~n15216 & ~n15217 ;
  assign n15219 = \wishbone_bd_ram_mem3_reg[2][24]/P0001  & n13975 ;
  assign n15220 = \wishbone_bd_ram_mem3_reg[75][24]/P0001  & n13605 ;
  assign n15221 = ~n15219 & ~n15220 ;
  assign n15222 = n15218 & n15221 ;
  assign n15223 = \wishbone_bd_ram_mem3_reg[181][24]/P0001  & n13587 ;
  assign n15224 = \wishbone_bd_ram_mem3_reg[244][24]/P0001  & n13474 ;
  assign n15225 = ~n15223 & ~n15224 ;
  assign n15226 = \wishbone_bd_ram_mem3_reg[109][24]/P0001  & n13306 ;
  assign n15227 = \wishbone_bd_ram_mem3_reg[88][24]/P0001  & n13347 ;
  assign n15228 = ~n15226 & ~n15227 ;
  assign n15229 = n15225 & n15228 ;
  assign n15230 = n15222 & n15229 ;
  assign n15231 = \wishbone_bd_ram_mem3_reg[120][24]/P0001  & n13550 ;
  assign n15232 = \wishbone_bd_ram_mem3_reg[250][24]/P0001  & n13677 ;
  assign n15233 = ~n15231 & ~n15232 ;
  assign n15234 = \wishbone_bd_ram_mem3_reg[215][24]/P0001  & n13901 ;
  assign n15235 = \wishbone_bd_ram_mem3_reg[67][24]/P0001  & n13663 ;
  assign n15236 = ~n15234 & ~n15235 ;
  assign n15237 = n15233 & n15236 ;
  assign n15238 = \wishbone_bd_ram_mem3_reg[80][24]/P0001  & n13516 ;
  assign n15239 = \wishbone_bd_ram_mem3_reg[140][24]/P0001  & n13287 ;
  assign n15240 = ~n15238 & ~n15239 ;
  assign n15241 = \wishbone_bd_ram_mem3_reg[160][24]/P0001  & n13271 ;
  assign n15242 = \wishbone_bd_ram_mem3_reg[219][24]/P0001  & n13577 ;
  assign n15243 = ~n15241 & ~n15242 ;
  assign n15244 = n15240 & n15243 ;
  assign n15245 = n15237 & n15244 ;
  assign n15246 = n15230 & n15245 ;
  assign n15247 = n15215 & n15246 ;
  assign n15248 = \wishbone_bd_ram_mem3_reg[212][24]/P0001  & n13634 ;
  assign n15249 = \wishbone_bd_ram_mem3_reg[10][24]/P0001  & n13837 ;
  assign n15250 = ~n15248 & ~n15249 ;
  assign n15251 = \wishbone_bd_ram_mem3_reg[139][24]/P0001  & n13566 ;
  assign n15252 = \wishbone_bd_ram_mem3_reg[30][24]/P0001  & n13713 ;
  assign n15253 = ~n15251 & ~n15252 ;
  assign n15254 = n15250 & n15253 ;
  assign n15255 = \wishbone_bd_ram_mem3_reg[247][24]/P0001  & n13571 ;
  assign n15256 = \wishbone_bd_ram_mem3_reg[29][24]/P0001  & n13412 ;
  assign n15257 = ~n15255 & ~n15256 ;
  assign n15258 = \wishbone_bd_ram_mem3_reg[216][24]/P0001  & n14005 ;
  assign n15259 = \wishbone_bd_ram_mem3_reg[145][24]/P0001  & n13715 ;
  assign n15260 = ~n15258 & ~n15259 ;
  assign n15261 = n15257 & n15260 ;
  assign n15262 = n15254 & n15261 ;
  assign n15263 = \wishbone_bd_ram_mem3_reg[192][24]/P0001  & n13390 ;
  assign n15264 = \wishbone_bd_ram_mem3_reg[162][24]/P0001  & n13726 ;
  assign n15265 = ~n15263 & ~n15264 ;
  assign n15266 = \wishbone_bd_ram_mem3_reg[36][24]/P0001  & n13639 ;
  assign n15267 = \wishbone_bd_ram_mem3_reg[9][24]/P0001  & n13580 ;
  assign n15268 = ~n15266 & ~n15267 ;
  assign n15269 = n15265 & n15268 ;
  assign n15270 = \wishbone_bd_ram_mem3_reg[132][24]/P0001  & n13927 ;
  assign n15271 = \wishbone_bd_ram_mem3_reg[187][24]/P0001  & n13756 ;
  assign n15272 = ~n15270 & ~n15271 ;
  assign n15273 = \wishbone_bd_ram_mem3_reg[43][24]/P0001  & n13761 ;
  assign n15274 = \wishbone_bd_ram_mem3_reg[239][24]/P0001  & n13349 ;
  assign n15275 = ~n15273 & ~n15274 ;
  assign n15276 = n15272 & n15275 ;
  assign n15277 = n15269 & n15276 ;
  assign n15278 = n15262 & n15277 ;
  assign n15279 = \wishbone_bd_ram_mem3_reg[168][24]/P0001  & n13795 ;
  assign n15280 = \wishbone_bd_ram_mem3_reg[182][24]/P0001  & n13598 ;
  assign n15281 = ~n15279 & ~n15280 ;
  assign n15282 = \wishbone_bd_ram_mem3_reg[230][24]/P0001  & n13994 ;
  assign n15283 = \wishbone_bd_ram_mem3_reg[21][24]/P0001  & n13438 ;
  assign n15284 = ~n15282 & ~n15283 ;
  assign n15285 = n15281 & n15284 ;
  assign n15286 = \wishbone_bd_ram_mem3_reg[178][24]/P0001  & n13301 ;
  assign n15287 = \wishbone_bd_ram_mem3_reg[127][24]/P0001  & n13803 ;
  assign n15288 = ~n15286 & ~n15287 ;
  assign n15289 = \wishbone_bd_ram_mem3_reg[60][24]/P0001  & n13790 ;
  assign n15290 = \wishbone_bd_ram_mem3_reg[18][24]/P0001  & n13532 ;
  assign n15291 = ~n15289 & ~n15290 ;
  assign n15292 = n15288 & n15291 ;
  assign n15293 = n15285 & n15292 ;
  assign n15294 = \wishbone_bd_ram_mem3_reg[41][24]/P0001  & n14017 ;
  assign n15295 = \wishbone_bd_ram_mem3_reg[52][24]/P0001  & n13988 ;
  assign n15296 = ~n15294 & ~n15295 ;
  assign n15297 = \wishbone_bd_ram_mem3_reg[147][24]/P0001  & n13702 ;
  assign n15298 = \wishbone_bd_ram_mem3_reg[20][24]/P0001  & n13839 ;
  assign n15299 = ~n15297 & ~n15298 ;
  assign n15300 = n15296 & n15299 ;
  assign n15301 = \wishbone_bd_ram_mem3_reg[22][24]/P0001  & n13744 ;
  assign n15302 = \wishbone_bd_ram_mem3_reg[97][24]/P0001  & n13724 ;
  assign n15303 = ~n15301 & ~n15302 ;
  assign n15304 = \wishbone_bd_ram_mem3_reg[255][24]/P0001  & n13952 ;
  assign n15305 = \wishbone_bd_ram_mem3_reg[164][24]/P0001  & n13236 ;
  assign n15306 = ~n15304 & ~n15305 ;
  assign n15307 = n15303 & n15306 ;
  assign n15308 = n15300 & n15307 ;
  assign n15309 = n15293 & n15308 ;
  assign n15310 = n15278 & n15309 ;
  assign n15311 = n15247 & n15310 ;
  assign n15312 = \wishbone_bd_ram_mem3_reg[201][24]/P0001  & n13600 ;
  assign n15313 = \wishbone_bd_ram_mem3_reg[91][24]/P0001  & n13954 ;
  assign n15314 = ~n15312 & ~n15313 ;
  assign n15315 = \wishbone_bd_ram_mem3_reg[211][24]/P0001  & n13805 ;
  assign n15316 = \wishbone_bd_ram_mem3_reg[149][24]/P0001  & n13469 ;
  assign n15317 = ~n15315 & ~n15316 ;
  assign n15318 = n15314 & n15317 ;
  assign n15319 = \wishbone_bd_ram_mem3_reg[205][24]/P0001  & n13947 ;
  assign n15320 = \wishbone_bd_ram_mem3_reg[176][24]/P0001  & n13262 ;
  assign n15321 = ~n15319 & ~n15320 ;
  assign n15322 = \wishbone_bd_ram_mem3_reg[131][24]/P0001  & n13358 ;
  assign n15323 = \wishbone_bd_ram_mem3_reg[39][24]/P0001  & n13893 ;
  assign n15324 = ~n15322 & ~n15323 ;
  assign n15325 = n15321 & n15324 ;
  assign n15326 = n15318 & n15325 ;
  assign n15327 = \wishbone_bd_ram_mem3_reg[35][24]/P0001  & n13523 ;
  assign n15328 = \wishbone_bd_ram_mem3_reg[218][24]/P0001  & n13792 ;
  assign n15329 = ~n15327 & ~n15328 ;
  assign n15330 = \wishbone_bd_ram_mem3_reg[241][24]/P0001  & n13854 ;
  assign n15331 = \wishbone_bd_ram_mem3_reg[170][24]/P0001  & n14007 ;
  assign n15332 = ~n15330 & ~n15331 ;
  assign n15333 = n15329 & n15332 ;
  assign n15334 = \wishbone_bd_ram_mem3_reg[196][24]/P0001  & n13977 ;
  assign n15335 = \wishbone_bd_ram_mem3_reg[84][24]/P0001  & n13385 ;
  assign n15336 = ~n15334 & ~n15335 ;
  assign n15337 = \wishbone_bd_ram_mem3_reg[121][24]/P0001  & n13983 ;
  assign n15338 = \wishbone_bd_ram_mem3_reg[83][24]/P0001  & n13454 ;
  assign n15339 = ~n15337 & ~n15338 ;
  assign n15340 = n15336 & n15339 ;
  assign n15341 = n15333 & n15340 ;
  assign n15342 = n15326 & n15341 ;
  assign n15343 = \wishbone_bd_ram_mem3_reg[3][24]/P0001  & n13354 ;
  assign n15344 = \wishbone_bd_ram_mem3_reg[126][24]/P0001  & n13786 ;
  assign n15345 = ~n15343 & ~n15344 ;
  assign n15346 = \wishbone_bd_ram_mem3_reg[34][24]/P0001  & n13450 ;
  assign n15347 = \wishbone_bd_ram_mem3_reg[55][24]/P0001  & n13618 ;
  assign n15348 = ~n15346 & ~n15347 ;
  assign n15349 = n15345 & n15348 ;
  assign n15350 = \wishbone_bd_ram_mem3_reg[78][24]/P0001  & n13277 ;
  assign n15351 = \wishbone_bd_ram_mem3_reg[157][24]/P0001  & n13445 ;
  assign n15352 = ~n15350 & ~n15351 ;
  assign n15353 = \wishbone_bd_ram_mem3_reg[17][24]/P0001  & n13324 ;
  assign n15354 = \wishbone_bd_ram_mem3_reg[0][24]/P0001  & n13539 ;
  assign n15355 = ~n15353 & ~n15354 ;
  assign n15356 = n15352 & n15355 ;
  assign n15357 = n15349 & n15356 ;
  assign n15358 = \wishbone_bd_ram_mem3_reg[144][24]/P0001  & n13508 ;
  assign n15359 = \wishbone_bd_ram_mem3_reg[227][24]/P0001  & n13388 ;
  assign n15360 = ~n15358 & ~n15359 ;
  assign n15361 = \wishbone_bd_ram_mem3_reg[57][24]/P0001  & n13731 ;
  assign n15362 = \wishbone_bd_ram_mem3_reg[188][24]/P0001  & n13407 ;
  assign n15363 = ~n15361 & ~n15362 ;
  assign n15364 = n15360 & n15363 ;
  assign n15365 = \wishbone_bd_ram_mem3_reg[104][24]/P0001  & n13684 ;
  assign n15366 = \wishbone_bd_ram_mem3_reg[252][24]/P0001  & n13986 ;
  assign n15367 = ~n15365 & ~n15366 ;
  assign n15368 = \wishbone_bd_ram_mem3_reg[197][24]/P0001  & n13594 ;
  assign n15369 = \wishbone_bd_ram_mem3_reg[137][24]/P0001  & n13808 ;
  assign n15370 = ~n15368 & ~n15369 ;
  assign n15371 = n15367 & n15370 ;
  assign n15372 = n15364 & n15371 ;
  assign n15373 = n15357 & n15372 ;
  assign n15374 = n15342 & n15373 ;
  assign n15375 = \wishbone_bd_ram_mem3_reg[66][24]/P0001  & n13603 ;
  assign n15376 = \wishbone_bd_ram_mem3_reg[105][24]/P0001  & n13503 ;
  assign n15377 = ~n15375 & ~n15376 ;
  assign n15378 = \wishbone_bd_ram_mem3_reg[89][24]/P0001  & n13910 ;
  assign n15379 = \wishbone_bd_ram_mem3_reg[224][24]/P0001  & n13433 ;
  assign n15380 = ~n15378 & ~n15379 ;
  assign n15381 = n15377 & n15380 ;
  assign n15382 = \wishbone_bd_ram_mem3_reg[173][24]/P0001  & n13360 ;
  assign n15383 = \wishbone_bd_ram_mem3_reg[226][24]/P0001  & n13668 ;
  assign n15384 = ~n15382 & ~n15383 ;
  assign n15385 = \wishbone_bd_ram_mem3_reg[204][24]/P0001  & n13821 ;
  assign n15386 = \wishbone_bd_ram_mem3_reg[24][24]/P0001  & n13970 ;
  assign n15387 = ~n15385 & ~n15386 ;
  assign n15388 = n15384 & n15387 ;
  assign n15389 = n15381 & n15388 ;
  assign n15390 = \wishbone_bd_ram_mem3_reg[158][24]/P0001  & n13294 ;
  assign n15391 = \wishbone_bd_ram_mem3_reg[26][24]/P0001  & n13521 ;
  assign n15392 = ~n15390 & ~n15391 ;
  assign n15393 = \wishbone_bd_ram_mem3_reg[165][24]/P0001  & n14028 ;
  assign n15394 = \wishbone_bd_ram_mem3_reg[209][24]/P0001  & n13689 ;
  assign n15395 = ~n15393 & ~n15394 ;
  assign n15396 = n15392 & n15395 ;
  assign n15397 = \wishbone_bd_ram_mem3_reg[90][24]/P0001  & n13906 ;
  assign n15398 = \wishbone_bd_ram_mem3_reg[184][24]/P0001  & n13960 ;
  assign n15399 = ~n15397 & ~n15398 ;
  assign n15400 = \wishbone_bd_ram_mem3_reg[73][24]/P0001  & n13456 ;
  assign n15401 = \wishbone_bd_ram_mem3_reg[31][24]/P0001  & n13758 ;
  assign n15402 = ~n15400 & ~n15401 ;
  assign n15403 = n15399 & n15402 ;
  assign n15404 = n15396 & n15403 ;
  assign n15405 = n15389 & n15404 ;
  assign n15406 = \wishbone_bd_ram_mem3_reg[130][24]/P0001  & n13427 ;
  assign n15407 = \wishbone_bd_ram_mem3_reg[133][24]/P0001  & n13492 ;
  assign n15408 = ~n15406 & ~n15407 ;
  assign n15409 = \wishbone_bd_ram_mem3_reg[152][24]/P0001  & n13912 ;
  assign n15410 = \wishbone_bd_ram_mem3_reg[25][24]/P0001  & n13742 ;
  assign n15411 = ~n15409 & ~n15410 ;
  assign n15412 = n15408 & n15411 ;
  assign n15413 = \wishbone_bd_ram_mem3_reg[100][24]/P0001  & n13401 ;
  assign n15414 = \wishbone_bd_ram_mem3_reg[229][24]/P0001  & n13552 ;
  assign n15415 = ~n15413 & ~n15414 ;
  assign n15416 = \wishbone_bd_ram_mem3_reg[110][24]/P0001  & n14030 ;
  assign n15417 = \wishbone_bd_ram_mem3_reg[99][24]/P0001  & n13996 ;
  assign n15418 = ~n15416 & ~n15417 ;
  assign n15419 = n15415 & n15418 ;
  assign n15420 = n15412 & n15419 ;
  assign n15421 = \wishbone_bd_ram_mem3_reg[114][24]/P0001  & n13763 ;
  assign n15422 = \wishbone_bd_ram_mem3_reg[93][24]/P0001  & n13891 ;
  assign n15423 = ~n15421 & ~n15422 ;
  assign n15424 = \wishbone_bd_ram_mem3_reg[141][24]/P0001  & n13852 ;
  assign n15425 = \wishbone_bd_ram_mem3_reg[146][24]/P0001  & n13958 ;
  assign n15426 = ~n15424 & ~n15425 ;
  assign n15427 = n15423 & n15426 ;
  assign n15428 = \wishbone_bd_ram_mem3_reg[220][24]/P0001  & n13965 ;
  assign n15429 = \wishbone_bd_ram_mem3_reg[245][24]/P0001  & n13877 ;
  assign n15430 = ~n15428 & ~n15429 ;
  assign n15431 = \wishbone_bd_ram_mem3_reg[33][24]/P0001  & n13933 ;
  assign n15432 = \wishbone_bd_ram_mem3_reg[61][24]/P0001  & n13544 ;
  assign n15433 = ~n15431 & ~n15432 ;
  assign n15434 = n15430 & n15433 ;
  assign n15435 = n15427 & n15434 ;
  assign n15436 = n15420 & n15435 ;
  assign n15437 = n15405 & n15436 ;
  assign n15438 = n15374 & n15437 ;
  assign n15439 = n15311 & n15438 ;
  assign n15440 = \wishbone_bd_ram_mem3_reg[153][24]/P0001  & n13309 ;
  assign n15441 = \wishbone_bd_ram_mem3_reg[44][24]/P0001  & n13291 ;
  assign n15442 = ~n15440 & ~n15441 ;
  assign n15443 = \wishbone_bd_ram_mem3_reg[191][24]/P0001  & n14012 ;
  assign n15444 = \wishbone_bd_ram_mem3_reg[217][24]/P0001  & n13767 ;
  assign n15445 = ~n15443 & ~n15444 ;
  assign n15446 = n15442 & n15445 ;
  assign n15447 = \wishbone_bd_ram_mem3_reg[68][24]/P0001  & n13379 ;
  assign n15448 = \wishbone_bd_ram_mem3_reg[38][24]/P0001  & n13828 ;
  assign n15449 = ~n15447 & ~n15448 ;
  assign n15450 = \wishbone_bd_ram_mem3_reg[233][24]/P0001  & n13332 ;
  assign n15451 = \wishbone_bd_ram_mem3_reg[117][24]/P0001  & n13557 ;
  assign n15452 = ~n15450 & ~n15451 ;
  assign n15453 = n15449 & n15452 ;
  assign n15454 = n15446 & n15453 ;
  assign n15455 = \wishbone_bd_ram_mem3_reg[189][24]/P0001  & n14001 ;
  assign n15456 = \wishbone_bd_ram_mem3_reg[180][24]/P0001  & n13650 ;
  assign n15457 = ~n15455 & ~n15456 ;
  assign n15458 = \wishbone_bd_ram_mem3_reg[243][24]/P0001  & n13575 ;
  assign n15459 = \wishbone_bd_ram_mem3_reg[116][24]/P0001  & n13865 ;
  assign n15460 = ~n15458 & ~n15459 ;
  assign n15461 = n15457 & n15460 ;
  assign n15462 = \wishbone_bd_ram_mem3_reg[77][24]/P0001  & n13935 ;
  assign n15463 = \wishbone_bd_ram_mem3_reg[125][24]/P0001  & n13396 ;
  assign n15464 = ~n15462 & ~n15463 ;
  assign n15465 = \wishbone_bd_ram_mem3_reg[237][24]/P0001  & n13924 ;
  assign n15466 = \wishbone_bd_ram_mem3_reg[195][24]/P0001  & n13700 ;
  assign n15467 = ~n15465 & ~n15466 ;
  assign n15468 = n15464 & n15467 ;
  assign n15469 = n15461 & n15468 ;
  assign n15470 = n15454 & n15469 ;
  assign n15471 = \wishbone_bd_ram_mem3_reg[214][24]/P0001  & n13938 ;
  assign n15472 = \wishbone_bd_ram_mem3_reg[177][24]/P0001  & n13863 ;
  assign n15473 = ~n15471 & ~n15472 ;
  assign n15474 = \wishbone_bd_ram_mem3_reg[166][24]/P0001  & n13999 ;
  assign n15475 = \wishbone_bd_ram_mem3_reg[102][24]/P0001  & n13534 ;
  assign n15476 = ~n15474 & ~n15475 ;
  assign n15477 = n15473 & n15476 ;
  assign n15478 = \wishbone_bd_ram_mem3_reg[238][24]/P0001  & n13819 ;
  assign n15479 = \wishbone_bd_ram_mem3_reg[124][24]/P0001  & n14024 ;
  assign n15480 = ~n15478 & ~n15479 ;
  assign n15481 = \wishbone_bd_ram_mem3_reg[234][24]/P0001  & n13781 ;
  assign n15482 = \wishbone_bd_ram_mem3_reg[232][24]/P0001  & n13510 ;
  assign n15483 = ~n15481 & ~n15482 ;
  assign n15484 = n15480 & n15483 ;
  assign n15485 = n15477 & n15484 ;
  assign n15486 = \wishbone_bd_ram_mem3_reg[118][24]/P0001  & n13589 ;
  assign n15487 = \wishbone_bd_ram_mem3_reg[50][24]/P0001  & n13686 ;
  assign n15488 = ~n15486 & ~n15487 ;
  assign n15489 = \wishbone_bd_ram_mem3_reg[81][24]/P0001  & n13409 ;
  assign n15490 = \wishbone_bd_ram_mem3_reg[82][24]/P0001  & n13374 ;
  assign n15491 = ~n15489 & ~n15490 ;
  assign n15492 = n15488 & n15491 ;
  assign n15493 = \wishbone_bd_ram_mem3_reg[11][24]/P0001  & n13774 ;
  assign n15494 = \wishbone_bd_ram_mem3_reg[53][24]/P0001  & n13875 ;
  assign n15495 = ~n15493 & ~n15494 ;
  assign n15496 = \wishbone_bd_ram_mem3_reg[169][24]/P0001  & n13541 ;
  assign n15497 = \wishbone_bd_ram_mem3_reg[59][24]/P0001  & n13613 ;
  assign n15498 = ~n15496 & ~n15497 ;
  assign n15499 = n15495 & n15498 ;
  assign n15500 = n15492 & n15499 ;
  assign n15501 = n15485 & n15500 ;
  assign n15502 = n15470 & n15501 ;
  assign n15503 = \wishbone_bd_ram_mem3_reg[213][24]/P0001  & n13870 ;
  assign n15504 = \wishbone_bd_ram_mem3_reg[76][24]/P0001  & n13831 ;
  assign n15505 = ~n15503 & ~n15504 ;
  assign n15506 = \wishbone_bd_ram_mem3_reg[16][24]/P0001  & n13695 ;
  assign n15507 = \wishbone_bd_ram_mem3_reg[175][24]/P0001  & n13674 ;
  assign n15508 = ~n15506 & ~n15507 ;
  assign n15509 = n15505 & n15508 ;
  assign n15510 = \wishbone_bd_ram_mem3_reg[253][24]/P0001  & n13708 ;
  assign n15511 = \wishbone_bd_ram_mem3_reg[62][24]/P0001  & n13529 ;
  assign n15512 = ~n15510 & ~n15511 ;
  assign n15513 = \wishbone_bd_ram_mem3_reg[122][24]/P0001  & n13679 ;
  assign n15514 = \wishbone_bd_ram_mem3_reg[6][24]/P0001  & n13915 ;
  assign n15515 = ~n15513 & ~n15514 ;
  assign n15516 = n15512 & n15515 ;
  assign n15517 = n15509 & n15516 ;
  assign n15518 = \wishbone_bd_ram_mem3_reg[13][24]/P0001  & n13844 ;
  assign n15519 = \wishbone_bd_ram_mem3_reg[193][24]/P0001  & n14022 ;
  assign n15520 = ~n15518 & ~n15519 ;
  assign n15521 = \wishbone_bd_ram_mem3_reg[4][24]/P0001  & n13527 ;
  assign n15522 = \wishbone_bd_ram_mem3_reg[236][24]/P0001  & n13480 ;
  assign n15523 = ~n15521 & ~n15522 ;
  assign n15524 = n15520 & n15523 ;
  assign n15525 = \wishbone_bd_ram_mem3_reg[27][24]/P0001  & n13251 ;
  assign n15526 = \wishbone_bd_ram_mem3_reg[159][24]/P0001  & n13627 ;
  assign n15527 = ~n15525 & ~n15526 ;
  assign n15528 = \wishbone_bd_ram_mem3_reg[32][24]/P0001  & n13736 ;
  assign n15529 = \wishbone_bd_ram_mem3_reg[14][24]/P0001  & n13972 ;
  assign n15530 = ~n15528 & ~n15529 ;
  assign n15531 = n15527 & n15530 ;
  assign n15532 = n15524 & n15531 ;
  assign n15533 = n15517 & n15532 ;
  assign n15534 = \wishbone_bd_ram_mem3_reg[128][24]/P0001  & n13652 ;
  assign n15535 = \wishbone_bd_ram_mem3_reg[113][24]/P0001  & n13882 ;
  assign n15536 = ~n15534 & ~n15535 ;
  assign n15537 = \wishbone_bd_ram_mem3_reg[123][24]/P0001  & n13749 ;
  assign n15538 = \wishbone_bd_ram_mem3_reg[206][24]/P0001  & n13414 ;
  assign n15539 = ~n15537 & ~n15538 ;
  assign n15540 = n15536 & n15539 ;
  assign n15541 = \wishbone_bd_ram_mem3_reg[174][24]/P0001  & n13899 ;
  assign n15542 = \wishbone_bd_ram_mem3_reg[242][24]/P0001  & n13383 ;
  assign n15543 = ~n15541 & ~n15542 ;
  assign n15544 = \wishbone_bd_ram_mem3_reg[194][24]/P0001  & n13624 ;
  assign n15545 = \wishbone_bd_ram_mem3_reg[223][24]/P0001  & n13335 ;
  assign n15546 = ~n15544 & ~n15545 ;
  assign n15547 = n15543 & n15546 ;
  assign n15548 = n15540 & n15547 ;
  assign n15549 = \wishbone_bd_ram_mem3_reg[221][24]/P0001  & n13641 ;
  assign n15550 = \wishbone_bd_ram_mem3_reg[85][24]/P0001  & n13784 ;
  assign n15551 = ~n15549 & ~n15550 ;
  assign n15552 = \wishbone_bd_ram_mem3_reg[63][24]/P0001  & n13327 ;
  assign n15553 = \wishbone_bd_ram_mem3_reg[71][24]/P0001  & n13636 ;
  assign n15554 = ~n15552 & ~n15553 ;
  assign n15555 = n15551 & n15554 ;
  assign n15556 = \wishbone_bd_ram_mem3_reg[74][24]/P0001  & n13564 ;
  assign n15557 = \wishbone_bd_ram_mem3_reg[56][24]/P0001  & n13611 ;
  assign n15558 = ~n15556 & ~n15557 ;
  assign n15559 = \wishbone_bd_ram_mem3_reg[95][24]/P0001  & n13317 ;
  assign n15560 = \wishbone_bd_ram_mem3_reg[49][24]/P0001  & n13929 ;
  assign n15561 = ~n15559 & ~n15560 ;
  assign n15562 = n15558 & n15561 ;
  assign n15563 = n15555 & n15562 ;
  assign n15564 = n15548 & n15563 ;
  assign n15565 = n15533 & n15564 ;
  assign n15566 = n15502 & n15565 ;
  assign n15567 = \wishbone_bd_ram_mem3_reg[37][24]/P0001  & n13710 ;
  assign n15568 = \wishbone_bd_ram_mem3_reg[222][24]/P0001  & n13721 ;
  assign n15569 = ~n15567 & ~n15568 ;
  assign n15570 = \wishbone_bd_ram_mem3_reg[92][24]/P0001  & n13859 ;
  assign n15571 = \wishbone_bd_ram_mem3_reg[208][24]/P0001  & n14010 ;
  assign n15572 = ~n15570 & ~n15571 ;
  assign n15573 = n15569 & n15572 ;
  assign n15574 = \wishbone_bd_ram_mem3_reg[231][24]/P0001  & n13363 ;
  assign n15575 = \wishbone_bd_ram_mem3_reg[48][24]/P0001  & n13917 ;
  assign n15576 = ~n15574 & ~n15575 ;
  assign n15577 = \wishbone_bd_ram_mem3_reg[12][24]/P0001  & n13733 ;
  assign n15578 = \wishbone_bd_ram_mem3_reg[240][24]/P0001  & n13352 ;
  assign n15579 = ~n15577 & ~n15578 ;
  assign n15580 = n15576 & n15579 ;
  assign n15581 = n15573 & n15580 ;
  assign n15582 = \wishbone_bd_ram_mem3_reg[138][24]/P0001  & n13398 ;
  assign n15583 = \wishbone_bd_ram_mem3_reg[246][24]/P0001  & n13981 ;
  assign n15584 = ~n15582 & ~n15583 ;
  assign n15585 = \wishbone_bd_ram_mem3_reg[210][24]/P0001  & n13443 ;
  assign n15586 = \wishbone_bd_ram_mem3_reg[107][24]/P0001  & n13476 ;
  assign n15587 = ~n15585 & ~n15586 ;
  assign n15588 = n15584 & n15587 ;
  assign n15589 = \wishbone_bd_ram_mem3_reg[51][24]/P0001  & n13880 ;
  assign n15590 = \wishbone_bd_ram_mem3_reg[5][24]/P0001  & n13243 ;
  assign n15591 = ~n15589 & ~n15590 ;
  assign n15592 = \wishbone_bd_ram_mem3_reg[155][24]/P0001  & n13738 ;
  assign n15593 = \wishbone_bd_ram_mem3_reg[72][24]/P0001  & n13582 ;
  assign n15594 = ~n15592 & ~n15593 ;
  assign n15595 = n15591 & n15594 ;
  assign n15596 = n15588 & n15595 ;
  assign n15597 = n15581 & n15596 ;
  assign n15598 = \wishbone_bd_ram_mem3_reg[98][24]/P0001  & n13569 ;
  assign n15599 = \wishbone_bd_ram_mem3_reg[45][24]/P0001  & n13420 ;
  assign n15600 = ~n15598 & ~n15599 ;
  assign n15601 = \wishbone_bd_ram_mem3_reg[86][24]/P0001  & n13485 ;
  assign n15602 = \wishbone_bd_ram_mem3_reg[64][24]/P0001  & n13904 ;
  assign n15603 = ~n15601 & ~n15602 ;
  assign n15604 = n15600 & n15603 ;
  assign n15605 = \wishbone_bd_ram_mem3_reg[108][24]/P0001  & n13814 ;
  assign n15606 = \wishbone_bd_ram_mem3_reg[19][24]/P0001  & n13886 ;
  assign n15607 = ~n15605 & ~n15606 ;
  assign n15608 = \wishbone_bd_ram_mem3_reg[15][24]/P0001  & n13797 ;
  assign n15609 = \wishbone_bd_ram_mem3_reg[23][24]/P0001  & n13857 ;
  assign n15610 = ~n15608 & ~n15609 ;
  assign n15611 = n15607 & n15610 ;
  assign n15612 = n15604 & n15611 ;
  assign n15613 = \wishbone_bd_ram_mem3_reg[179][24]/P0001  & n14035 ;
  assign n15614 = \wishbone_bd_ram_mem3_reg[167][24]/P0001  & n13940 ;
  assign n15615 = ~n15613 & ~n15614 ;
  assign n15616 = \wishbone_bd_ram_mem3_reg[202][24]/P0001  & n13268 ;
  assign n15617 = \wishbone_bd_ram_mem3_reg[119][24]/P0001  & n14033 ;
  assign n15618 = ~n15616 & ~n15617 ;
  assign n15619 = n15615 & n15618 ;
  assign n15620 = \wishbone_bd_ram_mem3_reg[183][24]/P0001  & n13645 ;
  assign n15621 = \wishbone_bd_ram_mem3_reg[161][24]/P0001  & n13505 ;
  assign n15622 = ~n15620 & ~n15621 ;
  assign n15623 = \wishbone_bd_ram_mem3_reg[190][24]/P0001  & n13365 ;
  assign n15624 = \wishbone_bd_ram_mem3_reg[54][24]/P0001  & n13622 ;
  assign n15625 = ~n15623 & ~n15624 ;
  assign n15626 = n15622 & n15625 ;
  assign n15627 = n15619 & n15626 ;
  assign n15628 = n15612 & n15627 ;
  assign n15629 = n15597 & n15628 ;
  assign n15630 = \wishbone_bd_ram_mem3_reg[235][24]/P0001  & n13518 ;
  assign n15631 = \wishbone_bd_ram_mem3_reg[42][24]/P0001  & n13341 ;
  assign n15632 = ~n15630 & ~n15631 ;
  assign n15633 = \wishbone_bd_ram_mem3_reg[200][24]/P0001  & n13922 ;
  assign n15634 = \wishbone_bd_ram_mem3_reg[112][24]/P0001  & n13482 ;
  assign n15635 = ~n15633 & ~n15634 ;
  assign n15636 = n15632 & n15635 ;
  assign n15637 = \wishbone_bd_ram_mem3_reg[148][24]/P0001  & n13868 ;
  assign n15638 = \wishbone_bd_ram_mem3_reg[134][24]/P0001  & n13494 ;
  assign n15639 = ~n15637 & ~n15638 ;
  assign n15640 = \wishbone_bd_ram_mem3_reg[163][24]/P0001  & n13255 ;
  assign n15641 = \wishbone_bd_ram_mem3_reg[186][24]/P0001  & n13616 ;
  assign n15642 = ~n15640 & ~n15641 ;
  assign n15643 = n15639 & n15642 ;
  assign n15644 = n15636 & n15643 ;
  assign n15645 = \wishbone_bd_ram_mem3_reg[69][24]/P0001  & n13487 ;
  assign n15646 = \wishbone_bd_ram_mem3_reg[225][24]/P0001  & n13719 ;
  assign n15647 = ~n15645 & ~n15646 ;
  assign n15648 = \wishbone_bd_ram_mem3_reg[1][24]/P0001  & n13888 ;
  assign n15649 = \wishbone_bd_ram_mem3_reg[70][24]/P0001  & n13339 ;
  assign n15650 = ~n15648 & ~n15649 ;
  assign n15651 = n15647 & n15650 ;
  assign n15652 = \wishbone_bd_ram_mem3_reg[251][24]/P0001  & n14019 ;
  assign n15653 = \wishbone_bd_ram_mem3_reg[151][24]/P0001  & n13697 ;
  assign n15654 = ~n15652 & ~n15653 ;
  assign n15655 = \wishbone_bd_ram_mem3_reg[254][24]/P0001  & n13283 ;
  assign n15656 = \wishbone_bd_ram_mem3_reg[103][24]/P0001  & n13320 ;
  assign n15657 = ~n15655 & ~n15656 ;
  assign n15658 = n15654 & n15657 ;
  assign n15659 = n15651 & n15658 ;
  assign n15660 = n15644 & n15659 ;
  assign n15661 = \wishbone_bd_ram_mem3_reg[79][24]/P0001  & n13779 ;
  assign n15662 = \wishbone_bd_ram_mem3_reg[101][24]/P0001  & n13772 ;
  assign n15663 = ~n15661 & ~n15662 ;
  assign n15664 = \wishbone_bd_ram_mem3_reg[199][24]/P0001  & n13499 ;
  assign n15665 = \wishbone_bd_ram_mem3_reg[58][24]/P0001  & n13949 ;
  assign n15666 = ~n15664 & ~n15665 ;
  assign n15667 = n15663 & n15666 ;
  assign n15668 = \wishbone_bd_ram_mem3_reg[136][24]/P0001  & n13963 ;
  assign n15669 = \wishbone_bd_ram_mem3_reg[135][24]/P0001  & n13672 ;
  assign n15670 = ~n15668 & ~n15669 ;
  assign n15671 = \wishbone_bd_ram_mem3_reg[87][24]/P0001  & n13691 ;
  assign n15672 = \wishbone_bd_ram_mem3_reg[156][24]/P0001  & n13769 ;
  assign n15673 = ~n15671 & ~n15672 ;
  assign n15674 = n15670 & n15673 ;
  assign n15675 = n15667 & n15674 ;
  assign n15676 = \wishbone_bd_ram_mem3_reg[207][24]/P0001  & n13826 ;
  assign n15677 = \wishbone_bd_ram_mem3_reg[248][24]/P0001  & n13647 ;
  assign n15678 = ~n15676 & ~n15677 ;
  assign n15679 = \wishbone_bd_ram_mem3_reg[94][24]/P0001  & n13833 ;
  assign n15680 = \wishbone_bd_ram_mem3_reg[7][24]/P0001  & n13546 ;
  assign n15681 = ~n15679 & ~n15680 ;
  assign n15682 = n15678 & n15681 ;
  assign n15683 = \wishbone_bd_ram_mem3_reg[198][24]/P0001  & n13592 ;
  assign n15684 = \wishbone_bd_ram_mem3_reg[46][24]/P0001  & n13298 ;
  assign n15685 = ~n15683 & ~n15684 ;
  assign n15686 = \wishbone_bd_ram_mem3_reg[96][24]/P0001  & n13425 ;
  assign n15687 = \wishbone_bd_ram_mem3_reg[203][24]/P0001  & n13816 ;
  assign n15688 = ~n15686 & ~n15687 ;
  assign n15689 = n15685 & n15688 ;
  assign n15690 = n15682 & n15689 ;
  assign n15691 = n15675 & n15690 ;
  assign n15692 = n15660 & n15691 ;
  assign n15693 = n15629 & n15692 ;
  assign n15694 = n15566 & n15693 ;
  assign n15695 = n15439 & n15694 ;
  assign n15696 = n14047 & ~n15695 ;
  assign n15697 = ~\wishbone_TxLength_reg[7]/NET0131  & n14056 ;
  assign n15698 = n14055 & n15697 ;
  assign n15699 = n14049 & n15698 ;
  assign n15700 = ~n14072 & n15699 ;
  assign n15701 = ~n14064 & n15700 ;
  assign n15702 = ~\wishbone_TxLength_reg[8]/NET0131  & ~n15701 ;
  assign n15703 = ~n14072 & n15698 ;
  assign n15704 = ~n14064 & ~n15703 ;
  assign n15705 = \wishbone_TxLength_reg[8]/NET0131  & n14049 ;
  assign n15706 = ~n15704 & n15705 ;
  assign n15707 = ~n14046 & ~n15706 ;
  assign n15708 = ~n15702 & n15707 ;
  assign n15709 = ~n15696 & ~n15708 ;
  assign n15710 = n13112 & n13114 ;
  assign n15711 = n13111 & n15710 ;
  assign n15712 = \m_wb_adr_o[25]_pad  & n15711 ;
  assign n15713 = ~\m_wb_adr_o[26]_pad  & ~n15712 ;
  assign n15714 = \wishbone_TxPointerMSB_reg[26]/NET0131  & ~n13166 ;
  assign n15715 = ~n13164 & n15714 ;
  assign n15716 = n15177 & ~n15715 ;
  assign n15717 = ~n13118 & ~n15716 ;
  assign n15718 = ~n15713 & n15717 ;
  assign n15719 = \m_wb_adr_o[26]_pad  & n13197 ;
  assign n15720 = \wishbone_TxPointerMSB_reg[26]/NET0131  & ~n13201 ;
  assign n15721 = \wishbone_RxPointerMSB_reg[26]/NET0131  & n13207 ;
  assign n15722 = ~n13196 & n15721 ;
  assign n15723 = ~n15720 & ~n15722 ;
  assign n15724 = ~n15719 & n15723 ;
  assign n15725 = ~n15718 & n15724 ;
  assign n15726 = \rxethmac1_RxStartFrm_reg/NET0131  & \rxethmac1_RxValid_reg/NET0131  ;
  assign n15727 = \wishbone_RxPointerLSB_rst_reg[0]/NET0131  & \wishbone_RxReady_reg/NET0131  ;
  assign n15728 = n15726 & n15727 ;
  assign n15729 = \wishbone_RxPointerLSB_rst_reg[1]/NET0131  & n15728 ;
  assign n15730 = ~\rxethmac1_RxStartFrm_reg/NET0131  & \rxethmac1_RxValid_reg/NET0131  ;
  assign n15731 = \wishbone_RxEnableWindow_reg/NET0131  & n15730 ;
  assign n15732 = \wishbone_RxByteCnt_reg[0]/NET0131  & \wishbone_RxByteCnt_reg[1]/NET0131  ;
  assign n15733 = \wishbone_RxReady_reg/NET0131  & n15732 ;
  assign n15734 = n15731 & n15733 ;
  assign n15735 = ~n15729 & ~n15734 ;
  assign n15736 = \wishbone_LastByteIn_reg/NET0131  & \wishbone_ShiftWillEnd_reg/NET0131  ;
  assign n15737 = n15732 & n15736 ;
  assign n15738 = \wishbone_RxDataLatched2_reg[10]/NET0131  & ~n15737 ;
  assign n15739 = n15735 & n15738 ;
  assign n15740 = ~\wishbone_ShiftWillEnd_reg/NET0131  & ~n15735 ;
  assign n15741 = ~\wishbone_RxValidBytes_reg[0]/NET0131  & ~\wishbone_RxValidBytes_reg[1]/NET0131  ;
  assign n15742 = \wishbone_RxValidBytes_reg[0]/NET0131  & \wishbone_RxValidBytes_reg[1]/NET0131  ;
  assign n15743 = ~n15741 & ~n15742 ;
  assign n15744 = ~n15740 & n15743 ;
  assign n15745 = n15735 & ~n15737 ;
  assign n15746 = \wishbone_RxDataLatched1_reg[10]/NET0131  & ~n15745 ;
  assign n15747 = ~n15744 & n15746 ;
  assign n15748 = ~n15739 & ~n15747 ;
  assign n15749 = \wishbone_RxDataLatched2_reg[11]/NET0131  & ~n15737 ;
  assign n15750 = n15735 & n15749 ;
  assign n15751 = \wishbone_RxDataLatched1_reg[11]/NET0131  & ~n15745 ;
  assign n15752 = ~n15744 & n15751 ;
  assign n15753 = ~n15750 & ~n15752 ;
  assign n15754 = \wishbone_RxDataLatched2_reg[12]/NET0131  & ~n15737 ;
  assign n15755 = n15735 & n15754 ;
  assign n15756 = \wishbone_RxDataLatched1_reg[12]/NET0131  & ~n15745 ;
  assign n15757 = ~n15744 & n15756 ;
  assign n15758 = ~n15755 & ~n15757 ;
  assign n15759 = \wishbone_RxDataLatched2_reg[13]/NET0131  & ~n15737 ;
  assign n15760 = n15735 & n15759 ;
  assign n15761 = \wishbone_RxDataLatched1_reg[13]/NET0131  & ~n15745 ;
  assign n15762 = ~n15744 & n15761 ;
  assign n15763 = ~n15760 & ~n15762 ;
  assign n15764 = \wishbone_RxDataLatched2_reg[14]/NET0131  & ~n15737 ;
  assign n15765 = n15735 & n15764 ;
  assign n15766 = \wishbone_RxDataLatched1_reg[14]/NET0131  & ~n15745 ;
  assign n15767 = ~n15744 & n15766 ;
  assign n15768 = ~n15765 & ~n15767 ;
  assign n15769 = \wishbone_RxDataLatched2_reg[15]/NET0131  & ~n15737 ;
  assign n15770 = n15735 & n15769 ;
  assign n15771 = \wishbone_RxDataLatched1_reg[15]/NET0131  & ~n15745 ;
  assign n15772 = ~n15744 & n15771 ;
  assign n15773 = ~n15770 & ~n15772 ;
  assign n15774 = \wishbone_RxDataLatched2_reg[8]/NET0131  & ~n15737 ;
  assign n15775 = n15735 & n15774 ;
  assign n15776 = \wishbone_RxDataLatched1_reg[8]/NET0131  & ~n15745 ;
  assign n15777 = ~n15744 & n15776 ;
  assign n15778 = ~n15775 & ~n15777 ;
  assign n15779 = \wishbone_RxEn_q_reg/NET0131  & \wishbone_RxEn_reg/NET0131  ;
  assign n15780 = \wishbone_RxBDRead_reg/NET0131  & n15779 ;
  assign n15781 = \wishbone_RxBDReady_reg/NET0131  & ~\wishbone_RxPointerRead_reg/NET0131  ;
  assign n15782 = \wishbone_RxBDRead_reg/NET0131  & ~\wishbone_RxPointerRead_reg/NET0131  ;
  assign n15783 = n15779 & n15782 ;
  assign n15784 = ~n15781 & ~n15783 ;
  assign n15785 = ~n15780 & ~n15784 ;
  assign n15786 = \wishbone_bd_ram_mem1_reg[44][15]/P0001  & n13291 ;
  assign n15787 = \wishbone_bd_ram_mem1_reg[243][15]/P0001  & n13575 ;
  assign n15788 = ~n15786 & ~n15787 ;
  assign n15789 = \wishbone_bd_ram_mem1_reg[118][15]/P0001  & n13589 ;
  assign n15790 = \wishbone_bd_ram_mem1_reg[193][15]/P0001  & n14022 ;
  assign n15791 = ~n15789 & ~n15790 ;
  assign n15792 = n15788 & n15791 ;
  assign n15793 = \wishbone_bd_ram_mem1_reg[234][15]/P0001  & n13781 ;
  assign n15794 = \wishbone_bd_ram_mem1_reg[162][15]/P0001  & n13726 ;
  assign n15795 = ~n15793 & ~n15794 ;
  assign n15796 = \wishbone_bd_ram_mem1_reg[145][15]/P0001  & n13715 ;
  assign n15797 = \wishbone_bd_ram_mem1_reg[72][15]/P0001  & n13582 ;
  assign n15798 = ~n15796 & ~n15797 ;
  assign n15799 = n15795 & n15798 ;
  assign n15800 = n15792 & n15799 ;
  assign n15801 = \wishbone_bd_ram_mem1_reg[105][15]/P0001  & n13503 ;
  assign n15802 = \wishbone_bd_ram_mem1_reg[141][15]/P0001  & n13852 ;
  assign n15803 = ~n15801 & ~n15802 ;
  assign n15804 = \wishbone_bd_ram_mem1_reg[149][15]/P0001  & n13469 ;
  assign n15805 = \wishbone_bd_ram_mem1_reg[194][15]/P0001  & n13624 ;
  assign n15806 = ~n15804 & ~n15805 ;
  assign n15807 = n15803 & n15806 ;
  assign n15808 = \wishbone_bd_ram_mem1_reg[132][15]/P0001  & n13927 ;
  assign n15809 = \wishbone_bd_ram_mem1_reg[83][15]/P0001  & n13454 ;
  assign n15810 = ~n15808 & ~n15809 ;
  assign n15811 = \wishbone_bd_ram_mem1_reg[167][15]/P0001  & n13940 ;
  assign n15812 = \wishbone_bd_ram_mem1_reg[151][15]/P0001  & n13697 ;
  assign n15813 = ~n15811 & ~n15812 ;
  assign n15814 = n15810 & n15813 ;
  assign n15815 = n15807 & n15814 ;
  assign n15816 = n15800 & n15815 ;
  assign n15817 = \wishbone_bd_ram_mem1_reg[47][15]/P0001  & n13436 ;
  assign n15818 = \wishbone_bd_ram_mem1_reg[21][15]/P0001  & n13438 ;
  assign n15819 = ~n15817 & ~n15818 ;
  assign n15820 = \wishbone_bd_ram_mem1_reg[77][15]/P0001  & n13935 ;
  assign n15821 = \wishbone_bd_ram_mem1_reg[206][15]/P0001  & n13414 ;
  assign n15822 = ~n15820 & ~n15821 ;
  assign n15823 = n15819 & n15822 ;
  assign n15824 = \wishbone_bd_ram_mem1_reg[15][15]/P0001  & n13797 ;
  assign n15825 = \wishbone_bd_ram_mem1_reg[26][15]/P0001  & n13521 ;
  assign n15826 = ~n15824 & ~n15825 ;
  assign n15827 = \wishbone_bd_ram_mem1_reg[97][15]/P0001  & n13724 ;
  assign n15828 = \wishbone_bd_ram_mem1_reg[160][15]/P0001  & n13271 ;
  assign n15829 = ~n15827 & ~n15828 ;
  assign n15830 = n15826 & n15829 ;
  assign n15831 = n15823 & n15830 ;
  assign n15832 = \wishbone_bd_ram_mem1_reg[4][15]/P0001  & n13527 ;
  assign n15833 = \wishbone_bd_ram_mem1_reg[117][15]/P0001  & n13557 ;
  assign n15834 = ~n15832 & ~n15833 ;
  assign n15835 = \wishbone_bd_ram_mem1_reg[152][15]/P0001  & n13912 ;
  assign n15836 = \wishbone_bd_ram_mem1_reg[103][15]/P0001  & n13320 ;
  assign n15837 = ~n15835 & ~n15836 ;
  assign n15838 = n15834 & n15837 ;
  assign n15839 = \wishbone_bd_ram_mem1_reg[153][15]/P0001  & n13309 ;
  assign n15840 = \wishbone_bd_ram_mem1_reg[98][15]/P0001  & n13569 ;
  assign n15841 = ~n15839 & ~n15840 ;
  assign n15842 = \wishbone_bd_ram_mem1_reg[192][15]/P0001  & n13390 ;
  assign n15843 = \wishbone_bd_ram_mem1_reg[142][15]/P0001  & n13448 ;
  assign n15844 = ~n15842 & ~n15843 ;
  assign n15845 = n15841 & n15844 ;
  assign n15846 = n15838 & n15845 ;
  assign n15847 = n15831 & n15846 ;
  assign n15848 = n15816 & n15847 ;
  assign n15849 = \wishbone_bd_ram_mem1_reg[50][15]/P0001  & n13686 ;
  assign n15850 = \wishbone_bd_ram_mem1_reg[213][15]/P0001  & n13870 ;
  assign n15851 = ~n15849 & ~n15850 ;
  assign n15852 = \wishbone_bd_ram_mem1_reg[32][15]/P0001  & n13736 ;
  assign n15853 = \wishbone_bd_ram_mem1_reg[182][15]/P0001  & n13598 ;
  assign n15854 = ~n15852 & ~n15853 ;
  assign n15855 = n15851 & n15854 ;
  assign n15856 = \wishbone_bd_ram_mem1_reg[29][15]/P0001  & n13412 ;
  assign n15857 = \wishbone_bd_ram_mem1_reg[39][15]/P0001  & n13893 ;
  assign n15858 = ~n15856 & ~n15857 ;
  assign n15859 = \wishbone_bd_ram_mem1_reg[134][15]/P0001  & n13494 ;
  assign n15860 = \wishbone_bd_ram_mem1_reg[43][15]/P0001  & n13761 ;
  assign n15861 = ~n15859 & ~n15860 ;
  assign n15862 = n15858 & n15861 ;
  assign n15863 = n15855 & n15862 ;
  assign n15864 = \wishbone_bd_ram_mem1_reg[13][15]/P0001  & n13844 ;
  assign n15865 = \wishbone_bd_ram_mem1_reg[46][15]/P0001  & n13298 ;
  assign n15866 = ~n15864 & ~n15865 ;
  assign n15867 = \wishbone_bd_ram_mem1_reg[101][15]/P0001  & n13772 ;
  assign n15868 = \wishbone_bd_ram_mem1_reg[202][15]/P0001  & n13268 ;
  assign n15869 = ~n15867 & ~n15868 ;
  assign n15870 = n15866 & n15869 ;
  assign n15871 = \wishbone_bd_ram_mem1_reg[163][15]/P0001  & n13255 ;
  assign n15872 = \wishbone_bd_ram_mem1_reg[75][15]/P0001  & n13605 ;
  assign n15873 = ~n15871 & ~n15872 ;
  assign n15874 = \wishbone_bd_ram_mem1_reg[9][15]/P0001  & n13580 ;
  assign n15875 = \wishbone_bd_ram_mem1_reg[14][15]/P0001  & n13972 ;
  assign n15876 = ~n15874 & ~n15875 ;
  assign n15877 = n15873 & n15876 ;
  assign n15878 = n15870 & n15877 ;
  assign n15879 = n15863 & n15878 ;
  assign n15880 = \wishbone_bd_ram_mem1_reg[218][15]/P0001  & n13792 ;
  assign n15881 = \wishbone_bd_ram_mem1_reg[90][15]/P0001  & n13906 ;
  assign n15882 = ~n15880 & ~n15881 ;
  assign n15883 = \wishbone_bd_ram_mem1_reg[126][15]/P0001  & n13786 ;
  assign n15884 = \wishbone_bd_ram_mem1_reg[119][15]/P0001  & n14033 ;
  assign n15885 = ~n15883 & ~n15884 ;
  assign n15886 = n15882 & n15885 ;
  assign n15887 = \wishbone_bd_ram_mem1_reg[109][15]/P0001  & n13306 ;
  assign n15888 = \wishbone_bd_ram_mem1_reg[42][15]/P0001  & n13341 ;
  assign n15889 = ~n15887 & ~n15888 ;
  assign n15890 = \wishbone_bd_ram_mem1_reg[144][15]/P0001  & n13508 ;
  assign n15891 = \wishbone_bd_ram_mem1_reg[166][15]/P0001  & n13999 ;
  assign n15892 = ~n15890 & ~n15891 ;
  assign n15893 = n15889 & n15892 ;
  assign n15894 = n15886 & n15893 ;
  assign n15895 = \wishbone_bd_ram_mem1_reg[123][15]/P0001  & n13749 ;
  assign n15896 = \wishbone_bd_ram_mem1_reg[247][15]/P0001  & n13571 ;
  assign n15897 = ~n15895 & ~n15896 ;
  assign n15898 = \wishbone_bd_ram_mem1_reg[133][15]/P0001  & n13492 ;
  assign n15899 = \wishbone_bd_ram_mem1_reg[49][15]/P0001  & n13929 ;
  assign n15900 = ~n15898 & ~n15899 ;
  assign n15901 = n15897 & n15900 ;
  assign n15902 = \wishbone_bd_ram_mem1_reg[240][15]/P0001  & n13352 ;
  assign n15903 = \wishbone_bd_ram_mem1_reg[76][15]/P0001  & n13831 ;
  assign n15904 = ~n15902 & ~n15903 ;
  assign n15905 = \wishbone_bd_ram_mem1_reg[84][15]/P0001  & n13385 ;
  assign n15906 = \wishbone_bd_ram_mem1_reg[177][15]/P0001  & n13863 ;
  assign n15907 = ~n15905 & ~n15906 ;
  assign n15908 = n15904 & n15907 ;
  assign n15909 = n15901 & n15908 ;
  assign n15910 = n15894 & n15909 ;
  assign n15911 = n15879 & n15910 ;
  assign n15912 = n15848 & n15911 ;
  assign n15913 = \wishbone_bd_ram_mem1_reg[203][15]/P0001  & n13816 ;
  assign n15914 = \wishbone_bd_ram_mem1_reg[147][15]/P0001  & n13702 ;
  assign n15915 = ~n15913 & ~n15914 ;
  assign n15916 = \wishbone_bd_ram_mem1_reg[1][15]/P0001  & n13888 ;
  assign n15917 = \wishbone_bd_ram_mem1_reg[179][15]/P0001  & n14035 ;
  assign n15918 = ~n15916 & ~n15917 ;
  assign n15919 = n15915 & n15918 ;
  assign n15920 = \wishbone_bd_ram_mem1_reg[80][15]/P0001  & n13516 ;
  assign n15921 = \wishbone_bd_ram_mem1_reg[237][15]/P0001  & n13924 ;
  assign n15922 = ~n15920 & ~n15921 ;
  assign n15923 = \wishbone_bd_ram_mem1_reg[235][15]/P0001  & n13518 ;
  assign n15924 = \wishbone_bd_ram_mem1_reg[86][15]/P0001  & n13485 ;
  assign n15925 = ~n15923 & ~n15924 ;
  assign n15926 = n15922 & n15925 ;
  assign n15927 = n15919 & n15926 ;
  assign n15928 = \wishbone_bd_ram_mem1_reg[138][15]/P0001  & n13398 ;
  assign n15929 = \wishbone_bd_ram_mem1_reg[252][15]/P0001  & n13986 ;
  assign n15930 = ~n15928 & ~n15929 ;
  assign n15931 = \wishbone_bd_ram_mem1_reg[22][15]/P0001  & n13744 ;
  assign n15932 = \wishbone_bd_ram_mem1_reg[62][15]/P0001  & n13529 ;
  assign n15933 = ~n15931 & ~n15932 ;
  assign n15934 = n15930 & n15933 ;
  assign n15935 = \wishbone_bd_ram_mem1_reg[45][15]/P0001  & n13420 ;
  assign n15936 = \wishbone_bd_ram_mem1_reg[180][15]/P0001  & n13650 ;
  assign n15937 = ~n15935 & ~n15936 ;
  assign n15938 = \wishbone_bd_ram_mem1_reg[68][15]/P0001  & n13379 ;
  assign n15939 = \wishbone_bd_ram_mem1_reg[233][15]/P0001  & n13332 ;
  assign n15940 = ~n15938 & ~n15939 ;
  assign n15941 = n15937 & n15940 ;
  assign n15942 = n15934 & n15941 ;
  assign n15943 = n15927 & n15942 ;
  assign n15944 = \wishbone_bd_ram_mem1_reg[212][15]/P0001  & n13634 ;
  assign n15945 = \wishbone_bd_ram_mem1_reg[85][15]/P0001  & n13784 ;
  assign n15946 = ~n15944 & ~n15945 ;
  assign n15947 = \wishbone_bd_ram_mem1_reg[120][15]/P0001  & n13550 ;
  assign n15948 = \wishbone_bd_ram_mem1_reg[169][15]/P0001  & n13541 ;
  assign n15949 = ~n15947 & ~n15948 ;
  assign n15950 = n15946 & n15949 ;
  assign n15951 = \wishbone_bd_ram_mem1_reg[156][15]/P0001  & n13769 ;
  assign n15952 = \wishbone_bd_ram_mem1_reg[242][15]/P0001  & n13383 ;
  assign n15953 = ~n15951 & ~n15952 ;
  assign n15954 = \wishbone_bd_ram_mem1_reg[199][15]/P0001  & n13499 ;
  assign n15955 = \wishbone_bd_ram_mem1_reg[173][15]/P0001  & n13360 ;
  assign n15956 = ~n15954 & ~n15955 ;
  assign n15957 = n15953 & n15956 ;
  assign n15958 = n15950 & n15957 ;
  assign n15959 = \wishbone_bd_ram_mem1_reg[197][15]/P0001  & n13594 ;
  assign n15960 = \wishbone_bd_ram_mem1_reg[155][15]/P0001  & n13738 ;
  assign n15961 = ~n15959 & ~n15960 ;
  assign n15962 = \wishbone_bd_ram_mem1_reg[164][15]/P0001  & n13236 ;
  assign n15963 = \wishbone_bd_ram_mem1_reg[226][15]/P0001  & n13668 ;
  assign n15964 = ~n15962 & ~n15963 ;
  assign n15965 = n15961 & n15964 ;
  assign n15966 = \wishbone_bd_ram_mem1_reg[191][15]/P0001  & n14012 ;
  assign n15967 = \wishbone_bd_ram_mem1_reg[217][15]/P0001  & n13767 ;
  assign n15968 = ~n15966 & ~n15967 ;
  assign n15969 = \wishbone_bd_ram_mem1_reg[108][15]/P0001  & n13814 ;
  assign n15970 = \wishbone_bd_ram_mem1_reg[139][15]/P0001  & n13566 ;
  assign n15971 = ~n15969 & ~n15970 ;
  assign n15972 = n15968 & n15971 ;
  assign n15973 = n15965 & n15972 ;
  assign n15974 = n15958 & n15973 ;
  assign n15975 = n15943 & n15974 ;
  assign n15976 = \wishbone_bd_ram_mem1_reg[73][15]/P0001  & n13456 ;
  assign n15977 = \wishbone_bd_ram_mem1_reg[201][15]/P0001  & n13600 ;
  assign n15978 = ~n15976 & ~n15977 ;
  assign n15979 = \wishbone_bd_ram_mem1_reg[37][15]/P0001  & n13710 ;
  assign n15980 = \wishbone_bd_ram_mem1_reg[104][15]/P0001  & n13684 ;
  assign n15981 = ~n15979 & ~n15980 ;
  assign n15982 = n15978 & n15981 ;
  assign n15983 = \wishbone_bd_ram_mem1_reg[52][15]/P0001  & n13988 ;
  assign n15984 = \wishbone_bd_ram_mem1_reg[112][15]/P0001  & n13482 ;
  assign n15985 = ~n15983 & ~n15984 ;
  assign n15986 = \wishbone_bd_ram_mem1_reg[255][15]/P0001  & n13952 ;
  assign n15987 = \wishbone_bd_ram_mem1_reg[175][15]/P0001  & n13674 ;
  assign n15988 = ~n15986 & ~n15987 ;
  assign n15989 = n15985 & n15988 ;
  assign n15990 = n15982 & n15989 ;
  assign n15991 = \wishbone_bd_ram_mem1_reg[238][15]/P0001  & n13819 ;
  assign n15992 = \wishbone_bd_ram_mem1_reg[58][15]/P0001  & n13949 ;
  assign n15993 = ~n15991 & ~n15992 ;
  assign n15994 = \wishbone_bd_ram_mem1_reg[195][15]/P0001  & n13700 ;
  assign n15995 = \wishbone_bd_ram_mem1_reg[60][15]/P0001  & n13790 ;
  assign n15996 = ~n15994 & ~n15995 ;
  assign n15997 = n15993 & n15996 ;
  assign n15998 = \wishbone_bd_ram_mem1_reg[27][15]/P0001  & n13251 ;
  assign n15999 = \wishbone_bd_ram_mem1_reg[7][15]/P0001  & n13546 ;
  assign n16000 = ~n15998 & ~n15999 ;
  assign n16001 = \wishbone_bd_ram_mem1_reg[150][15]/P0001  & n13666 ;
  assign n16002 = \wishbone_bd_ram_mem1_reg[215][15]/P0001  & n13901 ;
  assign n16003 = ~n16001 & ~n16002 ;
  assign n16004 = n16000 & n16003 ;
  assign n16005 = n15997 & n16004 ;
  assign n16006 = n15990 & n16005 ;
  assign n16007 = \wishbone_bd_ram_mem1_reg[88][15]/P0001  & n13347 ;
  assign n16008 = \wishbone_bd_ram_mem1_reg[172][15]/P0001  & n13377 ;
  assign n16009 = ~n16007 & ~n16008 ;
  assign n16010 = \wishbone_bd_ram_mem1_reg[129][15]/P0001  & n13629 ;
  assign n16011 = \wishbone_bd_ram_mem1_reg[227][15]/P0001  & n13388 ;
  assign n16012 = ~n16010 & ~n16011 ;
  assign n16013 = n16009 & n16012 ;
  assign n16014 = \wishbone_bd_ram_mem1_reg[188][15]/P0001  & n13407 ;
  assign n16015 = \wishbone_bd_ram_mem1_reg[198][15]/P0001  & n13592 ;
  assign n16016 = ~n16014 & ~n16015 ;
  assign n16017 = \wishbone_bd_ram_mem1_reg[249][15]/P0001  & n13431 ;
  assign n16018 = \wishbone_bd_ram_mem1_reg[196][15]/P0001  & n13977 ;
  assign n16019 = ~n16017 & ~n16018 ;
  assign n16020 = n16016 & n16019 ;
  assign n16021 = n16013 & n16020 ;
  assign n16022 = \wishbone_bd_ram_mem1_reg[67][15]/P0001  & n13663 ;
  assign n16023 = \wishbone_bd_ram_mem1_reg[41][15]/P0001  & n14017 ;
  assign n16024 = ~n16022 & ~n16023 ;
  assign n16025 = \wishbone_bd_ram_mem1_reg[122][15]/P0001  & n13679 ;
  assign n16026 = \wishbone_bd_ram_mem1_reg[25][15]/P0001  & n13742 ;
  assign n16027 = ~n16025 & ~n16026 ;
  assign n16028 = n16024 & n16027 ;
  assign n16029 = \wishbone_bd_ram_mem1_reg[18][15]/P0001  & n13532 ;
  assign n16030 = \wishbone_bd_ram_mem1_reg[181][15]/P0001  & n13587 ;
  assign n16031 = ~n16029 & ~n16030 ;
  assign n16032 = \wishbone_bd_ram_mem1_reg[20][15]/P0001  & n13839 ;
  assign n16033 = \wishbone_bd_ram_mem1_reg[189][15]/P0001  & n14001 ;
  assign n16034 = ~n16032 & ~n16033 ;
  assign n16035 = n16031 & n16034 ;
  assign n16036 = n16028 & n16035 ;
  assign n16037 = n16021 & n16036 ;
  assign n16038 = n16006 & n16037 ;
  assign n16039 = n15975 & n16038 ;
  assign n16040 = n15912 & n16039 ;
  assign n16041 = \wishbone_bd_ram_mem1_reg[121][15]/P0001  & n13983 ;
  assign n16042 = \wishbone_bd_ram_mem1_reg[65][15]/P0001  & n13842 ;
  assign n16043 = ~n16041 & ~n16042 ;
  assign n16044 = \wishbone_bd_ram_mem1_reg[229][15]/P0001  & n13552 ;
  assign n16045 = \wishbone_bd_ram_mem1_reg[100][15]/P0001  & n13401 ;
  assign n16046 = ~n16044 & ~n16045 ;
  assign n16047 = n16043 & n16046 ;
  assign n16048 = \wishbone_bd_ram_mem1_reg[223][15]/P0001  & n13335 ;
  assign n16049 = \wishbone_bd_ram_mem1_reg[89][15]/P0001  & n13910 ;
  assign n16050 = ~n16048 & ~n16049 ;
  assign n16051 = \wishbone_bd_ram_mem1_reg[6][15]/P0001  & n13915 ;
  assign n16052 = \wishbone_bd_ram_mem1_reg[70][15]/P0001  & n13339 ;
  assign n16053 = ~n16051 & ~n16052 ;
  assign n16054 = n16050 & n16053 ;
  assign n16055 = n16047 & n16054 ;
  assign n16056 = \wishbone_bd_ram_mem1_reg[38][15]/P0001  & n13828 ;
  assign n16057 = \wishbone_bd_ram_mem1_reg[34][15]/P0001  & n13450 ;
  assign n16058 = ~n16056 & ~n16057 ;
  assign n16059 = \wishbone_bd_ram_mem1_reg[3][15]/P0001  & n13354 ;
  assign n16060 = \wishbone_bd_ram_mem1_reg[63][15]/P0001  & n13327 ;
  assign n16061 = ~n16059 & ~n16060 ;
  assign n16062 = n16058 & n16061 ;
  assign n16063 = \wishbone_bd_ram_mem1_reg[183][15]/P0001  & n13645 ;
  assign n16064 = \wishbone_bd_ram_mem1_reg[96][15]/P0001  & n13425 ;
  assign n16065 = ~n16063 & ~n16064 ;
  assign n16066 = \wishbone_bd_ram_mem1_reg[228][15]/P0001  & n13497 ;
  assign n16067 = \wishbone_bd_ram_mem1_reg[59][15]/P0001  & n13613 ;
  assign n16068 = ~n16066 & ~n16067 ;
  assign n16069 = n16065 & n16068 ;
  assign n16070 = n16062 & n16069 ;
  assign n16071 = n16055 & n16070 ;
  assign n16072 = \wishbone_bd_ram_mem1_reg[159][15]/P0001  & n13627 ;
  assign n16073 = \wishbone_bd_ram_mem1_reg[56][15]/P0001  & n13611 ;
  assign n16074 = ~n16072 & ~n16073 ;
  assign n16075 = \wishbone_bd_ram_mem1_reg[12][15]/P0001  & n13733 ;
  assign n16076 = \wishbone_bd_ram_mem1_reg[161][15]/P0001  & n13505 ;
  assign n16077 = ~n16075 & ~n16076 ;
  assign n16078 = n16074 & n16077 ;
  assign n16079 = \wishbone_bd_ram_mem1_reg[23][15]/P0001  & n13857 ;
  assign n16080 = \wishbone_bd_ram_mem1_reg[208][15]/P0001  & n14010 ;
  assign n16081 = ~n16079 & ~n16080 ;
  assign n16082 = \wishbone_bd_ram_mem1_reg[54][15]/P0001  & n13622 ;
  assign n16083 = \wishbone_bd_ram_mem1_reg[248][15]/P0001  & n13647 ;
  assign n16084 = ~n16082 & ~n16083 ;
  assign n16085 = n16081 & n16084 ;
  assign n16086 = n16078 & n16085 ;
  assign n16087 = \wishbone_bd_ram_mem1_reg[135][15]/P0001  & n13672 ;
  assign n16088 = \wishbone_bd_ram_mem1_reg[2][15]/P0001  & n13975 ;
  assign n16089 = ~n16087 & ~n16088 ;
  assign n16090 = \wishbone_bd_ram_mem1_reg[184][15]/P0001  & n13960 ;
  assign n16091 = \wishbone_bd_ram_mem1_reg[154][15]/P0001  & n13403 ;
  assign n16092 = ~n16090 & ~n16091 ;
  assign n16093 = n16089 & n16092 ;
  assign n16094 = \wishbone_bd_ram_mem1_reg[92][15]/P0001  & n13859 ;
  assign n16095 = \wishbone_bd_ram_mem1_reg[186][15]/P0001  & n13616 ;
  assign n16096 = ~n16094 & ~n16095 ;
  assign n16097 = \wishbone_bd_ram_mem1_reg[19][15]/P0001  & n13886 ;
  assign n16098 = \wishbone_bd_ram_mem1_reg[232][15]/P0001  & n13510 ;
  assign n16099 = ~n16097 & ~n16098 ;
  assign n16100 = n16096 & n16099 ;
  assign n16101 = n16093 & n16100 ;
  assign n16102 = n16086 & n16101 ;
  assign n16103 = n16071 & n16102 ;
  assign n16104 = \wishbone_bd_ram_mem1_reg[51][15]/P0001  & n13880 ;
  assign n16105 = \wishbone_bd_ram_mem1_reg[250][15]/P0001  & n13677 ;
  assign n16106 = ~n16104 & ~n16105 ;
  assign n16107 = \wishbone_bd_ram_mem1_reg[185][15]/P0001  & n13372 ;
  assign n16108 = \wishbone_bd_ram_mem1_reg[148][15]/P0001  & n13868 ;
  assign n16109 = ~n16107 & ~n16108 ;
  assign n16110 = n16106 & n16109 ;
  assign n16111 = \wishbone_bd_ram_mem1_reg[10][15]/P0001  & n13837 ;
  assign n16112 = \wishbone_bd_ram_mem1_reg[102][15]/P0001  & n13534 ;
  assign n16113 = ~n16111 & ~n16112 ;
  assign n16114 = \wishbone_bd_ram_mem1_reg[136][15]/P0001  & n13963 ;
  assign n16115 = \wishbone_bd_ram_mem1_reg[190][15]/P0001  & n13365 ;
  assign n16116 = ~n16114 & ~n16115 ;
  assign n16117 = n16113 & n16116 ;
  assign n16118 = n16110 & n16117 ;
  assign n16119 = \wishbone_bd_ram_mem1_reg[114][15]/P0001  & n13763 ;
  assign n16120 = \wishbone_bd_ram_mem1_reg[94][15]/P0001  & n13833 ;
  assign n16121 = ~n16119 & ~n16120 ;
  assign n16122 = \wishbone_bd_ram_mem1_reg[236][15]/P0001  & n13480 ;
  assign n16123 = \wishbone_bd_ram_mem1_reg[113][15]/P0001  & n13882 ;
  assign n16124 = ~n16122 & ~n16123 ;
  assign n16125 = n16121 & n16124 ;
  assign n16126 = \wishbone_bd_ram_mem1_reg[57][15]/P0001  & n13731 ;
  assign n16127 = \wishbone_bd_ram_mem1_reg[254][15]/P0001  & n13283 ;
  assign n16128 = ~n16126 & ~n16127 ;
  assign n16129 = \wishbone_bd_ram_mem1_reg[245][15]/P0001  & n13877 ;
  assign n16130 = \wishbone_bd_ram_mem1_reg[253][15]/P0001  & n13708 ;
  assign n16131 = ~n16129 & ~n16130 ;
  assign n16132 = n16128 & n16131 ;
  assign n16133 = n16125 & n16132 ;
  assign n16134 = n16118 & n16133 ;
  assign n16135 = \wishbone_bd_ram_mem1_reg[79][15]/P0001  & n13779 ;
  assign n16136 = \wishbone_bd_ram_mem1_reg[5][15]/P0001  & n13243 ;
  assign n16137 = ~n16135 & ~n16136 ;
  assign n16138 = \wishbone_bd_ram_mem1_reg[53][15]/P0001  & n13875 ;
  assign n16139 = \wishbone_bd_ram_mem1_reg[225][15]/P0001  & n13719 ;
  assign n16140 = ~n16138 & ~n16139 ;
  assign n16141 = n16137 & n16140 ;
  assign n16142 = \wishbone_bd_ram_mem1_reg[231][15]/P0001  & n13363 ;
  assign n16143 = \wishbone_bd_ram_mem1_reg[209][15]/P0001  & n13689 ;
  assign n16144 = ~n16142 & ~n16143 ;
  assign n16145 = \wishbone_bd_ram_mem1_reg[216][15]/P0001  & n14005 ;
  assign n16146 = \wishbone_bd_ram_mem1_reg[8][15]/P0001  & n13459 ;
  assign n16147 = ~n16145 & ~n16146 ;
  assign n16148 = n16144 & n16147 ;
  assign n16149 = n16141 & n16148 ;
  assign n16150 = \wishbone_bd_ram_mem1_reg[55][15]/P0001  & n13618 ;
  assign n16151 = \wishbone_bd_ram_mem1_reg[157][15]/P0001  & n13445 ;
  assign n16152 = ~n16150 & ~n16151 ;
  assign n16153 = \wishbone_bd_ram_mem1_reg[93][15]/P0001  & n13891 ;
  assign n16154 = \wishbone_bd_ram_mem1_reg[176][15]/P0001  & n13262 ;
  assign n16155 = ~n16153 & ~n16154 ;
  assign n16156 = n16152 & n16155 ;
  assign n16157 = \wishbone_bd_ram_mem1_reg[110][15]/P0001  & n14030 ;
  assign n16158 = \wishbone_bd_ram_mem1_reg[230][15]/P0001  & n13994 ;
  assign n16159 = ~n16157 & ~n16158 ;
  assign n16160 = \wishbone_bd_ram_mem1_reg[69][15]/P0001  & n13487 ;
  assign n16161 = \wishbone_bd_ram_mem1_reg[146][15]/P0001  & n13958 ;
  assign n16162 = ~n16160 & ~n16161 ;
  assign n16163 = n16159 & n16162 ;
  assign n16164 = n16156 & n16163 ;
  assign n16165 = n16149 & n16164 ;
  assign n16166 = n16134 & n16165 ;
  assign n16167 = n16103 & n16166 ;
  assign n16168 = \wishbone_bd_ram_mem1_reg[130][15]/P0001  & n13427 ;
  assign n16169 = \wishbone_bd_ram_mem1_reg[48][15]/P0001  & n13917 ;
  assign n16170 = ~n16168 & ~n16169 ;
  assign n16171 = \wishbone_bd_ram_mem1_reg[207][15]/P0001  & n13826 ;
  assign n16172 = \wishbone_bd_ram_mem1_reg[71][15]/P0001  & n13636 ;
  assign n16173 = ~n16171 & ~n16172 ;
  assign n16174 = n16170 & n16173 ;
  assign n16175 = \wishbone_bd_ram_mem1_reg[125][15]/P0001  & n13396 ;
  assign n16176 = \wishbone_bd_ram_mem1_reg[28][15]/P0001  & n13810 ;
  assign n16177 = ~n16175 & ~n16176 ;
  assign n16178 = \wishbone_bd_ram_mem1_reg[127][15]/P0001  & n13803 ;
  assign n16179 = \wishbone_bd_ram_mem1_reg[74][15]/P0001  & n13564 ;
  assign n16180 = ~n16178 & ~n16179 ;
  assign n16181 = n16177 & n16180 ;
  assign n16182 = n16174 & n16181 ;
  assign n16183 = \wishbone_bd_ram_mem1_reg[31][15]/P0001  & n13758 ;
  assign n16184 = \wishbone_bd_ram_mem1_reg[82][15]/P0001  & n13374 ;
  assign n16185 = ~n16183 & ~n16184 ;
  assign n16186 = \wishbone_bd_ram_mem1_reg[137][15]/P0001  & n13808 ;
  assign n16187 = \wishbone_bd_ram_mem1_reg[200][15]/P0001  & n13922 ;
  assign n16188 = ~n16186 & ~n16187 ;
  assign n16189 = n16185 & n16188 ;
  assign n16190 = \wishbone_bd_ram_mem1_reg[11][15]/P0001  & n13774 ;
  assign n16191 = \wishbone_bd_ram_mem1_reg[106][15]/P0001  & n13555 ;
  assign n16192 = ~n16190 & ~n16191 ;
  assign n16193 = \wishbone_bd_ram_mem1_reg[251][15]/P0001  & n14019 ;
  assign n16194 = \wishbone_bd_ram_mem1_reg[204][15]/P0001  & n13821 ;
  assign n16195 = ~n16193 & ~n16194 ;
  assign n16196 = n16192 & n16195 ;
  assign n16197 = n16189 & n16196 ;
  assign n16198 = n16182 & n16197 ;
  assign n16199 = \wishbone_bd_ram_mem1_reg[171][15]/P0001  & n13422 ;
  assign n16200 = \wishbone_bd_ram_mem1_reg[91][15]/P0001  & n13954 ;
  assign n16201 = ~n16199 & ~n16200 ;
  assign n16202 = \wishbone_bd_ram_mem1_reg[33][15]/P0001  & n13933 ;
  assign n16203 = \wishbone_bd_ram_mem1_reg[174][15]/P0001  & n13899 ;
  assign n16204 = ~n16202 & ~n16203 ;
  assign n16205 = n16201 & n16204 ;
  assign n16206 = \wishbone_bd_ram_mem1_reg[78][15]/P0001  & n13277 ;
  assign n16207 = \wishbone_bd_ram_mem1_reg[178][15]/P0001  & n13301 ;
  assign n16208 = ~n16206 & ~n16207 ;
  assign n16209 = \wishbone_bd_ram_mem1_reg[219][15]/P0001  & n13577 ;
  assign n16210 = \wishbone_bd_ram_mem1_reg[187][15]/P0001  & n13756 ;
  assign n16211 = ~n16209 & ~n16210 ;
  assign n16212 = n16208 & n16211 ;
  assign n16213 = n16205 & n16212 ;
  assign n16214 = \wishbone_bd_ram_mem1_reg[170][15]/P0001  & n14007 ;
  assign n16215 = \wishbone_bd_ram_mem1_reg[241][15]/P0001  & n13854 ;
  assign n16216 = ~n16214 & ~n16215 ;
  assign n16217 = \wishbone_bd_ram_mem1_reg[115][15]/P0001  & n13747 ;
  assign n16218 = \wishbone_bd_ram_mem1_reg[24][15]/P0001  & n13970 ;
  assign n16219 = ~n16217 & ~n16218 ;
  assign n16220 = n16216 & n16219 ;
  assign n16221 = \wishbone_bd_ram_mem1_reg[61][15]/P0001  & n13544 ;
  assign n16222 = \wishbone_bd_ram_mem1_reg[64][15]/P0001  & n13904 ;
  assign n16223 = ~n16221 & ~n16222 ;
  assign n16224 = \wishbone_bd_ram_mem1_reg[111][15]/P0001  & n13471 ;
  assign n16225 = \wishbone_bd_ram_mem1_reg[222][15]/P0001  & n13721 ;
  assign n16226 = ~n16224 & ~n16225 ;
  assign n16227 = n16223 & n16226 ;
  assign n16228 = n16220 & n16227 ;
  assign n16229 = n16213 & n16228 ;
  assign n16230 = n16198 & n16229 ;
  assign n16231 = \wishbone_bd_ram_mem1_reg[220][15]/P0001  & n13965 ;
  assign n16232 = \wishbone_bd_ram_mem1_reg[95][15]/P0001  & n13317 ;
  assign n16233 = ~n16231 & ~n16232 ;
  assign n16234 = \wishbone_bd_ram_mem1_reg[16][15]/P0001  & n13695 ;
  assign n16235 = \wishbone_bd_ram_mem1_reg[81][15]/P0001  & n13409 ;
  assign n16236 = ~n16234 & ~n16235 ;
  assign n16237 = n16233 & n16236 ;
  assign n16238 = \wishbone_bd_ram_mem1_reg[128][15]/P0001  & n13652 ;
  assign n16239 = \wishbone_bd_ram_mem1_reg[124][15]/P0001  & n14024 ;
  assign n16240 = ~n16238 & ~n16239 ;
  assign n16241 = \wishbone_bd_ram_mem1_reg[239][15]/P0001  & n13349 ;
  assign n16242 = \wishbone_bd_ram_mem1_reg[17][15]/P0001  & n13324 ;
  assign n16243 = ~n16241 & ~n16242 ;
  assign n16244 = n16240 & n16243 ;
  assign n16245 = n16237 & n16244 ;
  assign n16246 = \wishbone_bd_ram_mem1_reg[244][15]/P0001  & n13474 ;
  assign n16247 = \wishbone_bd_ram_mem1_reg[87][15]/P0001  & n13691 ;
  assign n16248 = ~n16246 & ~n16247 ;
  assign n16249 = \wishbone_bd_ram_mem1_reg[140][15]/P0001  & n13287 ;
  assign n16250 = \wishbone_bd_ram_mem1_reg[158][15]/P0001  & n13294 ;
  assign n16251 = ~n16249 & ~n16250 ;
  assign n16252 = n16248 & n16251 ;
  assign n16253 = \wishbone_bd_ram_mem1_reg[221][15]/P0001  & n13641 ;
  assign n16254 = \wishbone_bd_ram_mem1_reg[30][15]/P0001  & n13713 ;
  assign n16255 = ~n16253 & ~n16254 ;
  assign n16256 = \wishbone_bd_ram_mem1_reg[116][15]/P0001  & n13865 ;
  assign n16257 = \wishbone_bd_ram_mem1_reg[224][15]/P0001  & n13433 ;
  assign n16258 = ~n16256 & ~n16257 ;
  assign n16259 = n16255 & n16258 ;
  assign n16260 = n16252 & n16259 ;
  assign n16261 = n16245 & n16260 ;
  assign n16262 = \wishbone_bd_ram_mem1_reg[211][15]/P0001  & n13805 ;
  assign n16263 = \wishbone_bd_ram_mem1_reg[165][15]/P0001  & n14028 ;
  assign n16264 = ~n16262 & ~n16263 ;
  assign n16265 = \wishbone_bd_ram_mem1_reg[131][15]/P0001  & n13358 ;
  assign n16266 = \wishbone_bd_ram_mem1_reg[107][15]/P0001  & n13476 ;
  assign n16267 = ~n16265 & ~n16266 ;
  assign n16268 = n16264 & n16267 ;
  assign n16269 = \wishbone_bd_ram_mem1_reg[246][15]/P0001  & n13981 ;
  assign n16270 = \wishbone_bd_ram_mem1_reg[205][15]/P0001  & n13947 ;
  assign n16271 = ~n16269 & ~n16270 ;
  assign n16272 = \wishbone_bd_ram_mem1_reg[210][15]/P0001  & n13443 ;
  assign n16273 = \wishbone_bd_ram_mem1_reg[0][15]/P0001  & n13539 ;
  assign n16274 = ~n16272 & ~n16273 ;
  assign n16275 = n16271 & n16274 ;
  assign n16276 = n16268 & n16275 ;
  assign n16277 = \wishbone_bd_ram_mem1_reg[99][15]/P0001  & n13996 ;
  assign n16278 = \wishbone_bd_ram_mem1_reg[168][15]/P0001  & n13795 ;
  assign n16279 = ~n16277 & ~n16278 ;
  assign n16280 = \wishbone_bd_ram_mem1_reg[36][15]/P0001  & n13639 ;
  assign n16281 = \wishbone_bd_ram_mem1_reg[214][15]/P0001  & n13938 ;
  assign n16282 = ~n16280 & ~n16281 ;
  assign n16283 = n16279 & n16282 ;
  assign n16284 = \wishbone_bd_ram_mem1_reg[66][15]/P0001  & n13603 ;
  assign n16285 = \wishbone_bd_ram_mem1_reg[35][15]/P0001  & n13523 ;
  assign n16286 = ~n16284 & ~n16285 ;
  assign n16287 = \wishbone_bd_ram_mem1_reg[40][15]/P0001  & n13661 ;
  assign n16288 = \wishbone_bd_ram_mem1_reg[143][15]/P0001  & n13461 ;
  assign n16289 = ~n16287 & ~n16288 ;
  assign n16290 = n16286 & n16289 ;
  assign n16291 = n16283 & n16290 ;
  assign n16292 = n16276 & n16291 ;
  assign n16293 = n16261 & n16292 ;
  assign n16294 = n16230 & n16293 ;
  assign n16295 = n16167 & n16294 ;
  assign n16296 = n16040 & n16295 ;
  assign n16297 = ~wb_rst_i_pad & ~n15784 ;
  assign n16298 = ~n16296 & n16297 ;
  assign n16299 = ~n15785 & ~n16298 ;
  assign n16300 = \wishbone_RxDataLatched2_reg[9]/NET0131  & ~n15737 ;
  assign n16301 = n15735 & n16300 ;
  assign n16302 = \wishbone_RxDataLatched1_reg[9]/NET0131  & ~n15745 ;
  assign n16303 = ~n15744 & n16302 ;
  assign n16304 = ~n16301 & ~n16303 ;
  assign n16305 = \wishbone_RxPointerRead_reg/NET0131  & n15779 ;
  assign n16306 = ~\wishbone_RxPointerLSB_rst_reg[1]/NET0131  & ~n16305 ;
  assign n16307 = m_wb_ack_i_pad & \wishbone_MasterWbRX_reg/NET0131  ;
  assign n16308 = ~n16306 & ~n16307 ;
  assign n16309 = ~n16305 & n16308 ;
  assign n16310 = \wishbone_bd_ram_mem0_reg[166][1]/P0001  & n13999 ;
  assign n16311 = \wishbone_bd_ram_mem0_reg[57][1]/P0001  & n13731 ;
  assign n16312 = ~n16310 & ~n16311 ;
  assign n16313 = \wishbone_bd_ram_mem0_reg[50][1]/P0001  & n13686 ;
  assign n16314 = \wishbone_bd_ram_mem0_reg[216][1]/P0001  & n14005 ;
  assign n16315 = ~n16313 & ~n16314 ;
  assign n16316 = n16312 & n16315 ;
  assign n16317 = \wishbone_bd_ram_mem0_reg[201][1]/P0001  & n13600 ;
  assign n16318 = \wishbone_bd_ram_mem0_reg[122][1]/P0001  & n13679 ;
  assign n16319 = ~n16317 & ~n16318 ;
  assign n16320 = \wishbone_bd_ram_mem0_reg[130][1]/P0001  & n13427 ;
  assign n16321 = \wishbone_bd_ram_mem0_reg[13][1]/P0001  & n13844 ;
  assign n16322 = ~n16320 & ~n16321 ;
  assign n16323 = n16319 & n16322 ;
  assign n16324 = n16316 & n16323 ;
  assign n16325 = \wishbone_bd_ram_mem0_reg[19][1]/P0001  & n13886 ;
  assign n16326 = \wishbone_bd_ram_mem0_reg[40][1]/P0001  & n13661 ;
  assign n16327 = ~n16325 & ~n16326 ;
  assign n16328 = \wishbone_bd_ram_mem0_reg[126][1]/P0001  & n13786 ;
  assign n16329 = \wishbone_bd_ram_mem0_reg[222][1]/P0001  & n13721 ;
  assign n16330 = ~n16328 & ~n16329 ;
  assign n16331 = n16327 & n16330 ;
  assign n16332 = \wishbone_bd_ram_mem0_reg[249][1]/P0001  & n13431 ;
  assign n16333 = \wishbone_bd_ram_mem0_reg[241][1]/P0001  & n13854 ;
  assign n16334 = ~n16332 & ~n16333 ;
  assign n16335 = \wishbone_bd_ram_mem0_reg[168][1]/P0001  & n13795 ;
  assign n16336 = \wishbone_bd_ram_mem0_reg[244][1]/P0001  & n13474 ;
  assign n16337 = ~n16335 & ~n16336 ;
  assign n16338 = n16334 & n16337 ;
  assign n16339 = n16331 & n16338 ;
  assign n16340 = n16324 & n16339 ;
  assign n16341 = \wishbone_bd_ram_mem0_reg[44][1]/P0001  & n13291 ;
  assign n16342 = \wishbone_bd_ram_mem0_reg[33][1]/P0001  & n13933 ;
  assign n16343 = ~n16341 & ~n16342 ;
  assign n16344 = \wishbone_bd_ram_mem0_reg[17][1]/P0001  & n13324 ;
  assign n16345 = \wishbone_bd_ram_mem0_reg[31][1]/P0001  & n13758 ;
  assign n16346 = ~n16344 & ~n16345 ;
  assign n16347 = n16343 & n16346 ;
  assign n16348 = \wishbone_bd_ram_mem0_reg[7][1]/P0001  & n13546 ;
  assign n16349 = \wishbone_bd_ram_mem0_reg[21][1]/P0001  & n13438 ;
  assign n16350 = ~n16348 & ~n16349 ;
  assign n16351 = \wishbone_bd_ram_mem0_reg[217][1]/P0001  & n13767 ;
  assign n16352 = \wishbone_bd_ram_mem0_reg[85][1]/P0001  & n13784 ;
  assign n16353 = ~n16351 & ~n16352 ;
  assign n16354 = n16350 & n16353 ;
  assign n16355 = n16347 & n16354 ;
  assign n16356 = \wishbone_bd_ram_mem0_reg[84][1]/P0001  & n13385 ;
  assign n16357 = \wishbone_bd_ram_mem0_reg[35][1]/P0001  & n13523 ;
  assign n16358 = ~n16356 & ~n16357 ;
  assign n16359 = \wishbone_bd_ram_mem0_reg[187][1]/P0001  & n13756 ;
  assign n16360 = \wishbone_bd_ram_mem0_reg[205][1]/P0001  & n13947 ;
  assign n16361 = ~n16359 & ~n16360 ;
  assign n16362 = n16358 & n16361 ;
  assign n16363 = \wishbone_bd_ram_mem0_reg[3][1]/P0001  & n13354 ;
  assign n16364 = \wishbone_bd_ram_mem0_reg[79][1]/P0001  & n13779 ;
  assign n16365 = ~n16363 & ~n16364 ;
  assign n16366 = \wishbone_bd_ram_mem0_reg[149][1]/P0001  & n13469 ;
  assign n16367 = \wishbone_bd_ram_mem0_reg[46][1]/P0001  & n13298 ;
  assign n16368 = ~n16366 & ~n16367 ;
  assign n16369 = n16365 & n16368 ;
  assign n16370 = n16362 & n16369 ;
  assign n16371 = n16355 & n16370 ;
  assign n16372 = n16340 & n16371 ;
  assign n16373 = \wishbone_bd_ram_mem0_reg[114][1]/P0001  & n13763 ;
  assign n16374 = \wishbone_bd_ram_mem0_reg[226][1]/P0001  & n13668 ;
  assign n16375 = ~n16373 & ~n16374 ;
  assign n16376 = \wishbone_bd_ram_mem0_reg[87][1]/P0001  & n13691 ;
  assign n16377 = \wishbone_bd_ram_mem0_reg[170][1]/P0001  & n14007 ;
  assign n16378 = ~n16376 & ~n16377 ;
  assign n16379 = n16375 & n16378 ;
  assign n16380 = \wishbone_bd_ram_mem0_reg[125][1]/P0001  & n13396 ;
  assign n16381 = \wishbone_bd_ram_mem0_reg[88][1]/P0001  & n13347 ;
  assign n16382 = ~n16380 & ~n16381 ;
  assign n16383 = \wishbone_bd_ram_mem0_reg[159][1]/P0001  & n13627 ;
  assign n16384 = \wishbone_bd_ram_mem0_reg[62][1]/P0001  & n13529 ;
  assign n16385 = ~n16383 & ~n16384 ;
  assign n16386 = n16382 & n16385 ;
  assign n16387 = n16379 & n16386 ;
  assign n16388 = \wishbone_bd_ram_mem0_reg[242][1]/P0001  & n13383 ;
  assign n16389 = \wishbone_bd_ram_mem0_reg[245][1]/P0001  & n13877 ;
  assign n16390 = ~n16388 & ~n16389 ;
  assign n16391 = \wishbone_bd_ram_mem0_reg[123][1]/P0001  & n13749 ;
  assign n16392 = \wishbone_bd_ram_mem0_reg[250][1]/P0001  & n13677 ;
  assign n16393 = ~n16391 & ~n16392 ;
  assign n16394 = n16390 & n16393 ;
  assign n16395 = \wishbone_bd_ram_mem0_reg[109][1]/P0001  & n13306 ;
  assign n16396 = \wishbone_bd_ram_mem0_reg[22][1]/P0001  & n13744 ;
  assign n16397 = ~n16395 & ~n16396 ;
  assign n16398 = \wishbone_bd_ram_mem0_reg[107][1]/P0001  & n13476 ;
  assign n16399 = \wishbone_bd_ram_mem0_reg[184][1]/P0001  & n13960 ;
  assign n16400 = ~n16398 & ~n16399 ;
  assign n16401 = n16397 & n16400 ;
  assign n16402 = n16394 & n16401 ;
  assign n16403 = n16387 & n16402 ;
  assign n16404 = \wishbone_bd_ram_mem0_reg[63][1]/P0001  & n13327 ;
  assign n16405 = \wishbone_bd_ram_mem0_reg[135][1]/P0001  & n13672 ;
  assign n16406 = ~n16404 & ~n16405 ;
  assign n16407 = \wishbone_bd_ram_mem0_reg[58][1]/P0001  & n13949 ;
  assign n16408 = \wishbone_bd_ram_mem0_reg[175][1]/P0001  & n13674 ;
  assign n16409 = ~n16407 & ~n16408 ;
  assign n16410 = n16406 & n16409 ;
  assign n16411 = \wishbone_bd_ram_mem0_reg[55][1]/P0001  & n13618 ;
  assign n16412 = \wishbone_bd_ram_mem0_reg[18][1]/P0001  & n13532 ;
  assign n16413 = ~n16411 & ~n16412 ;
  assign n16414 = \wishbone_bd_ram_mem0_reg[47][1]/P0001  & n13436 ;
  assign n16415 = \wishbone_bd_ram_mem0_reg[143][1]/P0001  & n13461 ;
  assign n16416 = ~n16414 & ~n16415 ;
  assign n16417 = n16413 & n16416 ;
  assign n16418 = n16410 & n16417 ;
  assign n16419 = \wishbone_bd_ram_mem0_reg[225][1]/P0001  & n13719 ;
  assign n16420 = \wishbone_bd_ram_mem0_reg[27][1]/P0001  & n13251 ;
  assign n16421 = ~n16419 & ~n16420 ;
  assign n16422 = \wishbone_bd_ram_mem0_reg[124][1]/P0001  & n14024 ;
  assign n16423 = \wishbone_bd_ram_mem0_reg[177][1]/P0001  & n13863 ;
  assign n16424 = ~n16422 & ~n16423 ;
  assign n16425 = n16421 & n16424 ;
  assign n16426 = \wishbone_bd_ram_mem0_reg[214][1]/P0001  & n13938 ;
  assign n16427 = \wishbone_bd_ram_mem0_reg[196][1]/P0001  & n13977 ;
  assign n16428 = ~n16426 & ~n16427 ;
  assign n16429 = \wishbone_bd_ram_mem0_reg[1][1]/P0001  & n13888 ;
  assign n16430 = \wishbone_bd_ram_mem0_reg[160][1]/P0001  & n13271 ;
  assign n16431 = ~n16429 & ~n16430 ;
  assign n16432 = n16428 & n16431 ;
  assign n16433 = n16425 & n16432 ;
  assign n16434 = n16418 & n16433 ;
  assign n16435 = n16403 & n16434 ;
  assign n16436 = n16372 & n16435 ;
  assign n16437 = \wishbone_bd_ram_mem0_reg[231][1]/P0001  & n13363 ;
  assign n16438 = \wishbone_bd_ram_mem0_reg[45][1]/P0001  & n13420 ;
  assign n16439 = ~n16437 & ~n16438 ;
  assign n16440 = \wishbone_bd_ram_mem0_reg[220][1]/P0001  & n13965 ;
  assign n16441 = \wishbone_bd_ram_mem0_reg[145][1]/P0001  & n13715 ;
  assign n16442 = ~n16440 & ~n16441 ;
  assign n16443 = n16439 & n16442 ;
  assign n16444 = \wishbone_bd_ram_mem0_reg[230][1]/P0001  & n13994 ;
  assign n16445 = \wishbone_bd_ram_mem0_reg[111][1]/P0001  & n13471 ;
  assign n16446 = ~n16444 & ~n16445 ;
  assign n16447 = \wishbone_bd_ram_mem0_reg[199][1]/P0001  & n13499 ;
  assign n16448 = \wishbone_bd_ram_mem0_reg[146][1]/P0001  & n13958 ;
  assign n16449 = ~n16447 & ~n16448 ;
  assign n16450 = n16446 & n16449 ;
  assign n16451 = n16443 & n16450 ;
  assign n16452 = \wishbone_bd_ram_mem0_reg[215][1]/P0001  & n13901 ;
  assign n16453 = \wishbone_bd_ram_mem0_reg[238][1]/P0001  & n13819 ;
  assign n16454 = ~n16452 & ~n16453 ;
  assign n16455 = \wishbone_bd_ram_mem0_reg[252][1]/P0001  & n13986 ;
  assign n16456 = \wishbone_bd_ram_mem0_reg[52][1]/P0001  & n13988 ;
  assign n16457 = ~n16455 & ~n16456 ;
  assign n16458 = n16454 & n16457 ;
  assign n16459 = \wishbone_bd_ram_mem0_reg[53][1]/P0001  & n13875 ;
  assign n16460 = \wishbone_bd_ram_mem0_reg[69][1]/P0001  & n13487 ;
  assign n16461 = ~n16459 & ~n16460 ;
  assign n16462 = \wishbone_bd_ram_mem0_reg[42][1]/P0001  & n13341 ;
  assign n16463 = \wishbone_bd_ram_mem0_reg[213][1]/P0001  & n13870 ;
  assign n16464 = ~n16462 & ~n16463 ;
  assign n16465 = n16461 & n16464 ;
  assign n16466 = n16458 & n16465 ;
  assign n16467 = n16451 & n16466 ;
  assign n16468 = \wishbone_bd_ram_mem0_reg[197][1]/P0001  & n13594 ;
  assign n16469 = \wishbone_bd_ram_mem0_reg[16][1]/P0001  & n13695 ;
  assign n16470 = ~n16468 & ~n16469 ;
  assign n16471 = \wishbone_bd_ram_mem0_reg[2][1]/P0001  & n13975 ;
  assign n16472 = \wishbone_bd_ram_mem0_reg[198][1]/P0001  & n13592 ;
  assign n16473 = ~n16471 & ~n16472 ;
  assign n16474 = n16470 & n16473 ;
  assign n16475 = \wishbone_bd_ram_mem0_reg[108][1]/P0001  & n13814 ;
  assign n16476 = \wishbone_bd_ram_mem0_reg[200][1]/P0001  & n13922 ;
  assign n16477 = ~n16475 & ~n16476 ;
  assign n16478 = \wishbone_bd_ram_mem0_reg[90][1]/P0001  & n13906 ;
  assign n16479 = \wishbone_bd_ram_mem0_reg[247][1]/P0001  & n13571 ;
  assign n16480 = ~n16478 & ~n16479 ;
  assign n16481 = n16477 & n16480 ;
  assign n16482 = n16474 & n16481 ;
  assign n16483 = \wishbone_bd_ram_mem0_reg[72][1]/P0001  & n13582 ;
  assign n16484 = \wishbone_bd_ram_mem0_reg[163][1]/P0001  & n13255 ;
  assign n16485 = ~n16483 & ~n16484 ;
  assign n16486 = \wishbone_bd_ram_mem0_reg[161][1]/P0001  & n13505 ;
  assign n16487 = \wishbone_bd_ram_mem0_reg[75][1]/P0001  & n13605 ;
  assign n16488 = ~n16486 & ~n16487 ;
  assign n16489 = n16485 & n16488 ;
  assign n16490 = \wishbone_bd_ram_mem0_reg[60][1]/P0001  & n13790 ;
  assign n16491 = \wishbone_bd_ram_mem0_reg[229][1]/P0001  & n13552 ;
  assign n16492 = ~n16490 & ~n16491 ;
  assign n16493 = \wishbone_bd_ram_mem0_reg[104][1]/P0001  & n13684 ;
  assign n16494 = \wishbone_bd_ram_mem0_reg[11][1]/P0001  & n13774 ;
  assign n16495 = ~n16493 & ~n16494 ;
  assign n16496 = n16492 & n16495 ;
  assign n16497 = n16489 & n16496 ;
  assign n16498 = n16482 & n16497 ;
  assign n16499 = n16467 & n16498 ;
  assign n16500 = \wishbone_bd_ram_mem0_reg[115][1]/P0001  & n13747 ;
  assign n16501 = \wishbone_bd_ram_mem0_reg[100][1]/P0001  & n13401 ;
  assign n16502 = ~n16500 & ~n16501 ;
  assign n16503 = \wishbone_bd_ram_mem0_reg[38][1]/P0001  & n13828 ;
  assign n16504 = \wishbone_bd_ram_mem0_reg[12][1]/P0001  & n13733 ;
  assign n16505 = ~n16503 & ~n16504 ;
  assign n16506 = n16502 & n16505 ;
  assign n16507 = \wishbone_bd_ram_mem0_reg[174][1]/P0001  & n13899 ;
  assign n16508 = \wishbone_bd_ram_mem0_reg[105][1]/P0001  & n13503 ;
  assign n16509 = ~n16507 & ~n16508 ;
  assign n16510 = \wishbone_bd_ram_mem0_reg[127][1]/P0001  & n13803 ;
  assign n16511 = \wishbone_bd_ram_mem0_reg[140][1]/P0001  & n13287 ;
  assign n16512 = ~n16510 & ~n16511 ;
  assign n16513 = n16509 & n16512 ;
  assign n16514 = n16506 & n16513 ;
  assign n16515 = \wishbone_bd_ram_mem0_reg[181][1]/P0001  & n13587 ;
  assign n16516 = \wishbone_bd_ram_mem0_reg[151][1]/P0001  & n13697 ;
  assign n16517 = ~n16515 & ~n16516 ;
  assign n16518 = \wishbone_bd_ram_mem0_reg[167][1]/P0001  & n13940 ;
  assign n16519 = \wishbone_bd_ram_mem0_reg[171][1]/P0001  & n13422 ;
  assign n16520 = ~n16518 & ~n16519 ;
  assign n16521 = n16517 & n16520 ;
  assign n16522 = \wishbone_bd_ram_mem0_reg[95][1]/P0001  & n13317 ;
  assign n16523 = \wishbone_bd_ram_mem0_reg[14][1]/P0001  & n13972 ;
  assign n16524 = ~n16522 & ~n16523 ;
  assign n16525 = \wishbone_bd_ram_mem0_reg[248][1]/P0001  & n13647 ;
  assign n16526 = \wishbone_bd_ram_mem0_reg[190][1]/P0001  & n13365 ;
  assign n16527 = ~n16525 & ~n16526 ;
  assign n16528 = n16524 & n16527 ;
  assign n16529 = n16521 & n16528 ;
  assign n16530 = n16514 & n16529 ;
  assign n16531 = \wishbone_bd_ram_mem0_reg[34][1]/P0001  & n13450 ;
  assign n16532 = \wishbone_bd_ram_mem0_reg[137][1]/P0001  & n13808 ;
  assign n16533 = ~n16531 & ~n16532 ;
  assign n16534 = \wishbone_bd_ram_mem0_reg[59][1]/P0001  & n13613 ;
  assign n16535 = \wishbone_bd_ram_mem0_reg[94][1]/P0001  & n13833 ;
  assign n16536 = ~n16534 & ~n16535 ;
  assign n16537 = n16533 & n16536 ;
  assign n16538 = \wishbone_bd_ram_mem0_reg[54][1]/P0001  & n13622 ;
  assign n16539 = \wishbone_bd_ram_mem0_reg[73][1]/P0001  & n13456 ;
  assign n16540 = ~n16538 & ~n16539 ;
  assign n16541 = \wishbone_bd_ram_mem0_reg[129][1]/P0001  & n13629 ;
  assign n16542 = \wishbone_bd_ram_mem0_reg[91][1]/P0001  & n13954 ;
  assign n16543 = ~n16541 & ~n16542 ;
  assign n16544 = n16540 & n16543 ;
  assign n16545 = n16537 & n16544 ;
  assign n16546 = \wishbone_bd_ram_mem0_reg[141][1]/P0001  & n13852 ;
  assign n16547 = \wishbone_bd_ram_mem0_reg[193][1]/P0001  & n14022 ;
  assign n16548 = ~n16546 & ~n16547 ;
  assign n16549 = \wishbone_bd_ram_mem0_reg[51][1]/P0001  & n13880 ;
  assign n16550 = \wishbone_bd_ram_mem0_reg[218][1]/P0001  & n13792 ;
  assign n16551 = ~n16549 & ~n16550 ;
  assign n16552 = n16548 & n16551 ;
  assign n16553 = \wishbone_bd_ram_mem0_reg[5][1]/P0001  & n13243 ;
  assign n16554 = \wishbone_bd_ram_mem0_reg[155][1]/P0001  & n13738 ;
  assign n16555 = ~n16553 & ~n16554 ;
  assign n16556 = \wishbone_bd_ram_mem0_reg[255][1]/P0001  & n13952 ;
  assign n16557 = \wishbone_bd_ram_mem0_reg[89][1]/P0001  & n13910 ;
  assign n16558 = ~n16556 & ~n16557 ;
  assign n16559 = n16555 & n16558 ;
  assign n16560 = n16552 & n16559 ;
  assign n16561 = n16545 & n16560 ;
  assign n16562 = n16530 & n16561 ;
  assign n16563 = n16499 & n16562 ;
  assign n16564 = n16436 & n16563 ;
  assign n16565 = \wishbone_bd_ram_mem0_reg[224][1]/P0001  & n13433 ;
  assign n16566 = \wishbone_bd_ram_mem0_reg[30][1]/P0001  & n13713 ;
  assign n16567 = ~n16565 & ~n16566 ;
  assign n16568 = \wishbone_bd_ram_mem0_reg[237][1]/P0001  & n13924 ;
  assign n16569 = \wishbone_bd_ram_mem0_reg[234][1]/P0001  & n13781 ;
  assign n16570 = ~n16568 & ~n16569 ;
  assign n16571 = n16567 & n16570 ;
  assign n16572 = \wishbone_bd_ram_mem0_reg[180][1]/P0001  & n13650 ;
  assign n16573 = \wishbone_bd_ram_mem0_reg[120][1]/P0001  & n13550 ;
  assign n16574 = ~n16572 & ~n16573 ;
  assign n16575 = \wishbone_bd_ram_mem0_reg[221][1]/P0001  & n13641 ;
  assign n16576 = \wishbone_bd_ram_mem0_reg[202][1]/P0001  & n13268 ;
  assign n16577 = ~n16575 & ~n16576 ;
  assign n16578 = n16574 & n16577 ;
  assign n16579 = n16571 & n16578 ;
  assign n16580 = \wishbone_bd_ram_mem0_reg[49][1]/P0001  & n13929 ;
  assign n16581 = \wishbone_bd_ram_mem0_reg[153][1]/P0001  & n13309 ;
  assign n16582 = ~n16580 & ~n16581 ;
  assign n16583 = \wishbone_bd_ram_mem0_reg[77][1]/P0001  & n13935 ;
  assign n16584 = \wishbone_bd_ram_mem0_reg[172][1]/P0001  & n13377 ;
  assign n16585 = ~n16583 & ~n16584 ;
  assign n16586 = n16582 & n16585 ;
  assign n16587 = \wishbone_bd_ram_mem0_reg[86][1]/P0001  & n13485 ;
  assign n16588 = \wishbone_bd_ram_mem0_reg[118][1]/P0001  & n13589 ;
  assign n16589 = ~n16587 & ~n16588 ;
  assign n16590 = \wishbone_bd_ram_mem0_reg[99][1]/P0001  & n13996 ;
  assign n16591 = \wishbone_bd_ram_mem0_reg[206][1]/P0001  & n13414 ;
  assign n16592 = ~n16590 & ~n16591 ;
  assign n16593 = n16589 & n16592 ;
  assign n16594 = n16586 & n16593 ;
  assign n16595 = n16579 & n16594 ;
  assign n16596 = \wishbone_bd_ram_mem0_reg[176][1]/P0001  & n13262 ;
  assign n16597 = \wishbone_bd_ram_mem0_reg[204][1]/P0001  & n13821 ;
  assign n16598 = ~n16596 & ~n16597 ;
  assign n16599 = \wishbone_bd_ram_mem0_reg[211][1]/P0001  & n13805 ;
  assign n16600 = \wishbone_bd_ram_mem0_reg[121][1]/P0001  & n13983 ;
  assign n16601 = ~n16599 & ~n16600 ;
  assign n16602 = n16598 & n16601 ;
  assign n16603 = \wishbone_bd_ram_mem0_reg[81][1]/P0001  & n13409 ;
  assign n16604 = \wishbone_bd_ram_mem0_reg[132][1]/P0001  & n13927 ;
  assign n16605 = ~n16603 & ~n16604 ;
  assign n16606 = \wishbone_bd_ram_mem0_reg[66][1]/P0001  & n13603 ;
  assign n16607 = \wishbone_bd_ram_mem0_reg[70][1]/P0001  & n13339 ;
  assign n16608 = ~n16606 & ~n16607 ;
  assign n16609 = n16605 & n16608 ;
  assign n16610 = n16602 & n16609 ;
  assign n16611 = \wishbone_bd_ram_mem0_reg[80][1]/P0001  & n13516 ;
  assign n16612 = \wishbone_bd_ram_mem0_reg[144][1]/P0001  & n13508 ;
  assign n16613 = ~n16611 & ~n16612 ;
  assign n16614 = \wishbone_bd_ram_mem0_reg[112][1]/P0001  & n13482 ;
  assign n16615 = \wishbone_bd_ram_mem0_reg[10][1]/P0001  & n13837 ;
  assign n16616 = ~n16614 & ~n16615 ;
  assign n16617 = n16613 & n16616 ;
  assign n16618 = \wishbone_bd_ram_mem0_reg[25][1]/P0001  & n13742 ;
  assign n16619 = \wishbone_bd_ram_mem0_reg[207][1]/P0001  & n13826 ;
  assign n16620 = ~n16618 & ~n16619 ;
  assign n16621 = \wishbone_bd_ram_mem0_reg[233][1]/P0001  & n13332 ;
  assign n16622 = \wishbone_bd_ram_mem0_reg[194][1]/P0001  & n13624 ;
  assign n16623 = ~n16621 & ~n16622 ;
  assign n16624 = n16620 & n16623 ;
  assign n16625 = n16617 & n16624 ;
  assign n16626 = n16610 & n16625 ;
  assign n16627 = n16595 & n16626 ;
  assign n16628 = \wishbone_bd_ram_mem0_reg[240][1]/P0001  & n13352 ;
  assign n16629 = \wishbone_bd_ram_mem0_reg[32][1]/P0001  & n13736 ;
  assign n16630 = ~n16628 & ~n16629 ;
  assign n16631 = \wishbone_bd_ram_mem0_reg[106][1]/P0001  & n13555 ;
  assign n16632 = \wishbone_bd_ram_mem0_reg[185][1]/P0001  & n13372 ;
  assign n16633 = ~n16631 & ~n16632 ;
  assign n16634 = n16630 & n16633 ;
  assign n16635 = \wishbone_bd_ram_mem0_reg[92][1]/P0001  & n13859 ;
  assign n16636 = \wishbone_bd_ram_mem0_reg[37][1]/P0001  & n13710 ;
  assign n16637 = ~n16635 & ~n16636 ;
  assign n16638 = \wishbone_bd_ram_mem0_reg[82][1]/P0001  & n13374 ;
  assign n16639 = \wishbone_bd_ram_mem0_reg[117][1]/P0001  & n13557 ;
  assign n16640 = ~n16638 & ~n16639 ;
  assign n16641 = n16637 & n16640 ;
  assign n16642 = n16634 & n16641 ;
  assign n16643 = \wishbone_bd_ram_mem0_reg[173][1]/P0001  & n13360 ;
  assign n16644 = \wishbone_bd_ram_mem0_reg[136][1]/P0001  & n13963 ;
  assign n16645 = ~n16643 & ~n16644 ;
  assign n16646 = \wishbone_bd_ram_mem0_reg[9][1]/P0001  & n13580 ;
  assign n16647 = \wishbone_bd_ram_mem0_reg[131][1]/P0001  & n13358 ;
  assign n16648 = ~n16646 & ~n16647 ;
  assign n16649 = n16645 & n16648 ;
  assign n16650 = \wishbone_bd_ram_mem0_reg[20][1]/P0001  & n13839 ;
  assign n16651 = \wishbone_bd_ram_mem0_reg[36][1]/P0001  & n13639 ;
  assign n16652 = ~n16650 & ~n16651 ;
  assign n16653 = \wishbone_bd_ram_mem0_reg[28][1]/P0001  & n13810 ;
  assign n16654 = \wishbone_bd_ram_mem0_reg[101][1]/P0001  & n13772 ;
  assign n16655 = ~n16653 & ~n16654 ;
  assign n16656 = n16652 & n16655 ;
  assign n16657 = n16649 & n16656 ;
  assign n16658 = n16642 & n16657 ;
  assign n16659 = \wishbone_bd_ram_mem0_reg[192][1]/P0001  & n13390 ;
  assign n16660 = \wishbone_bd_ram_mem0_reg[0][1]/P0001  & n13539 ;
  assign n16661 = ~n16659 & ~n16660 ;
  assign n16662 = \wishbone_bd_ram_mem0_reg[195][1]/P0001  & n13700 ;
  assign n16663 = \wishbone_bd_ram_mem0_reg[178][1]/P0001  & n13301 ;
  assign n16664 = ~n16662 & ~n16663 ;
  assign n16665 = n16661 & n16664 ;
  assign n16666 = \wishbone_bd_ram_mem0_reg[98][1]/P0001  & n13569 ;
  assign n16667 = \wishbone_bd_ram_mem0_reg[203][1]/P0001  & n13816 ;
  assign n16668 = ~n16666 & ~n16667 ;
  assign n16669 = \wishbone_bd_ram_mem0_reg[253][1]/P0001  & n13708 ;
  assign n16670 = \wishbone_bd_ram_mem0_reg[156][1]/P0001  & n13769 ;
  assign n16671 = ~n16669 & ~n16670 ;
  assign n16672 = n16668 & n16671 ;
  assign n16673 = n16665 & n16672 ;
  assign n16674 = \wishbone_bd_ram_mem0_reg[15][1]/P0001  & n13797 ;
  assign n16675 = \wishbone_bd_ram_mem0_reg[39][1]/P0001  & n13893 ;
  assign n16676 = ~n16674 & ~n16675 ;
  assign n16677 = \wishbone_bd_ram_mem0_reg[186][1]/P0001  & n13616 ;
  assign n16678 = \wishbone_bd_ram_mem0_reg[138][1]/P0001  & n13398 ;
  assign n16679 = ~n16677 & ~n16678 ;
  assign n16680 = n16676 & n16679 ;
  assign n16681 = \wishbone_bd_ram_mem0_reg[246][1]/P0001  & n13981 ;
  assign n16682 = \wishbone_bd_ram_mem0_reg[179][1]/P0001  & n14035 ;
  assign n16683 = ~n16681 & ~n16682 ;
  assign n16684 = \wishbone_bd_ram_mem0_reg[189][1]/P0001  & n14001 ;
  assign n16685 = \wishbone_bd_ram_mem0_reg[183][1]/P0001  & n13645 ;
  assign n16686 = ~n16684 & ~n16685 ;
  assign n16687 = n16683 & n16686 ;
  assign n16688 = n16680 & n16687 ;
  assign n16689 = n16673 & n16688 ;
  assign n16690 = n16658 & n16689 ;
  assign n16691 = n16627 & n16690 ;
  assign n16692 = \wishbone_bd_ram_mem0_reg[102][1]/P0001  & n13534 ;
  assign n16693 = \wishbone_bd_ram_mem0_reg[134][1]/P0001  & n13494 ;
  assign n16694 = ~n16692 & ~n16693 ;
  assign n16695 = \wishbone_bd_ram_mem0_reg[93][1]/P0001  & n13891 ;
  assign n16696 = \wishbone_bd_ram_mem0_reg[162][1]/P0001  & n13726 ;
  assign n16697 = ~n16695 & ~n16696 ;
  assign n16698 = n16694 & n16697 ;
  assign n16699 = \wishbone_bd_ram_mem0_reg[61][1]/P0001  & n13544 ;
  assign n16700 = \wishbone_bd_ram_mem0_reg[158][1]/P0001  & n13294 ;
  assign n16701 = ~n16699 & ~n16700 ;
  assign n16702 = \wishbone_bd_ram_mem0_reg[148][1]/P0001  & n13868 ;
  assign n16703 = \wishbone_bd_ram_mem0_reg[142][1]/P0001  & n13448 ;
  assign n16704 = ~n16702 & ~n16703 ;
  assign n16705 = n16701 & n16704 ;
  assign n16706 = n16698 & n16705 ;
  assign n16707 = \wishbone_bd_ram_mem0_reg[48][1]/P0001  & n13917 ;
  assign n16708 = \wishbone_bd_ram_mem0_reg[232][1]/P0001  & n13510 ;
  assign n16709 = ~n16707 & ~n16708 ;
  assign n16710 = \wishbone_bd_ram_mem0_reg[154][1]/P0001  & n13403 ;
  assign n16711 = \wishbone_bd_ram_mem0_reg[113][1]/P0001  & n13882 ;
  assign n16712 = ~n16710 & ~n16711 ;
  assign n16713 = n16709 & n16712 ;
  assign n16714 = \wishbone_bd_ram_mem0_reg[188][1]/P0001  & n13407 ;
  assign n16715 = \wishbone_bd_ram_mem0_reg[223][1]/P0001  & n13335 ;
  assign n16716 = ~n16714 & ~n16715 ;
  assign n16717 = \wishbone_bd_ram_mem0_reg[227][1]/P0001  & n13388 ;
  assign n16718 = \wishbone_bd_ram_mem0_reg[24][1]/P0001  & n13970 ;
  assign n16719 = ~n16717 & ~n16718 ;
  assign n16720 = n16716 & n16719 ;
  assign n16721 = n16713 & n16720 ;
  assign n16722 = n16706 & n16721 ;
  assign n16723 = \wishbone_bd_ram_mem0_reg[191][1]/P0001  & n14012 ;
  assign n16724 = \wishbone_bd_ram_mem0_reg[139][1]/P0001  & n13566 ;
  assign n16725 = ~n16723 & ~n16724 ;
  assign n16726 = \wishbone_bd_ram_mem0_reg[182][1]/P0001  & n13598 ;
  assign n16727 = \wishbone_bd_ram_mem0_reg[119][1]/P0001  & n14033 ;
  assign n16728 = ~n16726 & ~n16727 ;
  assign n16729 = n16725 & n16728 ;
  assign n16730 = \wishbone_bd_ram_mem0_reg[29][1]/P0001  & n13412 ;
  assign n16731 = \wishbone_bd_ram_mem0_reg[152][1]/P0001  & n13912 ;
  assign n16732 = ~n16730 & ~n16731 ;
  assign n16733 = \wishbone_bd_ram_mem0_reg[239][1]/P0001  & n13349 ;
  assign n16734 = \wishbone_bd_ram_mem0_reg[219][1]/P0001  & n13577 ;
  assign n16735 = ~n16733 & ~n16734 ;
  assign n16736 = n16732 & n16735 ;
  assign n16737 = n16729 & n16736 ;
  assign n16738 = \wishbone_bd_ram_mem0_reg[243][1]/P0001  & n13575 ;
  assign n16739 = \wishbone_bd_ram_mem0_reg[150][1]/P0001  & n13666 ;
  assign n16740 = ~n16738 & ~n16739 ;
  assign n16741 = \wishbone_bd_ram_mem0_reg[251][1]/P0001  & n14019 ;
  assign n16742 = \wishbone_bd_ram_mem0_reg[43][1]/P0001  & n13761 ;
  assign n16743 = ~n16741 & ~n16742 ;
  assign n16744 = n16740 & n16743 ;
  assign n16745 = \wishbone_bd_ram_mem0_reg[103][1]/P0001  & n13320 ;
  assign n16746 = \wishbone_bd_ram_mem0_reg[96][1]/P0001  & n13425 ;
  assign n16747 = ~n16745 & ~n16746 ;
  assign n16748 = \wishbone_bd_ram_mem0_reg[83][1]/P0001  & n13454 ;
  assign n16749 = \wishbone_bd_ram_mem0_reg[133][1]/P0001  & n13492 ;
  assign n16750 = ~n16748 & ~n16749 ;
  assign n16751 = n16747 & n16750 ;
  assign n16752 = n16744 & n16751 ;
  assign n16753 = n16737 & n16752 ;
  assign n16754 = n16722 & n16753 ;
  assign n16755 = \wishbone_bd_ram_mem0_reg[64][1]/P0001  & n13904 ;
  assign n16756 = \wishbone_bd_ram_mem0_reg[209][1]/P0001  & n13689 ;
  assign n16757 = ~n16755 & ~n16756 ;
  assign n16758 = \wishbone_bd_ram_mem0_reg[78][1]/P0001  & n13277 ;
  assign n16759 = \wishbone_bd_ram_mem0_reg[116][1]/P0001  & n13865 ;
  assign n16760 = ~n16758 & ~n16759 ;
  assign n16761 = n16757 & n16760 ;
  assign n16762 = \wishbone_bd_ram_mem0_reg[56][1]/P0001  & n13611 ;
  assign n16763 = \wishbone_bd_ram_mem0_reg[147][1]/P0001  & n13702 ;
  assign n16764 = ~n16762 & ~n16763 ;
  assign n16765 = \wishbone_bd_ram_mem0_reg[210][1]/P0001  & n13443 ;
  assign n16766 = \wishbone_bd_ram_mem0_reg[157][1]/P0001  & n13445 ;
  assign n16767 = ~n16765 & ~n16766 ;
  assign n16768 = n16764 & n16767 ;
  assign n16769 = n16761 & n16768 ;
  assign n16770 = \wishbone_bd_ram_mem0_reg[4][1]/P0001  & n13527 ;
  assign n16771 = \wishbone_bd_ram_mem0_reg[6][1]/P0001  & n13915 ;
  assign n16772 = ~n16770 & ~n16771 ;
  assign n16773 = \wishbone_bd_ram_mem0_reg[26][1]/P0001  & n13521 ;
  assign n16774 = \wishbone_bd_ram_mem0_reg[74][1]/P0001  & n13564 ;
  assign n16775 = ~n16773 & ~n16774 ;
  assign n16776 = n16772 & n16775 ;
  assign n16777 = \wishbone_bd_ram_mem0_reg[71][1]/P0001  & n13636 ;
  assign n16778 = \wishbone_bd_ram_mem0_reg[235][1]/P0001  & n13518 ;
  assign n16779 = ~n16777 & ~n16778 ;
  assign n16780 = \wishbone_bd_ram_mem0_reg[228][1]/P0001  & n13497 ;
  assign n16781 = \wishbone_bd_ram_mem0_reg[128][1]/P0001  & n13652 ;
  assign n16782 = ~n16780 & ~n16781 ;
  assign n16783 = n16779 & n16782 ;
  assign n16784 = n16776 & n16783 ;
  assign n16785 = n16769 & n16784 ;
  assign n16786 = \wishbone_bd_ram_mem0_reg[212][1]/P0001  & n13634 ;
  assign n16787 = \wishbone_bd_ram_mem0_reg[208][1]/P0001  & n14010 ;
  assign n16788 = ~n16786 & ~n16787 ;
  assign n16789 = \wishbone_bd_ram_mem0_reg[68][1]/P0001  & n13379 ;
  assign n16790 = \wishbone_bd_ram_mem0_reg[67][1]/P0001  & n13663 ;
  assign n16791 = ~n16789 & ~n16790 ;
  assign n16792 = n16788 & n16791 ;
  assign n16793 = \wishbone_bd_ram_mem0_reg[165][1]/P0001  & n14028 ;
  assign n16794 = \wishbone_bd_ram_mem0_reg[164][1]/P0001  & n13236 ;
  assign n16795 = ~n16793 & ~n16794 ;
  assign n16796 = \wishbone_bd_ram_mem0_reg[76][1]/P0001  & n13831 ;
  assign n16797 = \wishbone_bd_ram_mem0_reg[8][1]/P0001  & n13459 ;
  assign n16798 = ~n16796 & ~n16797 ;
  assign n16799 = n16795 & n16798 ;
  assign n16800 = n16792 & n16799 ;
  assign n16801 = \wishbone_bd_ram_mem0_reg[110][1]/P0001  & n14030 ;
  assign n16802 = \wishbone_bd_ram_mem0_reg[23][1]/P0001  & n13857 ;
  assign n16803 = ~n16801 & ~n16802 ;
  assign n16804 = \wishbone_bd_ram_mem0_reg[97][1]/P0001  & n13724 ;
  assign n16805 = \wishbone_bd_ram_mem0_reg[254][1]/P0001  & n13283 ;
  assign n16806 = ~n16804 & ~n16805 ;
  assign n16807 = n16803 & n16806 ;
  assign n16808 = \wishbone_bd_ram_mem0_reg[169][1]/P0001  & n13541 ;
  assign n16809 = \wishbone_bd_ram_mem0_reg[41][1]/P0001  & n14017 ;
  assign n16810 = ~n16808 & ~n16809 ;
  assign n16811 = \wishbone_bd_ram_mem0_reg[236][1]/P0001  & n13480 ;
  assign n16812 = \wishbone_bd_ram_mem0_reg[65][1]/P0001  & n13842 ;
  assign n16813 = ~n16811 & ~n16812 ;
  assign n16814 = n16810 & n16813 ;
  assign n16815 = n16807 & n16814 ;
  assign n16816 = n16800 & n16815 ;
  assign n16817 = n16785 & n16816 ;
  assign n16818 = n16754 & n16817 ;
  assign n16819 = n16691 & n16818 ;
  assign n16820 = n16564 & n16819 ;
  assign n16821 = ~wb_rst_i_pad & n16308 ;
  assign n16822 = ~n16820 & n16821 ;
  assign n16823 = ~n16309 & ~n16822 ;
  assign n16824 = ~\rxethmac1_crcrx_Crc_reg[21]/NET0131  & n12133 ;
  assign n16825 = n11353 & n16824 ;
  assign n16826 = ~\rxethmac1_crcrx_Crc_reg[21]/NET0131  & n10663 ;
  assign n16827 = ~n12257 & ~n16826 ;
  assign n16828 = ~n16825 & ~n16827 ;
  assign n16829 = ~\txethmac1_txcrc_Crc_reg[4]/NET0131  & n13011 ;
  assign n16830 = n12998 & n16829 ;
  assign n16831 = ~\txethmac1_txcrc_Crc_reg[4]/NET0131  & n11464 ;
  assign n16832 = ~n13016 & ~n16831 ;
  assign n16833 = ~n16830 & ~n16832 ;
  assign n16834 = \m_wb_adr_o[16]_pad  & \m_wb_adr_o[17]_pad  ;
  assign n16835 = n13107 & n16834 ;
  assign n16836 = ~\m_wb_adr_o[18]_pad  & ~n16835 ;
  assign n16837 = \m_wb_adr_o[16]_pad  & n13108 ;
  assign n16838 = n13107 & n16837 ;
  assign n16839 = ~n15177 & ~n16838 ;
  assign n16840 = ~n16836 & n16839 ;
  assign n16841 = \m_wb_adr_o[18]_pad  & n13197 ;
  assign n16842 = \wishbone_RxPointerMSB_reg[18]/NET0131  & n13207 ;
  assign n16843 = ~n13196 & n16842 ;
  assign n16844 = \wishbone_TxPointerMSB_reg[18]/NET0131  & ~n13201 ;
  assign n16845 = ~n16843 & ~n16844 ;
  assign n16846 = ~n16841 & n16845 ;
  assign n16847 = ~n16840 & n16846 ;
  assign n16848 = \wishbone_bd_ram_mem2_reg[67][20]/P0001  & n13663 ;
  assign n16849 = \wishbone_bd_ram_mem2_reg[113][20]/P0001  & n13882 ;
  assign n16850 = ~n16848 & ~n16849 ;
  assign n16851 = \wishbone_bd_ram_mem2_reg[140][20]/P0001  & n13287 ;
  assign n16852 = \wishbone_bd_ram_mem2_reg[245][20]/P0001  & n13877 ;
  assign n16853 = ~n16851 & ~n16852 ;
  assign n16854 = n16850 & n16853 ;
  assign n16855 = \wishbone_bd_ram_mem2_reg[99][20]/P0001  & n13996 ;
  assign n16856 = \wishbone_bd_ram_mem2_reg[133][20]/P0001  & n13492 ;
  assign n16857 = ~n16855 & ~n16856 ;
  assign n16858 = \wishbone_bd_ram_mem2_reg[43][20]/P0001  & n13761 ;
  assign n16859 = \wishbone_bd_ram_mem2_reg[34][20]/P0001  & n13450 ;
  assign n16860 = ~n16858 & ~n16859 ;
  assign n16861 = n16857 & n16860 ;
  assign n16862 = n16854 & n16861 ;
  assign n16863 = \wishbone_bd_ram_mem2_reg[252][20]/P0001  & n13986 ;
  assign n16864 = \wishbone_bd_ram_mem2_reg[3][20]/P0001  & n13354 ;
  assign n16865 = ~n16863 & ~n16864 ;
  assign n16866 = \wishbone_bd_ram_mem2_reg[180][20]/P0001  & n13650 ;
  assign n16867 = \wishbone_bd_ram_mem2_reg[83][20]/P0001  & n13454 ;
  assign n16868 = ~n16866 & ~n16867 ;
  assign n16869 = n16865 & n16868 ;
  assign n16870 = \wishbone_bd_ram_mem2_reg[87][20]/P0001  & n13691 ;
  assign n16871 = \wishbone_bd_ram_mem2_reg[194][20]/P0001  & n13624 ;
  assign n16872 = ~n16870 & ~n16871 ;
  assign n16873 = \wishbone_bd_ram_mem2_reg[32][20]/P0001  & n13736 ;
  assign n16874 = \wishbone_bd_ram_mem2_reg[29][20]/P0001  & n13412 ;
  assign n16875 = ~n16873 & ~n16874 ;
  assign n16876 = n16872 & n16875 ;
  assign n16877 = n16869 & n16876 ;
  assign n16878 = n16862 & n16877 ;
  assign n16879 = \wishbone_bd_ram_mem2_reg[9][20]/P0001  & n13580 ;
  assign n16880 = \wishbone_bd_ram_mem2_reg[135][20]/P0001  & n13672 ;
  assign n16881 = ~n16879 & ~n16880 ;
  assign n16882 = \wishbone_bd_ram_mem2_reg[0][20]/P0001  & n13539 ;
  assign n16883 = \wishbone_bd_ram_mem2_reg[19][20]/P0001  & n13886 ;
  assign n16884 = ~n16882 & ~n16883 ;
  assign n16885 = n16881 & n16884 ;
  assign n16886 = \wishbone_bd_ram_mem2_reg[53][20]/P0001  & n13875 ;
  assign n16887 = \wishbone_bd_ram_mem2_reg[164][20]/P0001  & n13236 ;
  assign n16888 = ~n16886 & ~n16887 ;
  assign n16889 = \wishbone_bd_ram_mem2_reg[215][20]/P0001  & n13901 ;
  assign n16890 = \wishbone_bd_ram_mem2_reg[4][20]/P0001  & n13527 ;
  assign n16891 = ~n16889 & ~n16890 ;
  assign n16892 = n16888 & n16891 ;
  assign n16893 = n16885 & n16892 ;
  assign n16894 = \wishbone_bd_ram_mem2_reg[65][20]/P0001  & n13842 ;
  assign n16895 = \wishbone_bd_ram_mem2_reg[165][20]/P0001  & n14028 ;
  assign n16896 = ~n16894 & ~n16895 ;
  assign n16897 = \wishbone_bd_ram_mem2_reg[134][20]/P0001  & n13494 ;
  assign n16898 = \wishbone_bd_ram_mem2_reg[146][20]/P0001  & n13958 ;
  assign n16899 = ~n16897 & ~n16898 ;
  assign n16900 = n16896 & n16899 ;
  assign n16901 = \wishbone_bd_ram_mem2_reg[211][20]/P0001  & n13805 ;
  assign n16902 = \wishbone_bd_ram_mem2_reg[235][20]/P0001  & n13518 ;
  assign n16903 = ~n16901 & ~n16902 ;
  assign n16904 = \wishbone_bd_ram_mem2_reg[119][20]/P0001  & n14033 ;
  assign n16905 = \wishbone_bd_ram_mem2_reg[10][20]/P0001  & n13837 ;
  assign n16906 = ~n16904 & ~n16905 ;
  assign n16907 = n16903 & n16906 ;
  assign n16908 = n16900 & n16907 ;
  assign n16909 = n16893 & n16908 ;
  assign n16910 = n16878 & n16909 ;
  assign n16911 = \wishbone_bd_ram_mem2_reg[40][20]/P0001  & n13661 ;
  assign n16912 = \wishbone_bd_ram_mem2_reg[229][20]/P0001  & n13552 ;
  assign n16913 = ~n16911 & ~n16912 ;
  assign n16914 = \wishbone_bd_ram_mem2_reg[73][20]/P0001  & n13456 ;
  assign n16915 = \wishbone_bd_ram_mem2_reg[236][20]/P0001  & n13480 ;
  assign n16916 = ~n16914 & ~n16915 ;
  assign n16917 = n16913 & n16916 ;
  assign n16918 = \wishbone_bd_ram_mem2_reg[157][20]/P0001  & n13445 ;
  assign n16919 = \wishbone_bd_ram_mem2_reg[90][20]/P0001  & n13906 ;
  assign n16920 = ~n16918 & ~n16919 ;
  assign n16921 = \wishbone_bd_ram_mem2_reg[45][20]/P0001  & n13420 ;
  assign n16922 = \wishbone_bd_ram_mem2_reg[125][20]/P0001  & n13396 ;
  assign n16923 = ~n16921 & ~n16922 ;
  assign n16924 = n16920 & n16923 ;
  assign n16925 = n16917 & n16924 ;
  assign n16926 = \wishbone_bd_ram_mem2_reg[244][20]/P0001  & n13474 ;
  assign n16927 = \wishbone_bd_ram_mem2_reg[193][20]/P0001  & n14022 ;
  assign n16928 = ~n16926 & ~n16927 ;
  assign n16929 = \wishbone_bd_ram_mem2_reg[172][20]/P0001  & n13377 ;
  assign n16930 = \wishbone_bd_ram_mem2_reg[116][20]/P0001  & n13865 ;
  assign n16931 = ~n16929 & ~n16930 ;
  assign n16932 = n16928 & n16931 ;
  assign n16933 = \wishbone_bd_ram_mem2_reg[222][20]/P0001  & n13721 ;
  assign n16934 = \wishbone_bd_ram_mem2_reg[137][20]/P0001  & n13808 ;
  assign n16935 = ~n16933 & ~n16934 ;
  assign n16936 = \wishbone_bd_ram_mem2_reg[126][20]/P0001  & n13786 ;
  assign n16937 = \wishbone_bd_ram_mem2_reg[109][20]/P0001  & n13306 ;
  assign n16938 = ~n16936 & ~n16937 ;
  assign n16939 = n16935 & n16938 ;
  assign n16940 = n16932 & n16939 ;
  assign n16941 = n16925 & n16940 ;
  assign n16942 = \wishbone_bd_ram_mem2_reg[158][20]/P0001  & n13294 ;
  assign n16943 = \wishbone_bd_ram_mem2_reg[8][20]/P0001  & n13459 ;
  assign n16944 = ~n16942 & ~n16943 ;
  assign n16945 = \wishbone_bd_ram_mem2_reg[89][20]/P0001  & n13910 ;
  assign n16946 = \wishbone_bd_ram_mem2_reg[204][20]/P0001  & n13821 ;
  assign n16947 = ~n16945 & ~n16946 ;
  assign n16948 = n16944 & n16947 ;
  assign n16949 = \wishbone_bd_ram_mem2_reg[41][20]/P0001  & n14017 ;
  assign n16950 = \wishbone_bd_ram_mem2_reg[33][20]/P0001  & n13933 ;
  assign n16951 = ~n16949 & ~n16950 ;
  assign n16952 = \wishbone_bd_ram_mem2_reg[30][20]/P0001  & n13713 ;
  assign n16953 = \wishbone_bd_ram_mem2_reg[5][20]/P0001  & n13243 ;
  assign n16954 = ~n16952 & ~n16953 ;
  assign n16955 = n16951 & n16954 ;
  assign n16956 = n16948 & n16955 ;
  assign n16957 = \wishbone_bd_ram_mem2_reg[219][20]/P0001  & n13577 ;
  assign n16958 = \wishbone_bd_ram_mem2_reg[189][20]/P0001  & n14001 ;
  assign n16959 = ~n16957 & ~n16958 ;
  assign n16960 = \wishbone_bd_ram_mem2_reg[217][20]/P0001  & n13767 ;
  assign n16961 = \wishbone_bd_ram_mem2_reg[26][20]/P0001  & n13521 ;
  assign n16962 = ~n16960 & ~n16961 ;
  assign n16963 = n16959 & n16962 ;
  assign n16964 = \wishbone_bd_ram_mem2_reg[82][20]/P0001  & n13374 ;
  assign n16965 = \wishbone_bd_ram_mem2_reg[202][20]/P0001  & n13268 ;
  assign n16966 = ~n16964 & ~n16965 ;
  assign n16967 = \wishbone_bd_ram_mem2_reg[18][20]/P0001  & n13532 ;
  assign n16968 = \wishbone_bd_ram_mem2_reg[108][20]/P0001  & n13814 ;
  assign n16969 = ~n16967 & ~n16968 ;
  assign n16970 = n16966 & n16969 ;
  assign n16971 = n16963 & n16970 ;
  assign n16972 = n16956 & n16971 ;
  assign n16973 = n16941 & n16972 ;
  assign n16974 = n16910 & n16973 ;
  assign n16975 = \wishbone_bd_ram_mem2_reg[120][20]/P0001  & n13550 ;
  assign n16976 = \wishbone_bd_ram_mem2_reg[239][20]/P0001  & n13349 ;
  assign n16977 = ~n16975 & ~n16976 ;
  assign n16978 = \wishbone_bd_ram_mem2_reg[16][20]/P0001  & n13695 ;
  assign n16979 = \wishbone_bd_ram_mem2_reg[79][20]/P0001  & n13779 ;
  assign n16980 = ~n16978 & ~n16979 ;
  assign n16981 = n16977 & n16980 ;
  assign n16982 = \wishbone_bd_ram_mem2_reg[56][20]/P0001  & n13611 ;
  assign n16983 = \wishbone_bd_ram_mem2_reg[100][20]/P0001  & n13401 ;
  assign n16984 = ~n16982 & ~n16983 ;
  assign n16985 = \wishbone_bd_ram_mem2_reg[127][20]/P0001  & n13803 ;
  assign n16986 = \wishbone_bd_ram_mem2_reg[144][20]/P0001  & n13508 ;
  assign n16987 = ~n16985 & ~n16986 ;
  assign n16988 = n16984 & n16987 ;
  assign n16989 = n16981 & n16988 ;
  assign n16990 = \wishbone_bd_ram_mem2_reg[206][20]/P0001  & n13414 ;
  assign n16991 = \wishbone_bd_ram_mem2_reg[169][20]/P0001  & n13541 ;
  assign n16992 = ~n16990 & ~n16991 ;
  assign n16993 = \wishbone_bd_ram_mem2_reg[250][20]/P0001  & n13677 ;
  assign n16994 = \wishbone_bd_ram_mem2_reg[38][20]/P0001  & n13828 ;
  assign n16995 = ~n16993 & ~n16994 ;
  assign n16996 = n16992 & n16995 ;
  assign n16997 = \wishbone_bd_ram_mem2_reg[76][20]/P0001  & n13831 ;
  assign n16998 = \wishbone_bd_ram_mem2_reg[39][20]/P0001  & n13893 ;
  assign n16999 = ~n16997 & ~n16998 ;
  assign n17000 = \wishbone_bd_ram_mem2_reg[145][20]/P0001  & n13715 ;
  assign n17001 = \wishbone_bd_ram_mem2_reg[111][20]/P0001  & n13471 ;
  assign n17002 = ~n17000 & ~n17001 ;
  assign n17003 = n16999 & n17002 ;
  assign n17004 = n16996 & n17003 ;
  assign n17005 = n16989 & n17004 ;
  assign n17006 = \wishbone_bd_ram_mem2_reg[203][20]/P0001  & n13816 ;
  assign n17007 = \wishbone_bd_ram_mem2_reg[118][20]/P0001  & n13589 ;
  assign n17008 = ~n17006 & ~n17007 ;
  assign n17009 = \wishbone_bd_ram_mem2_reg[231][20]/P0001  & n13363 ;
  assign n17010 = \wishbone_bd_ram_mem2_reg[15][20]/P0001  & n13797 ;
  assign n17011 = ~n17009 & ~n17010 ;
  assign n17012 = n17008 & n17011 ;
  assign n17013 = \wishbone_bd_ram_mem2_reg[177][20]/P0001  & n13863 ;
  assign n17014 = \wishbone_bd_ram_mem2_reg[166][20]/P0001  & n13999 ;
  assign n17015 = ~n17013 & ~n17014 ;
  assign n17016 = \wishbone_bd_ram_mem2_reg[149][20]/P0001  & n13469 ;
  assign n17017 = \wishbone_bd_ram_mem2_reg[121][20]/P0001  & n13983 ;
  assign n17018 = ~n17016 & ~n17017 ;
  assign n17019 = n17015 & n17018 ;
  assign n17020 = n17012 & n17019 ;
  assign n17021 = \wishbone_bd_ram_mem2_reg[37][20]/P0001  & n13710 ;
  assign n17022 = \wishbone_bd_ram_mem2_reg[234][20]/P0001  & n13781 ;
  assign n17023 = ~n17021 & ~n17022 ;
  assign n17024 = \wishbone_bd_ram_mem2_reg[20][20]/P0001  & n13839 ;
  assign n17025 = \wishbone_bd_ram_mem2_reg[147][20]/P0001  & n13702 ;
  assign n17026 = ~n17024 & ~n17025 ;
  assign n17027 = n17023 & n17026 ;
  assign n17028 = \wishbone_bd_ram_mem2_reg[64][20]/P0001  & n13904 ;
  assign n17029 = \wishbone_bd_ram_mem2_reg[225][20]/P0001  & n13719 ;
  assign n17030 = ~n17028 & ~n17029 ;
  assign n17031 = \wishbone_bd_ram_mem2_reg[85][20]/P0001  & n13784 ;
  assign n17032 = \wishbone_bd_ram_mem2_reg[237][20]/P0001  & n13924 ;
  assign n17033 = ~n17031 & ~n17032 ;
  assign n17034 = n17030 & n17033 ;
  assign n17035 = n17027 & n17034 ;
  assign n17036 = n17020 & n17035 ;
  assign n17037 = n17005 & n17036 ;
  assign n17038 = \wishbone_bd_ram_mem2_reg[124][20]/P0001  & n14024 ;
  assign n17039 = \wishbone_bd_ram_mem2_reg[71][20]/P0001  & n13636 ;
  assign n17040 = ~n17038 & ~n17039 ;
  assign n17041 = \wishbone_bd_ram_mem2_reg[223][20]/P0001  & n13335 ;
  assign n17042 = \wishbone_bd_ram_mem2_reg[242][20]/P0001  & n13383 ;
  assign n17043 = ~n17041 & ~n17042 ;
  assign n17044 = n17040 & n17043 ;
  assign n17045 = \wishbone_bd_ram_mem2_reg[114][20]/P0001  & n13763 ;
  assign n17046 = \wishbone_bd_ram_mem2_reg[168][20]/P0001  & n13795 ;
  assign n17047 = ~n17045 & ~n17046 ;
  assign n17048 = \wishbone_bd_ram_mem2_reg[96][20]/P0001  & n13425 ;
  assign n17049 = \wishbone_bd_ram_mem2_reg[247][20]/P0001  & n13571 ;
  assign n17050 = ~n17048 & ~n17049 ;
  assign n17051 = n17047 & n17050 ;
  assign n17052 = n17044 & n17051 ;
  assign n17053 = \wishbone_bd_ram_mem2_reg[198][20]/P0001  & n13592 ;
  assign n17054 = \wishbone_bd_ram_mem2_reg[128][20]/P0001  & n13652 ;
  assign n17055 = ~n17053 & ~n17054 ;
  assign n17056 = \wishbone_bd_ram_mem2_reg[112][20]/P0001  & n13482 ;
  assign n17057 = \wishbone_bd_ram_mem2_reg[44][20]/P0001  & n13291 ;
  assign n17058 = ~n17056 & ~n17057 ;
  assign n17059 = n17055 & n17058 ;
  assign n17060 = \wishbone_bd_ram_mem2_reg[160][20]/P0001  & n13271 ;
  assign n17061 = \wishbone_bd_ram_mem2_reg[92][20]/P0001  & n13859 ;
  assign n17062 = ~n17060 & ~n17061 ;
  assign n17063 = \wishbone_bd_ram_mem2_reg[210][20]/P0001  & n13443 ;
  assign n17064 = \wishbone_bd_ram_mem2_reg[254][20]/P0001  & n13283 ;
  assign n17065 = ~n17063 & ~n17064 ;
  assign n17066 = n17062 & n17065 ;
  assign n17067 = n17059 & n17066 ;
  assign n17068 = n17052 & n17067 ;
  assign n17069 = \wishbone_bd_ram_mem2_reg[57][20]/P0001  & n13731 ;
  assign n17070 = \wishbone_bd_ram_mem2_reg[101][20]/P0001  & n13772 ;
  assign n17071 = ~n17069 & ~n17070 ;
  assign n17072 = \wishbone_bd_ram_mem2_reg[70][20]/P0001  & n13339 ;
  assign n17073 = \wishbone_bd_ram_mem2_reg[150][20]/P0001  & n13666 ;
  assign n17074 = ~n17072 & ~n17073 ;
  assign n17075 = n17071 & n17074 ;
  assign n17076 = \wishbone_bd_ram_mem2_reg[115][20]/P0001  & n13747 ;
  assign n17077 = \wishbone_bd_ram_mem2_reg[154][20]/P0001  & n13403 ;
  assign n17078 = ~n17076 & ~n17077 ;
  assign n17079 = \wishbone_bd_ram_mem2_reg[105][20]/P0001  & n13503 ;
  assign n17080 = \wishbone_bd_ram_mem2_reg[152][20]/P0001  & n13912 ;
  assign n17081 = ~n17079 & ~n17080 ;
  assign n17082 = n17078 & n17081 ;
  assign n17083 = n17075 & n17082 ;
  assign n17084 = \wishbone_bd_ram_mem2_reg[21][20]/P0001  & n13438 ;
  assign n17085 = \wishbone_bd_ram_mem2_reg[201][20]/P0001  & n13600 ;
  assign n17086 = ~n17084 & ~n17085 ;
  assign n17087 = \wishbone_bd_ram_mem2_reg[190][20]/P0001  & n13365 ;
  assign n17088 = \wishbone_bd_ram_mem2_reg[22][20]/P0001  & n13744 ;
  assign n17089 = ~n17087 & ~n17088 ;
  assign n17090 = n17086 & n17089 ;
  assign n17091 = \wishbone_bd_ram_mem2_reg[173][20]/P0001  & n13360 ;
  assign n17092 = \wishbone_bd_ram_mem2_reg[142][20]/P0001  & n13448 ;
  assign n17093 = ~n17091 & ~n17092 ;
  assign n17094 = \wishbone_bd_ram_mem2_reg[106][20]/P0001  & n13555 ;
  assign n17095 = \wishbone_bd_ram_mem2_reg[148][20]/P0001  & n13868 ;
  assign n17096 = ~n17094 & ~n17095 ;
  assign n17097 = n17093 & n17096 ;
  assign n17098 = n17090 & n17097 ;
  assign n17099 = n17083 & n17098 ;
  assign n17100 = n17068 & n17099 ;
  assign n17101 = n17037 & n17100 ;
  assign n17102 = n16974 & n17101 ;
  assign n17103 = \wishbone_bd_ram_mem2_reg[84][20]/P0001  & n13385 ;
  assign n17104 = \wishbone_bd_ram_mem2_reg[102][20]/P0001  & n13534 ;
  assign n17105 = ~n17103 & ~n17104 ;
  assign n17106 = \wishbone_bd_ram_mem2_reg[139][20]/P0001  & n13566 ;
  assign n17107 = \wishbone_bd_ram_mem2_reg[66][20]/P0001  & n13603 ;
  assign n17108 = ~n17106 & ~n17107 ;
  assign n17109 = n17105 & n17108 ;
  assign n17110 = \wishbone_bd_ram_mem2_reg[185][20]/P0001  & n13372 ;
  assign n17111 = \wishbone_bd_ram_mem2_reg[1][20]/P0001  & n13888 ;
  assign n17112 = ~n17110 & ~n17111 ;
  assign n17113 = \wishbone_bd_ram_mem2_reg[23][20]/P0001  & n13857 ;
  assign n17114 = \wishbone_bd_ram_mem2_reg[129][20]/P0001  & n13629 ;
  assign n17115 = ~n17113 & ~n17114 ;
  assign n17116 = n17112 & n17115 ;
  assign n17117 = n17109 & n17116 ;
  assign n17118 = \wishbone_bd_ram_mem2_reg[69][20]/P0001  & n13487 ;
  assign n17119 = \wishbone_bd_ram_mem2_reg[197][20]/P0001  & n13594 ;
  assign n17120 = ~n17118 & ~n17119 ;
  assign n17121 = \wishbone_bd_ram_mem2_reg[72][20]/P0001  & n13582 ;
  assign n17122 = \wishbone_bd_ram_mem2_reg[94][20]/P0001  & n13833 ;
  assign n17123 = ~n17121 & ~n17122 ;
  assign n17124 = n17120 & n17123 ;
  assign n17125 = \wishbone_bd_ram_mem2_reg[205][20]/P0001  & n13947 ;
  assign n17126 = \wishbone_bd_ram_mem2_reg[130][20]/P0001  & n13427 ;
  assign n17127 = ~n17125 & ~n17126 ;
  assign n17128 = \wishbone_bd_ram_mem2_reg[163][20]/P0001  & n13255 ;
  assign n17129 = \wishbone_bd_ram_mem2_reg[253][20]/P0001  & n13708 ;
  assign n17130 = ~n17128 & ~n17129 ;
  assign n17131 = n17127 & n17130 ;
  assign n17132 = n17124 & n17131 ;
  assign n17133 = n17117 & n17132 ;
  assign n17134 = \wishbone_bd_ram_mem2_reg[240][20]/P0001  & n13352 ;
  assign n17135 = \wishbone_bd_ram_mem2_reg[243][20]/P0001  & n13575 ;
  assign n17136 = ~n17134 & ~n17135 ;
  assign n17137 = \wishbone_bd_ram_mem2_reg[24][20]/P0001  & n13970 ;
  assign n17138 = \wishbone_bd_ram_mem2_reg[103][20]/P0001  & n13320 ;
  assign n17139 = ~n17137 & ~n17138 ;
  assign n17140 = n17136 & n17139 ;
  assign n17141 = \wishbone_bd_ram_mem2_reg[184][20]/P0001  & n13960 ;
  assign n17142 = \wishbone_bd_ram_mem2_reg[110][20]/P0001  & n14030 ;
  assign n17143 = ~n17141 & ~n17142 ;
  assign n17144 = \wishbone_bd_ram_mem2_reg[28][20]/P0001  & n13810 ;
  assign n17145 = \wishbone_bd_ram_mem2_reg[91][20]/P0001  & n13954 ;
  assign n17146 = ~n17144 & ~n17145 ;
  assign n17147 = n17143 & n17146 ;
  assign n17148 = n17140 & n17147 ;
  assign n17149 = \wishbone_bd_ram_mem2_reg[27][20]/P0001  & n13251 ;
  assign n17150 = \wishbone_bd_ram_mem2_reg[170][20]/P0001  & n14007 ;
  assign n17151 = ~n17149 & ~n17150 ;
  assign n17152 = \wishbone_bd_ram_mem2_reg[195][20]/P0001  & n13700 ;
  assign n17153 = \wishbone_bd_ram_mem2_reg[233][20]/P0001  & n13332 ;
  assign n17154 = ~n17152 & ~n17153 ;
  assign n17155 = n17151 & n17154 ;
  assign n17156 = \wishbone_bd_ram_mem2_reg[7][20]/P0001  & n13546 ;
  assign n17157 = \wishbone_bd_ram_mem2_reg[97][20]/P0001  & n13724 ;
  assign n17158 = ~n17156 & ~n17157 ;
  assign n17159 = \wishbone_bd_ram_mem2_reg[31][20]/P0001  & n13758 ;
  assign n17160 = \wishbone_bd_ram_mem2_reg[54][20]/P0001  & n13622 ;
  assign n17161 = ~n17159 & ~n17160 ;
  assign n17162 = n17158 & n17161 ;
  assign n17163 = n17155 & n17162 ;
  assign n17164 = n17148 & n17163 ;
  assign n17165 = n17133 & n17164 ;
  assign n17166 = \wishbone_bd_ram_mem2_reg[46][20]/P0001  & n13298 ;
  assign n17167 = \wishbone_bd_ram_mem2_reg[207][20]/P0001  & n13826 ;
  assign n17168 = ~n17166 & ~n17167 ;
  assign n17169 = \wishbone_bd_ram_mem2_reg[212][20]/P0001  & n13634 ;
  assign n17170 = \wishbone_bd_ram_mem2_reg[62][20]/P0001  & n13529 ;
  assign n17171 = ~n17169 & ~n17170 ;
  assign n17172 = n17168 & n17171 ;
  assign n17173 = \wishbone_bd_ram_mem2_reg[75][20]/P0001  & n13605 ;
  assign n17174 = \wishbone_bd_ram_mem2_reg[161][20]/P0001  & n13505 ;
  assign n17175 = ~n17173 & ~n17174 ;
  assign n17176 = \wishbone_bd_ram_mem2_reg[36][20]/P0001  & n13639 ;
  assign n17177 = \wishbone_bd_ram_mem2_reg[51][20]/P0001  & n13880 ;
  assign n17178 = ~n17176 & ~n17177 ;
  assign n17179 = n17175 & n17178 ;
  assign n17180 = n17172 & n17179 ;
  assign n17181 = \wishbone_bd_ram_mem2_reg[80][20]/P0001  & n13516 ;
  assign n17182 = \wishbone_bd_ram_mem2_reg[14][20]/P0001  & n13972 ;
  assign n17183 = ~n17181 & ~n17182 ;
  assign n17184 = \wishbone_bd_ram_mem2_reg[200][20]/P0001  & n13922 ;
  assign n17185 = \wishbone_bd_ram_mem2_reg[141][20]/P0001  & n13852 ;
  assign n17186 = ~n17184 & ~n17185 ;
  assign n17187 = n17183 & n17186 ;
  assign n17188 = \wishbone_bd_ram_mem2_reg[88][20]/P0001  & n13347 ;
  assign n17189 = \wishbone_bd_ram_mem2_reg[196][20]/P0001  & n13977 ;
  assign n17190 = ~n17188 & ~n17189 ;
  assign n17191 = \wishbone_bd_ram_mem2_reg[238][20]/P0001  & n13819 ;
  assign n17192 = \wishbone_bd_ram_mem2_reg[181][20]/P0001  & n13587 ;
  assign n17193 = ~n17191 & ~n17192 ;
  assign n17194 = n17190 & n17193 ;
  assign n17195 = n17187 & n17194 ;
  assign n17196 = n17180 & n17195 ;
  assign n17197 = \wishbone_bd_ram_mem2_reg[179][20]/P0001  & n14035 ;
  assign n17198 = \wishbone_bd_ram_mem2_reg[49][20]/P0001  & n13929 ;
  assign n17199 = ~n17197 & ~n17198 ;
  assign n17200 = \wishbone_bd_ram_mem2_reg[117][20]/P0001  & n13557 ;
  assign n17201 = \wishbone_bd_ram_mem2_reg[162][20]/P0001  & n13726 ;
  assign n17202 = ~n17200 & ~n17201 ;
  assign n17203 = n17199 & n17202 ;
  assign n17204 = \wishbone_bd_ram_mem2_reg[60][20]/P0001  & n13790 ;
  assign n17205 = \wishbone_bd_ram_mem2_reg[255][20]/P0001  & n13952 ;
  assign n17206 = ~n17204 & ~n17205 ;
  assign n17207 = \wishbone_bd_ram_mem2_reg[249][20]/P0001  & n13431 ;
  assign n17208 = \wishbone_bd_ram_mem2_reg[42][20]/P0001  & n13341 ;
  assign n17209 = ~n17207 & ~n17208 ;
  assign n17210 = n17206 & n17209 ;
  assign n17211 = n17203 & n17210 ;
  assign n17212 = \wishbone_bd_ram_mem2_reg[214][20]/P0001  & n13938 ;
  assign n17213 = \wishbone_bd_ram_mem2_reg[107][20]/P0001  & n13476 ;
  assign n17214 = ~n17212 & ~n17213 ;
  assign n17215 = \wishbone_bd_ram_mem2_reg[188][20]/P0001  & n13407 ;
  assign n17216 = \wishbone_bd_ram_mem2_reg[25][20]/P0001  & n13742 ;
  assign n17217 = ~n17215 & ~n17216 ;
  assign n17218 = n17214 & n17217 ;
  assign n17219 = \wishbone_bd_ram_mem2_reg[186][20]/P0001  & n13616 ;
  assign n17220 = \wishbone_bd_ram_mem2_reg[47][20]/P0001  & n13436 ;
  assign n17221 = ~n17219 & ~n17220 ;
  assign n17222 = \wishbone_bd_ram_mem2_reg[151][20]/P0001  & n13697 ;
  assign n17223 = \wishbone_bd_ram_mem2_reg[95][20]/P0001  & n13317 ;
  assign n17224 = ~n17222 & ~n17223 ;
  assign n17225 = n17221 & n17224 ;
  assign n17226 = n17218 & n17225 ;
  assign n17227 = n17211 & n17226 ;
  assign n17228 = n17196 & n17227 ;
  assign n17229 = n17165 & n17228 ;
  assign n17230 = \wishbone_bd_ram_mem2_reg[209][20]/P0001  & n13689 ;
  assign n17231 = \wishbone_bd_ram_mem2_reg[228][20]/P0001  & n13497 ;
  assign n17232 = ~n17230 & ~n17231 ;
  assign n17233 = \wishbone_bd_ram_mem2_reg[246][20]/P0001  & n13981 ;
  assign n17234 = \wishbone_bd_ram_mem2_reg[81][20]/P0001  & n13409 ;
  assign n17235 = ~n17233 & ~n17234 ;
  assign n17236 = n17232 & n17235 ;
  assign n17237 = \wishbone_bd_ram_mem2_reg[68][20]/P0001  & n13379 ;
  assign n17238 = \wishbone_bd_ram_mem2_reg[248][20]/P0001  & n13647 ;
  assign n17239 = ~n17237 & ~n17238 ;
  assign n17240 = \wishbone_bd_ram_mem2_reg[230][20]/P0001  & n13994 ;
  assign n17241 = \wishbone_bd_ram_mem2_reg[35][20]/P0001  & n13523 ;
  assign n17242 = ~n17240 & ~n17241 ;
  assign n17243 = n17239 & n17242 ;
  assign n17244 = n17236 & n17243 ;
  assign n17245 = \wishbone_bd_ram_mem2_reg[176][20]/P0001  & n13262 ;
  assign n17246 = \wishbone_bd_ram_mem2_reg[59][20]/P0001  & n13613 ;
  assign n17247 = ~n17245 & ~n17246 ;
  assign n17248 = \wishbone_bd_ram_mem2_reg[226][20]/P0001  & n13668 ;
  assign n17249 = \wishbone_bd_ram_mem2_reg[143][20]/P0001  & n13461 ;
  assign n17250 = ~n17248 & ~n17249 ;
  assign n17251 = n17247 & n17250 ;
  assign n17252 = \wishbone_bd_ram_mem2_reg[216][20]/P0001  & n14005 ;
  assign n17253 = \wishbone_bd_ram_mem2_reg[2][20]/P0001  & n13975 ;
  assign n17254 = ~n17252 & ~n17253 ;
  assign n17255 = \wishbone_bd_ram_mem2_reg[178][20]/P0001  & n13301 ;
  assign n17256 = \wishbone_bd_ram_mem2_reg[12][20]/P0001  & n13733 ;
  assign n17257 = ~n17255 & ~n17256 ;
  assign n17258 = n17254 & n17257 ;
  assign n17259 = n17251 & n17258 ;
  assign n17260 = n17244 & n17259 ;
  assign n17261 = \wishbone_bd_ram_mem2_reg[61][20]/P0001  & n13544 ;
  assign n17262 = \wishbone_bd_ram_mem2_reg[6][20]/P0001  & n13915 ;
  assign n17263 = ~n17261 & ~n17262 ;
  assign n17264 = \wishbone_bd_ram_mem2_reg[191][20]/P0001  & n14012 ;
  assign n17265 = \wishbone_bd_ram_mem2_reg[17][20]/P0001  & n13324 ;
  assign n17266 = ~n17264 & ~n17265 ;
  assign n17267 = n17263 & n17266 ;
  assign n17268 = \wishbone_bd_ram_mem2_reg[192][20]/P0001  & n13390 ;
  assign n17269 = \wishbone_bd_ram_mem2_reg[232][20]/P0001  & n13510 ;
  assign n17270 = ~n17268 & ~n17269 ;
  assign n17271 = \wishbone_bd_ram_mem2_reg[11][20]/P0001  & n13774 ;
  assign n17272 = \wishbone_bd_ram_mem2_reg[213][20]/P0001  & n13870 ;
  assign n17273 = ~n17271 & ~n17272 ;
  assign n17274 = n17270 & n17273 ;
  assign n17275 = n17267 & n17274 ;
  assign n17276 = \wishbone_bd_ram_mem2_reg[224][20]/P0001  & n13433 ;
  assign n17277 = \wishbone_bd_ram_mem2_reg[138][20]/P0001  & n13398 ;
  assign n17278 = ~n17276 & ~n17277 ;
  assign n17279 = \wishbone_bd_ram_mem2_reg[221][20]/P0001  & n13641 ;
  assign n17280 = \wishbone_bd_ram_mem2_reg[174][20]/P0001  & n13899 ;
  assign n17281 = ~n17279 & ~n17280 ;
  assign n17282 = n17278 & n17281 ;
  assign n17283 = \wishbone_bd_ram_mem2_reg[199][20]/P0001  & n13499 ;
  assign n17284 = \wishbone_bd_ram_mem2_reg[78][20]/P0001  & n13277 ;
  assign n17285 = ~n17283 & ~n17284 ;
  assign n17286 = \wishbone_bd_ram_mem2_reg[251][20]/P0001  & n14019 ;
  assign n17287 = \wishbone_bd_ram_mem2_reg[48][20]/P0001  & n13917 ;
  assign n17288 = ~n17286 & ~n17287 ;
  assign n17289 = n17285 & n17288 ;
  assign n17290 = n17282 & n17289 ;
  assign n17291 = n17275 & n17290 ;
  assign n17292 = n17260 & n17291 ;
  assign n17293 = \wishbone_bd_ram_mem2_reg[52][20]/P0001  & n13988 ;
  assign n17294 = \wishbone_bd_ram_mem2_reg[175][20]/P0001  & n13674 ;
  assign n17295 = ~n17293 & ~n17294 ;
  assign n17296 = \wishbone_bd_ram_mem2_reg[156][20]/P0001  & n13769 ;
  assign n17297 = \wishbone_bd_ram_mem2_reg[241][20]/P0001  & n13854 ;
  assign n17298 = ~n17296 & ~n17297 ;
  assign n17299 = n17295 & n17298 ;
  assign n17300 = \wishbone_bd_ram_mem2_reg[58][20]/P0001  & n13949 ;
  assign n17301 = \wishbone_bd_ram_mem2_reg[208][20]/P0001  & n14010 ;
  assign n17302 = ~n17300 & ~n17301 ;
  assign n17303 = \wishbone_bd_ram_mem2_reg[187][20]/P0001  & n13756 ;
  assign n17304 = \wishbone_bd_ram_mem2_reg[13][20]/P0001  & n13844 ;
  assign n17305 = ~n17303 & ~n17304 ;
  assign n17306 = n17302 & n17305 ;
  assign n17307 = n17299 & n17306 ;
  assign n17308 = \wishbone_bd_ram_mem2_reg[183][20]/P0001  & n13645 ;
  assign n17309 = \wishbone_bd_ram_mem2_reg[55][20]/P0001  & n13618 ;
  assign n17310 = ~n17308 & ~n17309 ;
  assign n17311 = \wishbone_bd_ram_mem2_reg[50][20]/P0001  & n13686 ;
  assign n17312 = \wishbone_bd_ram_mem2_reg[155][20]/P0001  & n13738 ;
  assign n17313 = ~n17311 & ~n17312 ;
  assign n17314 = n17310 & n17313 ;
  assign n17315 = \wishbone_bd_ram_mem2_reg[159][20]/P0001  & n13627 ;
  assign n17316 = \wishbone_bd_ram_mem2_reg[220][20]/P0001  & n13965 ;
  assign n17317 = ~n17315 & ~n17316 ;
  assign n17318 = \wishbone_bd_ram_mem2_reg[218][20]/P0001  & n13792 ;
  assign n17319 = \wishbone_bd_ram_mem2_reg[104][20]/P0001  & n13684 ;
  assign n17320 = ~n17318 & ~n17319 ;
  assign n17321 = n17317 & n17320 ;
  assign n17322 = n17314 & n17321 ;
  assign n17323 = n17307 & n17322 ;
  assign n17324 = \wishbone_bd_ram_mem2_reg[98][20]/P0001  & n13569 ;
  assign n17325 = \wishbone_bd_ram_mem2_reg[123][20]/P0001  & n13749 ;
  assign n17326 = ~n17324 & ~n17325 ;
  assign n17327 = \wishbone_bd_ram_mem2_reg[171][20]/P0001  & n13422 ;
  assign n17328 = \wishbone_bd_ram_mem2_reg[131][20]/P0001  & n13358 ;
  assign n17329 = ~n17327 & ~n17328 ;
  assign n17330 = n17326 & n17329 ;
  assign n17331 = \wishbone_bd_ram_mem2_reg[93][20]/P0001  & n13891 ;
  assign n17332 = \wishbone_bd_ram_mem2_reg[86][20]/P0001  & n13485 ;
  assign n17333 = ~n17331 & ~n17332 ;
  assign n17334 = \wishbone_bd_ram_mem2_reg[63][20]/P0001  & n13327 ;
  assign n17335 = \wishbone_bd_ram_mem2_reg[77][20]/P0001  & n13935 ;
  assign n17336 = ~n17334 & ~n17335 ;
  assign n17337 = n17333 & n17336 ;
  assign n17338 = n17330 & n17337 ;
  assign n17339 = \wishbone_bd_ram_mem2_reg[227][20]/P0001  & n13388 ;
  assign n17340 = \wishbone_bd_ram_mem2_reg[122][20]/P0001  & n13679 ;
  assign n17341 = ~n17339 & ~n17340 ;
  assign n17342 = \wishbone_bd_ram_mem2_reg[167][20]/P0001  & n13940 ;
  assign n17343 = \wishbone_bd_ram_mem2_reg[132][20]/P0001  & n13927 ;
  assign n17344 = ~n17342 & ~n17343 ;
  assign n17345 = n17341 & n17344 ;
  assign n17346 = \wishbone_bd_ram_mem2_reg[74][20]/P0001  & n13564 ;
  assign n17347 = \wishbone_bd_ram_mem2_reg[136][20]/P0001  & n13963 ;
  assign n17348 = ~n17346 & ~n17347 ;
  assign n17349 = \wishbone_bd_ram_mem2_reg[182][20]/P0001  & n13598 ;
  assign n17350 = \wishbone_bd_ram_mem2_reg[153][20]/P0001  & n13309 ;
  assign n17351 = ~n17349 & ~n17350 ;
  assign n17352 = n17348 & n17351 ;
  assign n17353 = n17345 & n17352 ;
  assign n17354 = n17338 & n17353 ;
  assign n17355 = n17323 & n17354 ;
  assign n17356 = n17292 & n17355 ;
  assign n17357 = n17229 & n17356 ;
  assign n17358 = n17102 & n17357 ;
  assign n17359 = n14047 & ~n17358 ;
  assign n17360 = n14049 & ~n14064 ;
  assign n17361 = \wishbone_TxLength_reg[4]/NET0131  & ~n14049 ;
  assign n17362 = ~n17360 & ~n17361 ;
  assign n17363 = \wishbone_TxLength_reg[4]/NET0131  & ~n14054 ;
  assign n17364 = ~n14055 & ~n17363 ;
  assign n17365 = \wishbone_TxLength_reg[0]/NET0131  & \wishbone_TxLength_reg[1]/NET0131  ;
  assign n17366 = n17364 & ~n17365 ;
  assign n17367 = \wishbone_TxPointerLSB_rst_reg[0]/NET0131  & ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n17368 = ~\wishbone_TxLength_reg[4]/NET0131  & n17365 ;
  assign n17369 = n17367 & ~n17368 ;
  assign n17370 = ~n17366 & n17369 ;
  assign n17371 = \wishbone_TxPointerLSB_rst_reg[0]/NET0131  & \wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n17372 = ~\wishbone_TxLength_reg[0]/NET0131  & ~\wishbone_TxLength_reg[1]/NET0131  ;
  assign n17373 = n14054 & n17372 ;
  assign n17374 = \wishbone_TxLength_reg[4]/NET0131  & ~n17373 ;
  assign n17375 = n14055 & n17372 ;
  assign n17376 = ~n17374 & ~n17375 ;
  assign n17377 = n17371 & ~n17376 ;
  assign n17378 = ~n17370 & ~n17377 ;
  assign n17379 = ~\wishbone_TxPointerLSB_rst_reg[0]/NET0131  & ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n17380 = ~n17364 & n17379 ;
  assign n17381 = ~\wishbone_TxPointerLSB_rst_reg[0]/NET0131  & \wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n17382 = ~\wishbone_TxLength_reg[1]/NET0131  & ~\wishbone_TxLength_reg[4]/NET0131  ;
  assign n17383 = n14054 & n17382 ;
  assign n17384 = n17381 & n17383 ;
  assign n17385 = ~\wishbone_TxLength_reg[1]/NET0131  & n14054 ;
  assign n17386 = \wishbone_TxLength_reg[4]/NET0131  & n17381 ;
  assign n17387 = ~n17385 & n17386 ;
  assign n17388 = ~n17384 & ~n17387 ;
  assign n17389 = ~n17380 & n17388 ;
  assign n17390 = ~n17361 & n17389 ;
  assign n17391 = n17378 & n17390 ;
  assign n17392 = ~n17362 & ~n17391 ;
  assign n17393 = ~n14046 & n17392 ;
  assign n17394 = ~n17359 & ~n17393 ;
  assign n17395 = \wishbone_bd_ram_mem3_reg[57][26]/P0001  & n13731 ;
  assign n17396 = \wishbone_bd_ram_mem3_reg[185][26]/P0001  & n13372 ;
  assign n17397 = ~n17395 & ~n17396 ;
  assign n17398 = \wishbone_bd_ram_mem3_reg[189][26]/P0001  & n14001 ;
  assign n17399 = \wishbone_bd_ram_mem3_reg[55][26]/P0001  & n13618 ;
  assign n17400 = ~n17398 & ~n17399 ;
  assign n17401 = n17397 & n17400 ;
  assign n17402 = \wishbone_bd_ram_mem3_reg[36][26]/P0001  & n13639 ;
  assign n17403 = \wishbone_bd_ram_mem3_reg[159][26]/P0001  & n13627 ;
  assign n17404 = ~n17402 & ~n17403 ;
  assign n17405 = \wishbone_bd_ram_mem3_reg[64][26]/P0001  & n13904 ;
  assign n17406 = \wishbone_bd_ram_mem3_reg[204][26]/P0001  & n13821 ;
  assign n17407 = ~n17405 & ~n17406 ;
  assign n17408 = n17404 & n17407 ;
  assign n17409 = n17401 & n17408 ;
  assign n17410 = \wishbone_bd_ram_mem3_reg[201][26]/P0001  & n13600 ;
  assign n17411 = \wishbone_bd_ram_mem3_reg[127][26]/P0001  & n13803 ;
  assign n17412 = ~n17410 & ~n17411 ;
  assign n17413 = \wishbone_bd_ram_mem3_reg[86][26]/P0001  & n13485 ;
  assign n17414 = \wishbone_bd_ram_mem3_reg[111][26]/P0001  & n13471 ;
  assign n17415 = ~n17413 & ~n17414 ;
  assign n17416 = n17412 & n17415 ;
  assign n17417 = \wishbone_bd_ram_mem3_reg[63][26]/P0001  & n13327 ;
  assign n17418 = \wishbone_bd_ram_mem3_reg[207][26]/P0001  & n13826 ;
  assign n17419 = ~n17417 & ~n17418 ;
  assign n17420 = \wishbone_bd_ram_mem3_reg[254][26]/P0001  & n13283 ;
  assign n17421 = \wishbone_bd_ram_mem3_reg[119][26]/P0001  & n14033 ;
  assign n17422 = ~n17420 & ~n17421 ;
  assign n17423 = n17419 & n17422 ;
  assign n17424 = n17416 & n17423 ;
  assign n17425 = n17409 & n17424 ;
  assign n17426 = \wishbone_bd_ram_mem3_reg[90][26]/P0001  & n13906 ;
  assign n17427 = \wishbone_bd_ram_mem3_reg[143][26]/P0001  & n13461 ;
  assign n17428 = ~n17426 & ~n17427 ;
  assign n17429 = \wishbone_bd_ram_mem3_reg[160][26]/P0001  & n13271 ;
  assign n17430 = \wishbone_bd_ram_mem3_reg[75][26]/P0001  & n13605 ;
  assign n17431 = ~n17429 & ~n17430 ;
  assign n17432 = n17428 & n17431 ;
  assign n17433 = \wishbone_bd_ram_mem3_reg[248][26]/P0001  & n13647 ;
  assign n17434 = \wishbone_bd_ram_mem3_reg[209][26]/P0001  & n13689 ;
  assign n17435 = ~n17433 & ~n17434 ;
  assign n17436 = \wishbone_bd_ram_mem3_reg[15][26]/P0001  & n13797 ;
  assign n17437 = \wishbone_bd_ram_mem3_reg[247][26]/P0001  & n13571 ;
  assign n17438 = ~n17436 & ~n17437 ;
  assign n17439 = n17435 & n17438 ;
  assign n17440 = n17432 & n17439 ;
  assign n17441 = \wishbone_bd_ram_mem3_reg[125][26]/P0001  & n13396 ;
  assign n17442 = \wishbone_bd_ram_mem3_reg[217][26]/P0001  & n13767 ;
  assign n17443 = ~n17441 & ~n17442 ;
  assign n17444 = \wishbone_bd_ram_mem3_reg[215][26]/P0001  & n13901 ;
  assign n17445 = \wishbone_bd_ram_mem3_reg[65][26]/P0001  & n13842 ;
  assign n17446 = ~n17444 & ~n17445 ;
  assign n17447 = n17443 & n17446 ;
  assign n17448 = \wishbone_bd_ram_mem3_reg[67][26]/P0001  & n13663 ;
  assign n17449 = \wishbone_bd_ram_mem3_reg[242][26]/P0001  & n13383 ;
  assign n17450 = ~n17448 & ~n17449 ;
  assign n17451 = \wishbone_bd_ram_mem3_reg[120][26]/P0001  & n13550 ;
  assign n17452 = \wishbone_bd_ram_mem3_reg[178][26]/P0001  & n13301 ;
  assign n17453 = ~n17451 & ~n17452 ;
  assign n17454 = n17450 & n17453 ;
  assign n17455 = n17447 & n17454 ;
  assign n17456 = n17440 & n17455 ;
  assign n17457 = n17425 & n17456 ;
  assign n17458 = \wishbone_bd_ram_mem3_reg[212][26]/P0001  & n13634 ;
  assign n17459 = \wishbone_bd_ram_mem3_reg[54][26]/P0001  & n13622 ;
  assign n17460 = ~n17458 & ~n17459 ;
  assign n17461 = \wishbone_bd_ram_mem3_reg[228][26]/P0001  & n13497 ;
  assign n17462 = \wishbone_bd_ram_mem3_reg[18][26]/P0001  & n13532 ;
  assign n17463 = ~n17461 & ~n17462 ;
  assign n17464 = n17460 & n17463 ;
  assign n17465 = \wishbone_bd_ram_mem3_reg[205][26]/P0001  & n13947 ;
  assign n17466 = \wishbone_bd_ram_mem3_reg[26][26]/P0001  & n13521 ;
  assign n17467 = ~n17465 & ~n17466 ;
  assign n17468 = \wishbone_bd_ram_mem3_reg[229][26]/P0001  & n13552 ;
  assign n17469 = \wishbone_bd_ram_mem3_reg[146][26]/P0001  & n13958 ;
  assign n17470 = ~n17468 & ~n17469 ;
  assign n17471 = n17467 & n17470 ;
  assign n17472 = n17464 & n17471 ;
  assign n17473 = \wishbone_bd_ram_mem3_reg[182][26]/P0001  & n13598 ;
  assign n17474 = \wishbone_bd_ram_mem3_reg[188][26]/P0001  & n13407 ;
  assign n17475 = ~n17473 & ~n17474 ;
  assign n17476 = \wishbone_bd_ram_mem3_reg[32][26]/P0001  & n13736 ;
  assign n17477 = \wishbone_bd_ram_mem3_reg[138][26]/P0001  & n13398 ;
  assign n17478 = ~n17476 & ~n17477 ;
  assign n17479 = n17475 & n17478 ;
  assign n17480 = \wishbone_bd_ram_mem3_reg[239][26]/P0001  & n13349 ;
  assign n17481 = \wishbone_bd_ram_mem3_reg[206][26]/P0001  & n13414 ;
  assign n17482 = ~n17480 & ~n17481 ;
  assign n17483 = \wishbone_bd_ram_mem3_reg[56][26]/P0001  & n13611 ;
  assign n17484 = \wishbone_bd_ram_mem3_reg[253][26]/P0001  & n13708 ;
  assign n17485 = ~n17483 & ~n17484 ;
  assign n17486 = n17482 & n17485 ;
  assign n17487 = n17479 & n17486 ;
  assign n17488 = n17472 & n17487 ;
  assign n17489 = \wishbone_bd_ram_mem3_reg[76][26]/P0001  & n13831 ;
  assign n17490 = \wishbone_bd_ram_mem3_reg[157][26]/P0001  & n13445 ;
  assign n17491 = ~n17489 & ~n17490 ;
  assign n17492 = \wishbone_bd_ram_mem3_reg[145][26]/P0001  & n13715 ;
  assign n17493 = \wishbone_bd_ram_mem3_reg[104][26]/P0001  & n13684 ;
  assign n17494 = ~n17492 & ~n17493 ;
  assign n17495 = n17491 & n17494 ;
  assign n17496 = \wishbone_bd_ram_mem3_reg[112][26]/P0001  & n13482 ;
  assign n17497 = \wishbone_bd_ram_mem3_reg[108][26]/P0001  & n13814 ;
  assign n17498 = ~n17496 & ~n17497 ;
  assign n17499 = \wishbone_bd_ram_mem3_reg[135][26]/P0001  & n13672 ;
  assign n17500 = \wishbone_bd_ram_mem3_reg[12][26]/P0001  & n13733 ;
  assign n17501 = ~n17499 & ~n17500 ;
  assign n17502 = n17498 & n17501 ;
  assign n17503 = n17495 & n17502 ;
  assign n17504 = \wishbone_bd_ram_mem3_reg[10][26]/P0001  & n13837 ;
  assign n17505 = \wishbone_bd_ram_mem3_reg[29][26]/P0001  & n13412 ;
  assign n17506 = ~n17504 & ~n17505 ;
  assign n17507 = \wishbone_bd_ram_mem3_reg[87][26]/P0001  & n13691 ;
  assign n17508 = \wishbone_bd_ram_mem3_reg[141][26]/P0001  & n13852 ;
  assign n17509 = ~n17507 & ~n17508 ;
  assign n17510 = n17506 & n17509 ;
  assign n17511 = \wishbone_bd_ram_mem3_reg[11][26]/P0001  & n13774 ;
  assign n17512 = \wishbone_bd_ram_mem3_reg[41][26]/P0001  & n14017 ;
  assign n17513 = ~n17511 & ~n17512 ;
  assign n17514 = \wishbone_bd_ram_mem3_reg[40][26]/P0001  & n13661 ;
  assign n17515 = \wishbone_bd_ram_mem3_reg[151][26]/P0001  & n13697 ;
  assign n17516 = ~n17514 & ~n17515 ;
  assign n17517 = n17513 & n17516 ;
  assign n17518 = n17510 & n17517 ;
  assign n17519 = n17503 & n17518 ;
  assign n17520 = n17488 & n17519 ;
  assign n17521 = n17457 & n17520 ;
  assign n17522 = \wishbone_bd_ram_mem3_reg[16][26]/P0001  & n13695 ;
  assign n17523 = \wishbone_bd_ram_mem3_reg[81][26]/P0001  & n13409 ;
  assign n17524 = ~n17522 & ~n17523 ;
  assign n17525 = \wishbone_bd_ram_mem3_reg[140][26]/P0001  & n13287 ;
  assign n17526 = \wishbone_bd_ram_mem3_reg[98][26]/P0001  & n13569 ;
  assign n17527 = ~n17525 & ~n17526 ;
  assign n17528 = n17524 & n17527 ;
  assign n17529 = \wishbone_bd_ram_mem3_reg[231][26]/P0001  & n13363 ;
  assign n17530 = \wishbone_bd_ram_mem3_reg[176][26]/P0001  & n13262 ;
  assign n17531 = ~n17529 & ~n17530 ;
  assign n17532 = \wishbone_bd_ram_mem3_reg[50][26]/P0001  & n13686 ;
  assign n17533 = \wishbone_bd_ram_mem3_reg[153][26]/P0001  & n13309 ;
  assign n17534 = ~n17532 & ~n17533 ;
  assign n17535 = n17531 & n17534 ;
  assign n17536 = n17528 & n17535 ;
  assign n17537 = \wishbone_bd_ram_mem3_reg[105][26]/P0001  & n13503 ;
  assign n17538 = \wishbone_bd_ram_mem3_reg[92][26]/P0001  & n13859 ;
  assign n17539 = ~n17537 & ~n17538 ;
  assign n17540 = \wishbone_bd_ram_mem3_reg[193][26]/P0001  & n14022 ;
  assign n17541 = \wishbone_bd_ram_mem3_reg[203][26]/P0001  & n13816 ;
  assign n17542 = ~n17540 & ~n17541 ;
  assign n17543 = n17539 & n17542 ;
  assign n17544 = \wishbone_bd_ram_mem3_reg[133][26]/P0001  & n13492 ;
  assign n17545 = \wishbone_bd_ram_mem3_reg[1][26]/P0001  & n13888 ;
  assign n17546 = ~n17544 & ~n17545 ;
  assign n17547 = \wishbone_bd_ram_mem3_reg[223][26]/P0001  & n13335 ;
  assign n17548 = \wishbone_bd_ram_mem3_reg[137][26]/P0001  & n13808 ;
  assign n17549 = ~n17547 & ~n17548 ;
  assign n17550 = n17546 & n17549 ;
  assign n17551 = n17543 & n17550 ;
  assign n17552 = n17536 & n17551 ;
  assign n17553 = \wishbone_bd_ram_mem3_reg[47][26]/P0001  & n13436 ;
  assign n17554 = \wishbone_bd_ram_mem3_reg[113][26]/P0001  & n13882 ;
  assign n17555 = ~n17553 & ~n17554 ;
  assign n17556 = \wishbone_bd_ram_mem3_reg[131][26]/P0001  & n13358 ;
  assign n17557 = \wishbone_bd_ram_mem3_reg[19][26]/P0001  & n13886 ;
  assign n17558 = ~n17556 & ~n17557 ;
  assign n17559 = n17555 & n17558 ;
  assign n17560 = \wishbone_bd_ram_mem3_reg[89][26]/P0001  & n13910 ;
  assign n17561 = \wishbone_bd_ram_mem3_reg[77][26]/P0001  & n13935 ;
  assign n17562 = ~n17560 & ~n17561 ;
  assign n17563 = \wishbone_bd_ram_mem3_reg[166][26]/P0001  & n13999 ;
  assign n17564 = \wishbone_bd_ram_mem3_reg[107][26]/P0001  & n13476 ;
  assign n17565 = ~n17563 & ~n17564 ;
  assign n17566 = n17562 & n17565 ;
  assign n17567 = n17559 & n17566 ;
  assign n17568 = \wishbone_bd_ram_mem3_reg[43][26]/P0001  & n13761 ;
  assign n17569 = \wishbone_bd_ram_mem3_reg[132][26]/P0001  & n13927 ;
  assign n17570 = ~n17568 & ~n17569 ;
  assign n17571 = \wishbone_bd_ram_mem3_reg[62][26]/P0001  & n13529 ;
  assign n17572 = \wishbone_bd_ram_mem3_reg[48][26]/P0001  & n13917 ;
  assign n17573 = ~n17571 & ~n17572 ;
  assign n17574 = n17570 & n17573 ;
  assign n17575 = \wishbone_bd_ram_mem3_reg[102][26]/P0001  & n13534 ;
  assign n17576 = \wishbone_bd_ram_mem3_reg[233][26]/P0001  & n13332 ;
  assign n17577 = ~n17575 & ~n17576 ;
  assign n17578 = \wishbone_bd_ram_mem3_reg[255][26]/P0001  & n13952 ;
  assign n17579 = \wishbone_bd_ram_mem3_reg[155][26]/P0001  & n13738 ;
  assign n17580 = ~n17578 & ~n17579 ;
  assign n17581 = n17577 & n17580 ;
  assign n17582 = n17574 & n17581 ;
  assign n17583 = n17567 & n17582 ;
  assign n17584 = n17552 & n17583 ;
  assign n17585 = \wishbone_bd_ram_mem3_reg[250][26]/P0001  & n13677 ;
  assign n17586 = \wishbone_bd_ram_mem3_reg[124][26]/P0001  & n14024 ;
  assign n17587 = ~n17585 & ~n17586 ;
  assign n17588 = \wishbone_bd_ram_mem3_reg[78][26]/P0001  & n13277 ;
  assign n17589 = \wishbone_bd_ram_mem3_reg[191][26]/P0001  & n14012 ;
  assign n17590 = ~n17588 & ~n17589 ;
  assign n17591 = n17587 & n17590 ;
  assign n17592 = \wishbone_bd_ram_mem3_reg[192][26]/P0001  & n13390 ;
  assign n17593 = \wishbone_bd_ram_mem3_reg[225][26]/P0001  & n13719 ;
  assign n17594 = ~n17592 & ~n17593 ;
  assign n17595 = \wishbone_bd_ram_mem3_reg[88][26]/P0001  & n13347 ;
  assign n17596 = \wishbone_bd_ram_mem3_reg[148][26]/P0001  & n13868 ;
  assign n17597 = ~n17595 & ~n17596 ;
  assign n17598 = n17594 & n17597 ;
  assign n17599 = n17591 & n17598 ;
  assign n17600 = \wishbone_bd_ram_mem3_reg[227][26]/P0001  & n13388 ;
  assign n17601 = \wishbone_bd_ram_mem3_reg[180][26]/P0001  & n13650 ;
  assign n17602 = ~n17600 & ~n17601 ;
  assign n17603 = \wishbone_bd_ram_mem3_reg[202][26]/P0001  & n13268 ;
  assign n17604 = \wishbone_bd_ram_mem3_reg[200][26]/P0001  & n13922 ;
  assign n17605 = ~n17603 & ~n17604 ;
  assign n17606 = n17602 & n17605 ;
  assign n17607 = \wishbone_bd_ram_mem3_reg[171][26]/P0001  & n13422 ;
  assign n17608 = \wishbone_bd_ram_mem3_reg[214][26]/P0001  & n13938 ;
  assign n17609 = ~n17607 & ~n17608 ;
  assign n17610 = \wishbone_bd_ram_mem3_reg[93][26]/P0001  & n13891 ;
  assign n17611 = \wishbone_bd_ram_mem3_reg[152][26]/P0001  & n13912 ;
  assign n17612 = ~n17610 & ~n17611 ;
  assign n17613 = n17609 & n17612 ;
  assign n17614 = n17606 & n17613 ;
  assign n17615 = n17599 & n17614 ;
  assign n17616 = \wishbone_bd_ram_mem3_reg[60][26]/P0001  & n13790 ;
  assign n17617 = \wishbone_bd_ram_mem3_reg[100][26]/P0001  & n13401 ;
  assign n17618 = ~n17616 & ~n17617 ;
  assign n17619 = \wishbone_bd_ram_mem3_reg[83][26]/P0001  & n13454 ;
  assign n17620 = \wishbone_bd_ram_mem3_reg[169][26]/P0001  & n13541 ;
  assign n17621 = ~n17619 & ~n17620 ;
  assign n17622 = n17618 & n17621 ;
  assign n17623 = \wishbone_bd_ram_mem3_reg[136][26]/P0001  & n13963 ;
  assign n17624 = \wishbone_bd_ram_mem3_reg[216][26]/P0001  & n14005 ;
  assign n17625 = ~n17623 & ~n17624 ;
  assign n17626 = \wishbone_bd_ram_mem3_reg[97][26]/P0001  & n13724 ;
  assign n17627 = \wishbone_bd_ram_mem3_reg[53][26]/P0001  & n13875 ;
  assign n17628 = ~n17626 & ~n17627 ;
  assign n17629 = n17625 & n17628 ;
  assign n17630 = n17622 & n17629 ;
  assign n17631 = \wishbone_bd_ram_mem3_reg[220][26]/P0001  & n13965 ;
  assign n17632 = \wishbone_bd_ram_mem3_reg[82][26]/P0001  & n13374 ;
  assign n17633 = ~n17631 & ~n17632 ;
  assign n17634 = \wishbone_bd_ram_mem3_reg[196][26]/P0001  & n13977 ;
  assign n17635 = \wishbone_bd_ram_mem3_reg[226][26]/P0001  & n13668 ;
  assign n17636 = ~n17634 & ~n17635 ;
  assign n17637 = n17633 & n17636 ;
  assign n17638 = \wishbone_bd_ram_mem3_reg[114][26]/P0001  & n13763 ;
  assign n17639 = \wishbone_bd_ram_mem3_reg[251][26]/P0001  & n14019 ;
  assign n17640 = ~n17638 & ~n17639 ;
  assign n17641 = \wishbone_bd_ram_mem3_reg[3][26]/P0001  & n13354 ;
  assign n17642 = \wishbone_bd_ram_mem3_reg[49][26]/P0001  & n13929 ;
  assign n17643 = ~n17641 & ~n17642 ;
  assign n17644 = n17640 & n17643 ;
  assign n17645 = n17637 & n17644 ;
  assign n17646 = n17630 & n17645 ;
  assign n17647 = n17615 & n17646 ;
  assign n17648 = n17584 & n17647 ;
  assign n17649 = n17521 & n17648 ;
  assign n17650 = \wishbone_bd_ram_mem3_reg[39][26]/P0001  & n13893 ;
  assign n17651 = \wishbone_bd_ram_mem3_reg[244][26]/P0001  & n13474 ;
  assign n17652 = ~n17650 & ~n17651 ;
  assign n17653 = \wishbone_bd_ram_mem3_reg[23][26]/P0001  & n13857 ;
  assign n17654 = \wishbone_bd_ram_mem3_reg[238][26]/P0001  & n13819 ;
  assign n17655 = ~n17653 & ~n17654 ;
  assign n17656 = n17652 & n17655 ;
  assign n17657 = \wishbone_bd_ram_mem3_reg[118][26]/P0001  & n13589 ;
  assign n17658 = \wishbone_bd_ram_mem3_reg[37][26]/P0001  & n13710 ;
  assign n17659 = ~n17657 & ~n17658 ;
  assign n17660 = \wishbone_bd_ram_mem3_reg[190][26]/P0001  & n13365 ;
  assign n17661 = \wishbone_bd_ram_mem3_reg[210][26]/P0001  & n13443 ;
  assign n17662 = ~n17660 & ~n17661 ;
  assign n17663 = n17659 & n17662 ;
  assign n17664 = n17656 & n17663 ;
  assign n17665 = \wishbone_bd_ram_mem3_reg[130][26]/P0001  & n13427 ;
  assign n17666 = \wishbone_bd_ram_mem3_reg[13][26]/P0001  & n13844 ;
  assign n17667 = ~n17665 & ~n17666 ;
  assign n17668 = \wishbone_bd_ram_mem3_reg[224][26]/P0001  & n13433 ;
  assign n17669 = \wishbone_bd_ram_mem3_reg[117][26]/P0001  & n13557 ;
  assign n17670 = ~n17668 & ~n17669 ;
  assign n17671 = n17667 & n17670 ;
  assign n17672 = \wishbone_bd_ram_mem3_reg[61][26]/P0001  & n13544 ;
  assign n17673 = \wishbone_bd_ram_mem3_reg[52][26]/P0001  & n13988 ;
  assign n17674 = ~n17672 & ~n17673 ;
  assign n17675 = \wishbone_bd_ram_mem3_reg[162][26]/P0001  & n13726 ;
  assign n17676 = \wishbone_bd_ram_mem3_reg[109][26]/P0001  & n13306 ;
  assign n17677 = ~n17675 & ~n17676 ;
  assign n17678 = n17674 & n17677 ;
  assign n17679 = n17671 & n17678 ;
  assign n17680 = n17664 & n17679 ;
  assign n17681 = \wishbone_bd_ram_mem3_reg[241][26]/P0001  & n13854 ;
  assign n17682 = \wishbone_bd_ram_mem3_reg[42][26]/P0001  & n13341 ;
  assign n17683 = ~n17681 & ~n17682 ;
  assign n17684 = \wishbone_bd_ram_mem3_reg[17][26]/P0001  & n13324 ;
  assign n17685 = \wishbone_bd_ram_mem3_reg[38][26]/P0001  & n13828 ;
  assign n17686 = ~n17684 & ~n17685 ;
  assign n17687 = n17683 & n17686 ;
  assign n17688 = \wishbone_bd_ram_mem3_reg[219][26]/P0001  & n13577 ;
  assign n17689 = \wishbone_bd_ram_mem3_reg[45][26]/P0001  & n13420 ;
  assign n17690 = ~n17688 & ~n17689 ;
  assign n17691 = \wishbone_bd_ram_mem3_reg[94][26]/P0001  & n13833 ;
  assign n17692 = \wishbone_bd_ram_mem3_reg[222][26]/P0001  & n13721 ;
  assign n17693 = ~n17691 & ~n17692 ;
  assign n17694 = n17690 & n17693 ;
  assign n17695 = n17687 & n17694 ;
  assign n17696 = \wishbone_bd_ram_mem3_reg[68][26]/P0001  & n13379 ;
  assign n17697 = \wishbone_bd_ram_mem3_reg[58][26]/P0001  & n13949 ;
  assign n17698 = ~n17696 & ~n17697 ;
  assign n17699 = \wishbone_bd_ram_mem3_reg[91][26]/P0001  & n13954 ;
  assign n17700 = \wishbone_bd_ram_mem3_reg[74][26]/P0001  & n13564 ;
  assign n17701 = ~n17699 & ~n17700 ;
  assign n17702 = n17698 & n17701 ;
  assign n17703 = \wishbone_bd_ram_mem3_reg[167][26]/P0001  & n13940 ;
  assign n17704 = \wishbone_bd_ram_mem3_reg[14][26]/P0001  & n13972 ;
  assign n17705 = ~n17703 & ~n17704 ;
  assign n17706 = \wishbone_bd_ram_mem3_reg[25][26]/P0001  & n13742 ;
  assign n17707 = \wishbone_bd_ram_mem3_reg[31][26]/P0001  & n13758 ;
  assign n17708 = ~n17706 & ~n17707 ;
  assign n17709 = n17705 & n17708 ;
  assign n17710 = n17702 & n17709 ;
  assign n17711 = n17695 & n17710 ;
  assign n17712 = n17680 & n17711 ;
  assign n17713 = \wishbone_bd_ram_mem3_reg[213][26]/P0001  & n13870 ;
  assign n17714 = \wishbone_bd_ram_mem3_reg[168][26]/P0001  & n13795 ;
  assign n17715 = ~n17713 & ~n17714 ;
  assign n17716 = \wishbone_bd_ram_mem3_reg[0][26]/P0001  & n13539 ;
  assign n17717 = \wishbone_bd_ram_mem3_reg[175][26]/P0001  & n13674 ;
  assign n17718 = ~n17716 & ~n17717 ;
  assign n17719 = n17715 & n17718 ;
  assign n17720 = \wishbone_bd_ram_mem3_reg[249][26]/P0001  & n13431 ;
  assign n17721 = \wishbone_bd_ram_mem3_reg[230][26]/P0001  & n13994 ;
  assign n17722 = ~n17720 & ~n17721 ;
  assign n17723 = \wishbone_bd_ram_mem3_reg[163][26]/P0001  & n13255 ;
  assign n17724 = \wishbone_bd_ram_mem3_reg[66][26]/P0001  & n13603 ;
  assign n17725 = ~n17723 & ~n17724 ;
  assign n17726 = n17722 & n17725 ;
  assign n17727 = n17719 & n17726 ;
  assign n17728 = \wishbone_bd_ram_mem3_reg[2][26]/P0001  & n13975 ;
  assign n17729 = \wishbone_bd_ram_mem3_reg[218][26]/P0001  & n13792 ;
  assign n17730 = ~n17728 & ~n17729 ;
  assign n17731 = \wishbone_bd_ram_mem3_reg[149][26]/P0001  & n13469 ;
  assign n17732 = \wishbone_bd_ram_mem3_reg[235][26]/P0001  & n13518 ;
  assign n17733 = ~n17731 & ~n17732 ;
  assign n17734 = n17730 & n17733 ;
  assign n17735 = \wishbone_bd_ram_mem3_reg[4][26]/P0001  & n13527 ;
  assign n17736 = \wishbone_bd_ram_mem3_reg[116][26]/P0001  & n13865 ;
  assign n17737 = ~n17735 & ~n17736 ;
  assign n17738 = \wishbone_bd_ram_mem3_reg[150][26]/P0001  & n13666 ;
  assign n17739 = \wishbone_bd_ram_mem3_reg[187][26]/P0001  & n13756 ;
  assign n17740 = ~n17738 & ~n17739 ;
  assign n17741 = n17737 & n17740 ;
  assign n17742 = n17734 & n17741 ;
  assign n17743 = n17727 & n17742 ;
  assign n17744 = \wishbone_bd_ram_mem3_reg[183][26]/P0001  & n13645 ;
  assign n17745 = \wishbone_bd_ram_mem3_reg[126][26]/P0001  & n13786 ;
  assign n17746 = ~n17744 & ~n17745 ;
  assign n17747 = \wishbone_bd_ram_mem3_reg[142][26]/P0001  & n13448 ;
  assign n17748 = \wishbone_bd_ram_mem3_reg[172][26]/P0001  & n13377 ;
  assign n17749 = ~n17747 & ~n17748 ;
  assign n17750 = n17746 & n17749 ;
  assign n17751 = \wishbone_bd_ram_mem3_reg[174][26]/P0001  & n13899 ;
  assign n17752 = \wishbone_bd_ram_mem3_reg[211][26]/P0001  & n13805 ;
  assign n17753 = ~n17751 & ~n17752 ;
  assign n17754 = \wishbone_bd_ram_mem3_reg[195][26]/P0001  & n13700 ;
  assign n17755 = \wishbone_bd_ram_mem3_reg[243][26]/P0001  & n13575 ;
  assign n17756 = ~n17754 & ~n17755 ;
  assign n17757 = n17753 & n17756 ;
  assign n17758 = n17750 & n17757 ;
  assign n17759 = \wishbone_bd_ram_mem3_reg[240][26]/P0001  & n13352 ;
  assign n17760 = \wishbone_bd_ram_mem3_reg[69][26]/P0001  & n13487 ;
  assign n17761 = ~n17759 & ~n17760 ;
  assign n17762 = \wishbone_bd_ram_mem3_reg[154][26]/P0001  & n13403 ;
  assign n17763 = \wishbone_bd_ram_mem3_reg[110][26]/P0001  & n14030 ;
  assign n17764 = ~n17762 & ~n17763 ;
  assign n17765 = n17761 & n17764 ;
  assign n17766 = \wishbone_bd_ram_mem3_reg[73][26]/P0001  & n13456 ;
  assign n17767 = \wishbone_bd_ram_mem3_reg[24][26]/P0001  & n13970 ;
  assign n17768 = ~n17766 & ~n17767 ;
  assign n17769 = \wishbone_bd_ram_mem3_reg[33][26]/P0001  & n13933 ;
  assign n17770 = \wishbone_bd_ram_mem3_reg[8][26]/P0001  & n13459 ;
  assign n17771 = ~n17769 & ~n17770 ;
  assign n17772 = n17768 & n17771 ;
  assign n17773 = n17765 & n17772 ;
  assign n17774 = n17758 & n17773 ;
  assign n17775 = n17743 & n17774 ;
  assign n17776 = n17712 & n17775 ;
  assign n17777 = \wishbone_bd_ram_mem3_reg[84][26]/P0001  & n13385 ;
  assign n17778 = \wishbone_bd_ram_mem3_reg[186][26]/P0001  & n13616 ;
  assign n17779 = ~n17777 & ~n17778 ;
  assign n17780 = \wishbone_bd_ram_mem3_reg[99][26]/P0001  & n13996 ;
  assign n17781 = \wishbone_bd_ram_mem3_reg[123][26]/P0001  & n13749 ;
  assign n17782 = ~n17780 & ~n17781 ;
  assign n17783 = n17779 & n17782 ;
  assign n17784 = \wishbone_bd_ram_mem3_reg[96][26]/P0001  & n13425 ;
  assign n17785 = \wishbone_bd_ram_mem3_reg[59][26]/P0001  & n13613 ;
  assign n17786 = ~n17784 & ~n17785 ;
  assign n17787 = \wishbone_bd_ram_mem3_reg[161][26]/P0001  & n13505 ;
  assign n17788 = \wishbone_bd_ram_mem3_reg[221][26]/P0001  & n13641 ;
  assign n17789 = ~n17787 & ~n17788 ;
  assign n17790 = n17786 & n17789 ;
  assign n17791 = n17783 & n17790 ;
  assign n17792 = \wishbone_bd_ram_mem3_reg[129][26]/P0001  & n13629 ;
  assign n17793 = \wishbone_bd_ram_mem3_reg[237][26]/P0001  & n13924 ;
  assign n17794 = ~n17792 & ~n17793 ;
  assign n17795 = \wishbone_bd_ram_mem3_reg[22][26]/P0001  & n13744 ;
  assign n17796 = \wishbone_bd_ram_mem3_reg[199][26]/P0001  & n13499 ;
  assign n17797 = ~n17795 & ~n17796 ;
  assign n17798 = n17794 & n17797 ;
  assign n17799 = \wishbone_bd_ram_mem3_reg[70][26]/P0001  & n13339 ;
  assign n17800 = \wishbone_bd_ram_mem3_reg[9][26]/P0001  & n13580 ;
  assign n17801 = ~n17799 & ~n17800 ;
  assign n17802 = \wishbone_bd_ram_mem3_reg[51][26]/P0001  & n13880 ;
  assign n17803 = \wishbone_bd_ram_mem3_reg[72][26]/P0001  & n13582 ;
  assign n17804 = ~n17802 & ~n17803 ;
  assign n17805 = n17801 & n17804 ;
  assign n17806 = n17798 & n17805 ;
  assign n17807 = n17791 & n17806 ;
  assign n17808 = \wishbone_bd_ram_mem3_reg[27][26]/P0001  & n13251 ;
  assign n17809 = \wishbone_bd_ram_mem3_reg[147][26]/P0001  & n13702 ;
  assign n17810 = ~n17808 & ~n17809 ;
  assign n17811 = \wishbone_bd_ram_mem3_reg[80][26]/P0001  & n13516 ;
  assign n17812 = \wishbone_bd_ram_mem3_reg[103][26]/P0001  & n13320 ;
  assign n17813 = ~n17811 & ~n17812 ;
  assign n17814 = n17810 & n17813 ;
  assign n17815 = \wishbone_bd_ram_mem3_reg[156][26]/P0001  & n13769 ;
  assign n17816 = \wishbone_bd_ram_mem3_reg[208][26]/P0001  & n14010 ;
  assign n17817 = ~n17815 & ~n17816 ;
  assign n17818 = \wishbone_bd_ram_mem3_reg[28][26]/P0001  & n13810 ;
  assign n17819 = \wishbone_bd_ram_mem3_reg[7][26]/P0001  & n13546 ;
  assign n17820 = ~n17818 & ~n17819 ;
  assign n17821 = n17817 & n17820 ;
  assign n17822 = n17814 & n17821 ;
  assign n17823 = \wishbone_bd_ram_mem3_reg[177][26]/P0001  & n13863 ;
  assign n17824 = \wishbone_bd_ram_mem3_reg[139][26]/P0001  & n13566 ;
  assign n17825 = ~n17823 & ~n17824 ;
  assign n17826 = \wishbone_bd_ram_mem3_reg[165][26]/P0001  & n14028 ;
  assign n17827 = \wishbone_bd_ram_mem3_reg[128][26]/P0001  & n13652 ;
  assign n17828 = ~n17826 & ~n17827 ;
  assign n17829 = n17825 & n17828 ;
  assign n17830 = \wishbone_bd_ram_mem3_reg[30][26]/P0001  & n13713 ;
  assign n17831 = \wishbone_bd_ram_mem3_reg[20][26]/P0001  & n13839 ;
  assign n17832 = ~n17830 & ~n17831 ;
  assign n17833 = \wishbone_bd_ram_mem3_reg[252][26]/P0001  & n13986 ;
  assign n17834 = \wishbone_bd_ram_mem3_reg[71][26]/P0001  & n13636 ;
  assign n17835 = ~n17833 & ~n17834 ;
  assign n17836 = n17832 & n17835 ;
  assign n17837 = n17829 & n17836 ;
  assign n17838 = n17822 & n17837 ;
  assign n17839 = n17807 & n17838 ;
  assign n17840 = \wishbone_bd_ram_mem3_reg[236][26]/P0001  & n13480 ;
  assign n17841 = \wishbone_bd_ram_mem3_reg[5][26]/P0001  & n13243 ;
  assign n17842 = ~n17840 & ~n17841 ;
  assign n17843 = \wishbone_bd_ram_mem3_reg[106][26]/P0001  & n13555 ;
  assign n17844 = \wishbone_bd_ram_mem3_reg[184][26]/P0001  & n13960 ;
  assign n17845 = ~n17843 & ~n17844 ;
  assign n17846 = n17842 & n17845 ;
  assign n17847 = \wishbone_bd_ram_mem3_reg[79][26]/P0001  & n13779 ;
  assign n17848 = \wishbone_bd_ram_mem3_reg[232][26]/P0001  & n13510 ;
  assign n17849 = ~n17847 & ~n17848 ;
  assign n17850 = \wishbone_bd_ram_mem3_reg[122][26]/P0001  & n13679 ;
  assign n17851 = \wishbone_bd_ram_mem3_reg[197][26]/P0001  & n13594 ;
  assign n17852 = ~n17850 & ~n17851 ;
  assign n17853 = n17849 & n17852 ;
  assign n17854 = n17846 & n17853 ;
  assign n17855 = \wishbone_bd_ram_mem3_reg[85][26]/P0001  & n13784 ;
  assign n17856 = \wishbone_bd_ram_mem3_reg[46][26]/P0001  & n13298 ;
  assign n17857 = ~n17855 & ~n17856 ;
  assign n17858 = \wishbone_bd_ram_mem3_reg[44][26]/P0001  & n13291 ;
  assign n17859 = \wishbone_bd_ram_mem3_reg[35][26]/P0001  & n13523 ;
  assign n17860 = ~n17858 & ~n17859 ;
  assign n17861 = n17857 & n17860 ;
  assign n17862 = \wishbone_bd_ram_mem3_reg[245][26]/P0001  & n13877 ;
  assign n17863 = \wishbone_bd_ram_mem3_reg[164][26]/P0001  & n13236 ;
  assign n17864 = ~n17862 & ~n17863 ;
  assign n17865 = \wishbone_bd_ram_mem3_reg[246][26]/P0001  & n13981 ;
  assign n17866 = \wishbone_bd_ram_mem3_reg[95][26]/P0001  & n13317 ;
  assign n17867 = ~n17865 & ~n17866 ;
  assign n17868 = n17864 & n17867 ;
  assign n17869 = n17861 & n17868 ;
  assign n17870 = n17854 & n17869 ;
  assign n17871 = \wishbone_bd_ram_mem3_reg[34][26]/P0001  & n13450 ;
  assign n17872 = \wishbone_bd_ram_mem3_reg[134][26]/P0001  & n13494 ;
  assign n17873 = ~n17871 & ~n17872 ;
  assign n17874 = \wishbone_bd_ram_mem3_reg[121][26]/P0001  & n13983 ;
  assign n17875 = \wishbone_bd_ram_mem3_reg[21][26]/P0001  & n13438 ;
  assign n17876 = ~n17874 & ~n17875 ;
  assign n17877 = n17873 & n17876 ;
  assign n17878 = \wishbone_bd_ram_mem3_reg[194][26]/P0001  & n13624 ;
  assign n17879 = \wishbone_bd_ram_mem3_reg[179][26]/P0001  & n14035 ;
  assign n17880 = ~n17878 & ~n17879 ;
  assign n17881 = \wishbone_bd_ram_mem3_reg[6][26]/P0001  & n13915 ;
  assign n17882 = \wishbone_bd_ram_mem3_reg[173][26]/P0001  & n13360 ;
  assign n17883 = ~n17881 & ~n17882 ;
  assign n17884 = n17880 & n17883 ;
  assign n17885 = n17877 & n17884 ;
  assign n17886 = \wishbone_bd_ram_mem3_reg[115][26]/P0001  & n13747 ;
  assign n17887 = \wishbone_bd_ram_mem3_reg[181][26]/P0001  & n13587 ;
  assign n17888 = ~n17886 & ~n17887 ;
  assign n17889 = \wishbone_bd_ram_mem3_reg[234][26]/P0001  & n13781 ;
  assign n17890 = \wishbone_bd_ram_mem3_reg[158][26]/P0001  & n13294 ;
  assign n17891 = ~n17889 & ~n17890 ;
  assign n17892 = n17888 & n17891 ;
  assign n17893 = \wishbone_bd_ram_mem3_reg[101][26]/P0001  & n13772 ;
  assign n17894 = \wishbone_bd_ram_mem3_reg[198][26]/P0001  & n13592 ;
  assign n17895 = ~n17893 & ~n17894 ;
  assign n17896 = \wishbone_bd_ram_mem3_reg[144][26]/P0001  & n13508 ;
  assign n17897 = \wishbone_bd_ram_mem3_reg[170][26]/P0001  & n14007 ;
  assign n17898 = ~n17896 & ~n17897 ;
  assign n17899 = n17895 & n17898 ;
  assign n17900 = n17892 & n17899 ;
  assign n17901 = n17885 & n17900 ;
  assign n17902 = n17870 & n17901 ;
  assign n17903 = n17839 & n17902 ;
  assign n17904 = n17776 & n17903 ;
  assign n17905 = n17649 & n17904 ;
  assign n17906 = n14047 & ~n17905 ;
  assign n17907 = \wishbone_TxLength_reg[10]/NET0131  & n14069 ;
  assign n17908 = \wishbone_TxLength_reg[10]/NET0131  & ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n17909 = ~n14070 & n17908 ;
  assign n17910 = ~n17907 & ~n17909 ;
  assign n17911 = ~n14063 & n17910 ;
  assign n17912 = n14049 & n14053 ;
  assign n17913 = n14057 & n17912 ;
  assign n17914 = ~n17911 & n17913 ;
  assign n17915 = n14049 & n14069 ;
  assign n17916 = ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  & n14049 ;
  assign n17917 = ~n14070 & n17916 ;
  assign n17918 = ~n17915 & ~n17917 ;
  assign n17919 = n14058 & ~n17918 ;
  assign n17920 = ~\wishbone_TxLength_reg[10]/NET0131  & ~n17919 ;
  assign n17921 = ~n14046 & ~n17920 ;
  assign n17922 = ~n17914 & n17921 ;
  assign n17923 = ~n17906 & ~n17922 ;
  assign n17924 = \wishbone_bd_ram_mem3_reg[157][25]/P0001  & n13445 ;
  assign n17925 = \wishbone_bd_ram_mem3_reg[183][25]/P0001  & n13645 ;
  assign n17926 = ~n17924 & ~n17925 ;
  assign n17927 = \wishbone_bd_ram_mem3_reg[24][25]/P0001  & n13970 ;
  assign n17928 = \wishbone_bd_ram_mem3_reg[51][25]/P0001  & n13880 ;
  assign n17929 = ~n17927 & ~n17928 ;
  assign n17930 = n17926 & n17929 ;
  assign n17931 = \wishbone_bd_ram_mem3_reg[222][25]/P0001  & n13721 ;
  assign n17932 = \wishbone_bd_ram_mem3_reg[172][25]/P0001  & n13377 ;
  assign n17933 = ~n17931 & ~n17932 ;
  assign n17934 = \wishbone_bd_ram_mem3_reg[85][25]/P0001  & n13784 ;
  assign n17935 = \wishbone_bd_ram_mem3_reg[242][25]/P0001  & n13383 ;
  assign n17936 = ~n17934 & ~n17935 ;
  assign n17937 = n17933 & n17936 ;
  assign n17938 = n17930 & n17937 ;
  assign n17939 = \wishbone_bd_ram_mem3_reg[217][25]/P0001  & n13767 ;
  assign n17940 = \wishbone_bd_ram_mem3_reg[140][25]/P0001  & n13287 ;
  assign n17941 = ~n17939 & ~n17940 ;
  assign n17942 = \wishbone_bd_ram_mem3_reg[34][25]/P0001  & n13450 ;
  assign n17943 = \wishbone_bd_ram_mem3_reg[93][25]/P0001  & n13891 ;
  assign n17944 = ~n17942 & ~n17943 ;
  assign n17945 = n17941 & n17944 ;
  assign n17946 = \wishbone_bd_ram_mem3_reg[234][25]/P0001  & n13781 ;
  assign n17947 = \wishbone_bd_ram_mem3_reg[105][25]/P0001  & n13503 ;
  assign n17948 = ~n17946 & ~n17947 ;
  assign n17949 = \wishbone_bd_ram_mem3_reg[253][25]/P0001  & n13708 ;
  assign n17950 = \wishbone_bd_ram_mem3_reg[108][25]/P0001  & n13814 ;
  assign n17951 = ~n17949 & ~n17950 ;
  assign n17952 = n17948 & n17951 ;
  assign n17953 = n17945 & n17952 ;
  assign n17954 = n17938 & n17953 ;
  assign n17955 = \wishbone_bd_ram_mem3_reg[61][25]/P0001  & n13544 ;
  assign n17956 = \wishbone_bd_ram_mem3_reg[98][25]/P0001  & n13569 ;
  assign n17957 = ~n17955 & ~n17956 ;
  assign n17958 = \wishbone_bd_ram_mem3_reg[79][25]/P0001  & n13779 ;
  assign n17959 = \wishbone_bd_ram_mem3_reg[202][25]/P0001  & n13268 ;
  assign n17960 = ~n17958 & ~n17959 ;
  assign n17961 = n17957 & n17960 ;
  assign n17962 = \wishbone_bd_ram_mem3_reg[213][25]/P0001  & n13870 ;
  assign n17963 = \wishbone_bd_ram_mem3_reg[90][25]/P0001  & n13906 ;
  assign n17964 = ~n17962 & ~n17963 ;
  assign n17965 = \wishbone_bd_ram_mem3_reg[110][25]/P0001  & n14030 ;
  assign n17966 = \wishbone_bd_ram_mem3_reg[243][25]/P0001  & n13575 ;
  assign n17967 = ~n17965 & ~n17966 ;
  assign n17968 = n17964 & n17967 ;
  assign n17969 = n17961 & n17968 ;
  assign n17970 = \wishbone_bd_ram_mem3_reg[153][25]/P0001  & n13309 ;
  assign n17971 = \wishbone_bd_ram_mem3_reg[94][25]/P0001  & n13833 ;
  assign n17972 = ~n17970 & ~n17971 ;
  assign n17973 = \wishbone_bd_ram_mem3_reg[122][25]/P0001  & n13679 ;
  assign n17974 = \wishbone_bd_ram_mem3_reg[144][25]/P0001  & n13508 ;
  assign n17975 = ~n17973 & ~n17974 ;
  assign n17976 = n17972 & n17975 ;
  assign n17977 = \wishbone_bd_ram_mem3_reg[1][25]/P0001  & n13888 ;
  assign n17978 = \wishbone_bd_ram_mem3_reg[220][25]/P0001  & n13965 ;
  assign n17979 = ~n17977 & ~n17978 ;
  assign n17980 = \wishbone_bd_ram_mem3_reg[64][25]/P0001  & n13904 ;
  assign n17981 = \wishbone_bd_ram_mem3_reg[190][25]/P0001  & n13365 ;
  assign n17982 = ~n17980 & ~n17981 ;
  assign n17983 = n17979 & n17982 ;
  assign n17984 = n17976 & n17983 ;
  assign n17985 = n17969 & n17984 ;
  assign n17986 = n17954 & n17985 ;
  assign n17987 = \wishbone_bd_ram_mem3_reg[127][25]/P0001  & n13803 ;
  assign n17988 = \wishbone_bd_ram_mem3_reg[101][25]/P0001  & n13772 ;
  assign n17989 = ~n17987 & ~n17988 ;
  assign n17990 = \wishbone_bd_ram_mem3_reg[154][25]/P0001  & n13403 ;
  assign n17991 = \wishbone_bd_ram_mem3_reg[50][25]/P0001  & n13686 ;
  assign n17992 = ~n17990 & ~n17991 ;
  assign n17993 = n17989 & n17992 ;
  assign n17994 = \wishbone_bd_ram_mem3_reg[211][25]/P0001  & n13805 ;
  assign n17995 = \wishbone_bd_ram_mem3_reg[149][25]/P0001  & n13469 ;
  assign n17996 = ~n17994 & ~n17995 ;
  assign n17997 = \wishbone_bd_ram_mem3_reg[227][25]/P0001  & n13388 ;
  assign n17998 = \wishbone_bd_ram_mem3_reg[96][25]/P0001  & n13425 ;
  assign n17999 = ~n17997 & ~n17998 ;
  assign n18000 = n17996 & n17999 ;
  assign n18001 = n17993 & n18000 ;
  assign n18002 = \wishbone_bd_ram_mem3_reg[52][25]/P0001  & n13988 ;
  assign n18003 = \wishbone_bd_ram_mem3_reg[196][25]/P0001  & n13977 ;
  assign n18004 = ~n18002 & ~n18003 ;
  assign n18005 = \wishbone_bd_ram_mem3_reg[74][25]/P0001  & n13564 ;
  assign n18006 = \wishbone_bd_ram_mem3_reg[112][25]/P0001  & n13482 ;
  assign n18007 = ~n18005 & ~n18006 ;
  assign n18008 = n18004 & n18007 ;
  assign n18009 = \wishbone_bd_ram_mem3_reg[165][25]/P0001  & n14028 ;
  assign n18010 = \wishbone_bd_ram_mem3_reg[252][25]/P0001  & n13986 ;
  assign n18011 = ~n18009 & ~n18010 ;
  assign n18012 = \wishbone_bd_ram_mem3_reg[29][25]/P0001  & n13412 ;
  assign n18013 = \wishbone_bd_ram_mem3_reg[205][25]/P0001  & n13947 ;
  assign n18014 = ~n18012 & ~n18013 ;
  assign n18015 = n18011 & n18014 ;
  assign n18016 = n18008 & n18015 ;
  assign n18017 = n18001 & n18016 ;
  assign n18018 = \wishbone_bd_ram_mem3_reg[59][25]/P0001  & n13613 ;
  assign n18019 = \wishbone_bd_ram_mem3_reg[128][25]/P0001  & n13652 ;
  assign n18020 = ~n18018 & ~n18019 ;
  assign n18021 = \wishbone_bd_ram_mem3_reg[47][25]/P0001  & n13436 ;
  assign n18022 = \wishbone_bd_ram_mem3_reg[177][25]/P0001  & n13863 ;
  assign n18023 = ~n18021 & ~n18022 ;
  assign n18024 = n18020 & n18023 ;
  assign n18025 = \wishbone_bd_ram_mem3_reg[100][25]/P0001  & n13401 ;
  assign n18026 = \wishbone_bd_ram_mem3_reg[60][25]/P0001  & n13790 ;
  assign n18027 = ~n18025 & ~n18026 ;
  assign n18028 = \wishbone_bd_ram_mem3_reg[39][25]/P0001  & n13893 ;
  assign n18029 = \wishbone_bd_ram_mem3_reg[166][25]/P0001  & n13999 ;
  assign n18030 = ~n18028 & ~n18029 ;
  assign n18031 = n18027 & n18030 ;
  assign n18032 = n18024 & n18031 ;
  assign n18033 = \wishbone_bd_ram_mem3_reg[176][25]/P0001  & n13262 ;
  assign n18034 = \wishbone_bd_ram_mem3_reg[3][25]/P0001  & n13354 ;
  assign n18035 = ~n18033 & ~n18034 ;
  assign n18036 = \wishbone_bd_ram_mem3_reg[81][25]/P0001  & n13409 ;
  assign n18037 = \wishbone_bd_ram_mem3_reg[77][25]/P0001  & n13935 ;
  assign n18038 = ~n18036 & ~n18037 ;
  assign n18039 = n18035 & n18038 ;
  assign n18040 = \wishbone_bd_ram_mem3_reg[36][25]/P0001  & n13639 ;
  assign n18041 = \wishbone_bd_ram_mem3_reg[55][25]/P0001  & n13618 ;
  assign n18042 = ~n18040 & ~n18041 ;
  assign n18043 = \wishbone_bd_ram_mem3_reg[106][25]/P0001  & n13555 ;
  assign n18044 = \wishbone_bd_ram_mem3_reg[143][25]/P0001  & n13461 ;
  assign n18045 = ~n18043 & ~n18044 ;
  assign n18046 = n18042 & n18045 ;
  assign n18047 = n18039 & n18046 ;
  assign n18048 = n18032 & n18047 ;
  assign n18049 = n18017 & n18048 ;
  assign n18050 = n17986 & n18049 ;
  assign n18051 = \wishbone_bd_ram_mem3_reg[38][25]/P0001  & n13828 ;
  assign n18052 = \wishbone_bd_ram_mem3_reg[229][25]/P0001  & n13552 ;
  assign n18053 = ~n18051 & ~n18052 ;
  assign n18054 = \wishbone_bd_ram_mem3_reg[126][25]/P0001  & n13786 ;
  assign n18055 = \wishbone_bd_ram_mem3_reg[86][25]/P0001  & n13485 ;
  assign n18056 = ~n18054 & ~n18055 ;
  assign n18057 = n18053 & n18056 ;
  assign n18058 = \wishbone_bd_ram_mem3_reg[130][25]/P0001  & n13427 ;
  assign n18059 = \wishbone_bd_ram_mem3_reg[124][25]/P0001  & n14024 ;
  assign n18060 = ~n18058 & ~n18059 ;
  assign n18061 = \wishbone_bd_ram_mem3_reg[0][25]/P0001  & n13539 ;
  assign n18062 = \wishbone_bd_ram_mem3_reg[5][25]/P0001  & n13243 ;
  assign n18063 = ~n18061 & ~n18062 ;
  assign n18064 = n18060 & n18063 ;
  assign n18065 = n18057 & n18064 ;
  assign n18066 = \wishbone_bd_ram_mem3_reg[195][25]/P0001  & n13700 ;
  assign n18067 = \wishbone_bd_ram_mem3_reg[251][25]/P0001  & n14019 ;
  assign n18068 = ~n18066 & ~n18067 ;
  assign n18069 = \wishbone_bd_ram_mem3_reg[159][25]/P0001  & n13627 ;
  assign n18070 = \wishbone_bd_ram_mem3_reg[199][25]/P0001  & n13499 ;
  assign n18071 = ~n18069 & ~n18070 ;
  assign n18072 = n18068 & n18071 ;
  assign n18073 = \wishbone_bd_ram_mem3_reg[152][25]/P0001  & n13912 ;
  assign n18074 = \wishbone_bd_ram_mem3_reg[230][25]/P0001  & n13994 ;
  assign n18075 = ~n18073 & ~n18074 ;
  assign n18076 = \wishbone_bd_ram_mem3_reg[164][25]/P0001  & n13236 ;
  assign n18077 = \wishbone_bd_ram_mem3_reg[109][25]/P0001  & n13306 ;
  assign n18078 = ~n18076 & ~n18077 ;
  assign n18079 = n18075 & n18078 ;
  assign n18080 = n18072 & n18079 ;
  assign n18081 = n18065 & n18080 ;
  assign n18082 = \wishbone_bd_ram_mem3_reg[57][25]/P0001  & n13731 ;
  assign n18083 = \wishbone_bd_ram_mem3_reg[179][25]/P0001  & n14035 ;
  assign n18084 = ~n18082 & ~n18083 ;
  assign n18085 = \wishbone_bd_ram_mem3_reg[160][25]/P0001  & n13271 ;
  assign n18086 = \wishbone_bd_ram_mem3_reg[169][25]/P0001  & n13541 ;
  assign n18087 = ~n18085 & ~n18086 ;
  assign n18088 = n18084 & n18087 ;
  assign n18089 = \wishbone_bd_ram_mem3_reg[17][25]/P0001  & n13324 ;
  assign n18090 = \wishbone_bd_ram_mem3_reg[235][25]/P0001  & n13518 ;
  assign n18091 = ~n18089 & ~n18090 ;
  assign n18092 = \wishbone_bd_ram_mem3_reg[141][25]/P0001  & n13852 ;
  assign n18093 = \wishbone_bd_ram_mem3_reg[49][25]/P0001  & n13929 ;
  assign n18094 = ~n18092 & ~n18093 ;
  assign n18095 = n18091 & n18094 ;
  assign n18096 = n18088 & n18095 ;
  assign n18097 = \wishbone_bd_ram_mem3_reg[12][25]/P0001  & n13733 ;
  assign n18098 = \wishbone_bd_ram_mem3_reg[237][25]/P0001  & n13924 ;
  assign n18099 = ~n18097 & ~n18098 ;
  assign n18100 = \wishbone_bd_ram_mem3_reg[68][25]/P0001  & n13379 ;
  assign n18101 = \wishbone_bd_ram_mem3_reg[19][25]/P0001  & n13886 ;
  assign n18102 = ~n18100 & ~n18101 ;
  assign n18103 = n18099 & n18102 ;
  assign n18104 = \wishbone_bd_ram_mem3_reg[13][25]/P0001  & n13844 ;
  assign n18105 = \wishbone_bd_ram_mem3_reg[214][25]/P0001  & n13938 ;
  assign n18106 = ~n18104 & ~n18105 ;
  assign n18107 = \wishbone_bd_ram_mem3_reg[156][25]/P0001  & n13769 ;
  assign n18108 = \wishbone_bd_ram_mem3_reg[167][25]/P0001  & n13940 ;
  assign n18109 = ~n18107 & ~n18108 ;
  assign n18110 = n18106 & n18109 ;
  assign n18111 = n18103 & n18110 ;
  assign n18112 = n18096 & n18111 ;
  assign n18113 = n18081 & n18112 ;
  assign n18114 = \wishbone_bd_ram_mem3_reg[225][25]/P0001  & n13719 ;
  assign n18115 = \wishbone_bd_ram_mem3_reg[22][25]/P0001  & n13744 ;
  assign n18116 = ~n18114 & ~n18115 ;
  assign n18117 = \wishbone_bd_ram_mem3_reg[203][25]/P0001  & n13816 ;
  assign n18118 = \wishbone_bd_ram_mem3_reg[209][25]/P0001  & n13689 ;
  assign n18119 = ~n18117 & ~n18118 ;
  assign n18120 = n18116 & n18119 ;
  assign n18121 = \wishbone_bd_ram_mem3_reg[161][25]/P0001  & n13505 ;
  assign n18122 = \wishbone_bd_ram_mem3_reg[184][25]/P0001  & n13960 ;
  assign n18123 = ~n18121 & ~n18122 ;
  assign n18124 = \wishbone_bd_ram_mem3_reg[89][25]/P0001  & n13910 ;
  assign n18125 = \wishbone_bd_ram_mem3_reg[26][25]/P0001  & n13521 ;
  assign n18126 = ~n18124 & ~n18125 ;
  assign n18127 = n18123 & n18126 ;
  assign n18128 = n18120 & n18127 ;
  assign n18129 = \wishbone_bd_ram_mem3_reg[240][25]/P0001  & n13352 ;
  assign n18130 = \wishbone_bd_ram_mem3_reg[84][25]/P0001  & n13385 ;
  assign n18131 = ~n18129 & ~n18130 ;
  assign n18132 = \wishbone_bd_ram_mem3_reg[198][25]/P0001  & n13592 ;
  assign n18133 = \wishbone_bd_ram_mem3_reg[197][25]/P0001  & n13594 ;
  assign n18134 = ~n18132 & ~n18133 ;
  assign n18135 = n18131 & n18134 ;
  assign n18136 = \wishbone_bd_ram_mem3_reg[192][25]/P0001  & n13390 ;
  assign n18137 = \wishbone_bd_ram_mem3_reg[215][25]/P0001  & n13901 ;
  assign n18138 = ~n18136 & ~n18137 ;
  assign n18139 = \wishbone_bd_ram_mem3_reg[137][25]/P0001  & n13808 ;
  assign n18140 = \wishbone_bd_ram_mem3_reg[117][25]/P0001  & n13557 ;
  assign n18141 = ~n18139 & ~n18140 ;
  assign n18142 = n18138 & n18141 ;
  assign n18143 = n18135 & n18142 ;
  assign n18144 = n18128 & n18143 ;
  assign n18145 = \wishbone_bd_ram_mem3_reg[43][25]/P0001  & n13761 ;
  assign n18146 = \wishbone_bd_ram_mem3_reg[48][25]/P0001  & n13917 ;
  assign n18147 = ~n18145 & ~n18146 ;
  assign n18148 = \wishbone_bd_ram_mem3_reg[75][25]/P0001  & n13605 ;
  assign n18149 = \wishbone_bd_ram_mem3_reg[142][25]/P0001  & n13448 ;
  assign n18150 = ~n18148 & ~n18149 ;
  assign n18151 = n18147 & n18150 ;
  assign n18152 = \wishbone_bd_ram_mem3_reg[63][25]/P0001  & n13327 ;
  assign n18153 = \wishbone_bd_ram_mem3_reg[201][25]/P0001  & n13600 ;
  assign n18154 = ~n18152 & ~n18153 ;
  assign n18155 = \wishbone_bd_ram_mem3_reg[76][25]/P0001  & n13831 ;
  assign n18156 = \wishbone_bd_ram_mem3_reg[134][25]/P0001  & n13494 ;
  assign n18157 = ~n18155 & ~n18156 ;
  assign n18158 = n18154 & n18157 ;
  assign n18159 = n18151 & n18158 ;
  assign n18160 = \wishbone_bd_ram_mem3_reg[224][25]/P0001  & n13433 ;
  assign n18161 = \wishbone_bd_ram_mem3_reg[35][25]/P0001  & n13523 ;
  assign n18162 = ~n18160 & ~n18161 ;
  assign n18163 = \wishbone_bd_ram_mem3_reg[31][25]/P0001  & n13758 ;
  assign n18164 = \wishbone_bd_ram_mem3_reg[187][25]/P0001  & n13756 ;
  assign n18165 = ~n18163 & ~n18164 ;
  assign n18166 = n18162 & n18165 ;
  assign n18167 = \wishbone_bd_ram_mem3_reg[236][25]/P0001  & n13480 ;
  assign n18168 = \wishbone_bd_ram_mem3_reg[238][25]/P0001  & n13819 ;
  assign n18169 = ~n18167 & ~n18168 ;
  assign n18170 = \wishbone_bd_ram_mem3_reg[174][25]/P0001  & n13899 ;
  assign n18171 = \wishbone_bd_ram_mem3_reg[62][25]/P0001  & n13529 ;
  assign n18172 = ~n18170 & ~n18171 ;
  assign n18173 = n18169 & n18172 ;
  assign n18174 = n18166 & n18173 ;
  assign n18175 = n18159 & n18174 ;
  assign n18176 = n18144 & n18175 ;
  assign n18177 = n18113 & n18176 ;
  assign n18178 = n18050 & n18177 ;
  assign n18179 = \wishbone_bd_ram_mem3_reg[171][25]/P0001  & n13422 ;
  assign n18180 = \wishbone_bd_ram_mem3_reg[255][25]/P0001  & n13952 ;
  assign n18181 = ~n18179 & ~n18180 ;
  assign n18182 = \wishbone_bd_ram_mem3_reg[45][25]/P0001  & n13420 ;
  assign n18183 = \wishbone_bd_ram_mem3_reg[226][25]/P0001  & n13668 ;
  assign n18184 = ~n18182 & ~n18183 ;
  assign n18185 = n18181 & n18184 ;
  assign n18186 = \wishbone_bd_ram_mem3_reg[135][25]/P0001  & n13672 ;
  assign n18187 = \wishbone_bd_ram_mem3_reg[2][25]/P0001  & n13975 ;
  assign n18188 = ~n18186 & ~n18187 ;
  assign n18189 = \wishbone_bd_ram_mem3_reg[248][25]/P0001  & n13647 ;
  assign n18190 = \wishbone_bd_ram_mem3_reg[87][25]/P0001  & n13691 ;
  assign n18191 = ~n18189 & ~n18190 ;
  assign n18192 = n18188 & n18191 ;
  assign n18193 = n18185 & n18192 ;
  assign n18194 = \wishbone_bd_ram_mem3_reg[148][25]/P0001  & n13868 ;
  assign n18195 = \wishbone_bd_ram_mem3_reg[95][25]/P0001  & n13317 ;
  assign n18196 = ~n18194 & ~n18195 ;
  assign n18197 = \wishbone_bd_ram_mem3_reg[113][25]/P0001  & n13882 ;
  assign n18198 = \wishbone_bd_ram_mem3_reg[150][25]/P0001  & n13666 ;
  assign n18199 = ~n18197 & ~n18198 ;
  assign n18200 = n18196 & n18199 ;
  assign n18201 = \wishbone_bd_ram_mem3_reg[119][25]/P0001  & n14033 ;
  assign n18202 = \wishbone_bd_ram_mem3_reg[88][25]/P0001  & n13347 ;
  assign n18203 = ~n18201 & ~n18202 ;
  assign n18204 = \wishbone_bd_ram_mem3_reg[82][25]/P0001  & n13374 ;
  assign n18205 = \wishbone_bd_ram_mem3_reg[155][25]/P0001  & n13738 ;
  assign n18206 = ~n18204 & ~n18205 ;
  assign n18207 = n18203 & n18206 ;
  assign n18208 = n18200 & n18207 ;
  assign n18209 = n18193 & n18208 ;
  assign n18210 = \wishbone_bd_ram_mem3_reg[208][25]/P0001  & n14010 ;
  assign n18211 = \wishbone_bd_ram_mem3_reg[66][25]/P0001  & n13603 ;
  assign n18212 = ~n18210 & ~n18211 ;
  assign n18213 = \wishbone_bd_ram_mem3_reg[30][25]/P0001  & n13713 ;
  assign n18214 = \wishbone_bd_ram_mem3_reg[40][25]/P0001  & n13661 ;
  assign n18215 = ~n18213 & ~n18214 ;
  assign n18216 = n18212 & n18215 ;
  assign n18217 = \wishbone_bd_ram_mem3_reg[239][25]/P0001  & n13349 ;
  assign n18218 = \wishbone_bd_ram_mem3_reg[46][25]/P0001  & n13298 ;
  assign n18219 = ~n18217 & ~n18218 ;
  assign n18220 = \wishbone_bd_ram_mem3_reg[99][25]/P0001  & n13996 ;
  assign n18221 = \wishbone_bd_ram_mem3_reg[54][25]/P0001  & n13622 ;
  assign n18222 = ~n18220 & ~n18221 ;
  assign n18223 = n18219 & n18222 ;
  assign n18224 = n18216 & n18223 ;
  assign n18225 = \wishbone_bd_ram_mem3_reg[9][25]/P0001  & n13580 ;
  assign n18226 = \wishbone_bd_ram_mem3_reg[65][25]/P0001  & n13842 ;
  assign n18227 = ~n18225 & ~n18226 ;
  assign n18228 = \wishbone_bd_ram_mem3_reg[25][25]/P0001  & n13742 ;
  assign n18229 = \wishbone_bd_ram_mem3_reg[6][25]/P0001  & n13915 ;
  assign n18230 = ~n18228 & ~n18229 ;
  assign n18231 = n18227 & n18230 ;
  assign n18232 = \wishbone_bd_ram_mem3_reg[83][25]/P0001  & n13454 ;
  assign n18233 = \wishbone_bd_ram_mem3_reg[139][25]/P0001  & n13566 ;
  assign n18234 = ~n18232 & ~n18233 ;
  assign n18235 = \wishbone_bd_ram_mem3_reg[115][25]/P0001  & n13747 ;
  assign n18236 = \wishbone_bd_ram_mem3_reg[158][25]/P0001  & n13294 ;
  assign n18237 = ~n18235 & ~n18236 ;
  assign n18238 = n18234 & n18237 ;
  assign n18239 = n18231 & n18238 ;
  assign n18240 = n18224 & n18239 ;
  assign n18241 = n18209 & n18240 ;
  assign n18242 = \wishbone_bd_ram_mem3_reg[178][25]/P0001  & n13301 ;
  assign n18243 = \wishbone_bd_ram_mem3_reg[14][25]/P0001  & n13972 ;
  assign n18244 = ~n18242 & ~n18243 ;
  assign n18245 = \wishbone_bd_ram_mem3_reg[204][25]/P0001  & n13821 ;
  assign n18246 = \wishbone_bd_ram_mem3_reg[118][25]/P0001  & n13589 ;
  assign n18247 = ~n18245 & ~n18246 ;
  assign n18248 = n18244 & n18247 ;
  assign n18249 = \wishbone_bd_ram_mem3_reg[181][25]/P0001  & n13587 ;
  assign n18250 = \wishbone_bd_ram_mem3_reg[193][25]/P0001  & n14022 ;
  assign n18251 = ~n18249 & ~n18250 ;
  assign n18252 = \wishbone_bd_ram_mem3_reg[28][25]/P0001  & n13810 ;
  assign n18253 = \wishbone_bd_ram_mem3_reg[210][25]/P0001  & n13443 ;
  assign n18254 = ~n18252 & ~n18253 ;
  assign n18255 = n18251 & n18254 ;
  assign n18256 = n18248 & n18255 ;
  assign n18257 = \wishbone_bd_ram_mem3_reg[27][25]/P0001  & n13251 ;
  assign n18258 = \wishbone_bd_ram_mem3_reg[129][25]/P0001  & n13629 ;
  assign n18259 = ~n18257 & ~n18258 ;
  assign n18260 = \wishbone_bd_ram_mem3_reg[20][25]/P0001  & n13839 ;
  assign n18261 = \wishbone_bd_ram_mem3_reg[200][25]/P0001  & n13922 ;
  assign n18262 = ~n18260 & ~n18261 ;
  assign n18263 = n18259 & n18262 ;
  assign n18264 = \wishbone_bd_ram_mem3_reg[67][25]/P0001  & n13663 ;
  assign n18265 = \wishbone_bd_ram_mem3_reg[10][25]/P0001  & n13837 ;
  assign n18266 = ~n18264 & ~n18265 ;
  assign n18267 = \wishbone_bd_ram_mem3_reg[123][25]/P0001  & n13749 ;
  assign n18268 = \wishbone_bd_ram_mem3_reg[207][25]/P0001  & n13826 ;
  assign n18269 = ~n18267 & ~n18268 ;
  assign n18270 = n18266 & n18269 ;
  assign n18271 = n18263 & n18270 ;
  assign n18272 = n18256 & n18271 ;
  assign n18273 = \wishbone_bd_ram_mem3_reg[104][25]/P0001  & n13684 ;
  assign n18274 = \wishbone_bd_ram_mem3_reg[212][25]/P0001  & n13634 ;
  assign n18275 = ~n18273 & ~n18274 ;
  assign n18276 = \wishbone_bd_ram_mem3_reg[92][25]/P0001  & n13859 ;
  assign n18277 = \wishbone_bd_ram_mem3_reg[91][25]/P0001  & n13954 ;
  assign n18278 = ~n18276 & ~n18277 ;
  assign n18279 = n18275 & n18278 ;
  assign n18280 = \wishbone_bd_ram_mem3_reg[102][25]/P0001  & n13534 ;
  assign n18281 = \wishbone_bd_ram_mem3_reg[173][25]/P0001  & n13360 ;
  assign n18282 = ~n18280 & ~n18281 ;
  assign n18283 = \wishbone_bd_ram_mem3_reg[216][25]/P0001  & n14005 ;
  assign n18284 = \wishbone_bd_ram_mem3_reg[246][25]/P0001  & n13981 ;
  assign n18285 = ~n18283 & ~n18284 ;
  assign n18286 = n18282 & n18285 ;
  assign n18287 = n18279 & n18286 ;
  assign n18288 = \wishbone_bd_ram_mem3_reg[245][25]/P0001  & n13877 ;
  assign n18289 = \wishbone_bd_ram_mem3_reg[56][25]/P0001  & n13611 ;
  assign n18290 = ~n18288 & ~n18289 ;
  assign n18291 = \wishbone_bd_ram_mem3_reg[15][25]/P0001  & n13797 ;
  assign n18292 = \wishbone_bd_ram_mem3_reg[132][25]/P0001  & n13927 ;
  assign n18293 = ~n18291 & ~n18292 ;
  assign n18294 = n18290 & n18293 ;
  assign n18295 = \wishbone_bd_ram_mem3_reg[188][25]/P0001  & n13407 ;
  assign n18296 = \wishbone_bd_ram_mem3_reg[107][25]/P0001  & n13476 ;
  assign n18297 = ~n18295 & ~n18296 ;
  assign n18298 = \wishbone_bd_ram_mem3_reg[18][25]/P0001  & n13532 ;
  assign n18299 = \wishbone_bd_ram_mem3_reg[120][25]/P0001  & n13550 ;
  assign n18300 = ~n18298 & ~n18299 ;
  assign n18301 = n18297 & n18300 ;
  assign n18302 = n18294 & n18301 ;
  assign n18303 = n18287 & n18302 ;
  assign n18304 = n18272 & n18303 ;
  assign n18305 = n18241 & n18304 ;
  assign n18306 = \wishbone_bd_ram_mem3_reg[78][25]/P0001  & n13277 ;
  assign n18307 = \wishbone_bd_ram_mem3_reg[162][25]/P0001  & n13726 ;
  assign n18308 = ~n18306 & ~n18307 ;
  assign n18309 = \wishbone_bd_ram_mem3_reg[138][25]/P0001  & n13398 ;
  assign n18310 = \wishbone_bd_ram_mem3_reg[41][25]/P0001  & n14017 ;
  assign n18311 = ~n18309 & ~n18310 ;
  assign n18312 = n18308 & n18311 ;
  assign n18313 = \wishbone_bd_ram_mem3_reg[80][25]/P0001  & n13516 ;
  assign n18314 = \wishbone_bd_ram_mem3_reg[116][25]/P0001  & n13865 ;
  assign n18315 = ~n18313 & ~n18314 ;
  assign n18316 = \wishbone_bd_ram_mem3_reg[131][25]/P0001  & n13358 ;
  assign n18317 = \wishbone_bd_ram_mem3_reg[249][25]/P0001  & n13431 ;
  assign n18318 = ~n18316 & ~n18317 ;
  assign n18319 = n18315 & n18318 ;
  assign n18320 = n18312 & n18319 ;
  assign n18321 = \wishbone_bd_ram_mem3_reg[147][25]/P0001  & n13702 ;
  assign n18322 = \wishbone_bd_ram_mem3_reg[133][25]/P0001  & n13492 ;
  assign n18323 = ~n18321 & ~n18322 ;
  assign n18324 = \wishbone_bd_ram_mem3_reg[97][25]/P0001  & n13724 ;
  assign n18325 = \wishbone_bd_ram_mem3_reg[114][25]/P0001  & n13763 ;
  assign n18326 = ~n18324 & ~n18325 ;
  assign n18327 = n18323 & n18326 ;
  assign n18328 = \wishbone_bd_ram_mem3_reg[73][25]/P0001  & n13456 ;
  assign n18329 = \wishbone_bd_ram_mem3_reg[58][25]/P0001  & n13949 ;
  assign n18330 = ~n18328 & ~n18329 ;
  assign n18331 = \wishbone_bd_ram_mem3_reg[7][25]/P0001  & n13546 ;
  assign n18332 = \wishbone_bd_ram_mem3_reg[151][25]/P0001  & n13697 ;
  assign n18333 = ~n18331 & ~n18332 ;
  assign n18334 = n18330 & n18333 ;
  assign n18335 = n18327 & n18334 ;
  assign n18336 = n18320 & n18335 ;
  assign n18337 = \wishbone_bd_ram_mem3_reg[145][25]/P0001  & n13715 ;
  assign n18338 = \wishbone_bd_ram_mem3_reg[11][25]/P0001  & n13774 ;
  assign n18339 = ~n18337 & ~n18338 ;
  assign n18340 = \wishbone_bd_ram_mem3_reg[21][25]/P0001  & n13438 ;
  assign n18341 = \wishbone_bd_ram_mem3_reg[121][25]/P0001  & n13983 ;
  assign n18342 = ~n18340 & ~n18341 ;
  assign n18343 = n18339 & n18342 ;
  assign n18344 = \wishbone_bd_ram_mem3_reg[125][25]/P0001  & n13396 ;
  assign n18345 = \wishbone_bd_ram_mem3_reg[44][25]/P0001  & n13291 ;
  assign n18346 = ~n18344 & ~n18345 ;
  assign n18347 = \wishbone_bd_ram_mem3_reg[70][25]/P0001  & n13339 ;
  assign n18348 = \wishbone_bd_ram_mem3_reg[206][25]/P0001  & n13414 ;
  assign n18349 = ~n18347 & ~n18348 ;
  assign n18350 = n18346 & n18349 ;
  assign n18351 = n18343 & n18350 ;
  assign n18352 = \wishbone_bd_ram_mem3_reg[170][25]/P0001  & n14007 ;
  assign n18353 = \wishbone_bd_ram_mem3_reg[71][25]/P0001  & n13636 ;
  assign n18354 = ~n18352 & ~n18353 ;
  assign n18355 = \wishbone_bd_ram_mem3_reg[186][25]/P0001  & n13616 ;
  assign n18356 = \wishbone_bd_ram_mem3_reg[37][25]/P0001  & n13710 ;
  assign n18357 = ~n18355 & ~n18356 ;
  assign n18358 = n18354 & n18357 ;
  assign n18359 = \wishbone_bd_ram_mem3_reg[4][25]/P0001  & n13527 ;
  assign n18360 = \wishbone_bd_ram_mem3_reg[33][25]/P0001  & n13933 ;
  assign n18361 = ~n18359 & ~n18360 ;
  assign n18362 = \wishbone_bd_ram_mem3_reg[221][25]/P0001  & n13641 ;
  assign n18363 = \wishbone_bd_ram_mem3_reg[168][25]/P0001  & n13795 ;
  assign n18364 = ~n18362 & ~n18363 ;
  assign n18365 = n18361 & n18364 ;
  assign n18366 = n18358 & n18365 ;
  assign n18367 = n18351 & n18366 ;
  assign n18368 = n18336 & n18367 ;
  assign n18369 = \wishbone_bd_ram_mem3_reg[247][25]/P0001  & n13571 ;
  assign n18370 = \wishbone_bd_ram_mem3_reg[103][25]/P0001  & n13320 ;
  assign n18371 = ~n18369 & ~n18370 ;
  assign n18372 = \wishbone_bd_ram_mem3_reg[223][25]/P0001  & n13335 ;
  assign n18373 = \wishbone_bd_ram_mem3_reg[228][25]/P0001  & n13497 ;
  assign n18374 = ~n18372 & ~n18373 ;
  assign n18375 = n18371 & n18374 ;
  assign n18376 = \wishbone_bd_ram_mem3_reg[72][25]/P0001  & n13582 ;
  assign n18377 = \wishbone_bd_ram_mem3_reg[182][25]/P0001  & n13598 ;
  assign n18378 = ~n18376 & ~n18377 ;
  assign n18379 = \wishbone_bd_ram_mem3_reg[136][25]/P0001  & n13963 ;
  assign n18380 = \wishbone_bd_ram_mem3_reg[185][25]/P0001  & n13372 ;
  assign n18381 = ~n18379 & ~n18380 ;
  assign n18382 = n18378 & n18381 ;
  assign n18383 = n18375 & n18382 ;
  assign n18384 = \wishbone_bd_ram_mem3_reg[8][25]/P0001  & n13459 ;
  assign n18385 = \wishbone_bd_ram_mem3_reg[219][25]/P0001  & n13577 ;
  assign n18386 = ~n18384 & ~n18385 ;
  assign n18387 = \wishbone_bd_ram_mem3_reg[180][25]/P0001  & n13650 ;
  assign n18388 = \wishbone_bd_ram_mem3_reg[23][25]/P0001  & n13857 ;
  assign n18389 = ~n18387 & ~n18388 ;
  assign n18390 = n18386 & n18389 ;
  assign n18391 = \wishbone_bd_ram_mem3_reg[254][25]/P0001  & n13283 ;
  assign n18392 = \wishbone_bd_ram_mem3_reg[146][25]/P0001  & n13958 ;
  assign n18393 = ~n18391 & ~n18392 ;
  assign n18394 = \wishbone_bd_ram_mem3_reg[233][25]/P0001  & n13332 ;
  assign n18395 = \wishbone_bd_ram_mem3_reg[69][25]/P0001  & n13487 ;
  assign n18396 = ~n18394 & ~n18395 ;
  assign n18397 = n18393 & n18396 ;
  assign n18398 = n18390 & n18397 ;
  assign n18399 = n18383 & n18398 ;
  assign n18400 = \wishbone_bd_ram_mem3_reg[42][25]/P0001  & n13341 ;
  assign n18401 = \wishbone_bd_ram_mem3_reg[163][25]/P0001  & n13255 ;
  assign n18402 = ~n18400 & ~n18401 ;
  assign n18403 = \wishbone_bd_ram_mem3_reg[231][25]/P0001  & n13363 ;
  assign n18404 = \wishbone_bd_ram_mem3_reg[16][25]/P0001  & n13695 ;
  assign n18405 = ~n18403 & ~n18404 ;
  assign n18406 = n18402 & n18405 ;
  assign n18407 = \wishbone_bd_ram_mem3_reg[250][25]/P0001  & n13677 ;
  assign n18408 = \wishbone_bd_ram_mem3_reg[244][25]/P0001  & n13474 ;
  assign n18409 = ~n18407 & ~n18408 ;
  assign n18410 = \wishbone_bd_ram_mem3_reg[232][25]/P0001  & n13510 ;
  assign n18411 = \wishbone_bd_ram_mem3_reg[175][25]/P0001  & n13674 ;
  assign n18412 = ~n18410 & ~n18411 ;
  assign n18413 = n18409 & n18412 ;
  assign n18414 = n18406 & n18413 ;
  assign n18415 = \wishbone_bd_ram_mem3_reg[32][25]/P0001  & n13736 ;
  assign n18416 = \wishbone_bd_ram_mem3_reg[194][25]/P0001  & n13624 ;
  assign n18417 = ~n18415 & ~n18416 ;
  assign n18418 = \wishbone_bd_ram_mem3_reg[241][25]/P0001  & n13854 ;
  assign n18419 = \wishbone_bd_ram_mem3_reg[53][25]/P0001  & n13875 ;
  assign n18420 = ~n18418 & ~n18419 ;
  assign n18421 = n18417 & n18420 ;
  assign n18422 = \wishbone_bd_ram_mem3_reg[218][25]/P0001  & n13792 ;
  assign n18423 = \wishbone_bd_ram_mem3_reg[111][25]/P0001  & n13471 ;
  assign n18424 = ~n18422 & ~n18423 ;
  assign n18425 = \wishbone_bd_ram_mem3_reg[189][25]/P0001  & n14001 ;
  assign n18426 = \wishbone_bd_ram_mem3_reg[191][25]/P0001  & n14012 ;
  assign n18427 = ~n18425 & ~n18426 ;
  assign n18428 = n18424 & n18427 ;
  assign n18429 = n18421 & n18428 ;
  assign n18430 = n18414 & n18429 ;
  assign n18431 = n18399 & n18430 ;
  assign n18432 = n18368 & n18431 ;
  assign n18433 = n18305 & n18432 ;
  assign n18434 = n18178 & n18433 ;
  assign n18435 = n14047 & ~n18434 ;
  assign n18436 = \wishbone_TxLength_reg[9]/NET0131  & n14052 ;
  assign n18437 = n14057 & n18436 ;
  assign n18438 = ~n17918 & n18437 ;
  assign n18439 = ~\wishbone_TxLength_reg[9]/NET0131  & ~n14057 ;
  assign n18440 = ~\wishbone_TxLength_reg[9]/NET0131  & ~n14052 ;
  assign n18441 = ~n18439 & ~n18440 ;
  assign n18442 = ~n18438 & n18441 ;
  assign n18443 = ~\wishbone_TxLength_reg[9]/NET0131  & n17918 ;
  assign n18444 = n14046 & ~n14595 ;
  assign n18445 = n14063 & ~n14595 ;
  assign n18446 = n14058 & n18445 ;
  assign n18447 = ~n18444 & ~n18446 ;
  assign n18448 = ~n18443 & n18447 ;
  assign n18449 = n18442 & n18448 ;
  assign n18450 = ~n18435 & ~n18449 ;
  assign n18451 = \wishbone_RxDataLatched2_reg[0]/NET0131  & ~n15737 ;
  assign n18452 = n15735 & n18451 ;
  assign n18453 = \rxethmac1_RxData_reg[0]/NET0131  & n15740 ;
  assign n18454 = \rxethmac1_RxData_reg[0]/NET0131  & n15741 ;
  assign n18455 = ~n15745 & n18454 ;
  assign n18456 = ~n18453 & ~n18455 ;
  assign n18457 = ~n18452 & n18456 ;
  assign n18458 = \wishbone_RxDataLatched2_reg[1]/NET0131  & ~n15737 ;
  assign n18459 = n15735 & n18458 ;
  assign n18460 = \rxethmac1_RxData_reg[1]/NET0131  & n15740 ;
  assign n18461 = \rxethmac1_RxData_reg[1]/NET0131  & n15741 ;
  assign n18462 = ~n15745 & n18461 ;
  assign n18463 = ~n18460 & ~n18462 ;
  assign n18464 = ~n18459 & n18463 ;
  assign n18465 = \wishbone_RxDataLatched2_reg[2]/NET0131  & ~n15737 ;
  assign n18466 = n15735 & n18465 ;
  assign n18467 = \rxethmac1_RxData_reg[2]/NET0131  & n15740 ;
  assign n18468 = \rxethmac1_RxData_reg[2]/NET0131  & n15741 ;
  assign n18469 = ~n15745 & n18468 ;
  assign n18470 = ~n18467 & ~n18469 ;
  assign n18471 = ~n18466 & n18470 ;
  assign n18472 = \wishbone_RxDataLatched2_reg[3]/NET0131  & ~n15737 ;
  assign n18473 = n15735 & n18472 ;
  assign n18474 = \rxethmac1_RxData_reg[3]/NET0131  & n15740 ;
  assign n18475 = \rxethmac1_RxData_reg[3]/NET0131  & n15741 ;
  assign n18476 = ~n15745 & n18475 ;
  assign n18477 = ~n18474 & ~n18476 ;
  assign n18478 = ~n18473 & n18477 ;
  assign n18479 = \wishbone_RxDataLatched2_reg[5]/NET0131  & ~n15737 ;
  assign n18480 = n15735 & n18479 ;
  assign n18481 = \rxethmac1_RxData_reg[5]/NET0131  & n15740 ;
  assign n18482 = \rxethmac1_RxData_reg[5]/NET0131  & n15741 ;
  assign n18483 = ~n15745 & n18482 ;
  assign n18484 = ~n18481 & ~n18483 ;
  assign n18485 = ~n18480 & n18484 ;
  assign n18486 = \wishbone_RxDataLatched2_reg[4]/NET0131  & ~n15737 ;
  assign n18487 = n15735 & n18486 ;
  assign n18488 = \rxethmac1_RxData_reg[4]/NET0131  & n15740 ;
  assign n18489 = \rxethmac1_RxData_reg[4]/NET0131  & n15741 ;
  assign n18490 = ~n15745 & n18489 ;
  assign n18491 = ~n18488 & ~n18490 ;
  assign n18492 = ~n18487 & n18491 ;
  assign n18493 = \wishbone_RxDataLatched2_reg[6]/NET0131  & ~n15737 ;
  assign n18494 = n15735 & n18493 ;
  assign n18495 = \rxethmac1_RxData_reg[6]/NET0131  & n15740 ;
  assign n18496 = \rxethmac1_RxData_reg[6]/NET0131  & n15741 ;
  assign n18497 = ~n15745 & n18496 ;
  assign n18498 = ~n18495 & ~n18497 ;
  assign n18499 = ~n18494 & n18498 ;
  assign n18500 = \wishbone_RxDataLatched2_reg[7]/NET0131  & ~n15737 ;
  assign n18501 = n15735 & n18500 ;
  assign n18502 = \rxethmac1_RxData_reg[7]/NET0131  & n15740 ;
  assign n18503 = \rxethmac1_RxData_reg[7]/NET0131  & n15741 ;
  assign n18504 = ~n15745 & n18503 ;
  assign n18505 = ~n18502 & ~n18504 ;
  assign n18506 = ~n18501 & n18505 ;
  assign n18507 = ~wb_rst_i_pad & n16305 ;
  assign n18508 = ~n15114 & n18507 ;
  assign n18509 = \wishbone_RxPointerMSB_reg[2]/NET0131  & \wishbone_RxPointerMSB_reg[3]/NET0131  ;
  assign n18510 = n16307 & n18509 ;
  assign n18511 = \wishbone_RxPointerMSB_reg[4]/NET0131  & \wishbone_RxPointerMSB_reg[6]/NET0131  ;
  assign n18512 = \wishbone_RxPointerMSB_reg[5]/NET0131  & n18511 ;
  assign n18513 = n18510 & n18512 ;
  assign n18514 = \wishbone_RxPointerMSB_reg[8]/NET0131  & \wishbone_RxPointerMSB_reg[9]/NET0131  ;
  assign n18515 = \wishbone_RxPointerMSB_reg[10]/NET0131  & \wishbone_RxPointerMSB_reg[7]/NET0131  ;
  assign n18516 = n18514 & n18515 ;
  assign n18517 = n18513 & n18516 ;
  assign n18518 = \wishbone_RxPointerMSB_reg[12]/NET0131  & \wishbone_RxPointerMSB_reg[13]/NET0131  ;
  assign n18519 = \wishbone_RxPointerMSB_reg[11]/NET0131  & \wishbone_RxPointerMSB_reg[14]/NET0131  ;
  assign n18520 = n18518 & n18519 ;
  assign n18521 = n18517 & n18520 ;
  assign n18522 = \wishbone_RxPointerMSB_reg[16]/NET0131  & \wishbone_RxPointerMSB_reg[17]/NET0131  ;
  assign n18523 = \wishbone_RxPointerMSB_reg[18]/NET0131  & \wishbone_RxPointerMSB_reg[19]/NET0131  ;
  assign n18524 = n18522 & n18523 ;
  assign n18525 = \wishbone_RxPointerMSB_reg[15]/NET0131  & \wishbone_RxPointerMSB_reg[20]/NET0131  ;
  assign n18526 = n18524 & n18525 ;
  assign n18527 = n18521 & n18526 ;
  assign n18528 = \wishbone_RxPointerMSB_reg[21]/NET0131  & \wishbone_RxPointerMSB_reg[22]/NET0131  ;
  assign n18529 = \wishbone_RxPointerMSB_reg[23]/NET0131  & \wishbone_RxPointerMSB_reg[24]/NET0131  ;
  assign n18530 = n18528 & n18529 ;
  assign n18531 = n18527 & n18530 ;
  assign n18532 = \wishbone_RxPointerMSB_reg[26]/NET0131  & \wishbone_RxPointerMSB_reg[27]/NET0131  ;
  assign n18533 = \wishbone_RxPointerMSB_reg[28]/NET0131  & n18532 ;
  assign n18534 = \wishbone_RxPointerMSB_reg[25]/NET0131  & \wishbone_RxPointerMSB_reg[29]/NET0131  ;
  assign n18535 = n18533 & n18534 ;
  assign n18536 = n18531 & n18535 ;
  assign n18537 = ~\wishbone_RxPointerMSB_reg[30]/NET0131  & ~n18536 ;
  assign n18538 = \wishbone_RxPointerMSB_reg[29]/NET0131  & \wishbone_RxPointerMSB_reg[30]/NET0131  ;
  assign n18539 = \wishbone_RxPointerMSB_reg[25]/NET0131  & n18538 ;
  assign n18540 = n18533 & n18539 ;
  assign n18541 = n18531 & n18540 ;
  assign n18542 = ~n16305 & ~n18541 ;
  assign n18543 = ~n18537 & n18542 ;
  assign n18544 = ~n18508 & ~n18543 ;
  assign n18545 = \wishbone_TxPointerRead_reg/NET0131  & n14045 ;
  assign n18546 = ~\wishbone_BlockingIncrementTxPointer_reg/NET0131  & \wishbone_IncrTxPointer_reg/NET0131  ;
  assign n18547 = \wishbone_TxPointerMSB_reg[2]/NET0131  & \wishbone_TxPointerMSB_reg[3]/NET0131  ;
  assign n18548 = n18546 & n18547 ;
  assign n18549 = \wishbone_TxPointerMSB_reg[4]/NET0131  & \wishbone_TxPointerMSB_reg[6]/NET0131  ;
  assign n18550 = \wishbone_TxPointerMSB_reg[5]/NET0131  & n18549 ;
  assign n18551 = n18548 & n18550 ;
  assign n18552 = \wishbone_TxPointerMSB_reg[7]/NET0131  & \wishbone_TxPointerMSB_reg[9]/NET0131  ;
  assign n18553 = \wishbone_TxPointerMSB_reg[8]/NET0131  & n18552 ;
  assign n18554 = n18551 & n18553 ;
  assign n18555 = \wishbone_TxPointerMSB_reg[10]/NET0131  & \wishbone_TxPointerMSB_reg[12]/NET0131  ;
  assign n18556 = \wishbone_TxPointerMSB_reg[11]/NET0131  & n18555 ;
  assign n18557 = n18554 & n18556 ;
  assign n18558 = \wishbone_TxPointerMSB_reg[15]/NET0131  & \wishbone_TxPointerMSB_reg[16]/NET0131  ;
  assign n18559 = \wishbone_TxPointerMSB_reg[13]/NET0131  & \wishbone_TxPointerMSB_reg[14]/NET0131  ;
  assign n18560 = \wishbone_TxPointerMSB_reg[17]/NET0131  & n18559 ;
  assign n18561 = n18558 & n18560 ;
  assign n18562 = n18557 & n18561 ;
  assign n18563 = \wishbone_TxPointerMSB_reg[19]/NET0131  & \wishbone_TxPointerMSB_reg[20]/NET0131  ;
  assign n18564 = \wishbone_TxPointerMSB_reg[18]/NET0131  & n18563 ;
  assign n18565 = \wishbone_TxPointerMSB_reg[21]/NET0131  & \wishbone_TxPointerMSB_reg[22]/NET0131  ;
  assign n18566 = n18564 & n18565 ;
  assign n18567 = n18562 & n18566 ;
  assign n18568 = \wishbone_TxPointerMSB_reg[25]/NET0131  & \wishbone_TxPointerMSB_reg[26]/NET0131  ;
  assign n18569 = \wishbone_TxPointerMSB_reg[27]/NET0131  & \wishbone_TxPointerMSB_reg[28]/NET0131  ;
  assign n18570 = \wishbone_TxPointerMSB_reg[23]/NET0131  & \wishbone_TxPointerMSB_reg[24]/NET0131  ;
  assign n18571 = n18569 & n18570 ;
  assign n18572 = n18568 & n18571 ;
  assign n18573 = n18567 & n18572 ;
  assign n18574 = \wishbone_TxPointerMSB_reg[29]/NET0131  & \wishbone_TxPointerMSB_reg[30]/NET0131  ;
  assign n18575 = ~\wishbone_TxPointerMSB_reg[29]/NET0131  & ~\wishbone_TxPointerMSB_reg[30]/NET0131  ;
  assign n18576 = ~n18574 & ~n18575 ;
  assign n18577 = ~n18545 & ~n18576 ;
  assign n18578 = n18573 & n18577 ;
  assign n18579 = ~\wishbone_TxPointerMSB_reg[30]/NET0131  & ~n18545 ;
  assign n18580 = ~n18573 & n18579 ;
  assign n18581 = ~n18578 & ~n18580 ;
  assign n18582 = ~n18545 & n18581 ;
  assign n18583 = ~wb_rst_i_pad & n18581 ;
  assign n18584 = ~n15114 & n18583 ;
  assign n18585 = ~n18582 & ~n18584 ;
  assign n18586 = \wishbone_RxDataLatched2_reg[16]/NET0131  & ~n15737 ;
  assign n18587 = n15735 & n18586 ;
  assign n18588 = \wishbone_RxValidBytes_reg[0]/NET0131  & ~\wishbone_RxValidBytes_reg[1]/NET0131  ;
  assign n18589 = \wishbone_ShiftWillEnd_reg/NET0131  & n18588 ;
  assign n18590 = \wishbone_RxDataLatched1_reg[16]/NET0131  & ~n18589 ;
  assign n18591 = ~n15745 & n18590 ;
  assign n18592 = ~n18587 & ~n18591 ;
  assign n18593 = \wishbone_RxDataLatched2_reg[17]/NET0131  & ~n15737 ;
  assign n18594 = n15735 & n18593 ;
  assign n18595 = \wishbone_RxDataLatched1_reg[17]/NET0131  & ~n18589 ;
  assign n18596 = ~n15745 & n18595 ;
  assign n18597 = ~n18594 & ~n18596 ;
  assign n18598 = \wishbone_RxDataLatched2_reg[18]/NET0131  & ~n15737 ;
  assign n18599 = n15735 & n18598 ;
  assign n18600 = \wishbone_RxDataLatched1_reg[18]/NET0131  & ~n18589 ;
  assign n18601 = ~n15745 & n18600 ;
  assign n18602 = ~n18599 & ~n18601 ;
  assign n18603 = \wishbone_RxDataLatched2_reg[19]/NET0131  & ~n15737 ;
  assign n18604 = n15735 & n18603 ;
  assign n18605 = \wishbone_RxDataLatched1_reg[19]/NET0131  & ~n18589 ;
  assign n18606 = ~n15745 & n18605 ;
  assign n18607 = ~n18604 & ~n18606 ;
  assign n18608 = \wishbone_RxDataLatched2_reg[20]/NET0131  & ~n15737 ;
  assign n18609 = n15735 & n18608 ;
  assign n18610 = \wishbone_RxDataLatched1_reg[20]/NET0131  & ~n18589 ;
  assign n18611 = ~n15745 & n18610 ;
  assign n18612 = ~n18609 & ~n18611 ;
  assign n18613 = \wishbone_RxDataLatched2_reg[21]/NET0131  & ~n15737 ;
  assign n18614 = n15735 & n18613 ;
  assign n18615 = \wishbone_RxDataLatched1_reg[21]/NET0131  & ~n18589 ;
  assign n18616 = ~n15745 & n18615 ;
  assign n18617 = ~n18614 & ~n18616 ;
  assign n18618 = \wishbone_RxDataLatched2_reg[22]/NET0131  & ~n15737 ;
  assign n18619 = n15735 & n18618 ;
  assign n18620 = \wishbone_RxDataLatched1_reg[22]/NET0131  & ~n18589 ;
  assign n18621 = ~n15745 & n18620 ;
  assign n18622 = ~n18619 & ~n18621 ;
  assign n18623 = \wishbone_RxDataLatched2_reg[23]/NET0131  & ~n15737 ;
  assign n18624 = n15735 & n18623 ;
  assign n18625 = \wishbone_RxDataLatched1_reg[23]/NET0131  & ~n18589 ;
  assign n18626 = ~n15745 & n18625 ;
  assign n18627 = ~n18624 & ~n18626 ;
  assign n18628 = ~\wishbone_RxPointerMSB_reg[13]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n18629 = n13144 & n18628 ;
  assign n18630 = ~n13149 & ~n18629 ;
  assign n18631 = n13143 & n18630 ;
  assign n18632 = n13137 & n18631 ;
  assign n18633 = ~n13170 & ~n18632 ;
  assign n18634 = \m_wb_adr_o[12]_pad  & \m_wb_adr_o[13]_pad  ;
  assign n18635 = n13103 & n18634 ;
  assign n18636 = \m_wb_adr_o[12]_pad  & n13103 ;
  assign n18637 = ~\m_wb_adr_o[13]_pad  & ~n18636 ;
  assign n18638 = ~n18635 & ~n18637 ;
  assign n18639 = ~n18633 & n18638 ;
  assign n18640 = \m_wb_adr_o[13]_pad  & n13197 ;
  assign n18641 = \wishbone_TxPointerMSB_reg[13]/NET0131  & ~n13201 ;
  assign n18642 = \wishbone_RxPointerMSB_reg[13]/NET0131  & n13207 ;
  assign n18643 = ~n13196 & n18642 ;
  assign n18644 = ~n18641 & ~n18643 ;
  assign n18645 = ~n18640 & n18644 ;
  assign n18646 = ~n18639 & n18645 ;
  assign n18647 = \m_wb_adr_o[12]_pad  & n13104 ;
  assign n18648 = n13103 & n18647 ;
  assign n18649 = ~\m_wb_adr_o[14]_pad  & ~n18635 ;
  assign n18650 = ~n18648 & ~n18649 ;
  assign n18651 = ~n15177 & n18650 ;
  assign n18652 = \m_wb_adr_o[14]_pad  & n13197 ;
  assign n18653 = ~n18651 & ~n18652 ;
  assign n18654 = ~n13168 & n13188 ;
  assign n18655 = ~n18650 & n18654 ;
  assign n18656 = \wishbone_TxPointerMSB_reg[14]/NET0131  & ~n13189 ;
  assign n18657 = ~n18655 & n18656 ;
  assign n18658 = ~n13207 & ~n18650 ;
  assign n18659 = \wishbone_RxPointerMSB_reg[14]/NET0131  & ~n13196 ;
  assign n18660 = ~n18658 & n18659 ;
  assign n18661 = ~n18657 & ~n18660 ;
  assign n18662 = n18653 & n18661 ;
  assign n18663 = \m_wb_adr_o[8]_pad  & n13197 ;
  assign n18664 = \wishbone_RxPointerMSB_reg[8]/NET0131  & n13207 ;
  assign n18665 = ~n13196 & n18664 ;
  assign n18666 = ~n18663 & ~n18665 ;
  assign n18667 = \wishbone_TxPointerMSB_reg[8]/NET0131  & ~n13201 ;
  assign n18668 = \m_wb_adr_o[6]_pad  & \m_wb_adr_o[7]_pad  ;
  assign n18669 = n13097 & n18668 ;
  assign n18670 = ~\m_wb_adr_o[8]_pad  & ~n18669 ;
  assign n18671 = ~n13100 & ~n18670 ;
  assign n18672 = ~n15177 & n18671 ;
  assign n18673 = ~n18667 & ~n18672 ;
  assign n18674 = n18666 & n18673 ;
  assign n18675 = ~\wishbone_RxPointerMSB_reg[11]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n18676 = n13144 & n18675 ;
  assign n18677 = ~n13149 & ~n18676 ;
  assign n18678 = n13143 & n18677 ;
  assign n18679 = n13137 & n18678 ;
  assign n18680 = ~n13170 & ~n18679 ;
  assign n18681 = n13100 & n13101 ;
  assign n18682 = ~\m_wb_adr_o[11]_pad  & ~n18681 ;
  assign n18683 = ~n13103 & ~n18682 ;
  assign n18684 = ~n18680 & n18683 ;
  assign n18685 = \m_wb_adr_o[11]_pad  & n13197 ;
  assign n18686 = \wishbone_TxPointerMSB_reg[11]/NET0131  & ~n13201 ;
  assign n18687 = \wishbone_RxPointerMSB_reg[11]/NET0131  & n13207 ;
  assign n18688 = ~n13196 & n18687 ;
  assign n18689 = ~n18686 & ~n18688 ;
  assign n18690 = ~n18685 & n18689 ;
  assign n18691 = ~n18684 & n18690 ;
  assign n18692 = \wishbone_TxPointerMSB_reg[15]/NET0131  & ~n13166 ;
  assign n18693 = ~n13164 & n18692 ;
  assign n18694 = n15177 & ~n18693 ;
  assign n18695 = ~\m_wb_adr_o[15]_pad  & ~n18648 ;
  assign n18696 = ~n13107 & ~n18695 ;
  assign n18697 = ~n18694 & n18696 ;
  assign n18698 = \m_wb_adr_o[15]_pad  & n13197 ;
  assign n18699 = \wishbone_TxPointerMSB_reg[15]/NET0131  & ~n13201 ;
  assign n18700 = \wishbone_RxPointerMSB_reg[15]/NET0131  & n13207 ;
  assign n18701 = ~n13196 & n18700 ;
  assign n18702 = ~n18699 & ~n18701 ;
  assign n18703 = ~n18698 & n18702 ;
  assign n18704 = ~n18697 & n18703 ;
  assign n18705 = \m_wb_adr_o[4]_pad  & n13197 ;
  assign n18706 = \wishbone_RxPointerMSB_reg[4]/NET0131  & n13207 ;
  assign n18707 = ~n13196 & n18706 ;
  assign n18708 = ~n18705 & ~n18707 ;
  assign n18709 = \wishbone_TxPointerMSB_reg[4]/NET0131  & ~n13201 ;
  assign n18710 = \m_wb_adr_o[4]_pad  & n13095 ;
  assign n18711 = ~\m_wb_adr_o[4]_pad  & ~n13095 ;
  assign n18712 = ~n18710 & ~n18711 ;
  assign n18713 = ~n15177 & n18712 ;
  assign n18714 = ~n18709 & ~n18713 ;
  assign n18715 = n18708 & n18714 ;
  assign n18716 = \m_wb_adr_o[27]_pad  & n13118 ;
  assign n18717 = ~\m_wb_adr_o[27]_pad  & ~n13118 ;
  assign n18718 = \wishbone_TxPointerMSB_reg[27]/NET0131  & ~n13166 ;
  assign n18719 = ~n13164 & n18718 ;
  assign n18720 = n15177 & ~n18719 ;
  assign n18721 = ~n18717 & ~n18720 ;
  assign n18722 = ~n18716 & n18721 ;
  assign n18723 = \m_wb_adr_o[27]_pad  & n13197 ;
  assign n18724 = \wishbone_TxPointerMSB_reg[27]/NET0131  & ~n13201 ;
  assign n18725 = \wishbone_RxPointerMSB_reg[27]/NET0131  & n13207 ;
  assign n18726 = ~n13196 & n18725 ;
  assign n18727 = ~n18724 & ~n18726 ;
  assign n18728 = ~n18723 & n18727 ;
  assign n18729 = ~n18722 & n18728 ;
  assign n18730 = ~\wishbone_RxPointerMSB_reg[31]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n18731 = n13144 & n18730 ;
  assign n18732 = ~n13149 & ~n18731 ;
  assign n18733 = n13143 & n18732 ;
  assign n18734 = n13137 & n18733 ;
  assign n18735 = ~n13170 & ~n18734 ;
  assign n18736 = \m_wb_adr_o[31]_pad  & ~n18735 ;
  assign n18737 = ~n13125 & n18736 ;
  assign n18738 = ~\m_wb_adr_o[31]_pad  & ~n18735 ;
  assign n18739 = n13125 & n18738 ;
  assign n18740 = ~n18737 & ~n18739 ;
  assign n18741 = \m_wb_adr_o[31]_pad  & n13197 ;
  assign n18742 = \wishbone_RxPointerMSB_reg[31]/NET0131  & n13207 ;
  assign n18743 = ~n13196 & n18742 ;
  assign n18744 = \wishbone_TxPointerMSB_reg[31]/NET0131  & ~n13201 ;
  assign n18745 = ~n18743 & ~n18744 ;
  assign n18746 = ~n18741 & n18745 ;
  assign n18747 = n18740 & n18746 ;
  assign n18748 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  & \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n18749 = n12354 & n18748 ;
  assign n18750 = ~\macstatus1_ReceiveEnd_reg/NET0131  & ~n18749 ;
  assign n18751 = \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131  & n18750 ;
  assign n18752 = ~\rxethmac1_RxData_reg[0]/NET0131  & \rxethmac1_RxData_reg[3]/NET0131  ;
  assign n18753 = n12347 & n18752 ;
  assign n18754 = n12274 & n18753 ;
  assign n18755 = \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131  & n13224 ;
  assign n18756 = n18754 & n18755 ;
  assign n18757 = ~n18751 & ~n18756 ;
  assign n18758 = n12269 & n12272 ;
  assign n18759 = n18752 & n18758 ;
  assign n18760 = n12311 & n18759 ;
  assign n18761 = n13224 & n18760 ;
  assign n18762 = n18757 & ~n18761 ;
  assign n18763 = \wishbone_bd_ram_mem2_reg[85][18]/P0001  & n13784 ;
  assign n18764 = \wishbone_bd_ram_mem2_reg[106][18]/P0001  & n13555 ;
  assign n18765 = ~n18763 & ~n18764 ;
  assign n18766 = \wishbone_bd_ram_mem2_reg[197][18]/P0001  & n13594 ;
  assign n18767 = \wishbone_bd_ram_mem2_reg[176][18]/P0001  & n13262 ;
  assign n18768 = ~n18766 & ~n18767 ;
  assign n18769 = n18765 & n18768 ;
  assign n18770 = \wishbone_bd_ram_mem2_reg[221][18]/P0001  & n13641 ;
  assign n18771 = \wishbone_bd_ram_mem2_reg[55][18]/P0001  & n13618 ;
  assign n18772 = ~n18770 & ~n18771 ;
  assign n18773 = \wishbone_bd_ram_mem2_reg[102][18]/P0001  & n13534 ;
  assign n18774 = \wishbone_bd_ram_mem2_reg[157][18]/P0001  & n13445 ;
  assign n18775 = ~n18773 & ~n18774 ;
  assign n18776 = n18772 & n18775 ;
  assign n18777 = n18769 & n18776 ;
  assign n18778 = \wishbone_bd_ram_mem2_reg[7][18]/P0001  & n13546 ;
  assign n18779 = \wishbone_bd_ram_mem2_reg[3][18]/P0001  & n13354 ;
  assign n18780 = ~n18778 & ~n18779 ;
  assign n18781 = \wishbone_bd_ram_mem2_reg[191][18]/P0001  & n14012 ;
  assign n18782 = \wishbone_bd_ram_mem2_reg[254][18]/P0001  & n13283 ;
  assign n18783 = ~n18781 & ~n18782 ;
  assign n18784 = n18780 & n18783 ;
  assign n18785 = \wishbone_bd_ram_mem2_reg[6][18]/P0001  & n13915 ;
  assign n18786 = \wishbone_bd_ram_mem2_reg[222][18]/P0001  & n13721 ;
  assign n18787 = ~n18785 & ~n18786 ;
  assign n18788 = \wishbone_bd_ram_mem2_reg[32][18]/P0001  & n13736 ;
  assign n18789 = \wishbone_bd_ram_mem2_reg[119][18]/P0001  & n14033 ;
  assign n18790 = ~n18788 & ~n18789 ;
  assign n18791 = n18787 & n18790 ;
  assign n18792 = n18784 & n18791 ;
  assign n18793 = n18777 & n18792 ;
  assign n18794 = \wishbone_bd_ram_mem2_reg[40][18]/P0001  & n13661 ;
  assign n18795 = \wishbone_bd_ram_mem2_reg[42][18]/P0001  & n13341 ;
  assign n18796 = ~n18794 & ~n18795 ;
  assign n18797 = \wishbone_bd_ram_mem2_reg[179][18]/P0001  & n14035 ;
  assign n18798 = \wishbone_bd_ram_mem2_reg[210][18]/P0001  & n13443 ;
  assign n18799 = ~n18797 & ~n18798 ;
  assign n18800 = n18796 & n18799 ;
  assign n18801 = \wishbone_bd_ram_mem2_reg[14][18]/P0001  & n13972 ;
  assign n18802 = \wishbone_bd_ram_mem2_reg[61][18]/P0001  & n13544 ;
  assign n18803 = ~n18801 & ~n18802 ;
  assign n18804 = \wishbone_bd_ram_mem2_reg[234][18]/P0001  & n13781 ;
  assign n18805 = \wishbone_bd_ram_mem2_reg[4][18]/P0001  & n13527 ;
  assign n18806 = ~n18804 & ~n18805 ;
  assign n18807 = n18803 & n18806 ;
  assign n18808 = n18800 & n18807 ;
  assign n18809 = \wishbone_bd_ram_mem2_reg[80][18]/P0001  & n13516 ;
  assign n18810 = \wishbone_bd_ram_mem2_reg[99][18]/P0001  & n13996 ;
  assign n18811 = ~n18809 & ~n18810 ;
  assign n18812 = \wishbone_bd_ram_mem2_reg[159][18]/P0001  & n13627 ;
  assign n18813 = \wishbone_bd_ram_mem2_reg[107][18]/P0001  & n13476 ;
  assign n18814 = ~n18812 & ~n18813 ;
  assign n18815 = n18811 & n18814 ;
  assign n18816 = \wishbone_bd_ram_mem2_reg[146][18]/P0001  & n13958 ;
  assign n18817 = \wishbone_bd_ram_mem2_reg[65][18]/P0001  & n13842 ;
  assign n18818 = ~n18816 & ~n18817 ;
  assign n18819 = \wishbone_bd_ram_mem2_reg[13][18]/P0001  & n13844 ;
  assign n18820 = \wishbone_bd_ram_mem2_reg[10][18]/P0001  & n13837 ;
  assign n18821 = ~n18819 & ~n18820 ;
  assign n18822 = n18818 & n18821 ;
  assign n18823 = n18815 & n18822 ;
  assign n18824 = n18808 & n18823 ;
  assign n18825 = n18793 & n18824 ;
  assign n18826 = \wishbone_bd_ram_mem2_reg[12][18]/P0001  & n13733 ;
  assign n18827 = \wishbone_bd_ram_mem2_reg[184][18]/P0001  & n13960 ;
  assign n18828 = ~n18826 & ~n18827 ;
  assign n18829 = \wishbone_bd_ram_mem2_reg[82][18]/P0001  & n13374 ;
  assign n18830 = \wishbone_bd_ram_mem2_reg[174][18]/P0001  & n13899 ;
  assign n18831 = ~n18829 & ~n18830 ;
  assign n18832 = n18828 & n18831 ;
  assign n18833 = \wishbone_bd_ram_mem2_reg[79][18]/P0001  & n13779 ;
  assign n18834 = \wishbone_bd_ram_mem2_reg[90][18]/P0001  & n13906 ;
  assign n18835 = ~n18833 & ~n18834 ;
  assign n18836 = \wishbone_bd_ram_mem2_reg[45][18]/P0001  & n13420 ;
  assign n18837 = \wishbone_bd_ram_mem2_reg[128][18]/P0001  & n13652 ;
  assign n18838 = ~n18836 & ~n18837 ;
  assign n18839 = n18835 & n18838 ;
  assign n18840 = n18832 & n18839 ;
  assign n18841 = \wishbone_bd_ram_mem2_reg[84][18]/P0001  & n13385 ;
  assign n18842 = \wishbone_bd_ram_mem2_reg[193][18]/P0001  & n14022 ;
  assign n18843 = ~n18841 & ~n18842 ;
  assign n18844 = \wishbone_bd_ram_mem2_reg[241][18]/P0001  & n13854 ;
  assign n18845 = \wishbone_bd_ram_mem2_reg[138][18]/P0001  & n13398 ;
  assign n18846 = ~n18844 & ~n18845 ;
  assign n18847 = n18843 & n18846 ;
  assign n18848 = \wishbone_bd_ram_mem2_reg[11][18]/P0001  & n13774 ;
  assign n18849 = \wishbone_bd_ram_mem2_reg[218][18]/P0001  & n13792 ;
  assign n18850 = ~n18848 & ~n18849 ;
  assign n18851 = \wishbone_bd_ram_mem2_reg[126][18]/P0001  & n13786 ;
  assign n18852 = \wishbone_bd_ram_mem2_reg[115][18]/P0001  & n13747 ;
  assign n18853 = ~n18851 & ~n18852 ;
  assign n18854 = n18850 & n18853 ;
  assign n18855 = n18847 & n18854 ;
  assign n18856 = n18840 & n18855 ;
  assign n18857 = \wishbone_bd_ram_mem2_reg[195][18]/P0001  & n13700 ;
  assign n18858 = \wishbone_bd_ram_mem2_reg[103][18]/P0001  & n13320 ;
  assign n18859 = ~n18857 & ~n18858 ;
  assign n18860 = \wishbone_bd_ram_mem2_reg[86][18]/P0001  & n13485 ;
  assign n18861 = \wishbone_bd_ram_mem2_reg[170][18]/P0001  & n14007 ;
  assign n18862 = ~n18860 & ~n18861 ;
  assign n18863 = n18859 & n18862 ;
  assign n18864 = \wishbone_bd_ram_mem2_reg[48][18]/P0001  & n13917 ;
  assign n18865 = \wishbone_bd_ram_mem2_reg[43][18]/P0001  & n13761 ;
  assign n18866 = ~n18864 & ~n18865 ;
  assign n18867 = \wishbone_bd_ram_mem2_reg[230][18]/P0001  & n13994 ;
  assign n18868 = \wishbone_bd_ram_mem2_reg[242][18]/P0001  & n13383 ;
  assign n18869 = ~n18867 & ~n18868 ;
  assign n18870 = n18866 & n18869 ;
  assign n18871 = n18863 & n18870 ;
  assign n18872 = \wishbone_bd_ram_mem2_reg[178][18]/P0001  & n13301 ;
  assign n18873 = \wishbone_bd_ram_mem2_reg[29][18]/P0001  & n13412 ;
  assign n18874 = ~n18872 & ~n18873 ;
  assign n18875 = \wishbone_bd_ram_mem2_reg[229][18]/P0001  & n13552 ;
  assign n18876 = \wishbone_bd_ram_mem2_reg[130][18]/P0001  & n13427 ;
  assign n18877 = ~n18875 & ~n18876 ;
  assign n18878 = n18874 & n18877 ;
  assign n18879 = \wishbone_bd_ram_mem2_reg[251][18]/P0001  & n14019 ;
  assign n18880 = \wishbone_bd_ram_mem2_reg[206][18]/P0001  & n13414 ;
  assign n18881 = ~n18879 & ~n18880 ;
  assign n18882 = \wishbone_bd_ram_mem2_reg[224][18]/P0001  & n13433 ;
  assign n18883 = \wishbone_bd_ram_mem2_reg[185][18]/P0001  & n13372 ;
  assign n18884 = ~n18882 & ~n18883 ;
  assign n18885 = n18881 & n18884 ;
  assign n18886 = n18878 & n18885 ;
  assign n18887 = n18871 & n18886 ;
  assign n18888 = n18856 & n18887 ;
  assign n18889 = n18825 & n18888 ;
  assign n18890 = \wishbone_bd_ram_mem2_reg[16][18]/P0001  & n13695 ;
  assign n18891 = \wishbone_bd_ram_mem2_reg[167][18]/P0001  & n13940 ;
  assign n18892 = ~n18890 & ~n18891 ;
  assign n18893 = \wishbone_bd_ram_mem2_reg[120][18]/P0001  & n13550 ;
  assign n18894 = \wishbone_bd_ram_mem2_reg[247][18]/P0001  & n13571 ;
  assign n18895 = ~n18893 & ~n18894 ;
  assign n18896 = n18892 & n18895 ;
  assign n18897 = \wishbone_bd_ram_mem2_reg[113][18]/P0001  & n13882 ;
  assign n18898 = \wishbone_bd_ram_mem2_reg[134][18]/P0001  & n13494 ;
  assign n18899 = ~n18897 & ~n18898 ;
  assign n18900 = \wishbone_bd_ram_mem2_reg[47][18]/P0001  & n13436 ;
  assign n18901 = \wishbone_bd_ram_mem2_reg[153][18]/P0001  & n13309 ;
  assign n18902 = ~n18900 & ~n18901 ;
  assign n18903 = n18899 & n18902 ;
  assign n18904 = n18896 & n18903 ;
  assign n18905 = \wishbone_bd_ram_mem2_reg[216][18]/P0001  & n14005 ;
  assign n18906 = \wishbone_bd_ram_mem2_reg[238][18]/P0001  & n13819 ;
  assign n18907 = ~n18905 & ~n18906 ;
  assign n18908 = \wishbone_bd_ram_mem2_reg[87][18]/P0001  & n13691 ;
  assign n18909 = \wishbone_bd_ram_mem2_reg[38][18]/P0001  & n13828 ;
  assign n18910 = ~n18908 & ~n18909 ;
  assign n18911 = n18907 & n18910 ;
  assign n18912 = \wishbone_bd_ram_mem2_reg[75][18]/P0001  & n13605 ;
  assign n18913 = \wishbone_bd_ram_mem2_reg[39][18]/P0001  & n13893 ;
  assign n18914 = ~n18912 & ~n18913 ;
  assign n18915 = \wishbone_bd_ram_mem2_reg[2][18]/P0001  & n13975 ;
  assign n18916 = \wishbone_bd_ram_mem2_reg[111][18]/P0001  & n13471 ;
  assign n18917 = ~n18915 & ~n18916 ;
  assign n18918 = n18914 & n18917 ;
  assign n18919 = n18911 & n18918 ;
  assign n18920 = n18904 & n18919 ;
  assign n18921 = \wishbone_bd_ram_mem2_reg[156][18]/P0001  & n13769 ;
  assign n18922 = \wishbone_bd_ram_mem2_reg[37][18]/P0001  & n13710 ;
  assign n18923 = ~n18921 & ~n18922 ;
  assign n18924 = \wishbone_bd_ram_mem2_reg[88][18]/P0001  & n13347 ;
  assign n18925 = \wishbone_bd_ram_mem2_reg[252][18]/P0001  & n13986 ;
  assign n18926 = ~n18924 & ~n18925 ;
  assign n18927 = n18923 & n18926 ;
  assign n18928 = \wishbone_bd_ram_mem2_reg[211][18]/P0001  & n13805 ;
  assign n18929 = \wishbone_bd_ram_mem2_reg[200][18]/P0001  & n13922 ;
  assign n18930 = ~n18928 & ~n18929 ;
  assign n18931 = \wishbone_bd_ram_mem2_reg[96][18]/P0001  & n13425 ;
  assign n18932 = \wishbone_bd_ram_mem2_reg[5][18]/P0001  & n13243 ;
  assign n18933 = ~n18931 & ~n18932 ;
  assign n18934 = n18930 & n18933 ;
  assign n18935 = n18927 & n18934 ;
  assign n18936 = \wishbone_bd_ram_mem2_reg[68][18]/P0001  & n13379 ;
  assign n18937 = \wishbone_bd_ram_mem2_reg[76][18]/P0001  & n13831 ;
  assign n18938 = ~n18936 & ~n18937 ;
  assign n18939 = \wishbone_bd_ram_mem2_reg[125][18]/P0001  & n13396 ;
  assign n18940 = \wishbone_bd_ram_mem2_reg[163][18]/P0001  & n13255 ;
  assign n18941 = ~n18939 & ~n18940 ;
  assign n18942 = n18938 & n18941 ;
  assign n18943 = \wishbone_bd_ram_mem2_reg[95][18]/P0001  & n13317 ;
  assign n18944 = \wishbone_bd_ram_mem2_reg[101][18]/P0001  & n13772 ;
  assign n18945 = ~n18943 & ~n18944 ;
  assign n18946 = \wishbone_bd_ram_mem2_reg[89][18]/P0001  & n13910 ;
  assign n18947 = \wishbone_bd_ram_mem2_reg[172][18]/P0001  & n13377 ;
  assign n18948 = ~n18946 & ~n18947 ;
  assign n18949 = n18945 & n18948 ;
  assign n18950 = n18942 & n18949 ;
  assign n18951 = n18935 & n18950 ;
  assign n18952 = n18920 & n18951 ;
  assign n18953 = \wishbone_bd_ram_mem2_reg[41][18]/P0001  & n14017 ;
  assign n18954 = \wishbone_bd_ram_mem2_reg[97][18]/P0001  & n13724 ;
  assign n18955 = ~n18953 & ~n18954 ;
  assign n18956 = \wishbone_bd_ram_mem2_reg[160][18]/P0001  & n13271 ;
  assign n18957 = \wishbone_bd_ram_mem2_reg[0][18]/P0001  & n13539 ;
  assign n18958 = ~n18956 & ~n18957 ;
  assign n18959 = n18955 & n18958 ;
  assign n18960 = \wishbone_bd_ram_mem2_reg[114][18]/P0001  & n13763 ;
  assign n18961 = \wishbone_bd_ram_mem2_reg[91][18]/P0001  & n13954 ;
  assign n18962 = ~n18960 & ~n18961 ;
  assign n18963 = \wishbone_bd_ram_mem2_reg[151][18]/P0001  & n13697 ;
  assign n18964 = \wishbone_bd_ram_mem2_reg[244][18]/P0001  & n13474 ;
  assign n18965 = ~n18963 & ~n18964 ;
  assign n18966 = n18962 & n18965 ;
  assign n18967 = n18959 & n18966 ;
  assign n18968 = \wishbone_bd_ram_mem2_reg[208][18]/P0001  & n14010 ;
  assign n18969 = \wishbone_bd_ram_mem2_reg[121][18]/P0001  & n13983 ;
  assign n18970 = ~n18968 & ~n18969 ;
  assign n18971 = \wishbone_bd_ram_mem2_reg[187][18]/P0001  & n13756 ;
  assign n18972 = \wishbone_bd_ram_mem2_reg[131][18]/P0001  & n13358 ;
  assign n18973 = ~n18971 & ~n18972 ;
  assign n18974 = n18970 & n18973 ;
  assign n18975 = \wishbone_bd_ram_mem2_reg[9][18]/P0001  & n13580 ;
  assign n18976 = \wishbone_bd_ram_mem2_reg[25][18]/P0001  & n13742 ;
  assign n18977 = ~n18975 & ~n18976 ;
  assign n18978 = \wishbone_bd_ram_mem2_reg[201][18]/P0001  & n13600 ;
  assign n18979 = \wishbone_bd_ram_mem2_reg[250][18]/P0001  & n13677 ;
  assign n18980 = ~n18978 & ~n18979 ;
  assign n18981 = n18977 & n18980 ;
  assign n18982 = n18974 & n18981 ;
  assign n18983 = n18967 & n18982 ;
  assign n18984 = \wishbone_bd_ram_mem2_reg[20][18]/P0001  & n13839 ;
  assign n18985 = \wishbone_bd_ram_mem2_reg[123][18]/P0001  & n13749 ;
  assign n18986 = ~n18984 & ~n18985 ;
  assign n18987 = \wishbone_bd_ram_mem2_reg[122][18]/P0001  & n13679 ;
  assign n18988 = \wishbone_bd_ram_mem2_reg[162][18]/P0001  & n13726 ;
  assign n18989 = ~n18987 & ~n18988 ;
  assign n18990 = n18986 & n18989 ;
  assign n18991 = \wishbone_bd_ram_mem2_reg[232][18]/P0001  & n13510 ;
  assign n18992 = \wishbone_bd_ram_mem2_reg[70][18]/P0001  & n13339 ;
  assign n18993 = ~n18991 & ~n18992 ;
  assign n18994 = \wishbone_bd_ram_mem2_reg[59][18]/P0001  & n13613 ;
  assign n18995 = \wishbone_bd_ram_mem2_reg[169][18]/P0001  & n13541 ;
  assign n18996 = ~n18994 & ~n18995 ;
  assign n18997 = n18993 & n18996 ;
  assign n18998 = n18990 & n18997 ;
  assign n18999 = \wishbone_bd_ram_mem2_reg[149][18]/P0001  & n13469 ;
  assign n19000 = \wishbone_bd_ram_mem2_reg[100][18]/P0001  & n13401 ;
  assign n19001 = ~n18999 & ~n19000 ;
  assign n19002 = \wishbone_bd_ram_mem2_reg[226][18]/P0001  & n13668 ;
  assign n19003 = \wishbone_bd_ram_mem2_reg[196][18]/P0001  & n13977 ;
  assign n19004 = ~n19002 & ~n19003 ;
  assign n19005 = n19001 & n19004 ;
  assign n19006 = \wishbone_bd_ram_mem2_reg[34][18]/P0001  & n13450 ;
  assign n19007 = \wishbone_bd_ram_mem2_reg[207][18]/P0001  & n13826 ;
  assign n19008 = ~n19006 & ~n19007 ;
  assign n19009 = \wishbone_bd_ram_mem2_reg[127][18]/P0001  & n13803 ;
  assign n19010 = \wishbone_bd_ram_mem2_reg[166][18]/P0001  & n13999 ;
  assign n19011 = ~n19009 & ~n19010 ;
  assign n19012 = n19008 & n19011 ;
  assign n19013 = n19005 & n19012 ;
  assign n19014 = n18998 & n19013 ;
  assign n19015 = n18983 & n19014 ;
  assign n19016 = n18952 & n19015 ;
  assign n19017 = n18889 & n19016 ;
  assign n19018 = \wishbone_bd_ram_mem2_reg[1][18]/P0001  & n13888 ;
  assign n19019 = \wishbone_bd_ram_mem2_reg[33][18]/P0001  & n13933 ;
  assign n19020 = ~n19018 & ~n19019 ;
  assign n19021 = \wishbone_bd_ram_mem2_reg[23][18]/P0001  & n13857 ;
  assign n19022 = \wishbone_bd_ram_mem2_reg[155][18]/P0001  & n13738 ;
  assign n19023 = ~n19021 & ~n19022 ;
  assign n19024 = n19020 & n19023 ;
  assign n19025 = \wishbone_bd_ram_mem2_reg[108][18]/P0001  & n13814 ;
  assign n19026 = \wishbone_bd_ram_mem2_reg[50][18]/P0001  & n13686 ;
  assign n19027 = ~n19025 & ~n19026 ;
  assign n19028 = \wishbone_bd_ram_mem2_reg[139][18]/P0001  & n13566 ;
  assign n19029 = \wishbone_bd_ram_mem2_reg[132][18]/P0001  & n13927 ;
  assign n19030 = ~n19028 & ~n19029 ;
  assign n19031 = n19027 & n19030 ;
  assign n19032 = n19024 & n19031 ;
  assign n19033 = \wishbone_bd_ram_mem2_reg[72][18]/P0001  & n13582 ;
  assign n19034 = \wishbone_bd_ram_mem2_reg[140][18]/P0001  & n13287 ;
  assign n19035 = ~n19033 & ~n19034 ;
  assign n19036 = \wishbone_bd_ram_mem2_reg[67][18]/P0001  & n13663 ;
  assign n19037 = \wishbone_bd_ram_mem2_reg[94][18]/P0001  & n13833 ;
  assign n19038 = ~n19036 & ~n19037 ;
  assign n19039 = n19035 & n19038 ;
  assign n19040 = \wishbone_bd_ram_mem2_reg[205][18]/P0001  & n13947 ;
  assign n19041 = \wishbone_bd_ram_mem2_reg[18][18]/P0001  & n13532 ;
  assign n19042 = ~n19040 & ~n19041 ;
  assign n19043 = \wishbone_bd_ram_mem2_reg[188][18]/P0001  & n13407 ;
  assign n19044 = \wishbone_bd_ram_mem2_reg[198][18]/P0001  & n13592 ;
  assign n19045 = ~n19043 & ~n19044 ;
  assign n19046 = n19042 & n19045 ;
  assign n19047 = n19039 & n19046 ;
  assign n19048 = n19032 & n19047 ;
  assign n19049 = \wishbone_bd_ram_mem2_reg[240][18]/P0001  & n13352 ;
  assign n19050 = \wishbone_bd_ram_mem2_reg[143][18]/P0001  & n13461 ;
  assign n19051 = ~n19049 & ~n19050 ;
  assign n19052 = \wishbone_bd_ram_mem2_reg[24][18]/P0001  & n13970 ;
  assign n19053 = \wishbone_bd_ram_mem2_reg[104][18]/P0001  & n13684 ;
  assign n19054 = ~n19052 & ~n19053 ;
  assign n19055 = n19051 & n19054 ;
  assign n19056 = \wishbone_bd_ram_mem2_reg[165][18]/P0001  & n14028 ;
  assign n19057 = \wishbone_bd_ram_mem2_reg[105][18]/P0001  & n13503 ;
  assign n19058 = ~n19056 & ~n19057 ;
  assign n19059 = \wishbone_bd_ram_mem2_reg[46][18]/P0001  & n13298 ;
  assign n19060 = \wishbone_bd_ram_mem2_reg[93][18]/P0001  & n13891 ;
  assign n19061 = ~n19059 & ~n19060 ;
  assign n19062 = n19058 & n19061 ;
  assign n19063 = n19055 & n19062 ;
  assign n19064 = \wishbone_bd_ram_mem2_reg[209][18]/P0001  & n13689 ;
  assign n19065 = \wishbone_bd_ram_mem2_reg[21][18]/P0001  & n13438 ;
  assign n19066 = ~n19064 & ~n19065 ;
  assign n19067 = \wishbone_bd_ram_mem2_reg[233][18]/P0001  & n13332 ;
  assign n19068 = \wishbone_bd_ram_mem2_reg[186][18]/P0001  & n13616 ;
  assign n19069 = ~n19067 & ~n19068 ;
  assign n19070 = n19066 & n19069 ;
  assign n19071 = \wishbone_bd_ram_mem2_reg[194][18]/P0001  & n13624 ;
  assign n19072 = \wishbone_bd_ram_mem2_reg[71][18]/P0001  & n13636 ;
  assign n19073 = ~n19071 & ~n19072 ;
  assign n19074 = \wishbone_bd_ram_mem2_reg[31][18]/P0001  & n13758 ;
  assign n19075 = \wishbone_bd_ram_mem2_reg[53][18]/P0001  & n13875 ;
  assign n19076 = ~n19074 & ~n19075 ;
  assign n19077 = n19073 & n19076 ;
  assign n19078 = n19070 & n19077 ;
  assign n19079 = n19063 & n19078 ;
  assign n19080 = n19048 & n19079 ;
  assign n19081 = \wishbone_bd_ram_mem2_reg[19][18]/P0001  & n13886 ;
  assign n19082 = \wishbone_bd_ram_mem2_reg[239][18]/P0001  & n13349 ;
  assign n19083 = ~n19081 & ~n19082 ;
  assign n19084 = \wishbone_bd_ram_mem2_reg[78][18]/P0001  & n13277 ;
  assign n19085 = \wishbone_bd_ram_mem2_reg[52][18]/P0001  & n13988 ;
  assign n19086 = ~n19084 & ~n19085 ;
  assign n19087 = n19083 & n19086 ;
  assign n19088 = \wishbone_bd_ram_mem2_reg[74][18]/P0001  & n13564 ;
  assign n19089 = \wishbone_bd_ram_mem2_reg[199][18]/P0001  & n13499 ;
  assign n19090 = ~n19088 & ~n19089 ;
  assign n19091 = \wishbone_bd_ram_mem2_reg[217][18]/P0001  & n13767 ;
  assign n19092 = \wishbone_bd_ram_mem2_reg[214][18]/P0001  & n13938 ;
  assign n19093 = ~n19091 & ~n19092 ;
  assign n19094 = n19090 & n19093 ;
  assign n19095 = n19087 & n19094 ;
  assign n19096 = \wishbone_bd_ram_mem2_reg[235][18]/P0001  & n13518 ;
  assign n19097 = \wishbone_bd_ram_mem2_reg[110][18]/P0001  & n14030 ;
  assign n19098 = ~n19096 & ~n19097 ;
  assign n19099 = \wishbone_bd_ram_mem2_reg[27][18]/P0001  & n13251 ;
  assign n19100 = \wishbone_bd_ram_mem2_reg[183][18]/P0001  & n13645 ;
  assign n19101 = ~n19099 & ~n19100 ;
  assign n19102 = n19098 & n19101 ;
  assign n19103 = \wishbone_bd_ram_mem2_reg[192][18]/P0001  & n13390 ;
  assign n19104 = \wishbone_bd_ram_mem2_reg[116][18]/P0001  & n13865 ;
  assign n19105 = ~n19103 & ~n19104 ;
  assign n19106 = \wishbone_bd_ram_mem2_reg[36][18]/P0001  & n13639 ;
  assign n19107 = \wishbone_bd_ram_mem2_reg[219][18]/P0001  & n13577 ;
  assign n19108 = ~n19106 & ~n19107 ;
  assign n19109 = n19105 & n19108 ;
  assign n19110 = n19102 & n19109 ;
  assign n19111 = n19095 & n19110 ;
  assign n19112 = \wishbone_bd_ram_mem2_reg[145][18]/P0001  & n13715 ;
  assign n19113 = \wishbone_bd_ram_mem2_reg[8][18]/P0001  & n13459 ;
  assign n19114 = ~n19112 & ~n19113 ;
  assign n19115 = \wishbone_bd_ram_mem2_reg[133][18]/P0001  & n13492 ;
  assign n19116 = \wishbone_bd_ram_mem2_reg[202][18]/P0001  & n13268 ;
  assign n19117 = ~n19115 & ~n19116 ;
  assign n19118 = n19114 & n19117 ;
  assign n19119 = \wishbone_bd_ram_mem2_reg[62][18]/P0001  & n13529 ;
  assign n19120 = \wishbone_bd_ram_mem2_reg[57][18]/P0001  & n13731 ;
  assign n19121 = ~n19119 & ~n19120 ;
  assign n19122 = \wishbone_bd_ram_mem2_reg[117][18]/P0001  & n13557 ;
  assign n19123 = \wishbone_bd_ram_mem2_reg[30][18]/P0001  & n13713 ;
  assign n19124 = ~n19122 & ~n19123 ;
  assign n19125 = n19121 & n19124 ;
  assign n19126 = n19118 & n19125 ;
  assign n19127 = \wishbone_bd_ram_mem2_reg[137][18]/P0001  & n13808 ;
  assign n19128 = \wishbone_bd_ram_mem2_reg[177][18]/P0001  & n13863 ;
  assign n19129 = ~n19127 & ~n19128 ;
  assign n19130 = \wishbone_bd_ram_mem2_reg[154][18]/P0001  & n13403 ;
  assign n19131 = \wishbone_bd_ram_mem2_reg[152][18]/P0001  & n13912 ;
  assign n19132 = ~n19130 & ~n19131 ;
  assign n19133 = n19129 & n19132 ;
  assign n19134 = \wishbone_bd_ram_mem2_reg[158][18]/P0001  & n13294 ;
  assign n19135 = \wishbone_bd_ram_mem2_reg[49][18]/P0001  & n13929 ;
  assign n19136 = ~n19134 & ~n19135 ;
  assign n19137 = \wishbone_bd_ram_mem2_reg[204][18]/P0001  & n13821 ;
  assign n19138 = \wishbone_bd_ram_mem2_reg[64][18]/P0001  & n13904 ;
  assign n19139 = ~n19137 & ~n19138 ;
  assign n19140 = n19136 & n19139 ;
  assign n19141 = n19133 & n19140 ;
  assign n19142 = n19126 & n19141 ;
  assign n19143 = n19111 & n19142 ;
  assign n19144 = n19080 & n19143 ;
  assign n19145 = \wishbone_bd_ram_mem2_reg[203][18]/P0001  & n13816 ;
  assign n19146 = \wishbone_bd_ram_mem2_reg[129][18]/P0001  & n13629 ;
  assign n19147 = ~n19145 & ~n19146 ;
  assign n19148 = \wishbone_bd_ram_mem2_reg[246][18]/P0001  & n13981 ;
  assign n19149 = \wishbone_bd_ram_mem2_reg[245][18]/P0001  & n13877 ;
  assign n19150 = ~n19148 & ~n19149 ;
  assign n19151 = n19147 & n19150 ;
  assign n19152 = \wishbone_bd_ram_mem2_reg[144][18]/P0001  & n13508 ;
  assign n19153 = \wishbone_bd_ram_mem2_reg[248][18]/P0001  & n13647 ;
  assign n19154 = ~n19152 & ~n19153 ;
  assign n19155 = \wishbone_bd_ram_mem2_reg[135][18]/P0001  & n13672 ;
  assign n19156 = \wishbone_bd_ram_mem2_reg[150][18]/P0001  & n13666 ;
  assign n19157 = ~n19155 & ~n19156 ;
  assign n19158 = n19154 & n19157 ;
  assign n19159 = n19151 & n19158 ;
  assign n19160 = \wishbone_bd_ram_mem2_reg[215][18]/P0001  & n13901 ;
  assign n19161 = \wishbone_bd_ram_mem2_reg[181][18]/P0001  & n13587 ;
  assign n19162 = ~n19160 & ~n19161 ;
  assign n19163 = \wishbone_bd_ram_mem2_reg[190][18]/P0001  & n13365 ;
  assign n19164 = \wishbone_bd_ram_mem2_reg[161][18]/P0001  & n13505 ;
  assign n19165 = ~n19163 & ~n19164 ;
  assign n19166 = n19162 & n19165 ;
  assign n19167 = \wishbone_bd_ram_mem2_reg[35][18]/P0001  & n13523 ;
  assign n19168 = \wishbone_bd_ram_mem2_reg[255][18]/P0001  & n13952 ;
  assign n19169 = ~n19167 & ~n19168 ;
  assign n19170 = \wishbone_bd_ram_mem2_reg[54][18]/P0001  & n13622 ;
  assign n19171 = \wishbone_bd_ram_mem2_reg[180][18]/P0001  & n13650 ;
  assign n19172 = ~n19170 & ~n19171 ;
  assign n19173 = n19169 & n19172 ;
  assign n19174 = n19166 & n19173 ;
  assign n19175 = n19159 & n19174 ;
  assign n19176 = \wishbone_bd_ram_mem2_reg[220][18]/P0001  & n13965 ;
  assign n19177 = \wishbone_bd_ram_mem2_reg[51][18]/P0001  & n13880 ;
  assign n19178 = ~n19176 & ~n19177 ;
  assign n19179 = \wishbone_bd_ram_mem2_reg[60][18]/P0001  & n13790 ;
  assign n19180 = \wishbone_bd_ram_mem2_reg[148][18]/P0001  & n13868 ;
  assign n19181 = ~n19179 & ~n19180 ;
  assign n19182 = n19178 & n19181 ;
  assign n19183 = \wishbone_bd_ram_mem2_reg[231][18]/P0001  & n13363 ;
  assign n19184 = \wishbone_bd_ram_mem2_reg[136][18]/P0001  & n13963 ;
  assign n19185 = ~n19183 & ~n19184 ;
  assign n19186 = \wishbone_bd_ram_mem2_reg[225][18]/P0001  & n13719 ;
  assign n19187 = \wishbone_bd_ram_mem2_reg[81][18]/P0001  & n13409 ;
  assign n19188 = ~n19186 & ~n19187 ;
  assign n19189 = n19185 & n19188 ;
  assign n19190 = n19182 & n19189 ;
  assign n19191 = \wishbone_bd_ram_mem2_reg[26][18]/P0001  & n13521 ;
  assign n19192 = \wishbone_bd_ram_mem2_reg[22][18]/P0001  & n13744 ;
  assign n19193 = ~n19191 & ~n19192 ;
  assign n19194 = \wishbone_bd_ram_mem2_reg[92][18]/P0001  & n13859 ;
  assign n19195 = \wishbone_bd_ram_mem2_reg[175][18]/P0001  & n13674 ;
  assign n19196 = ~n19194 & ~n19195 ;
  assign n19197 = n19193 & n19196 ;
  assign n19198 = \wishbone_bd_ram_mem2_reg[243][18]/P0001  & n13575 ;
  assign n19199 = \wishbone_bd_ram_mem2_reg[236][18]/P0001  & n13480 ;
  assign n19200 = ~n19198 & ~n19199 ;
  assign n19201 = \wishbone_bd_ram_mem2_reg[73][18]/P0001  & n13456 ;
  assign n19202 = \wishbone_bd_ram_mem2_reg[124][18]/P0001  & n14024 ;
  assign n19203 = ~n19201 & ~n19202 ;
  assign n19204 = n19200 & n19203 ;
  assign n19205 = n19197 & n19204 ;
  assign n19206 = n19190 & n19205 ;
  assign n19207 = n19175 & n19206 ;
  assign n19208 = \wishbone_bd_ram_mem2_reg[141][18]/P0001  & n13852 ;
  assign n19209 = \wishbone_bd_ram_mem2_reg[171][18]/P0001  & n13422 ;
  assign n19210 = ~n19208 & ~n19209 ;
  assign n19211 = \wishbone_bd_ram_mem2_reg[164][18]/P0001  & n13236 ;
  assign n19212 = \wishbone_bd_ram_mem2_reg[237][18]/P0001  & n13924 ;
  assign n19213 = ~n19211 & ~n19212 ;
  assign n19214 = n19210 & n19213 ;
  assign n19215 = \wishbone_bd_ram_mem2_reg[118][18]/P0001  & n13589 ;
  assign n19216 = \wishbone_bd_ram_mem2_reg[227][18]/P0001  & n13388 ;
  assign n19217 = ~n19215 & ~n19216 ;
  assign n19218 = \wishbone_bd_ram_mem2_reg[112][18]/P0001  & n13482 ;
  assign n19219 = \wishbone_bd_ram_mem2_reg[189][18]/P0001  & n14001 ;
  assign n19220 = ~n19218 & ~n19219 ;
  assign n19221 = n19217 & n19220 ;
  assign n19222 = n19214 & n19221 ;
  assign n19223 = \wishbone_bd_ram_mem2_reg[223][18]/P0001  & n13335 ;
  assign n19224 = \wishbone_bd_ram_mem2_reg[249][18]/P0001  & n13431 ;
  assign n19225 = ~n19223 & ~n19224 ;
  assign n19226 = \wishbone_bd_ram_mem2_reg[173][18]/P0001  & n13360 ;
  assign n19227 = \wishbone_bd_ram_mem2_reg[66][18]/P0001  & n13603 ;
  assign n19228 = ~n19226 & ~n19227 ;
  assign n19229 = n19225 & n19228 ;
  assign n19230 = \wishbone_bd_ram_mem2_reg[142][18]/P0001  & n13448 ;
  assign n19231 = \wishbone_bd_ram_mem2_reg[77][18]/P0001  & n13935 ;
  assign n19232 = ~n19230 & ~n19231 ;
  assign n19233 = \wishbone_bd_ram_mem2_reg[83][18]/P0001  & n13454 ;
  assign n19234 = \wishbone_bd_ram_mem2_reg[56][18]/P0001  & n13611 ;
  assign n19235 = ~n19233 & ~n19234 ;
  assign n19236 = n19232 & n19235 ;
  assign n19237 = n19229 & n19236 ;
  assign n19238 = n19222 & n19237 ;
  assign n19239 = \wishbone_bd_ram_mem2_reg[98][18]/P0001  & n13569 ;
  assign n19240 = \wishbone_bd_ram_mem2_reg[228][18]/P0001  & n13497 ;
  assign n19241 = ~n19239 & ~n19240 ;
  assign n19242 = \wishbone_bd_ram_mem2_reg[69][18]/P0001  & n13487 ;
  assign n19243 = \wishbone_bd_ram_mem2_reg[44][18]/P0001  & n13291 ;
  assign n19244 = ~n19242 & ~n19243 ;
  assign n19245 = n19241 & n19244 ;
  assign n19246 = \wishbone_bd_ram_mem2_reg[213][18]/P0001  & n13870 ;
  assign n19247 = \wishbone_bd_ram_mem2_reg[212][18]/P0001  & n13634 ;
  assign n19248 = ~n19246 & ~n19247 ;
  assign n19249 = \wishbone_bd_ram_mem2_reg[63][18]/P0001  & n13327 ;
  assign n19250 = \wishbone_bd_ram_mem2_reg[17][18]/P0001  & n13324 ;
  assign n19251 = ~n19249 & ~n19250 ;
  assign n19252 = n19248 & n19251 ;
  assign n19253 = n19245 & n19252 ;
  assign n19254 = \wishbone_bd_ram_mem2_reg[253][18]/P0001  & n13708 ;
  assign n19255 = \wishbone_bd_ram_mem2_reg[147][18]/P0001  & n13702 ;
  assign n19256 = ~n19254 & ~n19255 ;
  assign n19257 = \wishbone_bd_ram_mem2_reg[28][18]/P0001  & n13810 ;
  assign n19258 = \wishbone_bd_ram_mem2_reg[15][18]/P0001  & n13797 ;
  assign n19259 = ~n19257 & ~n19258 ;
  assign n19260 = n19256 & n19259 ;
  assign n19261 = \wishbone_bd_ram_mem2_reg[168][18]/P0001  & n13795 ;
  assign n19262 = \wishbone_bd_ram_mem2_reg[109][18]/P0001  & n13306 ;
  assign n19263 = ~n19261 & ~n19262 ;
  assign n19264 = \wishbone_bd_ram_mem2_reg[182][18]/P0001  & n13598 ;
  assign n19265 = \wishbone_bd_ram_mem2_reg[58][18]/P0001  & n13949 ;
  assign n19266 = ~n19264 & ~n19265 ;
  assign n19267 = n19263 & n19266 ;
  assign n19268 = n19260 & n19267 ;
  assign n19269 = n19253 & n19268 ;
  assign n19270 = n19238 & n19269 ;
  assign n19271 = n19207 & n19270 ;
  assign n19272 = n19144 & n19271 ;
  assign n19273 = n19017 & n19272 ;
  assign n19274 = n14047 & ~n19273 ;
  assign n19275 = n14049 & n14063 ;
  assign n19276 = n14058 & n19275 ;
  assign n19277 = ~n14046 & ~n19276 ;
  assign n19278 = ~\wishbone_TxLength_reg[2]/NET0131  & n17918 ;
  assign n19279 = \wishbone_TxLength_reg[2]/NET0131  & ~n17918 ;
  assign n19280 = ~n19278 & ~n19279 ;
  assign n19281 = n19277 & n19280 ;
  assign n19282 = ~n19274 & ~n19281 ;
  assign n19283 = n10663 & ~n12137 ;
  assign n19284 = \wishbone_bd_ram_mem2_reg[128][16]/P0001  & n13652 ;
  assign n19285 = \wishbone_bd_ram_mem2_reg[55][16]/P0001  & n13618 ;
  assign n19286 = ~n19284 & ~n19285 ;
  assign n19287 = \wishbone_bd_ram_mem2_reg[34][16]/P0001  & n13450 ;
  assign n19288 = \wishbone_bd_ram_mem2_reg[125][16]/P0001  & n13396 ;
  assign n19289 = ~n19287 & ~n19288 ;
  assign n19290 = n19286 & n19289 ;
  assign n19291 = \wishbone_bd_ram_mem2_reg[220][16]/P0001  & n13965 ;
  assign n19292 = \wishbone_bd_ram_mem2_reg[118][16]/P0001  & n13589 ;
  assign n19293 = ~n19291 & ~n19292 ;
  assign n19294 = \wishbone_bd_ram_mem2_reg[138][16]/P0001  & n13398 ;
  assign n19295 = \wishbone_bd_ram_mem2_reg[127][16]/P0001  & n13803 ;
  assign n19296 = ~n19294 & ~n19295 ;
  assign n19297 = n19293 & n19296 ;
  assign n19298 = n19290 & n19297 ;
  assign n19299 = \wishbone_bd_ram_mem2_reg[103][16]/P0001  & n13320 ;
  assign n19300 = \wishbone_bd_ram_mem2_reg[69][16]/P0001  & n13487 ;
  assign n19301 = ~n19299 & ~n19300 ;
  assign n19302 = \wishbone_bd_ram_mem2_reg[254][16]/P0001  & n13283 ;
  assign n19303 = \wishbone_bd_ram_mem2_reg[39][16]/P0001  & n13893 ;
  assign n19304 = ~n19302 & ~n19303 ;
  assign n19305 = n19301 & n19304 ;
  assign n19306 = \wishbone_bd_ram_mem2_reg[137][16]/P0001  & n13808 ;
  assign n19307 = \wishbone_bd_ram_mem2_reg[20][16]/P0001  & n13839 ;
  assign n19308 = ~n19306 & ~n19307 ;
  assign n19309 = \wishbone_bd_ram_mem2_reg[31][16]/P0001  & n13758 ;
  assign n19310 = \wishbone_bd_ram_mem2_reg[237][16]/P0001  & n13924 ;
  assign n19311 = ~n19309 & ~n19310 ;
  assign n19312 = n19308 & n19311 ;
  assign n19313 = n19305 & n19312 ;
  assign n19314 = n19298 & n19313 ;
  assign n19315 = \wishbone_bd_ram_mem2_reg[204][16]/P0001  & n13821 ;
  assign n19316 = \wishbone_bd_ram_mem2_reg[120][16]/P0001  & n13550 ;
  assign n19317 = ~n19315 & ~n19316 ;
  assign n19318 = \wishbone_bd_ram_mem2_reg[79][16]/P0001  & n13779 ;
  assign n19319 = \wishbone_bd_ram_mem2_reg[6][16]/P0001  & n13915 ;
  assign n19320 = ~n19318 & ~n19319 ;
  assign n19321 = n19317 & n19320 ;
  assign n19322 = \wishbone_bd_ram_mem2_reg[221][16]/P0001  & n13641 ;
  assign n19323 = \wishbone_bd_ram_mem2_reg[0][16]/P0001  & n13539 ;
  assign n19324 = ~n19322 & ~n19323 ;
  assign n19325 = \wishbone_bd_ram_mem2_reg[8][16]/P0001  & n13459 ;
  assign n19326 = \wishbone_bd_ram_mem2_reg[100][16]/P0001  & n13401 ;
  assign n19327 = ~n19325 & ~n19326 ;
  assign n19328 = n19324 & n19327 ;
  assign n19329 = n19321 & n19328 ;
  assign n19330 = \wishbone_bd_ram_mem2_reg[164][16]/P0001  & n13236 ;
  assign n19331 = \wishbone_bd_ram_mem2_reg[188][16]/P0001  & n13407 ;
  assign n19332 = ~n19330 & ~n19331 ;
  assign n19333 = \wishbone_bd_ram_mem2_reg[241][16]/P0001  & n13854 ;
  assign n19334 = \wishbone_bd_ram_mem2_reg[197][16]/P0001  & n13594 ;
  assign n19335 = ~n19333 & ~n19334 ;
  assign n19336 = n19332 & n19335 ;
  assign n19337 = \wishbone_bd_ram_mem2_reg[122][16]/P0001  & n13679 ;
  assign n19338 = \wishbone_bd_ram_mem2_reg[33][16]/P0001  & n13933 ;
  assign n19339 = ~n19337 & ~n19338 ;
  assign n19340 = \wishbone_bd_ram_mem2_reg[91][16]/P0001  & n13954 ;
  assign n19341 = \wishbone_bd_ram_mem2_reg[161][16]/P0001  & n13505 ;
  assign n19342 = ~n19340 & ~n19341 ;
  assign n19343 = n19339 & n19342 ;
  assign n19344 = n19336 & n19343 ;
  assign n19345 = n19329 & n19344 ;
  assign n19346 = n19314 & n19345 ;
  assign n19347 = \wishbone_bd_ram_mem2_reg[170][16]/P0001  & n14007 ;
  assign n19348 = \wishbone_bd_ram_mem2_reg[71][16]/P0001  & n13636 ;
  assign n19349 = ~n19347 & ~n19348 ;
  assign n19350 = \wishbone_bd_ram_mem2_reg[52][16]/P0001  & n13988 ;
  assign n19351 = \wishbone_bd_ram_mem2_reg[40][16]/P0001  & n13661 ;
  assign n19352 = ~n19350 & ~n19351 ;
  assign n19353 = n19349 & n19352 ;
  assign n19354 = \wishbone_bd_ram_mem2_reg[244][16]/P0001  & n13474 ;
  assign n19355 = \wishbone_bd_ram_mem2_reg[129][16]/P0001  & n13629 ;
  assign n19356 = ~n19354 & ~n19355 ;
  assign n19357 = \wishbone_bd_ram_mem2_reg[242][16]/P0001  & n13383 ;
  assign n19358 = \wishbone_bd_ram_mem2_reg[11][16]/P0001  & n13774 ;
  assign n19359 = ~n19357 & ~n19358 ;
  assign n19360 = n19356 & n19359 ;
  assign n19361 = n19353 & n19360 ;
  assign n19362 = \wishbone_bd_ram_mem2_reg[41][16]/P0001  & n14017 ;
  assign n19363 = \wishbone_bd_ram_mem2_reg[240][16]/P0001  & n13352 ;
  assign n19364 = ~n19362 & ~n19363 ;
  assign n19365 = \wishbone_bd_ram_mem2_reg[143][16]/P0001  & n13461 ;
  assign n19366 = \wishbone_bd_ram_mem2_reg[139][16]/P0001  & n13566 ;
  assign n19367 = ~n19365 & ~n19366 ;
  assign n19368 = n19364 & n19367 ;
  assign n19369 = \wishbone_bd_ram_mem2_reg[19][16]/P0001  & n13886 ;
  assign n19370 = \wishbone_bd_ram_mem2_reg[247][16]/P0001  & n13571 ;
  assign n19371 = ~n19369 & ~n19370 ;
  assign n19372 = \wishbone_bd_ram_mem2_reg[192][16]/P0001  & n13390 ;
  assign n19373 = \wishbone_bd_ram_mem2_reg[81][16]/P0001  & n13409 ;
  assign n19374 = ~n19372 & ~n19373 ;
  assign n19375 = n19371 & n19374 ;
  assign n19376 = n19368 & n19375 ;
  assign n19377 = n19361 & n19376 ;
  assign n19378 = \wishbone_bd_ram_mem2_reg[121][16]/P0001  & n13983 ;
  assign n19379 = \wishbone_bd_ram_mem2_reg[102][16]/P0001  & n13534 ;
  assign n19380 = ~n19378 & ~n19379 ;
  assign n19381 = \wishbone_bd_ram_mem2_reg[93][16]/P0001  & n13891 ;
  assign n19382 = \wishbone_bd_ram_mem2_reg[158][16]/P0001  & n13294 ;
  assign n19383 = ~n19381 & ~n19382 ;
  assign n19384 = n19380 & n19383 ;
  assign n19385 = \wishbone_bd_ram_mem2_reg[202][16]/P0001  & n13268 ;
  assign n19386 = \wishbone_bd_ram_mem2_reg[99][16]/P0001  & n13996 ;
  assign n19387 = ~n19385 & ~n19386 ;
  assign n19388 = \wishbone_bd_ram_mem2_reg[13][16]/P0001  & n13844 ;
  assign n19389 = \wishbone_bd_ram_mem2_reg[193][16]/P0001  & n14022 ;
  assign n19390 = ~n19388 & ~n19389 ;
  assign n19391 = n19387 & n19390 ;
  assign n19392 = n19384 & n19391 ;
  assign n19393 = \wishbone_bd_ram_mem2_reg[229][16]/P0001  & n13552 ;
  assign n19394 = \wishbone_bd_ram_mem2_reg[206][16]/P0001  & n13414 ;
  assign n19395 = ~n19393 & ~n19394 ;
  assign n19396 = \wishbone_bd_ram_mem2_reg[239][16]/P0001  & n13349 ;
  assign n19397 = \wishbone_bd_ram_mem2_reg[48][16]/P0001  & n13917 ;
  assign n19398 = ~n19396 & ~n19397 ;
  assign n19399 = n19395 & n19398 ;
  assign n19400 = \wishbone_bd_ram_mem2_reg[28][16]/P0001  & n13810 ;
  assign n19401 = \wishbone_bd_ram_mem2_reg[105][16]/P0001  & n13503 ;
  assign n19402 = ~n19400 & ~n19401 ;
  assign n19403 = \wishbone_bd_ram_mem2_reg[252][16]/P0001  & n13986 ;
  assign n19404 = \wishbone_bd_ram_mem2_reg[149][16]/P0001  & n13469 ;
  assign n19405 = ~n19403 & ~n19404 ;
  assign n19406 = n19402 & n19405 ;
  assign n19407 = n19399 & n19406 ;
  assign n19408 = n19392 & n19407 ;
  assign n19409 = n19377 & n19408 ;
  assign n19410 = n19346 & n19409 ;
  assign n19411 = \wishbone_bd_ram_mem2_reg[182][16]/P0001  & n13598 ;
  assign n19412 = \wishbone_bd_ram_mem2_reg[42][16]/P0001  & n13341 ;
  assign n19413 = ~n19411 & ~n19412 ;
  assign n19414 = \wishbone_bd_ram_mem2_reg[23][16]/P0001  & n13857 ;
  assign n19415 = \wishbone_bd_ram_mem2_reg[213][16]/P0001  & n13870 ;
  assign n19416 = ~n19414 & ~n19415 ;
  assign n19417 = n19413 & n19416 ;
  assign n19418 = \wishbone_bd_ram_mem2_reg[74][16]/P0001  & n13564 ;
  assign n19419 = \wishbone_bd_ram_mem2_reg[116][16]/P0001  & n13865 ;
  assign n19420 = ~n19418 & ~n19419 ;
  assign n19421 = \wishbone_bd_ram_mem2_reg[101][16]/P0001  & n13772 ;
  assign n19422 = \wishbone_bd_ram_mem2_reg[58][16]/P0001  & n13949 ;
  assign n19423 = ~n19421 & ~n19422 ;
  assign n19424 = n19420 & n19423 ;
  assign n19425 = n19417 & n19424 ;
  assign n19426 = \wishbone_bd_ram_mem2_reg[196][16]/P0001  & n13977 ;
  assign n19427 = \wishbone_bd_ram_mem2_reg[1][16]/P0001  & n13888 ;
  assign n19428 = ~n19426 & ~n19427 ;
  assign n19429 = \wishbone_bd_ram_mem2_reg[17][16]/P0001  & n13324 ;
  assign n19430 = \wishbone_bd_ram_mem2_reg[2][16]/P0001  & n13975 ;
  assign n19431 = ~n19429 & ~n19430 ;
  assign n19432 = n19428 & n19431 ;
  assign n19433 = \wishbone_bd_ram_mem2_reg[218][16]/P0001  & n13792 ;
  assign n19434 = \wishbone_bd_ram_mem2_reg[10][16]/P0001  & n13837 ;
  assign n19435 = ~n19433 & ~n19434 ;
  assign n19436 = \wishbone_bd_ram_mem2_reg[75][16]/P0001  & n13605 ;
  assign n19437 = \wishbone_bd_ram_mem2_reg[184][16]/P0001  & n13960 ;
  assign n19438 = ~n19436 & ~n19437 ;
  assign n19439 = n19435 & n19438 ;
  assign n19440 = n19432 & n19439 ;
  assign n19441 = n19425 & n19440 ;
  assign n19442 = \wishbone_bd_ram_mem2_reg[126][16]/P0001  & n13786 ;
  assign n19443 = \wishbone_bd_ram_mem2_reg[235][16]/P0001  & n13518 ;
  assign n19444 = ~n19442 & ~n19443 ;
  assign n19445 = \wishbone_bd_ram_mem2_reg[32][16]/P0001  & n13736 ;
  assign n19446 = \wishbone_bd_ram_mem2_reg[185][16]/P0001  & n13372 ;
  assign n19447 = ~n19445 & ~n19446 ;
  assign n19448 = n19444 & n19447 ;
  assign n19449 = \wishbone_bd_ram_mem2_reg[24][16]/P0001  & n13970 ;
  assign n19450 = \wishbone_bd_ram_mem2_reg[108][16]/P0001  & n13814 ;
  assign n19451 = ~n19449 & ~n19450 ;
  assign n19452 = \wishbone_bd_ram_mem2_reg[77][16]/P0001  & n13935 ;
  assign n19453 = \wishbone_bd_ram_mem2_reg[147][16]/P0001  & n13702 ;
  assign n19454 = ~n19452 & ~n19453 ;
  assign n19455 = n19451 & n19454 ;
  assign n19456 = n19448 & n19455 ;
  assign n19457 = \wishbone_bd_ram_mem2_reg[219][16]/P0001  & n13577 ;
  assign n19458 = \wishbone_bd_ram_mem2_reg[47][16]/P0001  & n13436 ;
  assign n19459 = ~n19457 & ~n19458 ;
  assign n19460 = \wishbone_bd_ram_mem2_reg[30][16]/P0001  & n13713 ;
  assign n19461 = \wishbone_bd_ram_mem2_reg[7][16]/P0001  & n13546 ;
  assign n19462 = ~n19460 & ~n19461 ;
  assign n19463 = n19459 & n19462 ;
  assign n19464 = \wishbone_bd_ram_mem2_reg[148][16]/P0001  & n13868 ;
  assign n19465 = \wishbone_bd_ram_mem2_reg[117][16]/P0001  & n13557 ;
  assign n19466 = ~n19464 & ~n19465 ;
  assign n19467 = \wishbone_bd_ram_mem2_reg[59][16]/P0001  & n13613 ;
  assign n19468 = \wishbone_bd_ram_mem2_reg[160][16]/P0001  & n13271 ;
  assign n19469 = ~n19467 & ~n19468 ;
  assign n19470 = n19466 & n19469 ;
  assign n19471 = n19463 & n19470 ;
  assign n19472 = n19456 & n19471 ;
  assign n19473 = n19441 & n19472 ;
  assign n19474 = \wishbone_bd_ram_mem2_reg[124][16]/P0001  & n14024 ;
  assign n19475 = \wishbone_bd_ram_mem2_reg[57][16]/P0001  & n13731 ;
  assign n19476 = ~n19474 & ~n19475 ;
  assign n19477 = \wishbone_bd_ram_mem2_reg[45][16]/P0001  & n13420 ;
  assign n19478 = \wishbone_bd_ram_mem2_reg[190][16]/P0001  & n13365 ;
  assign n19479 = ~n19477 & ~n19478 ;
  assign n19480 = n19476 & n19479 ;
  assign n19481 = \wishbone_bd_ram_mem2_reg[134][16]/P0001  & n13494 ;
  assign n19482 = \wishbone_bd_ram_mem2_reg[234][16]/P0001  & n13781 ;
  assign n19483 = ~n19481 & ~n19482 ;
  assign n19484 = \wishbone_bd_ram_mem2_reg[203][16]/P0001  & n13816 ;
  assign n19485 = \wishbone_bd_ram_mem2_reg[49][16]/P0001  & n13929 ;
  assign n19486 = ~n19484 & ~n19485 ;
  assign n19487 = n19483 & n19486 ;
  assign n19488 = n19480 & n19487 ;
  assign n19489 = \wishbone_bd_ram_mem2_reg[36][16]/P0001  & n13639 ;
  assign n19490 = \wishbone_bd_ram_mem2_reg[150][16]/P0001  & n13666 ;
  assign n19491 = ~n19489 & ~n19490 ;
  assign n19492 = \wishbone_bd_ram_mem2_reg[115][16]/P0001  & n13747 ;
  assign n19493 = \wishbone_bd_ram_mem2_reg[163][16]/P0001  & n13255 ;
  assign n19494 = ~n19492 & ~n19493 ;
  assign n19495 = n19491 & n19494 ;
  assign n19496 = \wishbone_bd_ram_mem2_reg[200][16]/P0001  & n13922 ;
  assign n19497 = \wishbone_bd_ram_mem2_reg[44][16]/P0001  & n13291 ;
  assign n19498 = ~n19496 & ~n19497 ;
  assign n19499 = \wishbone_bd_ram_mem2_reg[96][16]/P0001  & n13425 ;
  assign n19500 = \wishbone_bd_ram_mem2_reg[38][16]/P0001  & n13828 ;
  assign n19501 = ~n19499 & ~n19500 ;
  assign n19502 = n19498 & n19501 ;
  assign n19503 = n19495 & n19502 ;
  assign n19504 = n19488 & n19503 ;
  assign n19505 = \wishbone_bd_ram_mem2_reg[62][16]/P0001  & n13529 ;
  assign n19506 = \wishbone_bd_ram_mem2_reg[21][16]/P0001  & n13438 ;
  assign n19507 = ~n19505 & ~n19506 ;
  assign n19508 = \wishbone_bd_ram_mem2_reg[67][16]/P0001  & n13663 ;
  assign n19509 = \wishbone_bd_ram_mem2_reg[159][16]/P0001  & n13627 ;
  assign n19510 = ~n19508 & ~n19509 ;
  assign n19511 = n19507 & n19510 ;
  assign n19512 = \wishbone_bd_ram_mem2_reg[191][16]/P0001  & n14012 ;
  assign n19513 = \wishbone_bd_ram_mem2_reg[80][16]/P0001  & n13516 ;
  assign n19514 = ~n19512 & ~n19513 ;
  assign n19515 = \wishbone_bd_ram_mem2_reg[214][16]/P0001  & n13938 ;
  assign n19516 = \wishbone_bd_ram_mem2_reg[194][16]/P0001  & n13624 ;
  assign n19517 = ~n19515 & ~n19516 ;
  assign n19518 = n19514 & n19517 ;
  assign n19519 = n19511 & n19518 ;
  assign n19520 = \wishbone_bd_ram_mem2_reg[246][16]/P0001  & n13981 ;
  assign n19521 = \wishbone_bd_ram_mem2_reg[151][16]/P0001  & n13697 ;
  assign n19522 = ~n19520 & ~n19521 ;
  assign n19523 = \wishbone_bd_ram_mem2_reg[172][16]/P0001  & n13377 ;
  assign n19524 = \wishbone_bd_ram_mem2_reg[86][16]/P0001  & n13485 ;
  assign n19525 = ~n19523 & ~n19524 ;
  assign n19526 = n19522 & n19525 ;
  assign n19527 = \wishbone_bd_ram_mem2_reg[231][16]/P0001  & n13363 ;
  assign n19528 = \wishbone_bd_ram_mem2_reg[183][16]/P0001  & n13645 ;
  assign n19529 = ~n19527 & ~n19528 ;
  assign n19530 = \wishbone_bd_ram_mem2_reg[112][16]/P0001  & n13482 ;
  assign n19531 = \wishbone_bd_ram_mem2_reg[88][16]/P0001  & n13347 ;
  assign n19532 = ~n19530 & ~n19531 ;
  assign n19533 = n19529 & n19532 ;
  assign n19534 = n19526 & n19533 ;
  assign n19535 = n19519 & n19534 ;
  assign n19536 = n19504 & n19535 ;
  assign n19537 = n19473 & n19536 ;
  assign n19538 = n19410 & n19537 ;
  assign n19539 = \wishbone_bd_ram_mem2_reg[3][16]/P0001  & n13354 ;
  assign n19540 = \wishbone_bd_ram_mem2_reg[98][16]/P0001  & n13569 ;
  assign n19541 = ~n19539 & ~n19540 ;
  assign n19542 = \wishbone_bd_ram_mem2_reg[168][16]/P0001  & n13795 ;
  assign n19543 = \wishbone_bd_ram_mem2_reg[64][16]/P0001  & n13904 ;
  assign n19544 = ~n19542 & ~n19543 ;
  assign n19545 = n19541 & n19544 ;
  assign n19546 = \wishbone_bd_ram_mem2_reg[18][16]/P0001  & n13532 ;
  assign n19547 = \wishbone_bd_ram_mem2_reg[136][16]/P0001  & n13963 ;
  assign n19548 = ~n19546 & ~n19547 ;
  assign n19549 = \wishbone_bd_ram_mem2_reg[152][16]/P0001  & n13912 ;
  assign n19550 = \wishbone_bd_ram_mem2_reg[146][16]/P0001  & n13958 ;
  assign n19551 = ~n19549 & ~n19550 ;
  assign n19552 = n19548 & n19551 ;
  assign n19553 = n19545 & n19552 ;
  assign n19554 = \wishbone_bd_ram_mem2_reg[51][16]/P0001  & n13880 ;
  assign n19555 = \wishbone_bd_ram_mem2_reg[223][16]/P0001  & n13335 ;
  assign n19556 = ~n19554 & ~n19555 ;
  assign n19557 = \wishbone_bd_ram_mem2_reg[9][16]/P0001  & n13580 ;
  assign n19558 = \wishbone_bd_ram_mem2_reg[70][16]/P0001  & n13339 ;
  assign n19559 = ~n19557 & ~n19558 ;
  assign n19560 = n19556 & n19559 ;
  assign n19561 = \wishbone_bd_ram_mem2_reg[215][16]/P0001  & n13901 ;
  assign n19562 = \wishbone_bd_ram_mem2_reg[176][16]/P0001  & n13262 ;
  assign n19563 = ~n19561 & ~n19562 ;
  assign n19564 = \wishbone_bd_ram_mem2_reg[37][16]/P0001  & n13710 ;
  assign n19565 = \wishbone_bd_ram_mem2_reg[54][16]/P0001  & n13622 ;
  assign n19566 = ~n19564 & ~n19565 ;
  assign n19567 = n19563 & n19566 ;
  assign n19568 = n19560 & n19567 ;
  assign n19569 = n19553 & n19568 ;
  assign n19570 = \wishbone_bd_ram_mem2_reg[50][16]/P0001  & n13686 ;
  assign n19571 = \wishbone_bd_ram_mem2_reg[162][16]/P0001  & n13726 ;
  assign n19572 = ~n19570 & ~n19571 ;
  assign n19573 = \wishbone_bd_ram_mem2_reg[157][16]/P0001  & n13445 ;
  assign n19574 = \wishbone_bd_ram_mem2_reg[253][16]/P0001  & n13708 ;
  assign n19575 = ~n19573 & ~n19574 ;
  assign n19576 = n19572 & n19575 ;
  assign n19577 = \wishbone_bd_ram_mem2_reg[22][16]/P0001  & n13744 ;
  assign n19578 = \wishbone_bd_ram_mem2_reg[236][16]/P0001  & n13480 ;
  assign n19579 = ~n19577 & ~n19578 ;
  assign n19580 = \wishbone_bd_ram_mem2_reg[255][16]/P0001  & n13952 ;
  assign n19581 = \wishbone_bd_ram_mem2_reg[211][16]/P0001  & n13805 ;
  assign n19582 = ~n19580 & ~n19581 ;
  assign n19583 = n19579 & n19582 ;
  assign n19584 = n19576 & n19583 ;
  assign n19585 = \wishbone_bd_ram_mem2_reg[72][16]/P0001  & n13582 ;
  assign n19586 = \wishbone_bd_ram_mem2_reg[174][16]/P0001  & n13899 ;
  assign n19587 = ~n19585 & ~n19586 ;
  assign n19588 = \wishbone_bd_ram_mem2_reg[27][16]/P0001  & n13251 ;
  assign n19589 = \wishbone_bd_ram_mem2_reg[154][16]/P0001  & n13403 ;
  assign n19590 = ~n19588 & ~n19589 ;
  assign n19591 = n19587 & n19590 ;
  assign n19592 = \wishbone_bd_ram_mem2_reg[156][16]/P0001  & n13769 ;
  assign n19593 = \wishbone_bd_ram_mem2_reg[166][16]/P0001  & n13999 ;
  assign n19594 = ~n19592 & ~n19593 ;
  assign n19595 = \wishbone_bd_ram_mem2_reg[53][16]/P0001  & n13875 ;
  assign n19596 = \wishbone_bd_ram_mem2_reg[123][16]/P0001  & n13749 ;
  assign n19597 = ~n19595 & ~n19596 ;
  assign n19598 = n19594 & n19597 ;
  assign n19599 = n19591 & n19598 ;
  assign n19600 = n19584 & n19599 ;
  assign n19601 = n19569 & n19600 ;
  assign n19602 = \wishbone_bd_ram_mem2_reg[4][16]/P0001  & n13527 ;
  assign n19603 = \wishbone_bd_ram_mem2_reg[224][16]/P0001  & n13433 ;
  assign n19604 = ~n19602 & ~n19603 ;
  assign n19605 = \wishbone_bd_ram_mem2_reg[107][16]/P0001  & n13476 ;
  assign n19606 = \wishbone_bd_ram_mem2_reg[145][16]/P0001  & n13715 ;
  assign n19607 = ~n19605 & ~n19606 ;
  assign n19608 = n19604 & n19607 ;
  assign n19609 = \wishbone_bd_ram_mem2_reg[84][16]/P0001  & n13385 ;
  assign n19610 = \wishbone_bd_ram_mem2_reg[83][16]/P0001  & n13454 ;
  assign n19611 = ~n19609 & ~n19610 ;
  assign n19612 = \wishbone_bd_ram_mem2_reg[179][16]/P0001  & n14035 ;
  assign n19613 = \wishbone_bd_ram_mem2_reg[130][16]/P0001  & n13427 ;
  assign n19614 = ~n19612 & ~n19613 ;
  assign n19615 = n19611 & n19614 ;
  assign n19616 = n19608 & n19615 ;
  assign n19617 = \wishbone_bd_ram_mem2_reg[94][16]/P0001  & n13833 ;
  assign n19618 = \wishbone_bd_ram_mem2_reg[217][16]/P0001  & n13767 ;
  assign n19619 = ~n19617 & ~n19618 ;
  assign n19620 = \wishbone_bd_ram_mem2_reg[144][16]/P0001  & n13508 ;
  assign n19621 = \wishbone_bd_ram_mem2_reg[73][16]/P0001  & n13456 ;
  assign n19622 = ~n19620 & ~n19621 ;
  assign n19623 = n19619 & n19622 ;
  assign n19624 = \wishbone_bd_ram_mem2_reg[210][16]/P0001  & n13443 ;
  assign n19625 = \wishbone_bd_ram_mem2_reg[198][16]/P0001  & n13592 ;
  assign n19626 = ~n19624 & ~n19625 ;
  assign n19627 = \wishbone_bd_ram_mem2_reg[153][16]/P0001  & n13309 ;
  assign n19628 = \wishbone_bd_ram_mem2_reg[131][16]/P0001  & n13358 ;
  assign n19629 = ~n19627 & ~n19628 ;
  assign n19630 = n19626 & n19629 ;
  assign n19631 = n19623 & n19630 ;
  assign n19632 = n19616 & n19631 ;
  assign n19633 = \wishbone_bd_ram_mem2_reg[187][16]/P0001  & n13756 ;
  assign n19634 = \wishbone_bd_ram_mem2_reg[68][16]/P0001  & n13379 ;
  assign n19635 = ~n19633 & ~n19634 ;
  assign n19636 = \wishbone_bd_ram_mem2_reg[66][16]/P0001  & n13603 ;
  assign n19637 = \wishbone_bd_ram_mem2_reg[14][16]/P0001  & n13972 ;
  assign n19638 = ~n19636 & ~n19637 ;
  assign n19639 = n19635 & n19638 ;
  assign n19640 = \wishbone_bd_ram_mem2_reg[222][16]/P0001  & n13721 ;
  assign n19641 = \wishbone_bd_ram_mem2_reg[155][16]/P0001  & n13738 ;
  assign n19642 = ~n19640 & ~n19641 ;
  assign n19643 = \wishbone_bd_ram_mem2_reg[78][16]/P0001  & n13277 ;
  assign n19644 = \wishbone_bd_ram_mem2_reg[177][16]/P0001  & n13863 ;
  assign n19645 = ~n19643 & ~n19644 ;
  assign n19646 = n19642 & n19645 ;
  assign n19647 = n19639 & n19646 ;
  assign n19648 = \wishbone_bd_ram_mem2_reg[238][16]/P0001  & n13819 ;
  assign n19649 = \wishbone_bd_ram_mem2_reg[5][16]/P0001  & n13243 ;
  assign n19650 = ~n19648 & ~n19649 ;
  assign n19651 = \wishbone_bd_ram_mem2_reg[133][16]/P0001  & n13492 ;
  assign n19652 = \wishbone_bd_ram_mem2_reg[114][16]/P0001  & n13763 ;
  assign n19653 = ~n19651 & ~n19652 ;
  assign n19654 = n19650 & n19653 ;
  assign n19655 = \wishbone_bd_ram_mem2_reg[232][16]/P0001  & n13510 ;
  assign n19656 = \wishbone_bd_ram_mem2_reg[16][16]/P0001  & n13695 ;
  assign n19657 = ~n19655 & ~n19656 ;
  assign n19658 = \wishbone_bd_ram_mem2_reg[109][16]/P0001  & n13306 ;
  assign n19659 = \wishbone_bd_ram_mem2_reg[216][16]/P0001  & n14005 ;
  assign n19660 = ~n19658 & ~n19659 ;
  assign n19661 = n19657 & n19660 ;
  assign n19662 = n19654 & n19661 ;
  assign n19663 = n19647 & n19662 ;
  assign n19664 = n19632 & n19663 ;
  assign n19665 = n19601 & n19664 ;
  assign n19666 = \wishbone_bd_ram_mem2_reg[65][16]/P0001  & n13842 ;
  assign n19667 = \wishbone_bd_ram_mem2_reg[207][16]/P0001  & n13826 ;
  assign n19668 = ~n19666 & ~n19667 ;
  assign n19669 = \wishbone_bd_ram_mem2_reg[142][16]/P0001  & n13448 ;
  assign n19670 = \wishbone_bd_ram_mem2_reg[181][16]/P0001  & n13587 ;
  assign n19671 = ~n19669 & ~n19670 ;
  assign n19672 = n19668 & n19671 ;
  assign n19673 = \wishbone_bd_ram_mem2_reg[15][16]/P0001  & n13797 ;
  assign n19674 = \wishbone_bd_ram_mem2_reg[230][16]/P0001  & n13994 ;
  assign n19675 = ~n19673 & ~n19674 ;
  assign n19676 = \wishbone_bd_ram_mem2_reg[189][16]/P0001  & n14001 ;
  assign n19677 = \wishbone_bd_ram_mem2_reg[243][16]/P0001  & n13575 ;
  assign n19678 = ~n19676 & ~n19677 ;
  assign n19679 = n19675 & n19678 ;
  assign n19680 = n19672 & n19679 ;
  assign n19681 = \wishbone_bd_ram_mem2_reg[25][16]/P0001  & n13742 ;
  assign n19682 = \wishbone_bd_ram_mem2_reg[97][16]/P0001  & n13724 ;
  assign n19683 = ~n19681 & ~n19682 ;
  assign n19684 = \wishbone_bd_ram_mem2_reg[251][16]/P0001  & n14019 ;
  assign n19685 = \wishbone_bd_ram_mem2_reg[61][16]/P0001  & n13544 ;
  assign n19686 = ~n19684 & ~n19685 ;
  assign n19687 = n19683 & n19686 ;
  assign n19688 = \wishbone_bd_ram_mem2_reg[249][16]/P0001  & n13431 ;
  assign n19689 = \wishbone_bd_ram_mem2_reg[110][16]/P0001  & n14030 ;
  assign n19690 = ~n19688 & ~n19689 ;
  assign n19691 = \wishbone_bd_ram_mem2_reg[63][16]/P0001  & n13327 ;
  assign n19692 = \wishbone_bd_ram_mem2_reg[104][16]/P0001  & n13684 ;
  assign n19693 = ~n19691 & ~n19692 ;
  assign n19694 = n19690 & n19693 ;
  assign n19695 = n19687 & n19694 ;
  assign n19696 = n19680 & n19695 ;
  assign n19697 = \wishbone_bd_ram_mem2_reg[225][16]/P0001  & n13719 ;
  assign n19698 = \wishbone_bd_ram_mem2_reg[135][16]/P0001  & n13672 ;
  assign n19699 = ~n19697 & ~n19698 ;
  assign n19700 = \wishbone_bd_ram_mem2_reg[199][16]/P0001  & n13499 ;
  assign n19701 = \wishbone_bd_ram_mem2_reg[186][16]/P0001  & n13616 ;
  assign n19702 = ~n19700 & ~n19701 ;
  assign n19703 = n19699 & n19702 ;
  assign n19704 = \wishbone_bd_ram_mem2_reg[180][16]/P0001  & n13650 ;
  assign n19705 = \wishbone_bd_ram_mem2_reg[167][16]/P0001  & n13940 ;
  assign n19706 = ~n19704 & ~n19705 ;
  assign n19707 = \wishbone_bd_ram_mem2_reg[113][16]/P0001  & n13882 ;
  assign n19708 = \wishbone_bd_ram_mem2_reg[95][16]/P0001  & n13317 ;
  assign n19709 = ~n19707 & ~n19708 ;
  assign n19710 = n19706 & n19709 ;
  assign n19711 = n19703 & n19710 ;
  assign n19712 = \wishbone_bd_ram_mem2_reg[26][16]/P0001  & n13521 ;
  assign n19713 = \wishbone_bd_ram_mem2_reg[250][16]/P0001  & n13677 ;
  assign n19714 = ~n19712 & ~n19713 ;
  assign n19715 = \wishbone_bd_ram_mem2_reg[82][16]/P0001  & n13374 ;
  assign n19716 = \wishbone_bd_ram_mem2_reg[248][16]/P0001  & n13647 ;
  assign n19717 = ~n19715 & ~n19716 ;
  assign n19718 = n19714 & n19717 ;
  assign n19719 = \wishbone_bd_ram_mem2_reg[60][16]/P0001  & n13790 ;
  assign n19720 = \wishbone_bd_ram_mem2_reg[35][16]/P0001  & n13523 ;
  assign n19721 = ~n19719 & ~n19720 ;
  assign n19722 = \wishbone_bd_ram_mem2_reg[89][16]/P0001  & n13910 ;
  assign n19723 = \wishbone_bd_ram_mem2_reg[165][16]/P0001  & n14028 ;
  assign n19724 = ~n19722 & ~n19723 ;
  assign n19725 = n19721 & n19724 ;
  assign n19726 = n19718 & n19725 ;
  assign n19727 = n19711 & n19726 ;
  assign n19728 = n19696 & n19727 ;
  assign n19729 = \wishbone_bd_ram_mem2_reg[201][16]/P0001  & n13600 ;
  assign n19730 = \wishbone_bd_ram_mem2_reg[208][16]/P0001  & n14010 ;
  assign n19731 = ~n19729 & ~n19730 ;
  assign n19732 = \wishbone_bd_ram_mem2_reg[29][16]/P0001  & n13412 ;
  assign n19733 = \wishbone_bd_ram_mem2_reg[132][16]/P0001  & n13927 ;
  assign n19734 = ~n19732 & ~n19733 ;
  assign n19735 = n19731 & n19734 ;
  assign n19736 = \wishbone_bd_ram_mem2_reg[92][16]/P0001  & n13859 ;
  assign n19737 = \wishbone_bd_ram_mem2_reg[227][16]/P0001  & n13388 ;
  assign n19738 = ~n19736 & ~n19737 ;
  assign n19739 = \wishbone_bd_ram_mem2_reg[245][16]/P0001  & n13877 ;
  assign n19740 = \wishbone_bd_ram_mem2_reg[111][16]/P0001  & n13471 ;
  assign n19741 = ~n19739 & ~n19740 ;
  assign n19742 = n19738 & n19741 ;
  assign n19743 = n19735 & n19742 ;
  assign n19744 = \wishbone_bd_ram_mem2_reg[12][16]/P0001  & n13733 ;
  assign n19745 = \wishbone_bd_ram_mem2_reg[90][16]/P0001  & n13906 ;
  assign n19746 = ~n19744 & ~n19745 ;
  assign n19747 = \wishbone_bd_ram_mem2_reg[85][16]/P0001  & n13784 ;
  assign n19748 = \wishbone_bd_ram_mem2_reg[87][16]/P0001  & n13691 ;
  assign n19749 = ~n19747 & ~n19748 ;
  assign n19750 = n19746 & n19749 ;
  assign n19751 = \wishbone_bd_ram_mem2_reg[212][16]/P0001  & n13634 ;
  assign n19752 = \wishbone_bd_ram_mem2_reg[173][16]/P0001  & n13360 ;
  assign n19753 = ~n19751 & ~n19752 ;
  assign n19754 = \wishbone_bd_ram_mem2_reg[43][16]/P0001  & n13761 ;
  assign n19755 = \wishbone_bd_ram_mem2_reg[233][16]/P0001  & n13332 ;
  assign n19756 = ~n19754 & ~n19755 ;
  assign n19757 = n19753 & n19756 ;
  assign n19758 = n19750 & n19757 ;
  assign n19759 = n19743 & n19758 ;
  assign n19760 = \wishbone_bd_ram_mem2_reg[76][16]/P0001  & n13831 ;
  assign n19761 = \wishbone_bd_ram_mem2_reg[106][16]/P0001  & n13555 ;
  assign n19762 = ~n19760 & ~n19761 ;
  assign n19763 = \wishbone_bd_ram_mem2_reg[228][16]/P0001  & n13497 ;
  assign n19764 = \wishbone_bd_ram_mem2_reg[169][16]/P0001  & n13541 ;
  assign n19765 = ~n19763 & ~n19764 ;
  assign n19766 = n19762 & n19765 ;
  assign n19767 = \wishbone_bd_ram_mem2_reg[209][16]/P0001  & n13689 ;
  assign n19768 = \wishbone_bd_ram_mem2_reg[178][16]/P0001  & n13301 ;
  assign n19769 = ~n19767 & ~n19768 ;
  assign n19770 = \wishbone_bd_ram_mem2_reg[205][16]/P0001  & n13947 ;
  assign n19771 = \wishbone_bd_ram_mem2_reg[141][16]/P0001  & n13852 ;
  assign n19772 = ~n19770 & ~n19771 ;
  assign n19773 = n19769 & n19772 ;
  assign n19774 = n19766 & n19773 ;
  assign n19775 = \wishbone_bd_ram_mem2_reg[140][16]/P0001  & n13287 ;
  assign n19776 = \wishbone_bd_ram_mem2_reg[56][16]/P0001  & n13611 ;
  assign n19777 = ~n19775 & ~n19776 ;
  assign n19778 = \wishbone_bd_ram_mem2_reg[175][16]/P0001  & n13674 ;
  assign n19779 = \wishbone_bd_ram_mem2_reg[46][16]/P0001  & n13298 ;
  assign n19780 = ~n19778 & ~n19779 ;
  assign n19781 = n19777 & n19780 ;
  assign n19782 = \wishbone_bd_ram_mem2_reg[195][16]/P0001  & n13700 ;
  assign n19783 = \wishbone_bd_ram_mem2_reg[119][16]/P0001  & n14033 ;
  assign n19784 = ~n19782 & ~n19783 ;
  assign n19785 = \wishbone_bd_ram_mem2_reg[171][16]/P0001  & n13422 ;
  assign n19786 = \wishbone_bd_ram_mem2_reg[226][16]/P0001  & n13668 ;
  assign n19787 = ~n19785 & ~n19786 ;
  assign n19788 = n19784 & n19787 ;
  assign n19789 = n19781 & n19788 ;
  assign n19790 = n19774 & n19789 ;
  assign n19791 = n19759 & n19790 ;
  assign n19792 = n19728 & n19791 ;
  assign n19793 = n19665 & n19792 ;
  assign n19794 = n19538 & n19793 ;
  assign n19795 = n14047 & ~n19794 ;
  assign n19796 = ~\wishbone_TxLength_reg[0]/NET0131  & ~\wishbone_TxPointerLSB_rst_reg[0]/NET0131  ;
  assign n19797 = ~n14068 & ~n19796 ;
  assign n19798 = n14065 & n19797 ;
  assign n19799 = ~n14064 & n19798 ;
  assign n19800 = \wishbone_TxLength_reg[0]/NET0131  & ~n14049 ;
  assign n19801 = ~n14046 & n19800 ;
  assign n19802 = ~n19799 & ~n19801 ;
  assign n19803 = ~n19795 & n19802 ;
  assign n19804 = \wishbone_bd_ram_mem3_reg[128][31]/P0001  & n13652 ;
  assign n19805 = \wishbone_bd_ram_mem3_reg[68][31]/P0001  & n13379 ;
  assign n19806 = ~n19804 & ~n19805 ;
  assign n19807 = \wishbone_bd_ram_mem3_reg[52][31]/P0001  & n13988 ;
  assign n19808 = \wishbone_bd_ram_mem3_reg[7][31]/P0001  & n13546 ;
  assign n19809 = ~n19807 & ~n19808 ;
  assign n19810 = n19806 & n19809 ;
  assign n19811 = \wishbone_bd_ram_mem3_reg[184][31]/P0001  & n13960 ;
  assign n19812 = \wishbone_bd_ram_mem3_reg[139][31]/P0001  & n13566 ;
  assign n19813 = ~n19811 & ~n19812 ;
  assign n19814 = \wishbone_bd_ram_mem3_reg[39][31]/P0001  & n13893 ;
  assign n19815 = \wishbone_bd_ram_mem3_reg[220][31]/P0001  & n13965 ;
  assign n19816 = ~n19814 & ~n19815 ;
  assign n19817 = n19813 & n19816 ;
  assign n19818 = n19810 & n19817 ;
  assign n19819 = \wishbone_bd_ram_mem3_reg[226][31]/P0001  & n13668 ;
  assign n19820 = \wishbone_bd_ram_mem3_reg[247][31]/P0001  & n13571 ;
  assign n19821 = ~n19819 & ~n19820 ;
  assign n19822 = \wishbone_bd_ram_mem3_reg[85][31]/P0001  & n13784 ;
  assign n19823 = \wishbone_bd_ram_mem3_reg[193][31]/P0001  & n14022 ;
  assign n19824 = ~n19822 & ~n19823 ;
  assign n19825 = n19821 & n19824 ;
  assign n19826 = \wishbone_bd_ram_mem3_reg[66][31]/P0001  & n13603 ;
  assign n19827 = \wishbone_bd_ram_mem3_reg[227][31]/P0001  & n13388 ;
  assign n19828 = ~n19826 & ~n19827 ;
  assign n19829 = \wishbone_bd_ram_mem3_reg[25][31]/P0001  & n13742 ;
  assign n19830 = \wishbone_bd_ram_mem3_reg[180][31]/P0001  & n13650 ;
  assign n19831 = ~n19829 & ~n19830 ;
  assign n19832 = n19828 & n19831 ;
  assign n19833 = n19825 & n19832 ;
  assign n19834 = n19818 & n19833 ;
  assign n19835 = \wishbone_bd_ram_mem3_reg[89][31]/P0001  & n13910 ;
  assign n19836 = \wishbone_bd_ram_mem3_reg[186][31]/P0001  & n13616 ;
  assign n19837 = ~n19835 & ~n19836 ;
  assign n19838 = \wishbone_bd_ram_mem3_reg[13][31]/P0001  & n13844 ;
  assign n19839 = \wishbone_bd_ram_mem3_reg[93][31]/P0001  & n13891 ;
  assign n19840 = ~n19838 & ~n19839 ;
  assign n19841 = n19837 & n19840 ;
  assign n19842 = \wishbone_bd_ram_mem3_reg[240][31]/P0001  & n13352 ;
  assign n19843 = \wishbone_bd_ram_mem3_reg[185][31]/P0001  & n13372 ;
  assign n19844 = ~n19842 & ~n19843 ;
  assign n19845 = \wishbone_bd_ram_mem3_reg[15][31]/P0001  & n13797 ;
  assign n19846 = \wishbone_bd_ram_mem3_reg[17][31]/P0001  & n13324 ;
  assign n19847 = ~n19845 & ~n19846 ;
  assign n19848 = n19844 & n19847 ;
  assign n19849 = n19841 & n19848 ;
  assign n19850 = \wishbone_bd_ram_mem3_reg[121][31]/P0001  & n13983 ;
  assign n19851 = \wishbone_bd_ram_mem3_reg[187][31]/P0001  & n13756 ;
  assign n19852 = ~n19850 & ~n19851 ;
  assign n19853 = \wishbone_bd_ram_mem3_reg[245][31]/P0001  & n13877 ;
  assign n19854 = \wishbone_bd_ram_mem3_reg[72][31]/P0001  & n13582 ;
  assign n19855 = ~n19853 & ~n19854 ;
  assign n19856 = n19852 & n19855 ;
  assign n19857 = \wishbone_bd_ram_mem3_reg[69][31]/P0001  & n13487 ;
  assign n19858 = \wishbone_bd_ram_mem3_reg[179][31]/P0001  & n14035 ;
  assign n19859 = ~n19857 & ~n19858 ;
  assign n19860 = \wishbone_bd_ram_mem3_reg[107][31]/P0001  & n13476 ;
  assign n19861 = \wishbone_bd_ram_mem3_reg[254][31]/P0001  & n13283 ;
  assign n19862 = ~n19860 & ~n19861 ;
  assign n19863 = n19859 & n19862 ;
  assign n19864 = n19856 & n19863 ;
  assign n19865 = n19849 & n19864 ;
  assign n19866 = n19834 & n19865 ;
  assign n19867 = \wishbone_bd_ram_mem3_reg[235][31]/P0001  & n13518 ;
  assign n19868 = \wishbone_bd_ram_mem3_reg[218][31]/P0001  & n13792 ;
  assign n19869 = ~n19867 & ~n19868 ;
  assign n19870 = \wishbone_bd_ram_mem3_reg[132][31]/P0001  & n13927 ;
  assign n19871 = \wishbone_bd_ram_mem3_reg[0][31]/P0001  & n13539 ;
  assign n19872 = ~n19870 & ~n19871 ;
  assign n19873 = n19869 & n19872 ;
  assign n19874 = \wishbone_bd_ram_mem3_reg[173][31]/P0001  & n13360 ;
  assign n19875 = \wishbone_bd_ram_mem3_reg[57][31]/P0001  & n13731 ;
  assign n19876 = ~n19874 & ~n19875 ;
  assign n19877 = \wishbone_bd_ram_mem3_reg[238][31]/P0001  & n13819 ;
  assign n19878 = \wishbone_bd_ram_mem3_reg[189][31]/P0001  & n14001 ;
  assign n19879 = ~n19877 & ~n19878 ;
  assign n19880 = n19876 & n19879 ;
  assign n19881 = n19873 & n19880 ;
  assign n19882 = \wishbone_bd_ram_mem3_reg[88][31]/P0001  & n13347 ;
  assign n19883 = \wishbone_bd_ram_mem3_reg[14][31]/P0001  & n13972 ;
  assign n19884 = ~n19882 & ~n19883 ;
  assign n19885 = \wishbone_bd_ram_mem3_reg[155][31]/P0001  & n13738 ;
  assign n19886 = \wishbone_bd_ram_mem3_reg[210][31]/P0001  & n13443 ;
  assign n19887 = ~n19885 & ~n19886 ;
  assign n19888 = n19884 & n19887 ;
  assign n19889 = \wishbone_bd_ram_mem3_reg[232][31]/P0001  & n13510 ;
  assign n19890 = \wishbone_bd_ram_mem3_reg[221][31]/P0001  & n13641 ;
  assign n19891 = ~n19889 & ~n19890 ;
  assign n19892 = \wishbone_bd_ram_mem3_reg[34][31]/P0001  & n13450 ;
  assign n19893 = \wishbone_bd_ram_mem3_reg[239][31]/P0001  & n13349 ;
  assign n19894 = ~n19892 & ~n19893 ;
  assign n19895 = n19891 & n19894 ;
  assign n19896 = n19888 & n19895 ;
  assign n19897 = n19881 & n19896 ;
  assign n19898 = \wishbone_bd_ram_mem3_reg[82][31]/P0001  & n13374 ;
  assign n19899 = \wishbone_bd_ram_mem3_reg[103][31]/P0001  & n13320 ;
  assign n19900 = ~n19898 & ~n19899 ;
  assign n19901 = \wishbone_bd_ram_mem3_reg[145][31]/P0001  & n13715 ;
  assign n19902 = \wishbone_bd_ram_mem3_reg[104][31]/P0001  & n13684 ;
  assign n19903 = ~n19901 & ~n19902 ;
  assign n19904 = n19900 & n19903 ;
  assign n19905 = \wishbone_bd_ram_mem3_reg[216][31]/P0001  & n14005 ;
  assign n19906 = \wishbone_bd_ram_mem3_reg[170][31]/P0001  & n14007 ;
  assign n19907 = ~n19905 & ~n19906 ;
  assign n19908 = \wishbone_bd_ram_mem3_reg[28][31]/P0001  & n13810 ;
  assign n19909 = \wishbone_bd_ram_mem3_reg[42][31]/P0001  & n13341 ;
  assign n19910 = ~n19908 & ~n19909 ;
  assign n19911 = n19907 & n19910 ;
  assign n19912 = n19904 & n19911 ;
  assign n19913 = \wishbone_bd_ram_mem3_reg[111][31]/P0001  & n13471 ;
  assign n19914 = \wishbone_bd_ram_mem3_reg[60][31]/P0001  & n13790 ;
  assign n19915 = ~n19913 & ~n19914 ;
  assign n19916 = \wishbone_bd_ram_mem3_reg[71][31]/P0001  & n13636 ;
  assign n19917 = \wishbone_bd_ram_mem3_reg[119][31]/P0001  & n14033 ;
  assign n19918 = ~n19916 & ~n19917 ;
  assign n19919 = n19915 & n19918 ;
  assign n19920 = \wishbone_bd_ram_mem3_reg[55][31]/P0001  & n13618 ;
  assign n19921 = \wishbone_bd_ram_mem3_reg[51][31]/P0001  & n13880 ;
  assign n19922 = ~n19920 & ~n19921 ;
  assign n19923 = \wishbone_bd_ram_mem3_reg[30][31]/P0001  & n13713 ;
  assign n19924 = \wishbone_bd_ram_mem3_reg[144][31]/P0001  & n13508 ;
  assign n19925 = ~n19923 & ~n19924 ;
  assign n19926 = n19922 & n19925 ;
  assign n19927 = n19919 & n19926 ;
  assign n19928 = n19912 & n19927 ;
  assign n19929 = n19897 & n19928 ;
  assign n19930 = n19866 & n19929 ;
  assign n19931 = \wishbone_bd_ram_mem3_reg[160][31]/P0001  & n13271 ;
  assign n19932 = \wishbone_bd_ram_mem3_reg[234][31]/P0001  & n13781 ;
  assign n19933 = ~n19931 & ~n19932 ;
  assign n19934 = \wishbone_bd_ram_mem3_reg[183][31]/P0001  & n13645 ;
  assign n19935 = \wishbone_bd_ram_mem3_reg[182][31]/P0001  & n13598 ;
  assign n19936 = ~n19934 & ~n19935 ;
  assign n19937 = n19933 & n19936 ;
  assign n19938 = \wishbone_bd_ram_mem3_reg[113][31]/P0001  & n13882 ;
  assign n19939 = \wishbone_bd_ram_mem3_reg[94][31]/P0001  & n13833 ;
  assign n19940 = ~n19938 & ~n19939 ;
  assign n19941 = \wishbone_bd_ram_mem3_reg[47][31]/P0001  & n13436 ;
  assign n19942 = \wishbone_bd_ram_mem3_reg[37][31]/P0001  & n13710 ;
  assign n19943 = ~n19941 & ~n19942 ;
  assign n19944 = n19940 & n19943 ;
  assign n19945 = n19937 & n19944 ;
  assign n19946 = \wishbone_bd_ram_mem3_reg[105][31]/P0001  & n13503 ;
  assign n19947 = \wishbone_bd_ram_mem3_reg[45][31]/P0001  & n13420 ;
  assign n19948 = ~n19946 & ~n19947 ;
  assign n19949 = \wishbone_bd_ram_mem3_reg[172][31]/P0001  & n13377 ;
  assign n19950 = \wishbone_bd_ram_mem3_reg[200][31]/P0001  & n13922 ;
  assign n19951 = ~n19949 & ~n19950 ;
  assign n19952 = n19948 & n19951 ;
  assign n19953 = \wishbone_bd_ram_mem3_reg[228][31]/P0001  & n13497 ;
  assign n19954 = \wishbone_bd_ram_mem3_reg[118][31]/P0001  & n13589 ;
  assign n19955 = ~n19953 & ~n19954 ;
  assign n19956 = \wishbone_bd_ram_mem3_reg[230][31]/P0001  & n13994 ;
  assign n19957 = \wishbone_bd_ram_mem3_reg[202][31]/P0001  & n13268 ;
  assign n19958 = ~n19956 & ~n19957 ;
  assign n19959 = n19955 & n19958 ;
  assign n19960 = n19952 & n19959 ;
  assign n19961 = n19945 & n19960 ;
  assign n19962 = \wishbone_bd_ram_mem3_reg[157][31]/P0001  & n13445 ;
  assign n19963 = \wishbone_bd_ram_mem3_reg[244][31]/P0001  & n13474 ;
  assign n19964 = ~n19962 & ~n19963 ;
  assign n19965 = \wishbone_bd_ram_mem3_reg[84][31]/P0001  & n13385 ;
  assign n19966 = \wishbone_bd_ram_mem3_reg[109][31]/P0001  & n13306 ;
  assign n19967 = ~n19965 & ~n19966 ;
  assign n19968 = n19964 & n19967 ;
  assign n19969 = \wishbone_bd_ram_mem3_reg[67][31]/P0001  & n13663 ;
  assign n19970 = \wishbone_bd_ram_mem3_reg[38][31]/P0001  & n13828 ;
  assign n19971 = ~n19969 & ~n19970 ;
  assign n19972 = \wishbone_bd_ram_mem3_reg[58][31]/P0001  & n13949 ;
  assign n19973 = \wishbone_bd_ram_mem3_reg[143][31]/P0001  & n13461 ;
  assign n19974 = ~n19972 & ~n19973 ;
  assign n19975 = n19971 & n19974 ;
  assign n19976 = n19968 & n19975 ;
  assign n19977 = \wishbone_bd_ram_mem3_reg[43][31]/P0001  & n13761 ;
  assign n19978 = \wishbone_bd_ram_mem3_reg[133][31]/P0001  & n13492 ;
  assign n19979 = ~n19977 & ~n19978 ;
  assign n19980 = \wishbone_bd_ram_mem3_reg[161][31]/P0001  & n13505 ;
  assign n19981 = \wishbone_bd_ram_mem3_reg[48][31]/P0001  & n13917 ;
  assign n19982 = ~n19980 & ~n19981 ;
  assign n19983 = n19979 & n19982 ;
  assign n19984 = \wishbone_bd_ram_mem3_reg[192][31]/P0001  & n13390 ;
  assign n19985 = \wishbone_bd_ram_mem3_reg[190][31]/P0001  & n13365 ;
  assign n19986 = ~n19984 & ~n19985 ;
  assign n19987 = \wishbone_bd_ram_mem3_reg[242][31]/P0001  & n13383 ;
  assign n19988 = \wishbone_bd_ram_mem3_reg[87][31]/P0001  & n13691 ;
  assign n19989 = ~n19987 & ~n19988 ;
  assign n19990 = n19986 & n19989 ;
  assign n19991 = n19983 & n19990 ;
  assign n19992 = n19976 & n19991 ;
  assign n19993 = n19961 & n19992 ;
  assign n19994 = \wishbone_bd_ram_mem3_reg[41][31]/P0001  & n14017 ;
  assign n19995 = \wishbone_bd_ram_mem3_reg[241][31]/P0001  & n13854 ;
  assign n19996 = ~n19994 & ~n19995 ;
  assign n19997 = \wishbone_bd_ram_mem3_reg[171][31]/P0001  & n13422 ;
  assign n19998 = \wishbone_bd_ram_mem3_reg[197][31]/P0001  & n13594 ;
  assign n19999 = ~n19997 & ~n19998 ;
  assign n20000 = n19996 & n19999 ;
  assign n20001 = \wishbone_bd_ram_mem3_reg[203][31]/P0001  & n13816 ;
  assign n20002 = \wishbone_bd_ram_mem3_reg[252][31]/P0001  & n13986 ;
  assign n20003 = ~n20001 & ~n20002 ;
  assign n20004 = \wishbone_bd_ram_mem3_reg[3][31]/P0001  & n13354 ;
  assign n20005 = \wishbone_bd_ram_mem3_reg[149][31]/P0001  & n13469 ;
  assign n20006 = ~n20004 & ~n20005 ;
  assign n20007 = n20003 & n20006 ;
  assign n20008 = n20000 & n20007 ;
  assign n20009 = \wishbone_bd_ram_mem3_reg[191][31]/P0001  & n14012 ;
  assign n20010 = \wishbone_bd_ram_mem3_reg[29][31]/P0001  & n13412 ;
  assign n20011 = ~n20009 & ~n20010 ;
  assign n20012 = \wishbone_bd_ram_mem3_reg[188][31]/P0001  & n13407 ;
  assign n20013 = \wishbone_bd_ram_mem3_reg[127][31]/P0001  & n13803 ;
  assign n20014 = ~n20012 & ~n20013 ;
  assign n20015 = n20011 & n20014 ;
  assign n20016 = \wishbone_bd_ram_mem3_reg[174][31]/P0001  & n13899 ;
  assign n20017 = \wishbone_bd_ram_mem3_reg[248][31]/P0001  & n13647 ;
  assign n20018 = ~n20016 & ~n20017 ;
  assign n20019 = \wishbone_bd_ram_mem3_reg[168][31]/P0001  & n13795 ;
  assign n20020 = \wishbone_bd_ram_mem3_reg[150][31]/P0001  & n13666 ;
  assign n20021 = ~n20019 & ~n20020 ;
  assign n20022 = n20018 & n20021 ;
  assign n20023 = n20015 & n20022 ;
  assign n20024 = n20008 & n20023 ;
  assign n20025 = \wishbone_bd_ram_mem3_reg[135][31]/P0001  & n13672 ;
  assign n20026 = \wishbone_bd_ram_mem3_reg[136][31]/P0001  & n13963 ;
  assign n20027 = ~n20025 & ~n20026 ;
  assign n20028 = \wishbone_bd_ram_mem3_reg[97][31]/P0001  & n13724 ;
  assign n20029 = \wishbone_bd_ram_mem3_reg[70][31]/P0001  & n13339 ;
  assign n20030 = ~n20028 & ~n20029 ;
  assign n20031 = n20027 & n20030 ;
  assign n20032 = \wishbone_bd_ram_mem3_reg[9][31]/P0001  & n13580 ;
  assign n20033 = \wishbone_bd_ram_mem3_reg[217][31]/P0001  & n13767 ;
  assign n20034 = ~n20032 & ~n20033 ;
  assign n20035 = \wishbone_bd_ram_mem3_reg[32][31]/P0001  & n13736 ;
  assign n20036 = \wishbone_bd_ram_mem3_reg[53][31]/P0001  & n13875 ;
  assign n20037 = ~n20035 & ~n20036 ;
  assign n20038 = n20034 & n20037 ;
  assign n20039 = n20031 & n20038 ;
  assign n20040 = \wishbone_bd_ram_mem3_reg[204][31]/P0001  & n13821 ;
  assign n20041 = \wishbone_bd_ram_mem3_reg[81][31]/P0001  & n13409 ;
  assign n20042 = ~n20040 & ~n20041 ;
  assign n20043 = \wishbone_bd_ram_mem3_reg[159][31]/P0001  & n13627 ;
  assign n20044 = \wishbone_bd_ram_mem3_reg[233][31]/P0001  & n13332 ;
  assign n20045 = ~n20043 & ~n20044 ;
  assign n20046 = n20042 & n20045 ;
  assign n20047 = \wishbone_bd_ram_mem3_reg[205][31]/P0001  & n13947 ;
  assign n20048 = \wishbone_bd_ram_mem3_reg[215][31]/P0001  & n13901 ;
  assign n20049 = ~n20047 & ~n20048 ;
  assign n20050 = \wishbone_bd_ram_mem3_reg[98][31]/P0001  & n13569 ;
  assign n20051 = \wishbone_bd_ram_mem3_reg[49][31]/P0001  & n13929 ;
  assign n20052 = ~n20050 & ~n20051 ;
  assign n20053 = n20049 & n20052 ;
  assign n20054 = n20046 & n20053 ;
  assign n20055 = n20039 & n20054 ;
  assign n20056 = n20024 & n20055 ;
  assign n20057 = n19993 & n20056 ;
  assign n20058 = n19930 & n20057 ;
  assign n20059 = \wishbone_bd_ram_mem3_reg[44][31]/P0001  & n13291 ;
  assign n20060 = \wishbone_bd_ram_mem3_reg[33][31]/P0001  & n13933 ;
  assign n20061 = ~n20059 & ~n20060 ;
  assign n20062 = \wishbone_bd_ram_mem3_reg[167][31]/P0001  & n13940 ;
  assign n20063 = \wishbone_bd_ram_mem3_reg[178][31]/P0001  & n13301 ;
  assign n20064 = ~n20062 & ~n20063 ;
  assign n20065 = n20061 & n20064 ;
  assign n20066 = \wishbone_bd_ram_mem3_reg[61][31]/P0001  & n13544 ;
  assign n20067 = \wishbone_bd_ram_mem3_reg[27][31]/P0001  & n13251 ;
  assign n20068 = ~n20066 & ~n20067 ;
  assign n20069 = \wishbone_bd_ram_mem3_reg[207][31]/P0001  & n13826 ;
  assign n20070 = \wishbone_bd_ram_mem3_reg[116][31]/P0001  & n13865 ;
  assign n20071 = ~n20069 & ~n20070 ;
  assign n20072 = n20068 & n20071 ;
  assign n20073 = n20065 & n20072 ;
  assign n20074 = \wishbone_bd_ram_mem3_reg[125][31]/P0001  & n13396 ;
  assign n20075 = \wishbone_bd_ram_mem3_reg[40][31]/P0001  & n13661 ;
  assign n20076 = ~n20074 & ~n20075 ;
  assign n20077 = \wishbone_bd_ram_mem3_reg[224][31]/P0001  & n13433 ;
  assign n20078 = \wishbone_bd_ram_mem3_reg[101][31]/P0001  & n13772 ;
  assign n20079 = ~n20077 & ~n20078 ;
  assign n20080 = n20076 & n20079 ;
  assign n20081 = \wishbone_bd_ram_mem3_reg[56][31]/P0001  & n13611 ;
  assign n20082 = \wishbone_bd_ram_mem3_reg[120][31]/P0001  & n13550 ;
  assign n20083 = ~n20081 & ~n20082 ;
  assign n20084 = \wishbone_bd_ram_mem3_reg[112][31]/P0001  & n13482 ;
  assign n20085 = \wishbone_bd_ram_mem3_reg[19][31]/P0001  & n13886 ;
  assign n20086 = ~n20084 & ~n20085 ;
  assign n20087 = n20083 & n20086 ;
  assign n20088 = n20080 & n20087 ;
  assign n20089 = n20073 & n20088 ;
  assign n20090 = \wishbone_bd_ram_mem3_reg[229][31]/P0001  & n13552 ;
  assign n20091 = \wishbone_bd_ram_mem3_reg[12][31]/P0001  & n13733 ;
  assign n20092 = ~n20090 & ~n20091 ;
  assign n20093 = \wishbone_bd_ram_mem3_reg[21][31]/P0001  & n13438 ;
  assign n20094 = \wishbone_bd_ram_mem3_reg[166][31]/P0001  & n13999 ;
  assign n20095 = ~n20093 & ~n20094 ;
  assign n20096 = n20092 & n20095 ;
  assign n20097 = \wishbone_bd_ram_mem3_reg[219][31]/P0001  & n13577 ;
  assign n20098 = \wishbone_bd_ram_mem3_reg[169][31]/P0001  & n13541 ;
  assign n20099 = ~n20097 & ~n20098 ;
  assign n20100 = \wishbone_bd_ram_mem3_reg[91][31]/P0001  & n13954 ;
  assign n20101 = \wishbone_bd_ram_mem3_reg[222][31]/P0001  & n13721 ;
  assign n20102 = ~n20100 & ~n20101 ;
  assign n20103 = n20099 & n20102 ;
  assign n20104 = n20096 & n20103 ;
  assign n20105 = \wishbone_bd_ram_mem3_reg[77][31]/P0001  & n13935 ;
  assign n20106 = \wishbone_bd_ram_mem3_reg[24][31]/P0001  & n13970 ;
  assign n20107 = ~n20105 & ~n20106 ;
  assign n20108 = \wishbone_bd_ram_mem3_reg[74][31]/P0001  & n13564 ;
  assign n20109 = \wishbone_bd_ram_mem3_reg[76][31]/P0001  & n13831 ;
  assign n20110 = ~n20108 & ~n20109 ;
  assign n20111 = n20107 & n20110 ;
  assign n20112 = \wishbone_bd_ram_mem3_reg[22][31]/P0001  & n13744 ;
  assign n20113 = \wishbone_bd_ram_mem3_reg[6][31]/P0001  & n13915 ;
  assign n20114 = ~n20112 & ~n20113 ;
  assign n20115 = \wishbone_bd_ram_mem3_reg[35][31]/P0001  & n13523 ;
  assign n20116 = \wishbone_bd_ram_mem3_reg[165][31]/P0001  & n14028 ;
  assign n20117 = ~n20115 & ~n20116 ;
  assign n20118 = n20114 & n20117 ;
  assign n20119 = n20111 & n20118 ;
  assign n20120 = n20104 & n20119 ;
  assign n20121 = n20089 & n20120 ;
  assign n20122 = \wishbone_bd_ram_mem3_reg[251][31]/P0001  & n14019 ;
  assign n20123 = \wishbone_bd_ram_mem3_reg[73][31]/P0001  & n13456 ;
  assign n20124 = ~n20122 & ~n20123 ;
  assign n20125 = \wishbone_bd_ram_mem3_reg[2][31]/P0001  & n13975 ;
  assign n20126 = \wishbone_bd_ram_mem3_reg[236][31]/P0001  & n13480 ;
  assign n20127 = ~n20125 & ~n20126 ;
  assign n20128 = n20124 & n20127 ;
  assign n20129 = \wishbone_bd_ram_mem3_reg[249][31]/P0001  & n13431 ;
  assign n20130 = \wishbone_bd_ram_mem3_reg[177][31]/P0001  & n13863 ;
  assign n20131 = ~n20129 & ~n20130 ;
  assign n20132 = \wishbone_bd_ram_mem3_reg[92][31]/P0001  & n13859 ;
  assign n20133 = \wishbone_bd_ram_mem3_reg[83][31]/P0001  & n13454 ;
  assign n20134 = ~n20132 & ~n20133 ;
  assign n20135 = n20131 & n20134 ;
  assign n20136 = n20128 & n20135 ;
  assign n20137 = \wishbone_bd_ram_mem3_reg[18][31]/P0001  & n13532 ;
  assign n20138 = \wishbone_bd_ram_mem3_reg[110][31]/P0001  & n14030 ;
  assign n20139 = ~n20137 & ~n20138 ;
  assign n20140 = \wishbone_bd_ram_mem3_reg[148][31]/P0001  & n13868 ;
  assign n20141 = \wishbone_bd_ram_mem3_reg[175][31]/P0001  & n13674 ;
  assign n20142 = ~n20140 & ~n20141 ;
  assign n20143 = n20139 & n20142 ;
  assign n20144 = \wishbone_bd_ram_mem3_reg[131][31]/P0001  & n13358 ;
  assign n20145 = \wishbone_bd_ram_mem3_reg[100][31]/P0001  & n13401 ;
  assign n20146 = ~n20144 & ~n20145 ;
  assign n20147 = \wishbone_bd_ram_mem3_reg[152][31]/P0001  & n13912 ;
  assign n20148 = \wishbone_bd_ram_mem3_reg[163][31]/P0001  & n13255 ;
  assign n20149 = ~n20147 & ~n20148 ;
  assign n20150 = n20146 & n20149 ;
  assign n20151 = n20143 & n20150 ;
  assign n20152 = n20136 & n20151 ;
  assign n20153 = \wishbone_bd_ram_mem3_reg[199][31]/P0001  & n13499 ;
  assign n20154 = \wishbone_bd_ram_mem3_reg[114][31]/P0001  & n13763 ;
  assign n20155 = ~n20153 & ~n20154 ;
  assign n20156 = \wishbone_bd_ram_mem3_reg[138][31]/P0001  & n13398 ;
  assign n20157 = \wishbone_bd_ram_mem3_reg[10][31]/P0001  & n13837 ;
  assign n20158 = ~n20156 & ~n20157 ;
  assign n20159 = n20155 & n20158 ;
  assign n20160 = \wishbone_bd_ram_mem3_reg[90][31]/P0001  & n13906 ;
  assign n20161 = \wishbone_bd_ram_mem3_reg[140][31]/P0001  & n13287 ;
  assign n20162 = ~n20160 & ~n20161 ;
  assign n20163 = \wishbone_bd_ram_mem3_reg[253][31]/P0001  & n13708 ;
  assign n20164 = \wishbone_bd_ram_mem3_reg[223][31]/P0001  & n13335 ;
  assign n20165 = ~n20163 & ~n20164 ;
  assign n20166 = n20162 & n20165 ;
  assign n20167 = n20159 & n20166 ;
  assign n20168 = \wishbone_bd_ram_mem3_reg[246][31]/P0001  & n13981 ;
  assign n20169 = \wishbone_bd_ram_mem3_reg[80][31]/P0001  & n13516 ;
  assign n20170 = ~n20168 & ~n20169 ;
  assign n20171 = \wishbone_bd_ram_mem3_reg[147][31]/P0001  & n13702 ;
  assign n20172 = \wishbone_bd_ram_mem3_reg[237][31]/P0001  & n13924 ;
  assign n20173 = ~n20171 & ~n20172 ;
  assign n20174 = n20170 & n20173 ;
  assign n20175 = \wishbone_bd_ram_mem3_reg[75][31]/P0001  & n13605 ;
  assign n20176 = \wishbone_bd_ram_mem3_reg[164][31]/P0001  & n13236 ;
  assign n20177 = ~n20175 & ~n20176 ;
  assign n20178 = \wishbone_bd_ram_mem3_reg[50][31]/P0001  & n13686 ;
  assign n20179 = \wishbone_bd_ram_mem3_reg[1][31]/P0001  & n13888 ;
  assign n20180 = ~n20178 & ~n20179 ;
  assign n20181 = n20177 & n20180 ;
  assign n20182 = n20174 & n20181 ;
  assign n20183 = n20167 & n20182 ;
  assign n20184 = n20152 & n20183 ;
  assign n20185 = n20121 & n20184 ;
  assign n20186 = \wishbone_bd_ram_mem3_reg[64][31]/P0001  & n13904 ;
  assign n20187 = \wishbone_bd_ram_mem3_reg[196][31]/P0001  & n13977 ;
  assign n20188 = ~n20186 & ~n20187 ;
  assign n20189 = \wishbone_bd_ram_mem3_reg[59][31]/P0001  & n13613 ;
  assign n20190 = \wishbone_bd_ram_mem3_reg[123][31]/P0001  & n13749 ;
  assign n20191 = ~n20189 & ~n20190 ;
  assign n20192 = n20188 & n20191 ;
  assign n20193 = \wishbone_bd_ram_mem3_reg[108][31]/P0001  & n13814 ;
  assign n20194 = \wishbone_bd_ram_mem3_reg[137][31]/P0001  & n13808 ;
  assign n20195 = ~n20193 & ~n20194 ;
  assign n20196 = \wishbone_bd_ram_mem3_reg[62][31]/P0001  & n13529 ;
  assign n20197 = \wishbone_bd_ram_mem3_reg[206][31]/P0001  & n13414 ;
  assign n20198 = ~n20196 & ~n20197 ;
  assign n20199 = n20195 & n20198 ;
  assign n20200 = n20192 & n20199 ;
  assign n20201 = \wishbone_bd_ram_mem3_reg[117][31]/P0001  & n13557 ;
  assign n20202 = \wishbone_bd_ram_mem3_reg[181][31]/P0001  & n13587 ;
  assign n20203 = ~n20201 & ~n20202 ;
  assign n20204 = \wishbone_bd_ram_mem3_reg[46][31]/P0001  & n13298 ;
  assign n20205 = \wishbone_bd_ram_mem3_reg[201][31]/P0001  & n13600 ;
  assign n20206 = ~n20204 & ~n20205 ;
  assign n20207 = n20203 & n20206 ;
  assign n20208 = \wishbone_bd_ram_mem3_reg[31][31]/P0001  & n13758 ;
  assign n20209 = \wishbone_bd_ram_mem3_reg[16][31]/P0001  & n13695 ;
  assign n20210 = ~n20208 & ~n20209 ;
  assign n20211 = \wishbone_bd_ram_mem3_reg[54][31]/P0001  & n13622 ;
  assign n20212 = \wishbone_bd_ram_mem3_reg[86][31]/P0001  & n13485 ;
  assign n20213 = ~n20211 & ~n20212 ;
  assign n20214 = n20210 & n20213 ;
  assign n20215 = n20207 & n20214 ;
  assign n20216 = n20200 & n20215 ;
  assign n20217 = \wishbone_bd_ram_mem3_reg[156][31]/P0001  & n13769 ;
  assign n20218 = \wishbone_bd_ram_mem3_reg[36][31]/P0001  & n13639 ;
  assign n20219 = ~n20217 & ~n20218 ;
  assign n20220 = \wishbone_bd_ram_mem3_reg[78][31]/P0001  & n13277 ;
  assign n20221 = \wishbone_bd_ram_mem3_reg[231][31]/P0001  & n13363 ;
  assign n20222 = ~n20220 & ~n20221 ;
  assign n20223 = n20219 & n20222 ;
  assign n20224 = \wishbone_bd_ram_mem3_reg[153][31]/P0001  & n13309 ;
  assign n20225 = \wishbone_bd_ram_mem3_reg[134][31]/P0001  & n13494 ;
  assign n20226 = ~n20224 & ~n20225 ;
  assign n20227 = \wishbone_bd_ram_mem3_reg[23][31]/P0001  & n13857 ;
  assign n20228 = \wishbone_bd_ram_mem3_reg[11][31]/P0001  & n13774 ;
  assign n20229 = ~n20227 & ~n20228 ;
  assign n20230 = n20226 & n20229 ;
  assign n20231 = n20223 & n20230 ;
  assign n20232 = \wishbone_bd_ram_mem3_reg[243][31]/P0001  & n13575 ;
  assign n20233 = \wishbone_bd_ram_mem3_reg[158][31]/P0001  & n13294 ;
  assign n20234 = ~n20232 & ~n20233 ;
  assign n20235 = \wishbone_bd_ram_mem3_reg[162][31]/P0001  & n13726 ;
  assign n20236 = \wishbone_bd_ram_mem3_reg[26][31]/P0001  & n13521 ;
  assign n20237 = ~n20235 & ~n20236 ;
  assign n20238 = n20234 & n20237 ;
  assign n20239 = \wishbone_bd_ram_mem3_reg[142][31]/P0001  & n13448 ;
  assign n20240 = \wishbone_bd_ram_mem3_reg[20][31]/P0001  & n13839 ;
  assign n20241 = ~n20239 & ~n20240 ;
  assign n20242 = \wishbone_bd_ram_mem3_reg[194][31]/P0001  & n13624 ;
  assign n20243 = \wishbone_bd_ram_mem3_reg[63][31]/P0001  & n13327 ;
  assign n20244 = ~n20242 & ~n20243 ;
  assign n20245 = n20241 & n20244 ;
  assign n20246 = n20238 & n20245 ;
  assign n20247 = n20231 & n20246 ;
  assign n20248 = n20216 & n20247 ;
  assign n20249 = \wishbone_bd_ram_mem3_reg[212][31]/P0001  & n13634 ;
  assign n20250 = \wishbone_bd_ram_mem3_reg[5][31]/P0001  & n13243 ;
  assign n20251 = ~n20249 & ~n20250 ;
  assign n20252 = \wishbone_bd_ram_mem3_reg[106][31]/P0001  & n13555 ;
  assign n20253 = \wishbone_bd_ram_mem3_reg[154][31]/P0001  & n13403 ;
  assign n20254 = ~n20252 & ~n20253 ;
  assign n20255 = n20251 & n20254 ;
  assign n20256 = \wishbone_bd_ram_mem3_reg[95][31]/P0001  & n13317 ;
  assign n20257 = \wishbone_bd_ram_mem3_reg[195][31]/P0001  & n13700 ;
  assign n20258 = ~n20256 & ~n20257 ;
  assign n20259 = \wishbone_bd_ram_mem3_reg[99][31]/P0001  & n13996 ;
  assign n20260 = \wishbone_bd_ram_mem3_reg[211][31]/P0001  & n13805 ;
  assign n20261 = ~n20259 & ~n20260 ;
  assign n20262 = n20258 & n20261 ;
  assign n20263 = n20255 & n20262 ;
  assign n20264 = \wishbone_bd_ram_mem3_reg[65][31]/P0001  & n13842 ;
  assign n20265 = \wishbone_bd_ram_mem3_reg[115][31]/P0001  & n13747 ;
  assign n20266 = ~n20264 & ~n20265 ;
  assign n20267 = \wishbone_bd_ram_mem3_reg[79][31]/P0001  & n13779 ;
  assign n20268 = \wishbone_bd_ram_mem3_reg[124][31]/P0001  & n14024 ;
  assign n20269 = ~n20267 & ~n20268 ;
  assign n20270 = n20266 & n20269 ;
  assign n20271 = \wishbone_bd_ram_mem3_reg[213][31]/P0001  & n13870 ;
  assign n20272 = \wishbone_bd_ram_mem3_reg[96][31]/P0001  & n13425 ;
  assign n20273 = ~n20271 & ~n20272 ;
  assign n20274 = \wishbone_bd_ram_mem3_reg[214][31]/P0001  & n13938 ;
  assign n20275 = \wishbone_bd_ram_mem3_reg[4][31]/P0001  & n13527 ;
  assign n20276 = ~n20274 & ~n20275 ;
  assign n20277 = n20273 & n20276 ;
  assign n20278 = n20270 & n20277 ;
  assign n20279 = n20263 & n20278 ;
  assign n20280 = \wishbone_bd_ram_mem3_reg[151][31]/P0001  & n13697 ;
  assign n20281 = \wishbone_bd_ram_mem3_reg[208][31]/P0001  & n14010 ;
  assign n20282 = ~n20280 & ~n20281 ;
  assign n20283 = \wishbone_bd_ram_mem3_reg[130][31]/P0001  & n13427 ;
  assign n20284 = \wishbone_bd_ram_mem3_reg[102][31]/P0001  & n13534 ;
  assign n20285 = ~n20283 & ~n20284 ;
  assign n20286 = n20282 & n20285 ;
  assign n20287 = \wishbone_bd_ram_mem3_reg[225][31]/P0001  & n13719 ;
  assign n20288 = \wishbone_bd_ram_mem3_reg[255][31]/P0001  & n13952 ;
  assign n20289 = ~n20287 & ~n20288 ;
  assign n20290 = \wishbone_bd_ram_mem3_reg[122][31]/P0001  & n13679 ;
  assign n20291 = \wishbone_bd_ram_mem3_reg[126][31]/P0001  & n13786 ;
  assign n20292 = ~n20290 & ~n20291 ;
  assign n20293 = n20289 & n20292 ;
  assign n20294 = n20286 & n20293 ;
  assign n20295 = \wishbone_bd_ram_mem3_reg[141][31]/P0001  & n13852 ;
  assign n20296 = \wishbone_bd_ram_mem3_reg[250][31]/P0001  & n13677 ;
  assign n20297 = ~n20295 & ~n20296 ;
  assign n20298 = \wishbone_bd_ram_mem3_reg[176][31]/P0001  & n13262 ;
  assign n20299 = \wishbone_bd_ram_mem3_reg[198][31]/P0001  & n13592 ;
  assign n20300 = ~n20298 & ~n20299 ;
  assign n20301 = n20297 & n20300 ;
  assign n20302 = \wishbone_bd_ram_mem3_reg[129][31]/P0001  & n13629 ;
  assign n20303 = \wishbone_bd_ram_mem3_reg[146][31]/P0001  & n13958 ;
  assign n20304 = ~n20302 & ~n20303 ;
  assign n20305 = \wishbone_bd_ram_mem3_reg[8][31]/P0001  & n13459 ;
  assign n20306 = \wishbone_bd_ram_mem3_reg[209][31]/P0001  & n13689 ;
  assign n20307 = ~n20305 & ~n20306 ;
  assign n20308 = n20304 & n20307 ;
  assign n20309 = n20301 & n20308 ;
  assign n20310 = n20294 & n20309 ;
  assign n20311 = n20279 & n20310 ;
  assign n20312 = n20248 & n20311 ;
  assign n20313 = n20185 & n20312 ;
  assign n20314 = n20058 & n20313 ;
  assign n20315 = ~wb_rst_i_pad & ~n20314 ;
  assign n20316 = n14046 & ~n20315 ;
  assign n20317 = ~\wishbone_TxLength_reg[15]/NET0131  & ~n14046 ;
  assign n20318 = n14060 & n14061 ;
  assign n20319 = ~n14046 & n20318 ;
  assign n20320 = n17919 & n20319 ;
  assign n20321 = ~n20317 & ~n20320 ;
  assign n20322 = ~n20316 & n20321 ;
  assign n20323 = \wishbone_bd_ram_mem2_reg[173][17]/P0001  & n13360 ;
  assign n20324 = \wishbone_bd_ram_mem2_reg[105][17]/P0001  & n13503 ;
  assign n20325 = ~n20323 & ~n20324 ;
  assign n20326 = \wishbone_bd_ram_mem2_reg[212][17]/P0001  & n13634 ;
  assign n20327 = \wishbone_bd_ram_mem2_reg[209][17]/P0001  & n13689 ;
  assign n20328 = ~n20326 & ~n20327 ;
  assign n20329 = n20325 & n20328 ;
  assign n20330 = \wishbone_bd_ram_mem2_reg[13][17]/P0001  & n13844 ;
  assign n20331 = \wishbone_bd_ram_mem2_reg[12][17]/P0001  & n13733 ;
  assign n20332 = ~n20330 & ~n20331 ;
  assign n20333 = \wishbone_bd_ram_mem2_reg[51][17]/P0001  & n13880 ;
  assign n20334 = \wishbone_bd_ram_mem2_reg[183][17]/P0001  & n13645 ;
  assign n20335 = ~n20333 & ~n20334 ;
  assign n20336 = n20332 & n20335 ;
  assign n20337 = n20329 & n20336 ;
  assign n20338 = \wishbone_bd_ram_mem2_reg[161][17]/P0001  & n13505 ;
  assign n20339 = \wishbone_bd_ram_mem2_reg[33][17]/P0001  & n13933 ;
  assign n20340 = ~n20338 & ~n20339 ;
  assign n20341 = \wishbone_bd_ram_mem2_reg[76][17]/P0001  & n13831 ;
  assign n20342 = \wishbone_bd_ram_mem2_reg[57][17]/P0001  & n13731 ;
  assign n20343 = ~n20341 & ~n20342 ;
  assign n20344 = n20340 & n20343 ;
  assign n20345 = \wishbone_bd_ram_mem2_reg[213][17]/P0001  & n13870 ;
  assign n20346 = \wishbone_bd_ram_mem2_reg[166][17]/P0001  & n13999 ;
  assign n20347 = ~n20345 & ~n20346 ;
  assign n20348 = \wishbone_bd_ram_mem2_reg[117][17]/P0001  & n13557 ;
  assign n20349 = \wishbone_bd_ram_mem2_reg[23][17]/P0001  & n13857 ;
  assign n20350 = ~n20348 & ~n20349 ;
  assign n20351 = n20347 & n20350 ;
  assign n20352 = n20344 & n20351 ;
  assign n20353 = n20337 & n20352 ;
  assign n20354 = \wishbone_bd_ram_mem2_reg[143][17]/P0001  & n13461 ;
  assign n20355 = \wishbone_bd_ram_mem2_reg[102][17]/P0001  & n13534 ;
  assign n20356 = ~n20354 & ~n20355 ;
  assign n20357 = \wishbone_bd_ram_mem2_reg[90][17]/P0001  & n13906 ;
  assign n20358 = \wishbone_bd_ram_mem2_reg[176][17]/P0001  & n13262 ;
  assign n20359 = ~n20357 & ~n20358 ;
  assign n20360 = n20356 & n20359 ;
  assign n20361 = \wishbone_bd_ram_mem2_reg[22][17]/P0001  & n13744 ;
  assign n20362 = \wishbone_bd_ram_mem2_reg[84][17]/P0001  & n13385 ;
  assign n20363 = ~n20361 & ~n20362 ;
  assign n20364 = \wishbone_bd_ram_mem2_reg[60][17]/P0001  & n13790 ;
  assign n20365 = \wishbone_bd_ram_mem2_reg[10][17]/P0001  & n13837 ;
  assign n20366 = ~n20364 & ~n20365 ;
  assign n20367 = n20363 & n20366 ;
  assign n20368 = n20360 & n20367 ;
  assign n20369 = \wishbone_bd_ram_mem2_reg[9][17]/P0001  & n13580 ;
  assign n20370 = \wishbone_bd_ram_mem2_reg[234][17]/P0001  & n13781 ;
  assign n20371 = ~n20369 & ~n20370 ;
  assign n20372 = \wishbone_bd_ram_mem2_reg[168][17]/P0001  & n13795 ;
  assign n20373 = \wishbone_bd_ram_mem2_reg[231][17]/P0001  & n13363 ;
  assign n20374 = ~n20372 & ~n20373 ;
  assign n20375 = n20371 & n20374 ;
  assign n20376 = \wishbone_bd_ram_mem2_reg[19][17]/P0001  & n13886 ;
  assign n20377 = \wishbone_bd_ram_mem2_reg[243][17]/P0001  & n13575 ;
  assign n20378 = ~n20376 & ~n20377 ;
  assign n20379 = \wishbone_bd_ram_mem2_reg[122][17]/P0001  & n13679 ;
  assign n20380 = \wishbone_bd_ram_mem2_reg[34][17]/P0001  & n13450 ;
  assign n20381 = ~n20379 & ~n20380 ;
  assign n20382 = n20378 & n20381 ;
  assign n20383 = n20375 & n20382 ;
  assign n20384 = n20368 & n20383 ;
  assign n20385 = n20353 & n20384 ;
  assign n20386 = \wishbone_bd_ram_mem2_reg[146][17]/P0001  & n13958 ;
  assign n20387 = \wishbone_bd_ram_mem2_reg[15][17]/P0001  & n13797 ;
  assign n20388 = ~n20386 & ~n20387 ;
  assign n20389 = \wishbone_bd_ram_mem2_reg[44][17]/P0001  & n13291 ;
  assign n20390 = \wishbone_bd_ram_mem2_reg[64][17]/P0001  & n13904 ;
  assign n20391 = ~n20389 & ~n20390 ;
  assign n20392 = n20388 & n20391 ;
  assign n20393 = \wishbone_bd_ram_mem2_reg[119][17]/P0001  & n14033 ;
  assign n20394 = \wishbone_bd_ram_mem2_reg[214][17]/P0001  & n13938 ;
  assign n20395 = ~n20393 & ~n20394 ;
  assign n20396 = \wishbone_bd_ram_mem2_reg[96][17]/P0001  & n13425 ;
  assign n20397 = \wishbone_bd_ram_mem2_reg[92][17]/P0001  & n13859 ;
  assign n20398 = ~n20396 & ~n20397 ;
  assign n20399 = n20395 & n20398 ;
  assign n20400 = n20392 & n20399 ;
  assign n20401 = \wishbone_bd_ram_mem2_reg[253][17]/P0001  & n13708 ;
  assign n20402 = \wishbone_bd_ram_mem2_reg[132][17]/P0001  & n13927 ;
  assign n20403 = ~n20401 & ~n20402 ;
  assign n20404 = \wishbone_bd_ram_mem2_reg[149][17]/P0001  & n13469 ;
  assign n20405 = \wishbone_bd_ram_mem2_reg[124][17]/P0001  & n14024 ;
  assign n20406 = ~n20404 & ~n20405 ;
  assign n20407 = n20403 & n20406 ;
  assign n20408 = \wishbone_bd_ram_mem2_reg[63][17]/P0001  & n13327 ;
  assign n20409 = \wishbone_bd_ram_mem2_reg[69][17]/P0001  & n13487 ;
  assign n20410 = ~n20408 & ~n20409 ;
  assign n20411 = \wishbone_bd_ram_mem2_reg[85][17]/P0001  & n13784 ;
  assign n20412 = \wishbone_bd_ram_mem2_reg[229][17]/P0001  & n13552 ;
  assign n20413 = ~n20411 & ~n20412 ;
  assign n20414 = n20410 & n20413 ;
  assign n20415 = n20407 & n20414 ;
  assign n20416 = n20400 & n20415 ;
  assign n20417 = \wishbone_bd_ram_mem2_reg[49][17]/P0001  & n13929 ;
  assign n20418 = \wishbone_bd_ram_mem2_reg[107][17]/P0001  & n13476 ;
  assign n20419 = ~n20417 & ~n20418 ;
  assign n20420 = \wishbone_bd_ram_mem2_reg[184][17]/P0001  & n13960 ;
  assign n20421 = \wishbone_bd_ram_mem2_reg[97][17]/P0001  & n13724 ;
  assign n20422 = ~n20420 & ~n20421 ;
  assign n20423 = n20419 & n20422 ;
  assign n20424 = \wishbone_bd_ram_mem2_reg[134][17]/P0001  & n13494 ;
  assign n20425 = \wishbone_bd_ram_mem2_reg[93][17]/P0001  & n13891 ;
  assign n20426 = ~n20424 & ~n20425 ;
  assign n20427 = \wishbone_bd_ram_mem2_reg[56][17]/P0001  & n13611 ;
  assign n20428 = \wishbone_bd_ram_mem2_reg[133][17]/P0001  & n13492 ;
  assign n20429 = ~n20427 & ~n20428 ;
  assign n20430 = n20426 & n20429 ;
  assign n20431 = n20423 & n20430 ;
  assign n20432 = \wishbone_bd_ram_mem2_reg[195][17]/P0001  & n13700 ;
  assign n20433 = \wishbone_bd_ram_mem2_reg[198][17]/P0001  & n13592 ;
  assign n20434 = ~n20432 & ~n20433 ;
  assign n20435 = \wishbone_bd_ram_mem2_reg[240][17]/P0001  & n13352 ;
  assign n20436 = \wishbone_bd_ram_mem2_reg[210][17]/P0001  & n13443 ;
  assign n20437 = ~n20435 & ~n20436 ;
  assign n20438 = n20434 & n20437 ;
  assign n20439 = \wishbone_bd_ram_mem2_reg[45][17]/P0001  & n13420 ;
  assign n20440 = \wishbone_bd_ram_mem2_reg[233][17]/P0001  & n13332 ;
  assign n20441 = ~n20439 & ~n20440 ;
  assign n20442 = \wishbone_bd_ram_mem2_reg[162][17]/P0001  & n13726 ;
  assign n20443 = \wishbone_bd_ram_mem2_reg[29][17]/P0001  & n13412 ;
  assign n20444 = ~n20442 & ~n20443 ;
  assign n20445 = n20441 & n20444 ;
  assign n20446 = n20438 & n20445 ;
  assign n20447 = n20431 & n20446 ;
  assign n20448 = n20416 & n20447 ;
  assign n20449 = n20385 & n20448 ;
  assign n20450 = \wishbone_bd_ram_mem2_reg[130][17]/P0001  & n13427 ;
  assign n20451 = \wishbone_bd_ram_mem2_reg[192][17]/P0001  & n13390 ;
  assign n20452 = ~n20450 & ~n20451 ;
  assign n20453 = \wishbone_bd_ram_mem2_reg[218][17]/P0001  & n13792 ;
  assign n20454 = \wishbone_bd_ram_mem2_reg[181][17]/P0001  & n13587 ;
  assign n20455 = ~n20453 & ~n20454 ;
  assign n20456 = n20452 & n20455 ;
  assign n20457 = \wishbone_bd_ram_mem2_reg[147][17]/P0001  & n13702 ;
  assign n20458 = \wishbone_bd_ram_mem2_reg[14][17]/P0001  & n13972 ;
  assign n20459 = ~n20457 & ~n20458 ;
  assign n20460 = \wishbone_bd_ram_mem2_reg[48][17]/P0001  & n13917 ;
  assign n20461 = \wishbone_bd_ram_mem2_reg[175][17]/P0001  & n13674 ;
  assign n20462 = ~n20460 & ~n20461 ;
  assign n20463 = n20459 & n20462 ;
  assign n20464 = n20456 & n20463 ;
  assign n20465 = \wishbone_bd_ram_mem2_reg[250][17]/P0001  & n13677 ;
  assign n20466 = \wishbone_bd_ram_mem2_reg[174][17]/P0001  & n13899 ;
  assign n20467 = ~n20465 & ~n20466 ;
  assign n20468 = \wishbone_bd_ram_mem2_reg[223][17]/P0001  & n13335 ;
  assign n20469 = \wishbone_bd_ram_mem2_reg[77][17]/P0001  & n13935 ;
  assign n20470 = ~n20468 & ~n20469 ;
  assign n20471 = n20467 & n20470 ;
  assign n20472 = \wishbone_bd_ram_mem2_reg[226][17]/P0001  & n13668 ;
  assign n20473 = \wishbone_bd_ram_mem2_reg[249][17]/P0001  & n13431 ;
  assign n20474 = ~n20472 & ~n20473 ;
  assign n20475 = \wishbone_bd_ram_mem2_reg[25][17]/P0001  & n13742 ;
  assign n20476 = \wishbone_bd_ram_mem2_reg[227][17]/P0001  & n13388 ;
  assign n20477 = ~n20475 & ~n20476 ;
  assign n20478 = n20474 & n20477 ;
  assign n20479 = n20471 & n20478 ;
  assign n20480 = n20464 & n20479 ;
  assign n20481 = \wishbone_bd_ram_mem2_reg[145][17]/P0001  & n13715 ;
  assign n20482 = \wishbone_bd_ram_mem2_reg[61][17]/P0001  & n13544 ;
  assign n20483 = ~n20481 & ~n20482 ;
  assign n20484 = \wishbone_bd_ram_mem2_reg[55][17]/P0001  & n13618 ;
  assign n20485 = \wishbone_bd_ram_mem2_reg[242][17]/P0001  & n13383 ;
  assign n20486 = ~n20484 & ~n20485 ;
  assign n20487 = n20483 & n20486 ;
  assign n20488 = \wishbone_bd_ram_mem2_reg[26][17]/P0001  & n13521 ;
  assign n20489 = \wishbone_bd_ram_mem2_reg[125][17]/P0001  & n13396 ;
  assign n20490 = ~n20488 & ~n20489 ;
  assign n20491 = \wishbone_bd_ram_mem2_reg[89][17]/P0001  & n13910 ;
  assign n20492 = \wishbone_bd_ram_mem2_reg[136][17]/P0001  & n13963 ;
  assign n20493 = ~n20491 & ~n20492 ;
  assign n20494 = n20490 & n20493 ;
  assign n20495 = n20487 & n20494 ;
  assign n20496 = \wishbone_bd_ram_mem2_reg[167][17]/P0001  & n13940 ;
  assign n20497 = \wishbone_bd_ram_mem2_reg[42][17]/P0001  & n13341 ;
  assign n20498 = ~n20496 & ~n20497 ;
  assign n20499 = \wishbone_bd_ram_mem2_reg[27][17]/P0001  & n13251 ;
  assign n20500 = \wishbone_bd_ram_mem2_reg[87][17]/P0001  & n13691 ;
  assign n20501 = ~n20499 & ~n20500 ;
  assign n20502 = n20498 & n20501 ;
  assign n20503 = \wishbone_bd_ram_mem2_reg[30][17]/P0001  & n13713 ;
  assign n20504 = \wishbone_bd_ram_mem2_reg[70][17]/P0001  & n13339 ;
  assign n20505 = ~n20503 & ~n20504 ;
  assign n20506 = \wishbone_bd_ram_mem2_reg[46][17]/P0001  & n13298 ;
  assign n20507 = \wishbone_bd_ram_mem2_reg[131][17]/P0001  & n13358 ;
  assign n20508 = ~n20506 & ~n20507 ;
  assign n20509 = n20505 & n20508 ;
  assign n20510 = n20502 & n20509 ;
  assign n20511 = n20495 & n20510 ;
  assign n20512 = n20480 & n20511 ;
  assign n20513 = \wishbone_bd_ram_mem2_reg[158][17]/P0001  & n13294 ;
  assign n20514 = \wishbone_bd_ram_mem2_reg[43][17]/P0001  & n13761 ;
  assign n20515 = ~n20513 & ~n20514 ;
  assign n20516 = \wishbone_bd_ram_mem2_reg[11][17]/P0001  & n13774 ;
  assign n20517 = \wishbone_bd_ram_mem2_reg[178][17]/P0001  & n13301 ;
  assign n20518 = ~n20516 & ~n20517 ;
  assign n20519 = n20515 & n20518 ;
  assign n20520 = \wishbone_bd_ram_mem2_reg[111][17]/P0001  & n13471 ;
  assign n20521 = \wishbone_bd_ram_mem2_reg[152][17]/P0001  & n13912 ;
  assign n20522 = ~n20520 & ~n20521 ;
  assign n20523 = \wishbone_bd_ram_mem2_reg[177][17]/P0001  & n13863 ;
  assign n20524 = \wishbone_bd_ram_mem2_reg[52][17]/P0001  & n13988 ;
  assign n20525 = ~n20523 & ~n20524 ;
  assign n20526 = n20522 & n20525 ;
  assign n20527 = n20519 & n20526 ;
  assign n20528 = \wishbone_bd_ram_mem2_reg[139][17]/P0001  & n13566 ;
  assign n20529 = \wishbone_bd_ram_mem2_reg[116][17]/P0001  & n13865 ;
  assign n20530 = ~n20528 & ~n20529 ;
  assign n20531 = \wishbone_bd_ram_mem2_reg[36][17]/P0001  & n13639 ;
  assign n20532 = \wishbone_bd_ram_mem2_reg[201][17]/P0001  & n13600 ;
  assign n20533 = ~n20531 & ~n20532 ;
  assign n20534 = n20530 & n20533 ;
  assign n20535 = \wishbone_bd_ram_mem2_reg[67][17]/P0001  & n13663 ;
  assign n20536 = \wishbone_bd_ram_mem2_reg[0][17]/P0001  & n13539 ;
  assign n20537 = ~n20535 & ~n20536 ;
  assign n20538 = \wishbone_bd_ram_mem2_reg[72][17]/P0001  & n13582 ;
  assign n20539 = \wishbone_bd_ram_mem2_reg[2][17]/P0001  & n13975 ;
  assign n20540 = ~n20538 & ~n20539 ;
  assign n20541 = n20537 & n20540 ;
  assign n20542 = n20534 & n20541 ;
  assign n20543 = n20527 & n20542 ;
  assign n20544 = \wishbone_bd_ram_mem2_reg[98][17]/P0001  & n13569 ;
  assign n20545 = \wishbone_bd_ram_mem2_reg[236][17]/P0001  & n13480 ;
  assign n20546 = ~n20544 & ~n20545 ;
  assign n20547 = \wishbone_bd_ram_mem2_reg[37][17]/P0001  & n13710 ;
  assign n20548 = \wishbone_bd_ram_mem2_reg[66][17]/P0001  & n13603 ;
  assign n20549 = ~n20547 & ~n20548 ;
  assign n20550 = n20546 & n20549 ;
  assign n20551 = \wishbone_bd_ram_mem2_reg[185][17]/P0001  & n13372 ;
  assign n20552 = \wishbone_bd_ram_mem2_reg[21][17]/P0001  & n13438 ;
  assign n20553 = ~n20551 & ~n20552 ;
  assign n20554 = \wishbone_bd_ram_mem2_reg[73][17]/P0001  & n13456 ;
  assign n20555 = \wishbone_bd_ram_mem2_reg[219][17]/P0001  & n13577 ;
  assign n20556 = ~n20554 & ~n20555 ;
  assign n20557 = n20553 & n20556 ;
  assign n20558 = n20550 & n20557 ;
  assign n20559 = \wishbone_bd_ram_mem2_reg[129][17]/P0001  & n13629 ;
  assign n20560 = \wishbone_bd_ram_mem2_reg[62][17]/P0001  & n13529 ;
  assign n20561 = ~n20559 & ~n20560 ;
  assign n20562 = \wishbone_bd_ram_mem2_reg[82][17]/P0001  & n13374 ;
  assign n20563 = \wishbone_bd_ram_mem2_reg[156][17]/P0001  & n13769 ;
  assign n20564 = ~n20562 & ~n20563 ;
  assign n20565 = n20561 & n20564 ;
  assign n20566 = \wishbone_bd_ram_mem2_reg[16][17]/P0001  & n13695 ;
  assign n20567 = \wishbone_bd_ram_mem2_reg[126][17]/P0001  & n13786 ;
  assign n20568 = ~n20566 & ~n20567 ;
  assign n20569 = \wishbone_bd_ram_mem2_reg[228][17]/P0001  & n13497 ;
  assign n20570 = \wishbone_bd_ram_mem2_reg[80][17]/P0001  & n13516 ;
  assign n20571 = ~n20569 & ~n20570 ;
  assign n20572 = n20568 & n20571 ;
  assign n20573 = n20565 & n20572 ;
  assign n20574 = n20558 & n20573 ;
  assign n20575 = n20543 & n20574 ;
  assign n20576 = n20512 & n20575 ;
  assign n20577 = n20449 & n20576 ;
  assign n20578 = \wishbone_bd_ram_mem2_reg[224][17]/P0001  & n13433 ;
  assign n20579 = \wishbone_bd_ram_mem2_reg[179][17]/P0001  & n14035 ;
  assign n20580 = ~n20578 & ~n20579 ;
  assign n20581 = \wishbone_bd_ram_mem2_reg[54][17]/P0001  & n13622 ;
  assign n20582 = \wishbone_bd_ram_mem2_reg[5][17]/P0001  & n13243 ;
  assign n20583 = ~n20581 & ~n20582 ;
  assign n20584 = n20580 & n20583 ;
  assign n20585 = \wishbone_bd_ram_mem2_reg[104][17]/P0001  & n13684 ;
  assign n20586 = \wishbone_bd_ram_mem2_reg[154][17]/P0001  & n13403 ;
  assign n20587 = ~n20585 & ~n20586 ;
  assign n20588 = \wishbone_bd_ram_mem2_reg[115][17]/P0001  & n13747 ;
  assign n20589 = \wishbone_bd_ram_mem2_reg[108][17]/P0001  & n13814 ;
  assign n20590 = ~n20588 & ~n20589 ;
  assign n20591 = n20587 & n20590 ;
  assign n20592 = n20584 & n20591 ;
  assign n20593 = \wishbone_bd_ram_mem2_reg[196][17]/P0001  & n13977 ;
  assign n20594 = \wishbone_bd_ram_mem2_reg[114][17]/P0001  & n13763 ;
  assign n20595 = ~n20593 & ~n20594 ;
  assign n20596 = \wishbone_bd_ram_mem2_reg[38][17]/P0001  & n13828 ;
  assign n20597 = \wishbone_bd_ram_mem2_reg[215][17]/P0001  & n13901 ;
  assign n20598 = ~n20596 & ~n20597 ;
  assign n20599 = n20595 & n20598 ;
  assign n20600 = \wishbone_bd_ram_mem2_reg[202][17]/P0001  & n13268 ;
  assign n20601 = \wishbone_bd_ram_mem2_reg[110][17]/P0001  & n14030 ;
  assign n20602 = ~n20600 & ~n20601 ;
  assign n20603 = \wishbone_bd_ram_mem2_reg[135][17]/P0001  & n13672 ;
  assign n20604 = \wishbone_bd_ram_mem2_reg[109][17]/P0001  & n13306 ;
  assign n20605 = ~n20603 & ~n20604 ;
  assign n20606 = n20602 & n20605 ;
  assign n20607 = n20599 & n20606 ;
  assign n20608 = n20592 & n20607 ;
  assign n20609 = \wishbone_bd_ram_mem2_reg[189][17]/P0001  & n14001 ;
  assign n20610 = \wishbone_bd_ram_mem2_reg[75][17]/P0001  & n13605 ;
  assign n20611 = ~n20609 & ~n20610 ;
  assign n20612 = \wishbone_bd_ram_mem2_reg[197][17]/P0001  & n13594 ;
  assign n20613 = \wishbone_bd_ram_mem2_reg[254][17]/P0001  & n13283 ;
  assign n20614 = ~n20612 & ~n20613 ;
  assign n20615 = n20611 & n20614 ;
  assign n20616 = \wishbone_bd_ram_mem2_reg[59][17]/P0001  & n13613 ;
  assign n20617 = \wishbone_bd_ram_mem2_reg[204][17]/P0001  & n13821 ;
  assign n20618 = ~n20616 & ~n20617 ;
  assign n20619 = \wishbone_bd_ram_mem2_reg[88][17]/P0001  & n13347 ;
  assign n20620 = \wishbone_bd_ram_mem2_reg[182][17]/P0001  & n13598 ;
  assign n20621 = ~n20619 & ~n20620 ;
  assign n20622 = n20618 & n20621 ;
  assign n20623 = n20615 & n20622 ;
  assign n20624 = \wishbone_bd_ram_mem2_reg[17][17]/P0001  & n13324 ;
  assign n20625 = \wishbone_bd_ram_mem2_reg[103][17]/P0001  & n13320 ;
  assign n20626 = ~n20624 & ~n20625 ;
  assign n20627 = \wishbone_bd_ram_mem2_reg[120][17]/P0001  & n13550 ;
  assign n20628 = \wishbone_bd_ram_mem2_reg[190][17]/P0001  & n13365 ;
  assign n20629 = ~n20627 & ~n20628 ;
  assign n20630 = n20626 & n20629 ;
  assign n20631 = \wishbone_bd_ram_mem2_reg[199][17]/P0001  & n13499 ;
  assign n20632 = \wishbone_bd_ram_mem2_reg[141][17]/P0001  & n13852 ;
  assign n20633 = ~n20631 & ~n20632 ;
  assign n20634 = \wishbone_bd_ram_mem2_reg[159][17]/P0001  & n13627 ;
  assign n20635 = \wishbone_bd_ram_mem2_reg[169][17]/P0001  & n13541 ;
  assign n20636 = ~n20634 & ~n20635 ;
  assign n20637 = n20633 & n20636 ;
  assign n20638 = n20630 & n20637 ;
  assign n20639 = n20623 & n20638 ;
  assign n20640 = n20608 & n20639 ;
  assign n20641 = \wishbone_bd_ram_mem2_reg[18][17]/P0001  & n13532 ;
  assign n20642 = \wishbone_bd_ram_mem2_reg[68][17]/P0001  & n13379 ;
  assign n20643 = ~n20641 & ~n20642 ;
  assign n20644 = \wishbone_bd_ram_mem2_reg[95][17]/P0001  & n13317 ;
  assign n20645 = \wishbone_bd_ram_mem2_reg[170][17]/P0001  & n14007 ;
  assign n20646 = ~n20644 & ~n20645 ;
  assign n20647 = n20643 & n20646 ;
  assign n20648 = \wishbone_bd_ram_mem2_reg[235][17]/P0001  & n13518 ;
  assign n20649 = \wishbone_bd_ram_mem2_reg[94][17]/P0001  & n13833 ;
  assign n20650 = ~n20648 & ~n20649 ;
  assign n20651 = \wishbone_bd_ram_mem2_reg[106][17]/P0001  & n13555 ;
  assign n20652 = \wishbone_bd_ram_mem2_reg[79][17]/P0001  & n13779 ;
  assign n20653 = ~n20651 & ~n20652 ;
  assign n20654 = n20650 & n20653 ;
  assign n20655 = n20647 & n20654 ;
  assign n20656 = \wishbone_bd_ram_mem2_reg[188][17]/P0001  & n13407 ;
  assign n20657 = \wishbone_bd_ram_mem2_reg[81][17]/P0001  & n13409 ;
  assign n20658 = ~n20656 & ~n20657 ;
  assign n20659 = \wishbone_bd_ram_mem2_reg[171][17]/P0001  & n13422 ;
  assign n20660 = \wishbone_bd_ram_mem2_reg[238][17]/P0001  & n13819 ;
  assign n20661 = ~n20659 & ~n20660 ;
  assign n20662 = n20658 & n20661 ;
  assign n20663 = \wishbone_bd_ram_mem2_reg[246][17]/P0001  & n13981 ;
  assign n20664 = \wishbone_bd_ram_mem2_reg[150][17]/P0001  & n13666 ;
  assign n20665 = ~n20663 & ~n20664 ;
  assign n20666 = \wishbone_bd_ram_mem2_reg[140][17]/P0001  & n13287 ;
  assign n20667 = \wishbone_bd_ram_mem2_reg[255][17]/P0001  & n13952 ;
  assign n20668 = ~n20666 & ~n20667 ;
  assign n20669 = n20665 & n20668 ;
  assign n20670 = n20662 & n20669 ;
  assign n20671 = n20655 & n20670 ;
  assign n20672 = \wishbone_bd_ram_mem2_reg[252][17]/P0001  & n13986 ;
  assign n20673 = \wishbone_bd_ram_mem2_reg[191][17]/P0001  & n14012 ;
  assign n20674 = ~n20672 & ~n20673 ;
  assign n20675 = \wishbone_bd_ram_mem2_reg[7][17]/P0001  & n13546 ;
  assign n20676 = \wishbone_bd_ram_mem2_reg[100][17]/P0001  & n13401 ;
  assign n20677 = ~n20675 & ~n20676 ;
  assign n20678 = n20674 & n20677 ;
  assign n20679 = \wishbone_bd_ram_mem2_reg[216][17]/P0001  & n14005 ;
  assign n20680 = \wishbone_bd_ram_mem2_reg[225][17]/P0001  & n13719 ;
  assign n20681 = ~n20679 & ~n20680 ;
  assign n20682 = \wishbone_bd_ram_mem2_reg[203][17]/P0001  & n13816 ;
  assign n20683 = \wishbone_bd_ram_mem2_reg[4][17]/P0001  & n13527 ;
  assign n20684 = ~n20682 & ~n20683 ;
  assign n20685 = n20681 & n20684 ;
  assign n20686 = n20678 & n20685 ;
  assign n20687 = \wishbone_bd_ram_mem2_reg[74][17]/P0001  & n13564 ;
  assign n20688 = \wishbone_bd_ram_mem2_reg[164][17]/P0001  & n13236 ;
  assign n20689 = ~n20687 & ~n20688 ;
  assign n20690 = \wishbone_bd_ram_mem2_reg[83][17]/P0001  & n13454 ;
  assign n20691 = \wishbone_bd_ram_mem2_reg[121][17]/P0001  & n13983 ;
  assign n20692 = ~n20690 & ~n20691 ;
  assign n20693 = n20689 & n20692 ;
  assign n20694 = \wishbone_bd_ram_mem2_reg[6][17]/P0001  & n13915 ;
  assign n20695 = \wishbone_bd_ram_mem2_reg[157][17]/P0001  & n13445 ;
  assign n20696 = ~n20694 & ~n20695 ;
  assign n20697 = \wishbone_bd_ram_mem2_reg[241][17]/P0001  & n13854 ;
  assign n20698 = \wishbone_bd_ram_mem2_reg[186][17]/P0001  & n13616 ;
  assign n20699 = ~n20697 & ~n20698 ;
  assign n20700 = n20696 & n20699 ;
  assign n20701 = n20693 & n20700 ;
  assign n20702 = n20686 & n20701 ;
  assign n20703 = n20671 & n20702 ;
  assign n20704 = n20640 & n20703 ;
  assign n20705 = \wishbone_bd_ram_mem2_reg[200][17]/P0001  & n13922 ;
  assign n20706 = \wishbone_bd_ram_mem2_reg[248][17]/P0001  & n13647 ;
  assign n20707 = ~n20705 & ~n20706 ;
  assign n20708 = \wishbone_bd_ram_mem2_reg[31][17]/P0001  & n13758 ;
  assign n20709 = \wishbone_bd_ram_mem2_reg[232][17]/P0001  & n13510 ;
  assign n20710 = ~n20708 & ~n20709 ;
  assign n20711 = n20707 & n20710 ;
  assign n20712 = \wishbone_bd_ram_mem2_reg[165][17]/P0001  & n14028 ;
  assign n20713 = \wishbone_bd_ram_mem2_reg[1][17]/P0001  & n13888 ;
  assign n20714 = ~n20712 & ~n20713 ;
  assign n20715 = \wishbone_bd_ram_mem2_reg[244][17]/P0001  & n13474 ;
  assign n20716 = \wishbone_bd_ram_mem2_reg[247][17]/P0001  & n13571 ;
  assign n20717 = ~n20715 & ~n20716 ;
  assign n20718 = n20714 & n20717 ;
  assign n20719 = n20711 & n20718 ;
  assign n20720 = \wishbone_bd_ram_mem2_reg[239][17]/P0001  & n13349 ;
  assign n20721 = \wishbone_bd_ram_mem2_reg[123][17]/P0001  & n13749 ;
  assign n20722 = ~n20720 & ~n20721 ;
  assign n20723 = \wishbone_bd_ram_mem2_reg[99][17]/P0001  & n13996 ;
  assign n20724 = \wishbone_bd_ram_mem2_reg[86][17]/P0001  & n13485 ;
  assign n20725 = ~n20723 & ~n20724 ;
  assign n20726 = n20722 & n20725 ;
  assign n20727 = \wishbone_bd_ram_mem2_reg[163][17]/P0001  & n13255 ;
  assign n20728 = \wishbone_bd_ram_mem2_reg[208][17]/P0001  & n14010 ;
  assign n20729 = ~n20727 & ~n20728 ;
  assign n20730 = \wishbone_bd_ram_mem2_reg[101][17]/P0001  & n13772 ;
  assign n20731 = \wishbone_bd_ram_mem2_reg[211][17]/P0001  & n13805 ;
  assign n20732 = ~n20730 & ~n20731 ;
  assign n20733 = n20729 & n20732 ;
  assign n20734 = n20726 & n20733 ;
  assign n20735 = n20719 & n20734 ;
  assign n20736 = \wishbone_bd_ram_mem2_reg[172][17]/P0001  & n13377 ;
  assign n20737 = \wishbone_bd_ram_mem2_reg[153][17]/P0001  & n13309 ;
  assign n20738 = ~n20736 & ~n20737 ;
  assign n20739 = \wishbone_bd_ram_mem2_reg[220][17]/P0001  & n13965 ;
  assign n20740 = \wishbone_bd_ram_mem2_reg[112][17]/P0001  & n13482 ;
  assign n20741 = ~n20739 & ~n20740 ;
  assign n20742 = n20738 & n20741 ;
  assign n20743 = \wishbone_bd_ram_mem2_reg[205][17]/P0001  & n13947 ;
  assign n20744 = \wishbone_bd_ram_mem2_reg[155][17]/P0001  & n13738 ;
  assign n20745 = ~n20743 & ~n20744 ;
  assign n20746 = \wishbone_bd_ram_mem2_reg[230][17]/P0001  & n13994 ;
  assign n20747 = \wishbone_bd_ram_mem2_reg[20][17]/P0001  & n13839 ;
  assign n20748 = ~n20746 & ~n20747 ;
  assign n20749 = n20745 & n20748 ;
  assign n20750 = n20742 & n20749 ;
  assign n20751 = \wishbone_bd_ram_mem2_reg[58][17]/P0001  & n13949 ;
  assign n20752 = \wishbone_bd_ram_mem2_reg[138][17]/P0001  & n13398 ;
  assign n20753 = ~n20751 & ~n20752 ;
  assign n20754 = \wishbone_bd_ram_mem2_reg[35][17]/P0001  & n13523 ;
  assign n20755 = \wishbone_bd_ram_mem2_reg[222][17]/P0001  & n13721 ;
  assign n20756 = ~n20754 & ~n20755 ;
  assign n20757 = n20753 & n20756 ;
  assign n20758 = \wishbone_bd_ram_mem2_reg[3][17]/P0001  & n13354 ;
  assign n20759 = \wishbone_bd_ram_mem2_reg[245][17]/P0001  & n13877 ;
  assign n20760 = ~n20758 & ~n20759 ;
  assign n20761 = \wishbone_bd_ram_mem2_reg[118][17]/P0001  & n13589 ;
  assign n20762 = \wishbone_bd_ram_mem2_reg[28][17]/P0001  & n13810 ;
  assign n20763 = ~n20761 & ~n20762 ;
  assign n20764 = n20760 & n20763 ;
  assign n20765 = n20757 & n20764 ;
  assign n20766 = n20750 & n20765 ;
  assign n20767 = n20735 & n20766 ;
  assign n20768 = \wishbone_bd_ram_mem2_reg[187][17]/P0001  & n13756 ;
  assign n20769 = \wishbone_bd_ram_mem2_reg[137][17]/P0001  & n13808 ;
  assign n20770 = ~n20768 & ~n20769 ;
  assign n20771 = \wishbone_bd_ram_mem2_reg[8][17]/P0001  & n13459 ;
  assign n20772 = \wishbone_bd_ram_mem2_reg[53][17]/P0001  & n13875 ;
  assign n20773 = ~n20771 & ~n20772 ;
  assign n20774 = n20770 & n20773 ;
  assign n20775 = \wishbone_bd_ram_mem2_reg[91][17]/P0001  & n13954 ;
  assign n20776 = \wishbone_bd_ram_mem2_reg[221][17]/P0001  & n13641 ;
  assign n20777 = ~n20775 & ~n20776 ;
  assign n20778 = \wishbone_bd_ram_mem2_reg[206][17]/P0001  & n13414 ;
  assign n20779 = \wishbone_bd_ram_mem2_reg[194][17]/P0001  & n13624 ;
  assign n20780 = ~n20778 & ~n20779 ;
  assign n20781 = n20777 & n20780 ;
  assign n20782 = n20774 & n20781 ;
  assign n20783 = \wishbone_bd_ram_mem2_reg[39][17]/P0001  & n13893 ;
  assign n20784 = \wishbone_bd_ram_mem2_reg[144][17]/P0001  & n13508 ;
  assign n20785 = ~n20783 & ~n20784 ;
  assign n20786 = \wishbone_bd_ram_mem2_reg[47][17]/P0001  & n13436 ;
  assign n20787 = \wishbone_bd_ram_mem2_reg[251][17]/P0001  & n14019 ;
  assign n20788 = ~n20786 & ~n20787 ;
  assign n20789 = n20785 & n20788 ;
  assign n20790 = \wishbone_bd_ram_mem2_reg[113][17]/P0001  & n13882 ;
  assign n20791 = \wishbone_bd_ram_mem2_reg[65][17]/P0001  & n13842 ;
  assign n20792 = ~n20790 & ~n20791 ;
  assign n20793 = \wishbone_bd_ram_mem2_reg[180][17]/P0001  & n13650 ;
  assign n20794 = \wishbone_bd_ram_mem2_reg[193][17]/P0001  & n14022 ;
  assign n20795 = ~n20793 & ~n20794 ;
  assign n20796 = n20792 & n20795 ;
  assign n20797 = n20789 & n20796 ;
  assign n20798 = n20782 & n20797 ;
  assign n20799 = \wishbone_bd_ram_mem2_reg[41][17]/P0001  & n14017 ;
  assign n20800 = \wishbone_bd_ram_mem2_reg[160][17]/P0001  & n13271 ;
  assign n20801 = ~n20799 & ~n20800 ;
  assign n20802 = \wishbone_bd_ram_mem2_reg[217][17]/P0001  & n13767 ;
  assign n20803 = \wishbone_bd_ram_mem2_reg[142][17]/P0001  & n13448 ;
  assign n20804 = ~n20802 & ~n20803 ;
  assign n20805 = n20801 & n20804 ;
  assign n20806 = \wishbone_bd_ram_mem2_reg[78][17]/P0001  & n13277 ;
  assign n20807 = \wishbone_bd_ram_mem2_reg[207][17]/P0001  & n13826 ;
  assign n20808 = ~n20806 & ~n20807 ;
  assign n20809 = \wishbone_bd_ram_mem2_reg[128][17]/P0001  & n13652 ;
  assign n20810 = \wishbone_bd_ram_mem2_reg[24][17]/P0001  & n13970 ;
  assign n20811 = ~n20809 & ~n20810 ;
  assign n20812 = n20808 & n20811 ;
  assign n20813 = n20805 & n20812 ;
  assign n20814 = \wishbone_bd_ram_mem2_reg[127][17]/P0001  & n13803 ;
  assign n20815 = \wishbone_bd_ram_mem2_reg[40][17]/P0001  & n13661 ;
  assign n20816 = ~n20814 & ~n20815 ;
  assign n20817 = \wishbone_bd_ram_mem2_reg[151][17]/P0001  & n13697 ;
  assign n20818 = \wishbone_bd_ram_mem2_reg[71][17]/P0001  & n13636 ;
  assign n20819 = ~n20817 & ~n20818 ;
  assign n20820 = n20816 & n20819 ;
  assign n20821 = \wishbone_bd_ram_mem2_reg[32][17]/P0001  & n13736 ;
  assign n20822 = \wishbone_bd_ram_mem2_reg[50][17]/P0001  & n13686 ;
  assign n20823 = ~n20821 & ~n20822 ;
  assign n20824 = \wishbone_bd_ram_mem2_reg[148][17]/P0001  & n13868 ;
  assign n20825 = \wishbone_bd_ram_mem2_reg[237][17]/P0001  & n13924 ;
  assign n20826 = ~n20824 & ~n20825 ;
  assign n20827 = n20823 & n20826 ;
  assign n20828 = n20820 & n20827 ;
  assign n20829 = n20813 & n20828 ;
  assign n20830 = n20798 & n20829 ;
  assign n20831 = n20767 & n20830 ;
  assign n20832 = n20704 & n20831 ;
  assign n20833 = n20577 & n20832 ;
  assign n20834 = n14047 & ~n20833 ;
  assign n20835 = \wishbone_TxLength_reg[1]/NET0131  & \wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n20836 = ~n14068 & n20835 ;
  assign n20837 = ~\wishbone_TxLength_reg[1]/NET0131  & \wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n20838 = n14068 & n20837 ;
  assign n20839 = ~n20836 & ~n20838 ;
  assign n20840 = ~\wishbone_TxLength_reg[1]/NET0131  & ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n20841 = ~n14068 & n20840 ;
  assign n20842 = \wishbone_TxLength_reg[1]/NET0131  & ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n20843 = n14068 & n20842 ;
  assign n20844 = ~n20841 & ~n20843 ;
  assign n20845 = n20839 & n20844 ;
  assign n20846 = n14065 & n20845 ;
  assign n20847 = ~n14064 & n20846 ;
  assign n20848 = \wishbone_TxLength_reg[1]/NET0131  & ~n14049 ;
  assign n20849 = ~n14046 & n20848 ;
  assign n20850 = ~n20847 & ~n20849 ;
  assign n20851 = ~n20834 & n20850 ;
  assign n20852 = \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  & n15157 ;
  assign n20853 = ~\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  & ~n20852 ;
  assign n20854 = n15142 & n15157 ;
  assign n20855 = n15162 & ~n20854 ;
  assign n20856 = ~n20853 & n20855 ;
  assign n20857 = ~\txethmac1_txcrc_Crc_reg[5]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n20858 = n11626 & n20857 ;
  assign n20859 = ~\txethmac1_txcrc_Crc_reg[5]/NET0131  & n11464 ;
  assign n20860 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n11464 ;
  assign n20861 = n11626 & n20860 ;
  assign n20862 = ~n20859 & ~n20861 ;
  assign n20863 = ~n20858 & ~n20862 ;
  assign n20864 = ~\wishbone_RxPointerMSB_reg[12]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n20865 = n13144 & n20864 ;
  assign n20866 = ~n13149 & ~n20865 ;
  assign n20867 = n13143 & n20866 ;
  assign n20868 = n13137 & n20867 ;
  assign n20869 = ~n13170 & ~n20868 ;
  assign n20870 = ~\m_wb_adr_o[12]_pad  & ~n13103 ;
  assign n20871 = ~n18636 & ~n20870 ;
  assign n20872 = ~n20869 & n20871 ;
  assign n20873 = \m_wb_adr_o[12]_pad  & n13197 ;
  assign n20874 = \wishbone_RxPointerMSB_reg[12]/NET0131  & n13207 ;
  assign n20875 = ~n13196 & n20874 ;
  assign n20876 = \wishbone_TxPointerMSB_reg[12]/NET0131  & ~n13201 ;
  assign n20877 = ~n20875 & ~n20876 ;
  assign n20878 = ~n20873 & n20877 ;
  assign n20879 = ~n20872 & n20878 ;
  assign n20880 = ~\wishbone_TxPointerMSB_reg[16]/NET0131  & ~\wishbone_tx_burst_cnt_reg[2]/NET0131  ;
  assign n20881 = n13167 & n20880 ;
  assign n20882 = ~n13166 & ~n20881 ;
  assign n20883 = ~n13164 & n20882 ;
  assign n20884 = ~n15176 & ~n20883 ;
  assign n20885 = \m_wb_adr_o[16]_pad  & n13107 ;
  assign n20886 = ~\m_wb_adr_o[16]_pad  & ~n13107 ;
  assign n20887 = ~n20885 & ~n20886 ;
  assign n20888 = ~n20884 & n20887 ;
  assign n20889 = \m_wb_adr_o[16]_pad  & n13197 ;
  assign n20890 = \wishbone_TxPointerMSB_reg[16]/NET0131  & ~n13201 ;
  assign n20891 = \wishbone_RxPointerMSB_reg[16]/NET0131  & n13207 ;
  assign n20892 = ~n13196 & n20891 ;
  assign n20893 = ~n20890 & ~n20892 ;
  assign n20894 = ~n20889 & n20893 ;
  assign n20895 = ~n20888 & n20894 ;
  assign n20896 = ~\m_wb_adr_o[17]_pad  & ~n20885 ;
  assign n20897 = ~\wishbone_TxPointerMSB_reg[17]/NET0131  & ~\wishbone_tx_burst_cnt_reg[2]/NET0131  ;
  assign n20898 = n13167 & n20897 ;
  assign n20899 = ~n13166 & ~n20898 ;
  assign n20900 = ~n13164 & n20899 ;
  assign n20901 = ~n15176 & ~n20900 ;
  assign n20902 = ~n16835 & ~n20901 ;
  assign n20903 = ~n20896 & n20902 ;
  assign n20904 = \m_wb_adr_o[17]_pad  & n13197 ;
  assign n20905 = \wishbone_TxPointerMSB_reg[17]/NET0131  & ~n13201 ;
  assign n20906 = \wishbone_RxPointerMSB_reg[17]/NET0131  & n13207 ;
  assign n20907 = ~n13196 & n20906 ;
  assign n20908 = ~n20905 & ~n20907 ;
  assign n20909 = ~n20904 & n20908 ;
  assign n20910 = ~n20903 & n20909 ;
  assign n20911 = ~\m_wb_adr_o[19]_pad  & ~n16838 ;
  assign n20912 = ~\wishbone_TxPointerMSB_reg[19]/NET0131  & ~\wishbone_tx_burst_cnt_reg[2]/NET0131  ;
  assign n20913 = n13167 & n20912 ;
  assign n20914 = ~n13166 & ~n20913 ;
  assign n20915 = ~n13164 & n20914 ;
  assign n20916 = ~n15176 & ~n20915 ;
  assign n20917 = ~n13111 & ~n20916 ;
  assign n20918 = ~n20911 & n20917 ;
  assign n20919 = \m_wb_adr_o[19]_pad  & n13197 ;
  assign n20920 = \wishbone_TxPointerMSB_reg[19]/NET0131  & ~n13201 ;
  assign n20921 = \wishbone_RxPointerMSB_reg[19]/NET0131  & n13207 ;
  assign n20922 = ~n13196 & n20921 ;
  assign n20923 = ~n20920 & ~n20922 ;
  assign n20924 = ~n20919 & n20923 ;
  assign n20925 = ~n20918 & n20924 ;
  assign n20926 = ~\m_wb_adr_o[20]_pad  & ~n13111 ;
  assign n20927 = \m_wb_adr_o[20]_pad  & n13111 ;
  assign n20928 = ~\wishbone_RxPointerMSB_reg[20]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n20929 = n13144 & n20928 ;
  assign n20930 = ~n13149 & ~n20929 ;
  assign n20931 = n13143 & n20930 ;
  assign n20932 = n13137 & n20931 ;
  assign n20933 = ~n13170 & ~n20932 ;
  assign n20934 = ~n20927 & ~n20933 ;
  assign n20935 = ~n20926 & n20934 ;
  assign n20936 = \m_wb_adr_o[20]_pad  & n13197 ;
  assign n20937 = \wishbone_TxPointerMSB_reg[20]/NET0131  & ~n13201 ;
  assign n20938 = \wishbone_RxPointerMSB_reg[20]/NET0131  & n13207 ;
  assign n20939 = ~n13196 & n20938 ;
  assign n20940 = ~n20937 & ~n20939 ;
  assign n20941 = ~n20936 & n20940 ;
  assign n20942 = ~n20935 & n20941 ;
  assign n20943 = ~\m_wb_adr_o[21]_pad  & ~n20927 ;
  assign n20944 = n13111 & n13112 ;
  assign n20945 = ~\wishbone_TxPointerMSB_reg[21]/NET0131  & ~\wishbone_tx_burst_cnt_reg[2]/NET0131  ;
  assign n20946 = n13167 & n20945 ;
  assign n20947 = ~n13166 & ~n20946 ;
  assign n20948 = ~n13164 & n20947 ;
  assign n20949 = ~n15176 & ~n20948 ;
  assign n20950 = ~n20944 & ~n20949 ;
  assign n20951 = ~n20943 & n20950 ;
  assign n20952 = \m_wb_adr_o[21]_pad  & n13197 ;
  assign n20953 = \wishbone_TxPointerMSB_reg[21]/NET0131  & ~n13201 ;
  assign n20954 = \wishbone_RxPointerMSB_reg[21]/NET0131  & n13207 ;
  assign n20955 = ~n13196 & n20954 ;
  assign n20956 = ~n20953 & ~n20955 ;
  assign n20957 = ~n20952 & n20956 ;
  assign n20958 = ~n20951 & n20957 ;
  assign n20959 = \m_wb_adr_o[3]_pad  & n13197 ;
  assign n20960 = \wishbone_RxPointerMSB_reg[3]/NET0131  & n13207 ;
  assign n20961 = ~n13196 & n20960 ;
  assign n20962 = ~n20959 & ~n20961 ;
  assign n20963 = \wishbone_TxPointerMSB_reg[3]/NET0131  & ~n13201 ;
  assign n20964 = ~\m_wb_adr_o[2]_pad  & ~\m_wb_adr_o[3]_pad  ;
  assign n20965 = ~n13095 & ~n20964 ;
  assign n20966 = ~n15177 & n20965 ;
  assign n20967 = ~n20963 & ~n20966 ;
  assign n20968 = n20962 & n20967 ;
  assign n20969 = ~\m_wb_adr_o[22]_pad  & ~n20944 ;
  assign n20970 = ~\wishbone_TxPointerMSB_reg[22]/NET0131  & ~\wishbone_tx_burst_cnt_reg[2]/NET0131  ;
  assign n20971 = n13167 & n20970 ;
  assign n20972 = ~n13166 & ~n20971 ;
  assign n20973 = ~n13164 & n20972 ;
  assign n20974 = ~n15176 & ~n20973 ;
  assign n20975 = \m_wb_adr_o[20]_pad  & \m_wb_adr_o[22]_pad  ;
  assign n20976 = \m_wb_adr_o[21]_pad  & n20975 ;
  assign n20977 = n13111 & n20976 ;
  assign n20978 = ~n20974 & ~n20977 ;
  assign n20979 = ~n20969 & n20978 ;
  assign n20980 = \m_wb_adr_o[22]_pad  & n13197 ;
  assign n20981 = \wishbone_TxPointerMSB_reg[22]/NET0131  & ~n13201 ;
  assign n20982 = \wishbone_RxPointerMSB_reg[22]/NET0131  & n13207 ;
  assign n20983 = ~n13196 & n20982 ;
  assign n20984 = ~n20981 & ~n20983 ;
  assign n20985 = ~n20980 & n20984 ;
  assign n20986 = ~n20979 & n20985 ;
  assign n20987 = \m_wb_adr_o[23]_pad  & n20977 ;
  assign n20988 = ~\m_wb_adr_o[23]_pad  & ~n20977 ;
  assign n20989 = ~n15177 & ~n20988 ;
  assign n20990 = ~n20987 & n20989 ;
  assign n20991 = \m_wb_adr_o[23]_pad  & n13197 ;
  assign n20992 = \wishbone_RxPointerMSB_reg[23]/NET0131  & n13207 ;
  assign n20993 = ~n13196 & n20992 ;
  assign n20994 = \wishbone_TxPointerMSB_reg[23]/NET0131  & ~n13201 ;
  assign n20995 = ~n20993 & ~n20994 ;
  assign n20996 = ~n20991 & n20995 ;
  assign n20997 = ~n20990 & n20996 ;
  assign n20998 = ~\m_wb_adr_o[24]_pad  & ~n20987 ;
  assign n20999 = ~\wishbone_RxPointerMSB_reg[24]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n21000 = n13144 & n20999 ;
  assign n21001 = ~n13149 & ~n21000 ;
  assign n21002 = n13143 & n21001 ;
  assign n21003 = n13137 & n21002 ;
  assign n21004 = ~n13170 & ~n21003 ;
  assign n21005 = ~n15711 & ~n21004 ;
  assign n21006 = ~n20998 & n21005 ;
  assign n21007 = \m_wb_adr_o[24]_pad  & n13197 ;
  assign n21008 = \wishbone_TxPointerMSB_reg[24]/NET0131  & ~n13201 ;
  assign n21009 = \wishbone_RxPointerMSB_reg[24]/NET0131  & n13207 ;
  assign n21010 = ~n13196 & n21009 ;
  assign n21011 = ~n21008 & ~n21010 ;
  assign n21012 = ~n21007 & n21011 ;
  assign n21013 = ~n21006 & n21012 ;
  assign n21014 = ~\m_wb_adr_o[25]_pad  & ~n13203 ;
  assign n21015 = ~n15711 & n21014 ;
  assign n21016 = \m_wb_adr_o[25]_pad  & ~n13203 ;
  assign n21017 = n15711 & n21016 ;
  assign n21018 = ~n21015 & ~n21017 ;
  assign n21019 = ~\wishbone_RxPointerMSB_reg[25]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n21020 = n13144 & n21019 ;
  assign n21021 = ~n13149 & ~n21020 ;
  assign n21022 = n13143 & n21021 ;
  assign n21023 = n13137 & n21022 ;
  assign n21024 = n21018 & n21023 ;
  assign n21025 = ~\m_wb_adr_o[25]_pad  & ~n13168 ;
  assign n21026 = ~n15711 & n21025 ;
  assign n21027 = \m_wb_adr_o[25]_pad  & ~n13168 ;
  assign n21028 = n15711 & n21027 ;
  assign n21029 = ~n21026 & ~n21028 ;
  assign n21030 = ~\wishbone_TxPointerMSB_reg[25]/NET0131  & ~\wishbone_tx_burst_cnt_reg[2]/NET0131  ;
  assign n21031 = n13167 & n21030 ;
  assign n21032 = ~n13166 & ~n21031 ;
  assign n21033 = ~n13164 & n21032 ;
  assign n21034 = n21029 & n21033 ;
  assign n21035 = \m_wb_adr_o[25]_pad  & n13197 ;
  assign n21036 = \wishbone_RxPointerMSB_reg[25]/NET0131  & n13192 ;
  assign n21037 = ~n13194 & n21036 ;
  assign n21038 = \wishbone_TxPointerMSB_reg[25]/NET0131  & ~n13188 ;
  assign n21039 = ~n21037 & ~n21038 ;
  assign n21040 = ~n21035 & n21039 ;
  assign n21041 = ~n21034 & n21040 ;
  assign n21042 = ~n21024 & n21041 ;
  assign n21043 = ~\m_wb_adr_o[28]_pad  & ~n18716 ;
  assign n21044 = n13118 & n13119 ;
  assign n21045 = ~\wishbone_RxPointerMSB_reg[28]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n21046 = n13144 & n21045 ;
  assign n21047 = ~n13149 & ~n21046 ;
  assign n21048 = n13143 & n21047 ;
  assign n21049 = n13137 & n21048 ;
  assign n21050 = ~n13170 & ~n21049 ;
  assign n21051 = ~n21044 & ~n21050 ;
  assign n21052 = ~n21043 & n21051 ;
  assign n21053 = \m_wb_adr_o[28]_pad  & n13197 ;
  assign n21054 = \wishbone_TxPointerMSB_reg[28]/NET0131  & ~n13201 ;
  assign n21055 = \wishbone_RxPointerMSB_reg[28]/NET0131  & n13207 ;
  assign n21056 = ~n13196 & n21055 ;
  assign n21057 = ~n21054 & ~n21056 ;
  assign n21058 = ~n21053 & n21057 ;
  assign n21059 = ~n21052 & n21058 ;
  assign n21060 = ~\m_wb_adr_o[29]_pad  & ~n21044 ;
  assign n21061 = ~\wishbone_RxPointerMSB_reg[29]/NET0131  & ~\wishbone_rx_burst_cnt_reg[2]/NET0131  ;
  assign n21062 = n13144 & n21061 ;
  assign n21063 = ~n13149 & ~n21062 ;
  assign n21064 = n13143 & n21063 ;
  assign n21065 = n13137 & n21064 ;
  assign n21066 = ~n13170 & ~n21065 ;
  assign n21067 = ~n13121 & ~n21066 ;
  assign n21068 = ~n21060 & n21067 ;
  assign n21069 = \m_wb_adr_o[29]_pad  & n13197 ;
  assign n21070 = \wishbone_RxPointerMSB_reg[29]/NET0131  & n13207 ;
  assign n21071 = ~n13196 & n21070 ;
  assign n21072 = \wishbone_TxPointerMSB_reg[29]/NET0131  & ~n13201 ;
  assign n21073 = ~n21071 & ~n21072 ;
  assign n21074 = ~n21069 & n21073 ;
  assign n21075 = ~n21068 & n21074 ;
  assign n21076 = \m_wb_adr_o[5]_pad  & n13197 ;
  assign n21077 = \wishbone_RxPointerMSB_reg[5]/NET0131  & n13207 ;
  assign n21078 = ~n13196 & n21077 ;
  assign n21079 = ~n21076 & ~n21078 ;
  assign n21080 = \wishbone_TxPointerMSB_reg[5]/NET0131  & ~n13201 ;
  assign n21081 = ~\m_wb_adr_o[5]_pad  & ~n18710 ;
  assign n21082 = ~n13097 & ~n21081 ;
  assign n21083 = ~n15177 & n21082 ;
  assign n21084 = ~n21080 & ~n21083 ;
  assign n21085 = n21079 & n21084 ;
  assign n21086 = \m_wb_adr_o[6]_pad  & n13197 ;
  assign n21087 = \wishbone_RxPointerMSB_reg[6]/NET0131  & n13207 ;
  assign n21088 = ~n13196 & n21087 ;
  assign n21089 = ~n21086 & ~n21088 ;
  assign n21090 = \wishbone_TxPointerMSB_reg[6]/NET0131  & ~n13201 ;
  assign n21091 = \m_wb_adr_o[6]_pad  & n13097 ;
  assign n21092 = ~\m_wb_adr_o[6]_pad  & ~n13097 ;
  assign n21093 = ~n21091 & ~n21092 ;
  assign n21094 = ~n15177 & n21093 ;
  assign n21095 = ~n21090 & ~n21094 ;
  assign n21096 = n21089 & n21095 ;
  assign n21097 = \m_wb_adr_o[7]_pad  & n13197 ;
  assign n21098 = \wishbone_RxPointerMSB_reg[7]/NET0131  & n13207 ;
  assign n21099 = ~n13196 & n21098 ;
  assign n21100 = ~n21097 & ~n21099 ;
  assign n21101 = \wishbone_TxPointerMSB_reg[7]/NET0131  & ~n13201 ;
  assign n21102 = ~\m_wb_adr_o[7]_pad  & ~n21091 ;
  assign n21103 = ~n18669 & ~n21102 ;
  assign n21104 = ~n15177 & n21103 ;
  assign n21105 = ~n21101 & ~n21104 ;
  assign n21106 = n21100 & n21105 ;
  assign n21107 = \wishbone_TxPointerMSB_reg[9]/NET0131  & ~n13201 ;
  assign n21108 = \wishbone_RxPointerMSB_reg[9]/NET0131  & n13207 ;
  assign n21109 = ~n13196 & n21108 ;
  assign n21110 = ~n21107 & ~n21109 ;
  assign n21111 = \m_wb_adr_o[9]_pad  & n13197 ;
  assign n21112 = \m_wb_adr_o[9]_pad  & n13100 ;
  assign n21113 = ~\m_wb_adr_o[9]_pad  & ~n13100 ;
  assign n21114 = ~n21112 & ~n21113 ;
  assign n21115 = ~n15177 & n21114 ;
  assign n21116 = ~n21111 & ~n21115 ;
  assign n21117 = n21110 & n21116 ;
  assign n21118 = \wishbone_TxPointerMSB_reg[10]/NET0131  & ~n13201 ;
  assign n21119 = \wishbone_RxPointerMSB_reg[10]/NET0131  & n13207 ;
  assign n21120 = ~n13196 & n21119 ;
  assign n21121 = ~n21118 & ~n21120 ;
  assign n21122 = \m_wb_adr_o[10]_pad  & n13197 ;
  assign n21123 = ~\m_wb_adr_o[10]_pad  & ~n21112 ;
  assign n21124 = ~n18681 & ~n21123 ;
  assign n21125 = ~n15177 & n21124 ;
  assign n21126 = ~n21122 & ~n21125 ;
  assign n21127 = n21121 & n21126 ;
  assign n21128 = \wishbone_LatchedTxLength_reg[0]/NET0131  & ~n14046 ;
  assign n21129 = ~n19795 & ~n21128 ;
  assign n21130 = \wishbone_LatchedTxLength_reg[10]/NET0131  & ~n14046 ;
  assign n21131 = ~n17906 & ~n21130 ;
  assign n21132 = \wishbone_LatchedTxLength_reg[11]/NET0131  & ~n14046 ;
  assign n21133 = \wishbone_bd_ram_mem3_reg[80][27]/P0001  & n13516 ;
  assign n21134 = \wishbone_bd_ram_mem3_reg[3][27]/P0001  & n13354 ;
  assign n21135 = ~n21133 & ~n21134 ;
  assign n21136 = \wishbone_bd_ram_mem3_reg[52][27]/P0001  & n13988 ;
  assign n21137 = \wishbone_bd_ram_mem3_reg[73][27]/P0001  & n13456 ;
  assign n21138 = ~n21136 & ~n21137 ;
  assign n21139 = n21135 & n21138 ;
  assign n21140 = \wishbone_bd_ram_mem3_reg[124][27]/P0001  & n14024 ;
  assign n21141 = \wishbone_bd_ram_mem3_reg[169][27]/P0001  & n13541 ;
  assign n21142 = ~n21140 & ~n21141 ;
  assign n21143 = \wishbone_bd_ram_mem3_reg[128][27]/P0001  & n13652 ;
  assign n21144 = \wishbone_bd_ram_mem3_reg[200][27]/P0001  & n13922 ;
  assign n21145 = ~n21143 & ~n21144 ;
  assign n21146 = n21142 & n21145 ;
  assign n21147 = n21139 & n21146 ;
  assign n21148 = \wishbone_bd_ram_mem3_reg[214][27]/P0001  & n13938 ;
  assign n21149 = \wishbone_bd_ram_mem3_reg[113][27]/P0001  & n13882 ;
  assign n21150 = ~n21148 & ~n21149 ;
  assign n21151 = \wishbone_bd_ram_mem3_reg[119][27]/P0001  & n14033 ;
  assign n21152 = \wishbone_bd_ram_mem3_reg[132][27]/P0001  & n13927 ;
  assign n21153 = ~n21151 & ~n21152 ;
  assign n21154 = n21150 & n21153 ;
  assign n21155 = \wishbone_bd_ram_mem3_reg[55][27]/P0001  & n13618 ;
  assign n21156 = \wishbone_bd_ram_mem3_reg[219][27]/P0001  & n13577 ;
  assign n21157 = ~n21155 & ~n21156 ;
  assign n21158 = \wishbone_bd_ram_mem3_reg[147][27]/P0001  & n13702 ;
  assign n21159 = \wishbone_bd_ram_mem3_reg[180][27]/P0001  & n13650 ;
  assign n21160 = ~n21158 & ~n21159 ;
  assign n21161 = n21157 & n21160 ;
  assign n21162 = n21154 & n21161 ;
  assign n21163 = n21147 & n21162 ;
  assign n21164 = \wishbone_bd_ram_mem3_reg[120][27]/P0001  & n13550 ;
  assign n21165 = \wishbone_bd_ram_mem3_reg[177][27]/P0001  & n13863 ;
  assign n21166 = ~n21164 & ~n21165 ;
  assign n21167 = \wishbone_bd_ram_mem3_reg[68][27]/P0001  & n13379 ;
  assign n21168 = \wishbone_bd_ram_mem3_reg[136][27]/P0001  & n13963 ;
  assign n21169 = ~n21167 & ~n21168 ;
  assign n21170 = n21166 & n21169 ;
  assign n21171 = \wishbone_bd_ram_mem3_reg[225][27]/P0001  & n13719 ;
  assign n21172 = \wishbone_bd_ram_mem3_reg[242][27]/P0001  & n13383 ;
  assign n21173 = ~n21171 & ~n21172 ;
  assign n21174 = \wishbone_bd_ram_mem3_reg[74][27]/P0001  & n13564 ;
  assign n21175 = \wishbone_bd_ram_mem3_reg[37][27]/P0001  & n13710 ;
  assign n21176 = ~n21174 & ~n21175 ;
  assign n21177 = n21173 & n21176 ;
  assign n21178 = n21170 & n21177 ;
  assign n21179 = \wishbone_bd_ram_mem3_reg[89][27]/P0001  & n13910 ;
  assign n21180 = \wishbone_bd_ram_mem3_reg[252][27]/P0001  & n13986 ;
  assign n21181 = ~n21179 & ~n21180 ;
  assign n21182 = \wishbone_bd_ram_mem3_reg[227][27]/P0001  & n13388 ;
  assign n21183 = \wishbone_bd_ram_mem3_reg[13][27]/P0001  & n13844 ;
  assign n21184 = ~n21182 & ~n21183 ;
  assign n21185 = n21181 & n21184 ;
  assign n21186 = \wishbone_bd_ram_mem3_reg[16][27]/P0001  & n13695 ;
  assign n21187 = \wishbone_bd_ram_mem3_reg[175][27]/P0001  & n13674 ;
  assign n21188 = ~n21186 & ~n21187 ;
  assign n21189 = \wishbone_bd_ram_mem3_reg[107][27]/P0001  & n13476 ;
  assign n21190 = \wishbone_bd_ram_mem3_reg[181][27]/P0001  & n13587 ;
  assign n21191 = ~n21189 & ~n21190 ;
  assign n21192 = n21188 & n21191 ;
  assign n21193 = n21185 & n21192 ;
  assign n21194 = n21178 & n21193 ;
  assign n21195 = n21163 & n21194 ;
  assign n21196 = \wishbone_bd_ram_mem3_reg[243][27]/P0001  & n13575 ;
  assign n21197 = \wishbone_bd_ram_mem3_reg[122][27]/P0001  & n13679 ;
  assign n21198 = ~n21196 & ~n21197 ;
  assign n21199 = \wishbone_bd_ram_mem3_reg[91][27]/P0001  & n13954 ;
  assign n21200 = \wishbone_bd_ram_mem3_reg[65][27]/P0001  & n13842 ;
  assign n21201 = ~n21199 & ~n21200 ;
  assign n21202 = n21198 & n21201 ;
  assign n21203 = \wishbone_bd_ram_mem3_reg[205][27]/P0001  & n13947 ;
  assign n21204 = \wishbone_bd_ram_mem3_reg[78][27]/P0001  & n13277 ;
  assign n21205 = ~n21203 & ~n21204 ;
  assign n21206 = \wishbone_bd_ram_mem3_reg[221][27]/P0001  & n13641 ;
  assign n21207 = \wishbone_bd_ram_mem3_reg[88][27]/P0001  & n13347 ;
  assign n21208 = ~n21206 & ~n21207 ;
  assign n21209 = n21205 & n21208 ;
  assign n21210 = n21202 & n21209 ;
  assign n21211 = \wishbone_bd_ram_mem3_reg[182][27]/P0001  & n13598 ;
  assign n21212 = \wishbone_bd_ram_mem3_reg[51][27]/P0001  & n13880 ;
  assign n21213 = ~n21211 & ~n21212 ;
  assign n21214 = \wishbone_bd_ram_mem3_reg[101][27]/P0001  & n13772 ;
  assign n21215 = \wishbone_bd_ram_mem3_reg[210][27]/P0001  & n13443 ;
  assign n21216 = ~n21214 & ~n21215 ;
  assign n21217 = n21213 & n21216 ;
  assign n21218 = \wishbone_bd_ram_mem3_reg[162][27]/P0001  & n13726 ;
  assign n21219 = \wishbone_bd_ram_mem3_reg[238][27]/P0001  & n13819 ;
  assign n21220 = ~n21218 & ~n21219 ;
  assign n21221 = \wishbone_bd_ram_mem3_reg[47][27]/P0001  & n13436 ;
  assign n21222 = \wishbone_bd_ram_mem3_reg[201][27]/P0001  & n13600 ;
  assign n21223 = ~n21221 & ~n21222 ;
  assign n21224 = n21220 & n21223 ;
  assign n21225 = n21217 & n21224 ;
  assign n21226 = n21210 & n21225 ;
  assign n21227 = \wishbone_bd_ram_mem3_reg[208][27]/P0001  & n14010 ;
  assign n21228 = \wishbone_bd_ram_mem3_reg[192][27]/P0001  & n13390 ;
  assign n21229 = ~n21227 & ~n21228 ;
  assign n21230 = \wishbone_bd_ram_mem3_reg[171][27]/P0001  & n13422 ;
  assign n21231 = \wishbone_bd_ram_mem3_reg[98][27]/P0001  & n13569 ;
  assign n21232 = ~n21230 & ~n21231 ;
  assign n21233 = n21229 & n21232 ;
  assign n21234 = \wishbone_bd_ram_mem3_reg[248][27]/P0001  & n13647 ;
  assign n21235 = \wishbone_bd_ram_mem3_reg[126][27]/P0001  & n13786 ;
  assign n21236 = ~n21234 & ~n21235 ;
  assign n21237 = \wishbone_bd_ram_mem3_reg[62][27]/P0001  & n13529 ;
  assign n21238 = \wishbone_bd_ram_mem3_reg[58][27]/P0001  & n13949 ;
  assign n21239 = ~n21237 & ~n21238 ;
  assign n21240 = n21236 & n21239 ;
  assign n21241 = n21233 & n21240 ;
  assign n21242 = \wishbone_bd_ram_mem3_reg[133][27]/P0001  & n13492 ;
  assign n21243 = \wishbone_bd_ram_mem3_reg[60][27]/P0001  & n13790 ;
  assign n21244 = ~n21242 & ~n21243 ;
  assign n21245 = \wishbone_bd_ram_mem3_reg[123][27]/P0001  & n13749 ;
  assign n21246 = \wishbone_bd_ram_mem3_reg[84][27]/P0001  & n13385 ;
  assign n21247 = ~n21245 & ~n21246 ;
  assign n21248 = n21244 & n21247 ;
  assign n21249 = \wishbone_bd_ram_mem3_reg[75][27]/P0001  & n13605 ;
  assign n21250 = \wishbone_bd_ram_mem3_reg[25][27]/P0001  & n13742 ;
  assign n21251 = ~n21249 & ~n21250 ;
  assign n21252 = \wishbone_bd_ram_mem3_reg[43][27]/P0001  & n13761 ;
  assign n21253 = \wishbone_bd_ram_mem3_reg[153][27]/P0001  & n13309 ;
  assign n21254 = ~n21252 & ~n21253 ;
  assign n21255 = n21251 & n21254 ;
  assign n21256 = n21248 & n21255 ;
  assign n21257 = n21241 & n21256 ;
  assign n21258 = n21226 & n21257 ;
  assign n21259 = n21195 & n21258 ;
  assign n21260 = \wishbone_bd_ram_mem3_reg[160][27]/P0001  & n13271 ;
  assign n21261 = \wishbone_bd_ram_mem3_reg[198][27]/P0001  & n13592 ;
  assign n21262 = ~n21260 & ~n21261 ;
  assign n21263 = \wishbone_bd_ram_mem3_reg[183][27]/P0001  & n13645 ;
  assign n21264 = \wishbone_bd_ram_mem3_reg[121][27]/P0001  & n13983 ;
  assign n21265 = ~n21263 & ~n21264 ;
  assign n21266 = n21262 & n21265 ;
  assign n21267 = \wishbone_bd_ram_mem3_reg[247][27]/P0001  & n13571 ;
  assign n21268 = \wishbone_bd_ram_mem3_reg[232][27]/P0001  & n13510 ;
  assign n21269 = ~n21267 & ~n21268 ;
  assign n21270 = \wishbone_bd_ram_mem3_reg[34][27]/P0001  & n13450 ;
  assign n21271 = \wishbone_bd_ram_mem3_reg[8][27]/P0001  & n13459 ;
  assign n21272 = ~n21270 & ~n21271 ;
  assign n21273 = n21269 & n21272 ;
  assign n21274 = n21266 & n21273 ;
  assign n21275 = \wishbone_bd_ram_mem3_reg[111][27]/P0001  & n13471 ;
  assign n21276 = \wishbone_bd_ram_mem3_reg[117][27]/P0001  & n13557 ;
  assign n21277 = ~n21275 & ~n21276 ;
  assign n21278 = \wishbone_bd_ram_mem3_reg[193][27]/P0001  & n14022 ;
  assign n21279 = \wishbone_bd_ram_mem3_reg[220][27]/P0001  & n13965 ;
  assign n21280 = ~n21278 & ~n21279 ;
  assign n21281 = n21277 & n21280 ;
  assign n21282 = \wishbone_bd_ram_mem3_reg[176][27]/P0001  & n13262 ;
  assign n21283 = \wishbone_bd_ram_mem3_reg[148][27]/P0001  & n13868 ;
  assign n21284 = ~n21282 & ~n21283 ;
  assign n21285 = \wishbone_bd_ram_mem3_reg[96][27]/P0001  & n13425 ;
  assign n21286 = \wishbone_bd_ram_mem3_reg[184][27]/P0001  & n13960 ;
  assign n21287 = ~n21285 & ~n21286 ;
  assign n21288 = n21284 & n21287 ;
  assign n21289 = n21281 & n21288 ;
  assign n21290 = n21274 & n21289 ;
  assign n21291 = \wishbone_bd_ram_mem3_reg[118][27]/P0001  & n13589 ;
  assign n21292 = \wishbone_bd_ram_mem3_reg[203][27]/P0001  & n13816 ;
  assign n21293 = ~n21291 & ~n21292 ;
  assign n21294 = \wishbone_bd_ram_mem3_reg[131][27]/P0001  & n13358 ;
  assign n21295 = \wishbone_bd_ram_mem3_reg[70][27]/P0001  & n13339 ;
  assign n21296 = ~n21294 & ~n21295 ;
  assign n21297 = n21293 & n21296 ;
  assign n21298 = \wishbone_bd_ram_mem3_reg[30][27]/P0001  & n13713 ;
  assign n21299 = \wishbone_bd_ram_mem3_reg[26][27]/P0001  & n13521 ;
  assign n21300 = ~n21298 & ~n21299 ;
  assign n21301 = \wishbone_bd_ram_mem3_reg[24][27]/P0001  & n13970 ;
  assign n21302 = \wishbone_bd_ram_mem3_reg[104][27]/P0001  & n13684 ;
  assign n21303 = ~n21301 & ~n21302 ;
  assign n21304 = n21300 & n21303 ;
  assign n21305 = n21297 & n21304 ;
  assign n21306 = \wishbone_bd_ram_mem3_reg[4][27]/P0001  & n13527 ;
  assign n21307 = \wishbone_bd_ram_mem3_reg[94][27]/P0001  & n13833 ;
  assign n21308 = ~n21306 & ~n21307 ;
  assign n21309 = \wishbone_bd_ram_mem3_reg[77][27]/P0001  & n13935 ;
  assign n21310 = \wishbone_bd_ram_mem3_reg[32][27]/P0001  & n13736 ;
  assign n21311 = ~n21309 & ~n21310 ;
  assign n21312 = n21308 & n21311 ;
  assign n21313 = \wishbone_bd_ram_mem3_reg[103][27]/P0001  & n13320 ;
  assign n21314 = \wishbone_bd_ram_mem3_reg[216][27]/P0001  & n14005 ;
  assign n21315 = ~n21313 & ~n21314 ;
  assign n21316 = \wishbone_bd_ram_mem3_reg[212][27]/P0001  & n13634 ;
  assign n21317 = \wishbone_bd_ram_mem3_reg[155][27]/P0001  & n13738 ;
  assign n21318 = ~n21316 & ~n21317 ;
  assign n21319 = n21315 & n21318 ;
  assign n21320 = n21312 & n21319 ;
  assign n21321 = n21305 & n21320 ;
  assign n21322 = n21290 & n21321 ;
  assign n21323 = \wishbone_bd_ram_mem3_reg[6][27]/P0001  & n13915 ;
  assign n21324 = \wishbone_bd_ram_mem3_reg[110][27]/P0001  & n14030 ;
  assign n21325 = ~n21323 & ~n21324 ;
  assign n21326 = \wishbone_bd_ram_mem3_reg[143][27]/P0001  & n13461 ;
  assign n21327 = \wishbone_bd_ram_mem3_reg[173][27]/P0001  & n13360 ;
  assign n21328 = ~n21326 & ~n21327 ;
  assign n21329 = n21325 & n21328 ;
  assign n21330 = \wishbone_bd_ram_mem3_reg[204][27]/P0001  & n13821 ;
  assign n21331 = \wishbone_bd_ram_mem3_reg[213][27]/P0001  & n13870 ;
  assign n21332 = ~n21330 & ~n21331 ;
  assign n21333 = \wishbone_bd_ram_mem3_reg[5][27]/P0001  & n13243 ;
  assign n21334 = \wishbone_bd_ram_mem3_reg[61][27]/P0001  & n13544 ;
  assign n21335 = ~n21333 & ~n21334 ;
  assign n21336 = n21332 & n21335 ;
  assign n21337 = n21329 & n21336 ;
  assign n21338 = \wishbone_bd_ram_mem3_reg[239][27]/P0001  & n13349 ;
  assign n21339 = \wishbone_bd_ram_mem3_reg[164][27]/P0001  & n13236 ;
  assign n21340 = ~n21338 & ~n21339 ;
  assign n21341 = \wishbone_bd_ram_mem3_reg[154][27]/P0001  & n13403 ;
  assign n21342 = \wishbone_bd_ram_mem3_reg[244][27]/P0001  & n13474 ;
  assign n21343 = ~n21341 & ~n21342 ;
  assign n21344 = n21340 & n21343 ;
  assign n21345 = \wishbone_bd_ram_mem3_reg[189][27]/P0001  & n14001 ;
  assign n21346 = \wishbone_bd_ram_mem3_reg[249][27]/P0001  & n13431 ;
  assign n21347 = ~n21345 & ~n21346 ;
  assign n21348 = \wishbone_bd_ram_mem3_reg[138][27]/P0001  & n13398 ;
  assign n21349 = \wishbone_bd_ram_mem3_reg[99][27]/P0001  & n13996 ;
  assign n21350 = ~n21348 & ~n21349 ;
  assign n21351 = n21347 & n21350 ;
  assign n21352 = n21344 & n21351 ;
  assign n21353 = n21337 & n21352 ;
  assign n21354 = \wishbone_bd_ram_mem3_reg[49][27]/P0001  & n13929 ;
  assign n21355 = \wishbone_bd_ram_mem3_reg[53][27]/P0001  & n13875 ;
  assign n21356 = ~n21354 & ~n21355 ;
  assign n21357 = \wishbone_bd_ram_mem3_reg[222][27]/P0001  & n13721 ;
  assign n21358 = \wishbone_bd_ram_mem3_reg[31][27]/P0001  & n13758 ;
  assign n21359 = ~n21357 & ~n21358 ;
  assign n21360 = n21356 & n21359 ;
  assign n21361 = \wishbone_bd_ram_mem3_reg[134][27]/P0001  & n13494 ;
  assign n21362 = \wishbone_bd_ram_mem3_reg[187][27]/P0001  & n13756 ;
  assign n21363 = ~n21361 & ~n21362 ;
  assign n21364 = \wishbone_bd_ram_mem3_reg[7][27]/P0001  & n13546 ;
  assign n21365 = \wishbone_bd_ram_mem3_reg[63][27]/P0001  & n13327 ;
  assign n21366 = ~n21364 & ~n21365 ;
  assign n21367 = n21363 & n21366 ;
  assign n21368 = n21360 & n21367 ;
  assign n21369 = \wishbone_bd_ram_mem3_reg[127][27]/P0001  & n13803 ;
  assign n21370 = \wishbone_bd_ram_mem3_reg[116][27]/P0001  & n13865 ;
  assign n21371 = ~n21369 & ~n21370 ;
  assign n21372 = \wishbone_bd_ram_mem3_reg[159][27]/P0001  & n13627 ;
  assign n21373 = \wishbone_bd_ram_mem3_reg[233][27]/P0001  & n13332 ;
  assign n21374 = ~n21372 & ~n21373 ;
  assign n21375 = n21371 & n21374 ;
  assign n21376 = \wishbone_bd_ram_mem3_reg[179][27]/P0001  & n14035 ;
  assign n21377 = \wishbone_bd_ram_mem3_reg[190][27]/P0001  & n13365 ;
  assign n21378 = ~n21376 & ~n21377 ;
  assign n21379 = \wishbone_bd_ram_mem3_reg[130][27]/P0001  & n13427 ;
  assign n21380 = \wishbone_bd_ram_mem3_reg[39][27]/P0001  & n13893 ;
  assign n21381 = ~n21379 & ~n21380 ;
  assign n21382 = n21378 & n21381 ;
  assign n21383 = n21375 & n21382 ;
  assign n21384 = n21368 & n21383 ;
  assign n21385 = n21353 & n21384 ;
  assign n21386 = n21322 & n21385 ;
  assign n21387 = n21259 & n21386 ;
  assign n21388 = \wishbone_bd_ram_mem3_reg[18][27]/P0001  & n13532 ;
  assign n21389 = \wishbone_bd_ram_mem3_reg[1][27]/P0001  & n13888 ;
  assign n21390 = ~n21388 & ~n21389 ;
  assign n21391 = \wishbone_bd_ram_mem3_reg[167][27]/P0001  & n13940 ;
  assign n21392 = \wishbone_bd_ram_mem3_reg[250][27]/P0001  & n13677 ;
  assign n21393 = ~n21391 & ~n21392 ;
  assign n21394 = n21390 & n21393 ;
  assign n21395 = \wishbone_bd_ram_mem3_reg[149][27]/P0001  & n13469 ;
  assign n21396 = \wishbone_bd_ram_mem3_reg[21][27]/P0001  & n13438 ;
  assign n21397 = ~n21395 & ~n21396 ;
  assign n21398 = \wishbone_bd_ram_mem3_reg[207][27]/P0001  & n13826 ;
  assign n21399 = \wishbone_bd_ram_mem3_reg[165][27]/P0001  & n14028 ;
  assign n21400 = ~n21398 & ~n21399 ;
  assign n21401 = n21397 & n21400 ;
  assign n21402 = n21394 & n21401 ;
  assign n21403 = \wishbone_bd_ram_mem3_reg[174][27]/P0001  & n13899 ;
  assign n21404 = \wishbone_bd_ram_mem3_reg[40][27]/P0001  & n13661 ;
  assign n21405 = ~n21403 & ~n21404 ;
  assign n21406 = \wishbone_bd_ram_mem3_reg[236][27]/P0001  & n13480 ;
  assign n21407 = \wishbone_bd_ram_mem3_reg[81][27]/P0001  & n13409 ;
  assign n21408 = ~n21406 & ~n21407 ;
  assign n21409 = n21405 & n21408 ;
  assign n21410 = \wishbone_bd_ram_mem3_reg[157][27]/P0001  & n13445 ;
  assign n21411 = \wishbone_bd_ram_mem3_reg[166][27]/P0001  & n13999 ;
  assign n21412 = ~n21410 & ~n21411 ;
  assign n21413 = \wishbone_bd_ram_mem3_reg[228][27]/P0001  & n13497 ;
  assign n21414 = \wishbone_bd_ram_mem3_reg[28][27]/P0001  & n13810 ;
  assign n21415 = ~n21413 & ~n21414 ;
  assign n21416 = n21412 & n21415 ;
  assign n21417 = n21409 & n21416 ;
  assign n21418 = n21402 & n21417 ;
  assign n21419 = \wishbone_bd_ram_mem3_reg[206][27]/P0001  & n13414 ;
  assign n21420 = \wishbone_bd_ram_mem3_reg[9][27]/P0001  & n13580 ;
  assign n21421 = ~n21419 & ~n21420 ;
  assign n21422 = \wishbone_bd_ram_mem3_reg[27][27]/P0001  & n13251 ;
  assign n21423 = \wishbone_bd_ram_mem3_reg[95][27]/P0001  & n13317 ;
  assign n21424 = ~n21422 & ~n21423 ;
  assign n21425 = n21421 & n21424 ;
  assign n21426 = \wishbone_bd_ram_mem3_reg[240][27]/P0001  & n13352 ;
  assign n21427 = \wishbone_bd_ram_mem3_reg[97][27]/P0001  & n13724 ;
  assign n21428 = ~n21426 & ~n21427 ;
  assign n21429 = \wishbone_bd_ram_mem3_reg[139][27]/P0001  & n13566 ;
  assign n21430 = \wishbone_bd_ram_mem3_reg[234][27]/P0001  & n13781 ;
  assign n21431 = ~n21429 & ~n21430 ;
  assign n21432 = n21428 & n21431 ;
  assign n21433 = n21425 & n21432 ;
  assign n21434 = \wishbone_bd_ram_mem3_reg[38][27]/P0001  & n13828 ;
  assign n21435 = \wishbone_bd_ram_mem3_reg[2][27]/P0001  & n13975 ;
  assign n21436 = ~n21434 & ~n21435 ;
  assign n21437 = \wishbone_bd_ram_mem3_reg[115][27]/P0001  & n13747 ;
  assign n21438 = \wishbone_bd_ram_mem3_reg[23][27]/P0001  & n13857 ;
  assign n21439 = ~n21437 & ~n21438 ;
  assign n21440 = n21436 & n21439 ;
  assign n21441 = \wishbone_bd_ram_mem3_reg[163][27]/P0001  & n13255 ;
  assign n21442 = \wishbone_bd_ram_mem3_reg[41][27]/P0001  & n14017 ;
  assign n21443 = ~n21441 & ~n21442 ;
  assign n21444 = \wishbone_bd_ram_mem3_reg[36][27]/P0001  & n13639 ;
  assign n21445 = \wishbone_bd_ram_mem3_reg[71][27]/P0001  & n13636 ;
  assign n21446 = ~n21444 & ~n21445 ;
  assign n21447 = n21443 & n21446 ;
  assign n21448 = n21440 & n21447 ;
  assign n21449 = n21433 & n21448 ;
  assign n21450 = n21418 & n21449 ;
  assign n21451 = \wishbone_bd_ram_mem3_reg[253][27]/P0001  & n13708 ;
  assign n21452 = \wishbone_bd_ram_mem3_reg[109][27]/P0001  & n13306 ;
  assign n21453 = ~n21451 & ~n21452 ;
  assign n21454 = \wishbone_bd_ram_mem3_reg[69][27]/P0001  & n13487 ;
  assign n21455 = \wishbone_bd_ram_mem3_reg[199][27]/P0001  & n13499 ;
  assign n21456 = ~n21454 & ~n21455 ;
  assign n21457 = n21453 & n21456 ;
  assign n21458 = \wishbone_bd_ram_mem3_reg[245][27]/P0001  & n13877 ;
  assign n21459 = \wishbone_bd_ram_mem3_reg[146][27]/P0001  & n13958 ;
  assign n21460 = ~n21458 & ~n21459 ;
  assign n21461 = \wishbone_bd_ram_mem3_reg[45][27]/P0001  & n13420 ;
  assign n21462 = \wishbone_bd_ram_mem3_reg[66][27]/P0001  & n13603 ;
  assign n21463 = ~n21461 & ~n21462 ;
  assign n21464 = n21460 & n21463 ;
  assign n21465 = n21457 & n21464 ;
  assign n21466 = \wishbone_bd_ram_mem3_reg[72][27]/P0001  & n13582 ;
  assign n21467 = \wishbone_bd_ram_mem3_reg[241][27]/P0001  & n13854 ;
  assign n21468 = ~n21466 & ~n21467 ;
  assign n21469 = \wishbone_bd_ram_mem3_reg[56][27]/P0001  & n13611 ;
  assign n21470 = \wishbone_bd_ram_mem3_reg[140][27]/P0001  & n13287 ;
  assign n21471 = ~n21469 & ~n21470 ;
  assign n21472 = n21468 & n21471 ;
  assign n21473 = \wishbone_bd_ram_mem3_reg[57][27]/P0001  & n13731 ;
  assign n21474 = \wishbone_bd_ram_mem3_reg[100][27]/P0001  & n13401 ;
  assign n21475 = ~n21473 & ~n21474 ;
  assign n21476 = \wishbone_bd_ram_mem3_reg[59][27]/P0001  & n13613 ;
  assign n21477 = \wishbone_bd_ram_mem3_reg[10][27]/P0001  & n13837 ;
  assign n21478 = ~n21476 & ~n21477 ;
  assign n21479 = n21475 & n21478 ;
  assign n21480 = n21472 & n21479 ;
  assign n21481 = n21465 & n21480 ;
  assign n21482 = \wishbone_bd_ram_mem3_reg[106][27]/P0001  & n13555 ;
  assign n21483 = \wishbone_bd_ram_mem3_reg[255][27]/P0001  & n13952 ;
  assign n21484 = ~n21482 & ~n21483 ;
  assign n21485 = \wishbone_bd_ram_mem3_reg[87][27]/P0001  & n13691 ;
  assign n21486 = \wishbone_bd_ram_mem3_reg[15][27]/P0001  & n13797 ;
  assign n21487 = ~n21485 & ~n21486 ;
  assign n21488 = n21484 & n21487 ;
  assign n21489 = \wishbone_bd_ram_mem3_reg[230][27]/P0001  & n13994 ;
  assign n21490 = \wishbone_bd_ram_mem3_reg[170][27]/P0001  & n14007 ;
  assign n21491 = ~n21489 & ~n21490 ;
  assign n21492 = \wishbone_bd_ram_mem3_reg[217][27]/P0001  & n13767 ;
  assign n21493 = \wishbone_bd_ram_mem3_reg[191][27]/P0001  & n14012 ;
  assign n21494 = ~n21492 & ~n21493 ;
  assign n21495 = n21491 & n21494 ;
  assign n21496 = n21488 & n21495 ;
  assign n21497 = \wishbone_bd_ram_mem3_reg[194][27]/P0001  & n13624 ;
  assign n21498 = \wishbone_bd_ram_mem3_reg[161][27]/P0001  & n13505 ;
  assign n21499 = ~n21497 & ~n21498 ;
  assign n21500 = \wishbone_bd_ram_mem3_reg[14][27]/P0001  & n13972 ;
  assign n21501 = \wishbone_bd_ram_mem3_reg[202][27]/P0001  & n13268 ;
  assign n21502 = ~n21500 & ~n21501 ;
  assign n21503 = n21499 & n21502 ;
  assign n21504 = \wishbone_bd_ram_mem3_reg[22][27]/P0001  & n13744 ;
  assign n21505 = \wishbone_bd_ram_mem3_reg[64][27]/P0001  & n13904 ;
  assign n21506 = ~n21504 & ~n21505 ;
  assign n21507 = \wishbone_bd_ram_mem3_reg[17][27]/P0001  & n13324 ;
  assign n21508 = \wishbone_bd_ram_mem3_reg[33][27]/P0001  & n13933 ;
  assign n21509 = ~n21507 & ~n21508 ;
  assign n21510 = n21506 & n21509 ;
  assign n21511 = n21503 & n21510 ;
  assign n21512 = n21496 & n21511 ;
  assign n21513 = n21481 & n21512 ;
  assign n21514 = n21450 & n21513 ;
  assign n21515 = \wishbone_bd_ram_mem3_reg[20][27]/P0001  & n13839 ;
  assign n21516 = \wishbone_bd_ram_mem3_reg[172][27]/P0001  & n13377 ;
  assign n21517 = ~n21515 & ~n21516 ;
  assign n21518 = \wishbone_bd_ram_mem3_reg[218][27]/P0001  & n13792 ;
  assign n21519 = \wishbone_bd_ram_mem3_reg[93][27]/P0001  & n13891 ;
  assign n21520 = ~n21518 & ~n21519 ;
  assign n21521 = n21517 & n21520 ;
  assign n21522 = \wishbone_bd_ram_mem3_reg[125][27]/P0001  & n13396 ;
  assign n21523 = \wishbone_bd_ram_mem3_reg[54][27]/P0001  & n13622 ;
  assign n21524 = ~n21522 & ~n21523 ;
  assign n21525 = \wishbone_bd_ram_mem3_reg[141][27]/P0001  & n13852 ;
  assign n21526 = \wishbone_bd_ram_mem3_reg[178][27]/P0001  & n13301 ;
  assign n21527 = ~n21525 & ~n21526 ;
  assign n21528 = n21524 & n21527 ;
  assign n21529 = n21521 & n21528 ;
  assign n21530 = \wishbone_bd_ram_mem3_reg[168][27]/P0001  & n13795 ;
  assign n21531 = \wishbone_bd_ram_mem3_reg[254][27]/P0001  & n13283 ;
  assign n21532 = ~n21530 & ~n21531 ;
  assign n21533 = \wishbone_bd_ram_mem3_reg[46][27]/P0001  & n13298 ;
  assign n21534 = \wishbone_bd_ram_mem3_reg[223][27]/P0001  & n13335 ;
  assign n21535 = ~n21533 & ~n21534 ;
  assign n21536 = n21532 & n21535 ;
  assign n21537 = \wishbone_bd_ram_mem3_reg[11][27]/P0001  & n13774 ;
  assign n21538 = \wishbone_bd_ram_mem3_reg[79][27]/P0001  & n13779 ;
  assign n21539 = ~n21537 & ~n21538 ;
  assign n21540 = \wishbone_bd_ram_mem3_reg[137][27]/P0001  & n13808 ;
  assign n21541 = \wishbone_bd_ram_mem3_reg[135][27]/P0001  & n13672 ;
  assign n21542 = ~n21540 & ~n21541 ;
  assign n21543 = n21539 & n21542 ;
  assign n21544 = n21536 & n21543 ;
  assign n21545 = n21529 & n21544 ;
  assign n21546 = \wishbone_bd_ram_mem3_reg[102][27]/P0001  & n13534 ;
  assign n21547 = \wishbone_bd_ram_mem3_reg[35][27]/P0001  & n13523 ;
  assign n21548 = ~n21546 & ~n21547 ;
  assign n21549 = \wishbone_bd_ram_mem3_reg[29][27]/P0001  & n13412 ;
  assign n21550 = \wishbone_bd_ram_mem3_reg[151][27]/P0001  & n13697 ;
  assign n21551 = ~n21549 & ~n21550 ;
  assign n21552 = n21548 & n21551 ;
  assign n21553 = \wishbone_bd_ram_mem3_reg[144][27]/P0001  & n13508 ;
  assign n21554 = \wishbone_bd_ram_mem3_reg[142][27]/P0001  & n13448 ;
  assign n21555 = ~n21553 & ~n21554 ;
  assign n21556 = \wishbone_bd_ram_mem3_reg[83][27]/P0001  & n13454 ;
  assign n21557 = \wishbone_bd_ram_mem3_reg[76][27]/P0001  & n13831 ;
  assign n21558 = ~n21556 & ~n21557 ;
  assign n21559 = n21555 & n21558 ;
  assign n21560 = n21552 & n21559 ;
  assign n21561 = \wishbone_bd_ram_mem3_reg[209][27]/P0001  & n13689 ;
  assign n21562 = \wishbone_bd_ram_mem3_reg[158][27]/P0001  & n13294 ;
  assign n21563 = ~n21561 & ~n21562 ;
  assign n21564 = \wishbone_bd_ram_mem3_reg[112][27]/P0001  & n13482 ;
  assign n21565 = \wishbone_bd_ram_mem3_reg[85][27]/P0001  & n13784 ;
  assign n21566 = ~n21564 & ~n21565 ;
  assign n21567 = n21563 & n21566 ;
  assign n21568 = \wishbone_bd_ram_mem3_reg[12][27]/P0001  & n13733 ;
  assign n21569 = \wishbone_bd_ram_mem3_reg[86][27]/P0001  & n13485 ;
  assign n21570 = ~n21568 & ~n21569 ;
  assign n21571 = \wishbone_bd_ram_mem3_reg[215][27]/P0001  & n13901 ;
  assign n21572 = \wishbone_bd_ram_mem3_reg[129][27]/P0001  & n13629 ;
  assign n21573 = ~n21571 & ~n21572 ;
  assign n21574 = n21570 & n21573 ;
  assign n21575 = n21567 & n21574 ;
  assign n21576 = n21560 & n21575 ;
  assign n21577 = n21545 & n21576 ;
  assign n21578 = \wishbone_bd_ram_mem3_reg[197][27]/P0001  & n13594 ;
  assign n21579 = \wishbone_bd_ram_mem3_reg[67][27]/P0001  & n13663 ;
  assign n21580 = ~n21578 & ~n21579 ;
  assign n21581 = \wishbone_bd_ram_mem3_reg[114][27]/P0001  & n13763 ;
  assign n21582 = \wishbone_bd_ram_mem3_reg[188][27]/P0001  & n13407 ;
  assign n21583 = ~n21581 & ~n21582 ;
  assign n21584 = n21580 & n21583 ;
  assign n21585 = \wishbone_bd_ram_mem3_reg[145][27]/P0001  & n13715 ;
  assign n21586 = \wishbone_bd_ram_mem3_reg[186][27]/P0001  & n13616 ;
  assign n21587 = ~n21585 & ~n21586 ;
  assign n21588 = \wishbone_bd_ram_mem3_reg[150][27]/P0001  & n13666 ;
  assign n21589 = \wishbone_bd_ram_mem3_reg[211][27]/P0001  & n13805 ;
  assign n21590 = ~n21588 & ~n21589 ;
  assign n21591 = n21587 & n21590 ;
  assign n21592 = n21584 & n21591 ;
  assign n21593 = \wishbone_bd_ram_mem3_reg[42][27]/P0001  & n13341 ;
  assign n21594 = \wishbone_bd_ram_mem3_reg[48][27]/P0001  & n13917 ;
  assign n21595 = ~n21593 & ~n21594 ;
  assign n21596 = \wishbone_bd_ram_mem3_reg[44][27]/P0001  & n13291 ;
  assign n21597 = \wishbone_bd_ram_mem3_reg[237][27]/P0001  & n13924 ;
  assign n21598 = ~n21596 & ~n21597 ;
  assign n21599 = n21595 & n21598 ;
  assign n21600 = \wishbone_bd_ram_mem3_reg[226][27]/P0001  & n13668 ;
  assign n21601 = \wishbone_bd_ram_mem3_reg[108][27]/P0001  & n13814 ;
  assign n21602 = ~n21600 & ~n21601 ;
  assign n21603 = \wishbone_bd_ram_mem3_reg[246][27]/P0001  & n13981 ;
  assign n21604 = \wishbone_bd_ram_mem3_reg[0][27]/P0001  & n13539 ;
  assign n21605 = ~n21603 & ~n21604 ;
  assign n21606 = n21602 & n21605 ;
  assign n21607 = n21599 & n21606 ;
  assign n21608 = n21592 & n21607 ;
  assign n21609 = \wishbone_bd_ram_mem3_reg[156][27]/P0001  & n13769 ;
  assign n21610 = \wishbone_bd_ram_mem3_reg[92][27]/P0001  & n13859 ;
  assign n21611 = ~n21609 & ~n21610 ;
  assign n21612 = \wishbone_bd_ram_mem3_reg[90][27]/P0001  & n13906 ;
  assign n21613 = \wishbone_bd_ram_mem3_reg[231][27]/P0001  & n13363 ;
  assign n21614 = ~n21612 & ~n21613 ;
  assign n21615 = n21611 & n21614 ;
  assign n21616 = \wishbone_bd_ram_mem3_reg[251][27]/P0001  & n14019 ;
  assign n21617 = \wishbone_bd_ram_mem3_reg[235][27]/P0001  & n13518 ;
  assign n21618 = ~n21616 & ~n21617 ;
  assign n21619 = \wishbone_bd_ram_mem3_reg[152][27]/P0001  & n13912 ;
  assign n21620 = \wishbone_bd_ram_mem3_reg[224][27]/P0001  & n13433 ;
  assign n21621 = ~n21619 & ~n21620 ;
  assign n21622 = n21618 & n21621 ;
  assign n21623 = n21615 & n21622 ;
  assign n21624 = \wishbone_bd_ram_mem3_reg[19][27]/P0001  & n13886 ;
  assign n21625 = \wishbone_bd_ram_mem3_reg[229][27]/P0001  & n13552 ;
  assign n21626 = ~n21624 & ~n21625 ;
  assign n21627 = \wishbone_bd_ram_mem3_reg[196][27]/P0001  & n13977 ;
  assign n21628 = \wishbone_bd_ram_mem3_reg[105][27]/P0001  & n13503 ;
  assign n21629 = ~n21627 & ~n21628 ;
  assign n21630 = n21626 & n21629 ;
  assign n21631 = \wishbone_bd_ram_mem3_reg[82][27]/P0001  & n13374 ;
  assign n21632 = \wishbone_bd_ram_mem3_reg[195][27]/P0001  & n13700 ;
  assign n21633 = ~n21631 & ~n21632 ;
  assign n21634 = \wishbone_bd_ram_mem3_reg[50][27]/P0001  & n13686 ;
  assign n21635 = \wishbone_bd_ram_mem3_reg[185][27]/P0001  & n13372 ;
  assign n21636 = ~n21634 & ~n21635 ;
  assign n21637 = n21633 & n21636 ;
  assign n21638 = n21630 & n21637 ;
  assign n21639 = n21623 & n21638 ;
  assign n21640 = n21608 & n21639 ;
  assign n21641 = n21577 & n21640 ;
  assign n21642 = n21514 & n21641 ;
  assign n21643 = n21387 & n21642 ;
  assign n21644 = n14047 & ~n21643 ;
  assign n21645 = ~n21132 & ~n21644 ;
  assign n21646 = \wishbone_LatchedTxLength_reg[12]/NET0131  & ~n14046 ;
  assign n21647 = ~n14048 & ~n21646 ;
  assign n21648 = \wishbone_LatchedTxLength_reg[13]/NET0131  & ~n14046 ;
  assign n21649 = ~n14594 & ~n21648 ;
  assign n21650 = \wishbone_LatchedTxLength_reg[14]/NET0131  & ~n14046 ;
  assign n21651 = ~n15115 & ~n21650 ;
  assign n21652 = ~\wishbone_LatchedTxLength_reg[15]/NET0131  & ~n14046 ;
  assign n21653 = ~n14046 & ~n21652 ;
  assign n21654 = ~wb_rst_i_pad & ~n21652 ;
  assign n21655 = ~n20314 & n21654 ;
  assign n21656 = ~n21653 & ~n21655 ;
  assign n21657 = \wishbone_LatchedTxLength_reg[1]/NET0131  & ~n14046 ;
  assign n21658 = ~n20834 & ~n21657 ;
  assign n21659 = \wishbone_LatchedTxLength_reg[2]/NET0131  & ~n14046 ;
  assign n21660 = ~n19274 & ~n21659 ;
  assign n21661 = \wishbone_LatchedTxLength_reg[3]/NET0131  & ~n14046 ;
  assign n21662 = \wishbone_bd_ram_mem2_reg[103][19]/P0001  & n13320 ;
  assign n21663 = \wishbone_bd_ram_mem2_reg[223][19]/P0001  & n13335 ;
  assign n21664 = ~n21662 & ~n21663 ;
  assign n21665 = \wishbone_bd_ram_mem2_reg[203][19]/P0001  & n13816 ;
  assign n21666 = \wishbone_bd_ram_mem2_reg[181][19]/P0001  & n13587 ;
  assign n21667 = ~n21665 & ~n21666 ;
  assign n21668 = n21664 & n21667 ;
  assign n21669 = \wishbone_bd_ram_mem2_reg[73][19]/P0001  & n13456 ;
  assign n21670 = \wishbone_bd_ram_mem2_reg[187][19]/P0001  & n13756 ;
  assign n21671 = ~n21669 & ~n21670 ;
  assign n21672 = \wishbone_bd_ram_mem2_reg[26][19]/P0001  & n13521 ;
  assign n21673 = \wishbone_bd_ram_mem2_reg[67][19]/P0001  & n13663 ;
  assign n21674 = ~n21672 & ~n21673 ;
  assign n21675 = n21671 & n21674 ;
  assign n21676 = n21668 & n21675 ;
  assign n21677 = \wishbone_bd_ram_mem2_reg[193][19]/P0001  & n14022 ;
  assign n21678 = \wishbone_bd_ram_mem2_reg[42][19]/P0001  & n13341 ;
  assign n21679 = ~n21677 & ~n21678 ;
  assign n21680 = \wishbone_bd_ram_mem2_reg[106][19]/P0001  & n13555 ;
  assign n21681 = \wishbone_bd_ram_mem2_reg[15][19]/P0001  & n13797 ;
  assign n21682 = ~n21680 & ~n21681 ;
  assign n21683 = n21679 & n21682 ;
  assign n21684 = \wishbone_bd_ram_mem2_reg[249][19]/P0001  & n13431 ;
  assign n21685 = \wishbone_bd_ram_mem2_reg[32][19]/P0001  & n13736 ;
  assign n21686 = ~n21684 & ~n21685 ;
  assign n21687 = \wishbone_bd_ram_mem2_reg[136][19]/P0001  & n13963 ;
  assign n21688 = \wishbone_bd_ram_mem2_reg[118][19]/P0001  & n13589 ;
  assign n21689 = ~n21687 & ~n21688 ;
  assign n21690 = n21686 & n21689 ;
  assign n21691 = n21683 & n21690 ;
  assign n21692 = n21676 & n21691 ;
  assign n21693 = \wishbone_bd_ram_mem2_reg[164][19]/P0001  & n13236 ;
  assign n21694 = \wishbone_bd_ram_mem2_reg[56][19]/P0001  & n13611 ;
  assign n21695 = ~n21693 & ~n21694 ;
  assign n21696 = \wishbone_bd_ram_mem2_reg[108][19]/P0001  & n13814 ;
  assign n21697 = \wishbone_bd_ram_mem2_reg[217][19]/P0001  & n13767 ;
  assign n21698 = ~n21696 & ~n21697 ;
  assign n21699 = n21695 & n21698 ;
  assign n21700 = \wishbone_bd_ram_mem2_reg[11][19]/P0001  & n13774 ;
  assign n21701 = \wishbone_bd_ram_mem2_reg[18][19]/P0001  & n13532 ;
  assign n21702 = ~n21700 & ~n21701 ;
  assign n21703 = \wishbone_bd_ram_mem2_reg[237][19]/P0001  & n13924 ;
  assign n21704 = \wishbone_bd_ram_mem2_reg[135][19]/P0001  & n13672 ;
  assign n21705 = ~n21703 & ~n21704 ;
  assign n21706 = n21702 & n21705 ;
  assign n21707 = n21699 & n21706 ;
  assign n21708 = \wishbone_bd_ram_mem2_reg[37][19]/P0001  & n13710 ;
  assign n21709 = \wishbone_bd_ram_mem2_reg[55][19]/P0001  & n13618 ;
  assign n21710 = ~n21708 & ~n21709 ;
  assign n21711 = \wishbone_bd_ram_mem2_reg[70][19]/P0001  & n13339 ;
  assign n21712 = \wishbone_bd_ram_mem2_reg[170][19]/P0001  & n14007 ;
  assign n21713 = ~n21711 & ~n21712 ;
  assign n21714 = n21710 & n21713 ;
  assign n21715 = \wishbone_bd_ram_mem2_reg[104][19]/P0001  & n13684 ;
  assign n21716 = \wishbone_bd_ram_mem2_reg[156][19]/P0001  & n13769 ;
  assign n21717 = ~n21715 & ~n21716 ;
  assign n21718 = \wishbone_bd_ram_mem2_reg[61][19]/P0001  & n13544 ;
  assign n21719 = \wishbone_bd_ram_mem2_reg[109][19]/P0001  & n13306 ;
  assign n21720 = ~n21718 & ~n21719 ;
  assign n21721 = n21717 & n21720 ;
  assign n21722 = n21714 & n21721 ;
  assign n21723 = n21707 & n21722 ;
  assign n21724 = n21692 & n21723 ;
  assign n21725 = \wishbone_bd_ram_mem2_reg[79][19]/P0001  & n13779 ;
  assign n21726 = \wishbone_bd_ram_mem2_reg[91][19]/P0001  & n13954 ;
  assign n21727 = ~n21725 & ~n21726 ;
  assign n21728 = \wishbone_bd_ram_mem2_reg[147][19]/P0001  & n13702 ;
  assign n21729 = \wishbone_bd_ram_mem2_reg[113][19]/P0001  & n13882 ;
  assign n21730 = ~n21728 & ~n21729 ;
  assign n21731 = n21727 & n21730 ;
  assign n21732 = \wishbone_bd_ram_mem2_reg[160][19]/P0001  & n13271 ;
  assign n21733 = \wishbone_bd_ram_mem2_reg[148][19]/P0001  & n13868 ;
  assign n21734 = ~n21732 & ~n21733 ;
  assign n21735 = \wishbone_bd_ram_mem2_reg[23][19]/P0001  & n13857 ;
  assign n21736 = \wishbone_bd_ram_mem2_reg[131][19]/P0001  & n13358 ;
  assign n21737 = ~n21735 & ~n21736 ;
  assign n21738 = n21734 & n21737 ;
  assign n21739 = n21731 & n21738 ;
  assign n21740 = \wishbone_bd_ram_mem2_reg[52][19]/P0001  & n13988 ;
  assign n21741 = \wishbone_bd_ram_mem2_reg[190][19]/P0001  & n13365 ;
  assign n21742 = ~n21740 & ~n21741 ;
  assign n21743 = \wishbone_bd_ram_mem2_reg[222][19]/P0001  & n13721 ;
  assign n21744 = \wishbone_bd_ram_mem2_reg[122][19]/P0001  & n13679 ;
  assign n21745 = ~n21743 & ~n21744 ;
  assign n21746 = n21742 & n21745 ;
  assign n21747 = \wishbone_bd_ram_mem2_reg[10][19]/P0001  & n13837 ;
  assign n21748 = \wishbone_bd_ram_mem2_reg[74][19]/P0001  & n13564 ;
  assign n21749 = ~n21747 & ~n21748 ;
  assign n21750 = \wishbone_bd_ram_mem2_reg[230][19]/P0001  & n13994 ;
  assign n21751 = \wishbone_bd_ram_mem2_reg[6][19]/P0001  & n13915 ;
  assign n21752 = ~n21750 & ~n21751 ;
  assign n21753 = n21749 & n21752 ;
  assign n21754 = n21746 & n21753 ;
  assign n21755 = n21739 & n21754 ;
  assign n21756 = \wishbone_bd_ram_mem2_reg[172][19]/P0001  & n13377 ;
  assign n21757 = \wishbone_bd_ram_mem2_reg[212][19]/P0001  & n13634 ;
  assign n21758 = ~n21756 & ~n21757 ;
  assign n21759 = \wishbone_bd_ram_mem2_reg[157][19]/P0001  & n13445 ;
  assign n21760 = \wishbone_bd_ram_mem2_reg[183][19]/P0001  & n13645 ;
  assign n21761 = ~n21759 & ~n21760 ;
  assign n21762 = n21758 & n21761 ;
  assign n21763 = \wishbone_bd_ram_mem2_reg[134][19]/P0001  & n13494 ;
  assign n21764 = \wishbone_bd_ram_mem2_reg[62][19]/P0001  & n13529 ;
  assign n21765 = ~n21763 & ~n21764 ;
  assign n21766 = \wishbone_bd_ram_mem2_reg[102][19]/P0001  & n13534 ;
  assign n21767 = \wishbone_bd_ram_mem2_reg[126][19]/P0001  & n13786 ;
  assign n21768 = ~n21766 & ~n21767 ;
  assign n21769 = n21765 & n21768 ;
  assign n21770 = n21762 & n21769 ;
  assign n21771 = \wishbone_bd_ram_mem2_reg[252][19]/P0001  & n13986 ;
  assign n21772 = \wishbone_bd_ram_mem2_reg[21][19]/P0001  & n13438 ;
  assign n21773 = ~n21771 & ~n21772 ;
  assign n21774 = \wishbone_bd_ram_mem2_reg[225][19]/P0001  & n13719 ;
  assign n21775 = \wishbone_bd_ram_mem2_reg[205][19]/P0001  & n13947 ;
  assign n21776 = ~n21774 & ~n21775 ;
  assign n21777 = n21773 & n21776 ;
  assign n21778 = \wishbone_bd_ram_mem2_reg[206][19]/P0001  & n13414 ;
  assign n21779 = \wishbone_bd_ram_mem2_reg[215][19]/P0001  & n13901 ;
  assign n21780 = ~n21778 & ~n21779 ;
  assign n21781 = \wishbone_bd_ram_mem2_reg[114][19]/P0001  & n13763 ;
  assign n21782 = \wishbone_bd_ram_mem2_reg[119][19]/P0001  & n14033 ;
  assign n21783 = ~n21781 & ~n21782 ;
  assign n21784 = n21780 & n21783 ;
  assign n21785 = n21777 & n21784 ;
  assign n21786 = n21770 & n21785 ;
  assign n21787 = n21755 & n21786 ;
  assign n21788 = n21724 & n21787 ;
  assign n21789 = \wishbone_bd_ram_mem2_reg[151][19]/P0001  & n13697 ;
  assign n21790 = \wishbone_bd_ram_mem2_reg[92][19]/P0001  & n13859 ;
  assign n21791 = ~n21789 & ~n21790 ;
  assign n21792 = \wishbone_bd_ram_mem2_reg[144][19]/P0001  & n13508 ;
  assign n21793 = \wishbone_bd_ram_mem2_reg[5][19]/P0001  & n13243 ;
  assign n21794 = ~n21792 & ~n21793 ;
  assign n21795 = n21791 & n21794 ;
  assign n21796 = \wishbone_bd_ram_mem2_reg[69][19]/P0001  & n13487 ;
  assign n21797 = \wishbone_bd_ram_mem2_reg[87][19]/P0001  & n13691 ;
  assign n21798 = ~n21796 & ~n21797 ;
  assign n21799 = \wishbone_bd_ram_mem2_reg[85][19]/P0001  & n13784 ;
  assign n21800 = \wishbone_bd_ram_mem2_reg[235][19]/P0001  & n13518 ;
  assign n21801 = ~n21799 & ~n21800 ;
  assign n21802 = n21798 & n21801 ;
  assign n21803 = n21795 & n21802 ;
  assign n21804 = \wishbone_bd_ram_mem2_reg[207][19]/P0001  & n13826 ;
  assign n21805 = \wishbone_bd_ram_mem2_reg[132][19]/P0001  & n13927 ;
  assign n21806 = ~n21804 & ~n21805 ;
  assign n21807 = \wishbone_bd_ram_mem2_reg[159][19]/P0001  & n13627 ;
  assign n21808 = \wishbone_bd_ram_mem2_reg[16][19]/P0001  & n13695 ;
  assign n21809 = ~n21807 & ~n21808 ;
  assign n21810 = n21806 & n21809 ;
  assign n21811 = \wishbone_bd_ram_mem2_reg[150][19]/P0001  & n13666 ;
  assign n21812 = \wishbone_bd_ram_mem2_reg[143][19]/P0001  & n13461 ;
  assign n21813 = ~n21811 & ~n21812 ;
  assign n21814 = \wishbone_bd_ram_mem2_reg[3][19]/P0001  & n13354 ;
  assign n21815 = \wishbone_bd_ram_mem2_reg[227][19]/P0001  & n13388 ;
  assign n21816 = ~n21814 & ~n21815 ;
  assign n21817 = n21813 & n21816 ;
  assign n21818 = n21810 & n21817 ;
  assign n21819 = n21803 & n21818 ;
  assign n21820 = \wishbone_bd_ram_mem2_reg[89][19]/P0001  & n13910 ;
  assign n21821 = \wishbone_bd_ram_mem2_reg[72][19]/P0001  & n13582 ;
  assign n21822 = ~n21820 & ~n21821 ;
  assign n21823 = \wishbone_bd_ram_mem2_reg[180][19]/P0001  & n13650 ;
  assign n21824 = \wishbone_bd_ram_mem2_reg[248][19]/P0001  & n13647 ;
  assign n21825 = ~n21823 & ~n21824 ;
  assign n21826 = n21822 & n21825 ;
  assign n21827 = \wishbone_bd_ram_mem2_reg[96][19]/P0001  & n13425 ;
  assign n21828 = \wishbone_bd_ram_mem2_reg[121][19]/P0001  & n13983 ;
  assign n21829 = ~n21827 & ~n21828 ;
  assign n21830 = \wishbone_bd_ram_mem2_reg[191][19]/P0001  & n14012 ;
  assign n21831 = \wishbone_bd_ram_mem2_reg[98][19]/P0001  & n13569 ;
  assign n21832 = ~n21830 & ~n21831 ;
  assign n21833 = n21829 & n21832 ;
  assign n21834 = n21826 & n21833 ;
  assign n21835 = \wishbone_bd_ram_mem2_reg[107][19]/P0001  & n13476 ;
  assign n21836 = \wishbone_bd_ram_mem2_reg[54][19]/P0001  & n13622 ;
  assign n21837 = ~n21835 & ~n21836 ;
  assign n21838 = \wishbone_bd_ram_mem2_reg[64][19]/P0001  & n13904 ;
  assign n21839 = \wishbone_bd_ram_mem2_reg[158][19]/P0001  & n13294 ;
  assign n21840 = ~n21838 & ~n21839 ;
  assign n21841 = n21837 & n21840 ;
  assign n21842 = \wishbone_bd_ram_mem2_reg[161][19]/P0001  & n13505 ;
  assign n21843 = \wishbone_bd_ram_mem2_reg[31][19]/P0001  & n13758 ;
  assign n21844 = ~n21842 & ~n21843 ;
  assign n21845 = \wishbone_bd_ram_mem2_reg[27][19]/P0001  & n13251 ;
  assign n21846 = \wishbone_bd_ram_mem2_reg[210][19]/P0001  & n13443 ;
  assign n21847 = ~n21845 & ~n21846 ;
  assign n21848 = n21844 & n21847 ;
  assign n21849 = n21841 & n21848 ;
  assign n21850 = n21834 & n21849 ;
  assign n21851 = n21819 & n21850 ;
  assign n21852 = \wishbone_bd_ram_mem2_reg[176][19]/P0001  & n13262 ;
  assign n21853 = \wishbone_bd_ram_mem2_reg[208][19]/P0001  & n14010 ;
  assign n21854 = ~n21852 & ~n21853 ;
  assign n21855 = \wishbone_bd_ram_mem2_reg[77][19]/P0001  & n13935 ;
  assign n21856 = \wishbone_bd_ram_mem2_reg[182][19]/P0001  & n13598 ;
  assign n21857 = ~n21855 & ~n21856 ;
  assign n21858 = n21854 & n21857 ;
  assign n21859 = \wishbone_bd_ram_mem2_reg[30][19]/P0001  & n13713 ;
  assign n21860 = \wishbone_bd_ram_mem2_reg[36][19]/P0001  & n13639 ;
  assign n21861 = ~n21859 & ~n21860 ;
  assign n21862 = \wishbone_bd_ram_mem2_reg[130][19]/P0001  & n13427 ;
  assign n21863 = \wishbone_bd_ram_mem2_reg[236][19]/P0001  & n13480 ;
  assign n21864 = ~n21862 & ~n21863 ;
  assign n21865 = n21861 & n21864 ;
  assign n21866 = n21858 & n21865 ;
  assign n21867 = \wishbone_bd_ram_mem2_reg[14][19]/P0001  & n13972 ;
  assign n21868 = \wishbone_bd_ram_mem2_reg[38][19]/P0001  & n13828 ;
  assign n21869 = ~n21867 & ~n21868 ;
  assign n21870 = \wishbone_bd_ram_mem2_reg[138][19]/P0001  & n13398 ;
  assign n21871 = \wishbone_bd_ram_mem2_reg[13][19]/P0001  & n13844 ;
  assign n21872 = ~n21870 & ~n21871 ;
  assign n21873 = n21869 & n21872 ;
  assign n21874 = \wishbone_bd_ram_mem2_reg[49][19]/P0001  & n13929 ;
  assign n21875 = \wishbone_bd_ram_mem2_reg[7][19]/P0001  & n13546 ;
  assign n21876 = ~n21874 & ~n21875 ;
  assign n21877 = \wishbone_bd_ram_mem2_reg[219][19]/P0001  & n13577 ;
  assign n21878 = \wishbone_bd_ram_mem2_reg[245][19]/P0001  & n13877 ;
  assign n21879 = ~n21877 & ~n21878 ;
  assign n21880 = n21876 & n21879 ;
  assign n21881 = n21873 & n21880 ;
  assign n21882 = n21866 & n21881 ;
  assign n21883 = \wishbone_bd_ram_mem2_reg[39][19]/P0001  & n13893 ;
  assign n21884 = \wishbone_bd_ram_mem2_reg[63][19]/P0001  & n13327 ;
  assign n21885 = ~n21883 & ~n21884 ;
  assign n21886 = \wishbone_bd_ram_mem2_reg[129][19]/P0001  & n13629 ;
  assign n21887 = \wishbone_bd_ram_mem2_reg[201][19]/P0001  & n13600 ;
  assign n21888 = ~n21886 & ~n21887 ;
  assign n21889 = n21885 & n21888 ;
  assign n21890 = \wishbone_bd_ram_mem2_reg[124][19]/P0001  & n14024 ;
  assign n21891 = \wishbone_bd_ram_mem2_reg[28][19]/P0001  & n13810 ;
  assign n21892 = ~n21890 & ~n21891 ;
  assign n21893 = \wishbone_bd_ram_mem2_reg[228][19]/P0001  & n13497 ;
  assign n21894 = \wishbone_bd_ram_mem2_reg[100][19]/P0001  & n13401 ;
  assign n21895 = ~n21893 & ~n21894 ;
  assign n21896 = n21892 & n21895 ;
  assign n21897 = n21889 & n21896 ;
  assign n21898 = \wishbone_bd_ram_mem2_reg[80][19]/P0001  & n13516 ;
  assign n21899 = \wishbone_bd_ram_mem2_reg[169][19]/P0001  & n13541 ;
  assign n21900 = ~n21898 & ~n21899 ;
  assign n21901 = \wishbone_bd_ram_mem2_reg[229][19]/P0001  & n13552 ;
  assign n21902 = \wishbone_bd_ram_mem2_reg[25][19]/P0001  & n13742 ;
  assign n21903 = ~n21901 & ~n21902 ;
  assign n21904 = n21900 & n21903 ;
  assign n21905 = \wishbone_bd_ram_mem2_reg[20][19]/P0001  & n13839 ;
  assign n21906 = \wishbone_bd_ram_mem2_reg[163][19]/P0001  & n13255 ;
  assign n21907 = ~n21905 & ~n21906 ;
  assign n21908 = \wishbone_bd_ram_mem2_reg[242][19]/P0001  & n13383 ;
  assign n21909 = \wishbone_bd_ram_mem2_reg[60][19]/P0001  & n13790 ;
  assign n21910 = ~n21908 & ~n21909 ;
  assign n21911 = n21907 & n21910 ;
  assign n21912 = n21904 & n21911 ;
  assign n21913 = n21897 & n21912 ;
  assign n21914 = n21882 & n21913 ;
  assign n21915 = n21851 & n21914 ;
  assign n21916 = n21788 & n21915 ;
  assign n21917 = \wishbone_bd_ram_mem2_reg[224][19]/P0001  & n13433 ;
  assign n21918 = \wishbone_bd_ram_mem2_reg[174][19]/P0001  & n13899 ;
  assign n21919 = ~n21917 & ~n21918 ;
  assign n21920 = \wishbone_bd_ram_mem2_reg[202][19]/P0001  & n13268 ;
  assign n21921 = \wishbone_bd_ram_mem2_reg[22][19]/P0001  & n13744 ;
  assign n21922 = ~n21920 & ~n21921 ;
  assign n21923 = n21919 & n21922 ;
  assign n21924 = \wishbone_bd_ram_mem2_reg[189][19]/P0001  & n14001 ;
  assign n21925 = \wishbone_bd_ram_mem2_reg[171][19]/P0001  & n13422 ;
  assign n21926 = ~n21924 & ~n21925 ;
  assign n21927 = \wishbone_bd_ram_mem2_reg[188][19]/P0001  & n13407 ;
  assign n21928 = \wishbone_bd_ram_mem2_reg[45][19]/P0001  & n13420 ;
  assign n21929 = ~n21927 & ~n21928 ;
  assign n21930 = n21926 & n21929 ;
  assign n21931 = n21923 & n21930 ;
  assign n21932 = \wishbone_bd_ram_mem2_reg[149][19]/P0001  & n13469 ;
  assign n21933 = \wishbone_bd_ram_mem2_reg[200][19]/P0001  & n13922 ;
  assign n21934 = ~n21932 & ~n21933 ;
  assign n21935 = \wishbone_bd_ram_mem2_reg[50][19]/P0001  & n13686 ;
  assign n21936 = \wishbone_bd_ram_mem2_reg[152][19]/P0001  & n13912 ;
  assign n21937 = ~n21935 & ~n21936 ;
  assign n21938 = n21934 & n21937 ;
  assign n21939 = \wishbone_bd_ram_mem2_reg[120][19]/P0001  & n13550 ;
  assign n21940 = \wishbone_bd_ram_mem2_reg[185][19]/P0001  & n13372 ;
  assign n21941 = ~n21939 & ~n21940 ;
  assign n21942 = \wishbone_bd_ram_mem2_reg[101][19]/P0001  & n13772 ;
  assign n21943 = \wishbone_bd_ram_mem2_reg[241][19]/P0001  & n13854 ;
  assign n21944 = ~n21942 & ~n21943 ;
  assign n21945 = n21941 & n21944 ;
  assign n21946 = n21938 & n21945 ;
  assign n21947 = n21931 & n21946 ;
  assign n21948 = \wishbone_bd_ram_mem2_reg[115][19]/P0001  & n13747 ;
  assign n21949 = \wishbone_bd_ram_mem2_reg[192][19]/P0001  & n13390 ;
  assign n21950 = ~n21948 & ~n21949 ;
  assign n21951 = \wishbone_bd_ram_mem2_reg[197][19]/P0001  & n13594 ;
  assign n21952 = \wishbone_bd_ram_mem2_reg[12][19]/P0001  & n13733 ;
  assign n21953 = ~n21951 & ~n21952 ;
  assign n21954 = n21950 & n21953 ;
  assign n21955 = \wishbone_bd_ram_mem2_reg[46][19]/P0001  & n13298 ;
  assign n21956 = \wishbone_bd_ram_mem2_reg[19][19]/P0001  & n13886 ;
  assign n21957 = ~n21955 & ~n21956 ;
  assign n21958 = \wishbone_bd_ram_mem2_reg[165][19]/P0001  & n14028 ;
  assign n21959 = \wishbone_bd_ram_mem2_reg[218][19]/P0001  & n13792 ;
  assign n21960 = ~n21958 & ~n21959 ;
  assign n21961 = n21957 & n21960 ;
  assign n21962 = n21954 & n21961 ;
  assign n21963 = \wishbone_bd_ram_mem2_reg[146][19]/P0001  & n13958 ;
  assign n21964 = \wishbone_bd_ram_mem2_reg[179][19]/P0001  & n14035 ;
  assign n21965 = ~n21963 & ~n21964 ;
  assign n21966 = \wishbone_bd_ram_mem2_reg[162][19]/P0001  & n13726 ;
  assign n21967 = \wishbone_bd_ram_mem2_reg[105][19]/P0001  & n13503 ;
  assign n21968 = ~n21966 & ~n21967 ;
  assign n21969 = n21965 & n21968 ;
  assign n21970 = \wishbone_bd_ram_mem2_reg[112][19]/P0001  & n13482 ;
  assign n21971 = \wishbone_bd_ram_mem2_reg[253][19]/P0001  & n13708 ;
  assign n21972 = ~n21970 & ~n21971 ;
  assign n21973 = \wishbone_bd_ram_mem2_reg[226][19]/P0001  & n13668 ;
  assign n21974 = \wishbone_bd_ram_mem2_reg[195][19]/P0001  & n13700 ;
  assign n21975 = ~n21973 & ~n21974 ;
  assign n21976 = n21972 & n21975 ;
  assign n21977 = n21969 & n21976 ;
  assign n21978 = n21962 & n21977 ;
  assign n21979 = n21947 & n21978 ;
  assign n21980 = \wishbone_bd_ram_mem2_reg[83][19]/P0001  & n13454 ;
  assign n21981 = \wishbone_bd_ram_mem2_reg[214][19]/P0001  & n13938 ;
  assign n21982 = ~n21980 & ~n21981 ;
  assign n21983 = \wishbone_bd_ram_mem2_reg[220][19]/P0001  & n13965 ;
  assign n21984 = \wishbone_bd_ram_mem2_reg[58][19]/P0001  & n13949 ;
  assign n21985 = ~n21983 & ~n21984 ;
  assign n21986 = n21982 & n21985 ;
  assign n21987 = \wishbone_bd_ram_mem2_reg[51][19]/P0001  & n13880 ;
  assign n21988 = \wishbone_bd_ram_mem2_reg[247][19]/P0001  & n13571 ;
  assign n21989 = ~n21987 & ~n21988 ;
  assign n21990 = \wishbone_bd_ram_mem2_reg[186][19]/P0001  & n13616 ;
  assign n21991 = \wishbone_bd_ram_mem2_reg[233][19]/P0001  & n13332 ;
  assign n21992 = ~n21990 & ~n21991 ;
  assign n21993 = n21989 & n21992 ;
  assign n21994 = n21986 & n21993 ;
  assign n21995 = \wishbone_bd_ram_mem2_reg[204][19]/P0001  & n13821 ;
  assign n21996 = \wishbone_bd_ram_mem2_reg[213][19]/P0001  & n13870 ;
  assign n21997 = ~n21995 & ~n21996 ;
  assign n21998 = \wishbone_bd_ram_mem2_reg[90][19]/P0001  & n13906 ;
  assign n21999 = \wishbone_bd_ram_mem2_reg[68][19]/P0001  & n13379 ;
  assign n22000 = ~n21998 & ~n21999 ;
  assign n22001 = n21997 & n22000 ;
  assign n22002 = \wishbone_bd_ram_mem2_reg[145][19]/P0001  & n13715 ;
  assign n22003 = \wishbone_bd_ram_mem2_reg[35][19]/P0001  & n13523 ;
  assign n22004 = ~n22002 & ~n22003 ;
  assign n22005 = \wishbone_bd_ram_mem2_reg[94][19]/P0001  & n13833 ;
  assign n22006 = \wishbone_bd_ram_mem2_reg[239][19]/P0001  & n13349 ;
  assign n22007 = ~n22005 & ~n22006 ;
  assign n22008 = n22004 & n22007 ;
  assign n22009 = n22001 & n22008 ;
  assign n22010 = n21994 & n22009 ;
  assign n22011 = \wishbone_bd_ram_mem2_reg[4][19]/P0001  & n13527 ;
  assign n22012 = \wishbone_bd_ram_mem2_reg[2][19]/P0001  & n13975 ;
  assign n22013 = ~n22011 & ~n22012 ;
  assign n22014 = \wishbone_bd_ram_mem2_reg[246][19]/P0001  & n13981 ;
  assign n22015 = \wishbone_bd_ram_mem2_reg[133][19]/P0001  & n13492 ;
  assign n22016 = ~n22014 & ~n22015 ;
  assign n22017 = n22013 & n22016 ;
  assign n22018 = \wishbone_bd_ram_mem2_reg[84][19]/P0001  & n13385 ;
  assign n22019 = \wishbone_bd_ram_mem2_reg[24][19]/P0001  & n13970 ;
  assign n22020 = ~n22018 & ~n22019 ;
  assign n22021 = \wishbone_bd_ram_mem2_reg[97][19]/P0001  & n13724 ;
  assign n22022 = \wishbone_bd_ram_mem2_reg[1][19]/P0001  & n13888 ;
  assign n22023 = ~n22021 & ~n22022 ;
  assign n22024 = n22020 & n22023 ;
  assign n22025 = n22017 & n22024 ;
  assign n22026 = \wishbone_bd_ram_mem2_reg[123][19]/P0001  & n13749 ;
  assign n22027 = \wishbone_bd_ram_mem2_reg[88][19]/P0001  & n13347 ;
  assign n22028 = ~n22026 & ~n22027 ;
  assign n22029 = \wishbone_bd_ram_mem2_reg[251][19]/P0001  & n14019 ;
  assign n22030 = \wishbone_bd_ram_mem2_reg[81][19]/P0001  & n13409 ;
  assign n22031 = ~n22029 & ~n22030 ;
  assign n22032 = n22028 & n22031 ;
  assign n22033 = \wishbone_bd_ram_mem2_reg[216][19]/P0001  & n14005 ;
  assign n22034 = \wishbone_bd_ram_mem2_reg[177][19]/P0001  & n13863 ;
  assign n22035 = ~n22033 & ~n22034 ;
  assign n22036 = \wishbone_bd_ram_mem2_reg[175][19]/P0001  & n13674 ;
  assign n22037 = \wishbone_bd_ram_mem2_reg[243][19]/P0001  & n13575 ;
  assign n22038 = ~n22036 & ~n22037 ;
  assign n22039 = n22035 & n22038 ;
  assign n22040 = n22032 & n22039 ;
  assign n22041 = n22025 & n22040 ;
  assign n22042 = n22010 & n22041 ;
  assign n22043 = n21979 & n22042 ;
  assign n22044 = \wishbone_bd_ram_mem2_reg[255][19]/P0001  & n13952 ;
  assign n22045 = \wishbone_bd_ram_mem2_reg[155][19]/P0001  & n13738 ;
  assign n22046 = ~n22044 & ~n22045 ;
  assign n22047 = \wishbone_bd_ram_mem2_reg[139][19]/P0001  & n13566 ;
  assign n22048 = \wishbone_bd_ram_mem2_reg[250][19]/P0001  & n13677 ;
  assign n22049 = ~n22047 & ~n22048 ;
  assign n22050 = n22046 & n22049 ;
  assign n22051 = \wishbone_bd_ram_mem2_reg[57][19]/P0001  & n13731 ;
  assign n22052 = \wishbone_bd_ram_mem2_reg[232][19]/P0001  & n13510 ;
  assign n22053 = ~n22051 & ~n22052 ;
  assign n22054 = \wishbone_bd_ram_mem2_reg[34][19]/P0001  & n13450 ;
  assign n22055 = \wishbone_bd_ram_mem2_reg[82][19]/P0001  & n13374 ;
  assign n22056 = ~n22054 & ~n22055 ;
  assign n22057 = n22053 & n22056 ;
  assign n22058 = n22050 & n22057 ;
  assign n22059 = \wishbone_bd_ram_mem2_reg[154][19]/P0001  & n13403 ;
  assign n22060 = \wishbone_bd_ram_mem2_reg[76][19]/P0001  & n13831 ;
  assign n22061 = ~n22059 & ~n22060 ;
  assign n22062 = \wishbone_bd_ram_mem2_reg[238][19]/P0001  & n13819 ;
  assign n22063 = \wishbone_bd_ram_mem2_reg[8][19]/P0001  & n13459 ;
  assign n22064 = ~n22062 & ~n22063 ;
  assign n22065 = n22061 & n22064 ;
  assign n22066 = \wishbone_bd_ram_mem2_reg[194][19]/P0001  & n13624 ;
  assign n22067 = \wishbone_bd_ram_mem2_reg[44][19]/P0001  & n13291 ;
  assign n22068 = ~n22066 & ~n22067 ;
  assign n22069 = \wishbone_bd_ram_mem2_reg[168][19]/P0001  & n13795 ;
  assign n22070 = \wishbone_bd_ram_mem2_reg[209][19]/P0001  & n13689 ;
  assign n22071 = ~n22069 & ~n22070 ;
  assign n22072 = n22068 & n22071 ;
  assign n22073 = n22065 & n22072 ;
  assign n22074 = n22058 & n22073 ;
  assign n22075 = \wishbone_bd_ram_mem2_reg[65][19]/P0001  & n13842 ;
  assign n22076 = \wishbone_bd_ram_mem2_reg[234][19]/P0001  & n13781 ;
  assign n22077 = ~n22075 & ~n22076 ;
  assign n22078 = \wishbone_bd_ram_mem2_reg[166][19]/P0001  & n13999 ;
  assign n22079 = \wishbone_bd_ram_mem2_reg[78][19]/P0001  & n13277 ;
  assign n22080 = ~n22078 & ~n22079 ;
  assign n22081 = n22077 & n22080 ;
  assign n22082 = \wishbone_bd_ram_mem2_reg[86][19]/P0001  & n13485 ;
  assign n22083 = \wishbone_bd_ram_mem2_reg[137][19]/P0001  & n13808 ;
  assign n22084 = ~n22082 & ~n22083 ;
  assign n22085 = \wishbone_bd_ram_mem2_reg[66][19]/P0001  & n13603 ;
  assign n22086 = \wishbone_bd_ram_mem2_reg[221][19]/P0001  & n13641 ;
  assign n22087 = ~n22085 & ~n22086 ;
  assign n22088 = n22084 & n22087 ;
  assign n22089 = n22081 & n22088 ;
  assign n22090 = \wishbone_bd_ram_mem2_reg[95][19]/P0001  & n13317 ;
  assign n22091 = \wishbone_bd_ram_mem2_reg[99][19]/P0001  & n13996 ;
  assign n22092 = ~n22090 & ~n22091 ;
  assign n22093 = \wishbone_bd_ram_mem2_reg[142][19]/P0001  & n13448 ;
  assign n22094 = \wishbone_bd_ram_mem2_reg[153][19]/P0001  & n13309 ;
  assign n22095 = ~n22093 & ~n22094 ;
  assign n22096 = n22092 & n22095 ;
  assign n22097 = \wishbone_bd_ram_mem2_reg[127][19]/P0001  & n13803 ;
  assign n22098 = \wishbone_bd_ram_mem2_reg[244][19]/P0001  & n13474 ;
  assign n22099 = ~n22097 & ~n22098 ;
  assign n22100 = \wishbone_bd_ram_mem2_reg[184][19]/P0001  & n13960 ;
  assign n22101 = \wishbone_bd_ram_mem2_reg[117][19]/P0001  & n13557 ;
  assign n22102 = ~n22100 & ~n22101 ;
  assign n22103 = n22099 & n22102 ;
  assign n22104 = n22096 & n22103 ;
  assign n22105 = n22089 & n22104 ;
  assign n22106 = n22074 & n22105 ;
  assign n22107 = \wishbone_bd_ram_mem2_reg[43][19]/P0001  & n13761 ;
  assign n22108 = \wishbone_bd_ram_mem2_reg[231][19]/P0001  & n13363 ;
  assign n22109 = ~n22107 & ~n22108 ;
  assign n22110 = \wishbone_bd_ram_mem2_reg[40][19]/P0001  & n13661 ;
  assign n22111 = \wishbone_bd_ram_mem2_reg[93][19]/P0001  & n13891 ;
  assign n22112 = ~n22110 & ~n22111 ;
  assign n22113 = n22109 & n22112 ;
  assign n22114 = \wishbone_bd_ram_mem2_reg[128][19]/P0001  & n13652 ;
  assign n22115 = \wishbone_bd_ram_mem2_reg[254][19]/P0001  & n13283 ;
  assign n22116 = ~n22114 & ~n22115 ;
  assign n22117 = \wishbone_bd_ram_mem2_reg[196][19]/P0001  & n13977 ;
  assign n22118 = \wishbone_bd_ram_mem2_reg[17][19]/P0001  & n13324 ;
  assign n22119 = ~n22117 & ~n22118 ;
  assign n22120 = n22116 & n22119 ;
  assign n22121 = n22113 & n22120 ;
  assign n22122 = \wishbone_bd_ram_mem2_reg[173][19]/P0001  & n13360 ;
  assign n22123 = \wishbone_bd_ram_mem2_reg[240][19]/P0001  & n13352 ;
  assign n22124 = ~n22122 & ~n22123 ;
  assign n22125 = \wishbone_bd_ram_mem2_reg[211][19]/P0001  & n13805 ;
  assign n22126 = \wishbone_bd_ram_mem2_reg[116][19]/P0001  & n13865 ;
  assign n22127 = ~n22125 & ~n22126 ;
  assign n22128 = n22124 & n22127 ;
  assign n22129 = \wishbone_bd_ram_mem2_reg[48][19]/P0001  & n13917 ;
  assign n22130 = \wishbone_bd_ram_mem2_reg[141][19]/P0001  & n13852 ;
  assign n22131 = ~n22129 & ~n22130 ;
  assign n22132 = \wishbone_bd_ram_mem2_reg[167][19]/P0001  & n13940 ;
  assign n22133 = \wishbone_bd_ram_mem2_reg[125][19]/P0001  & n13396 ;
  assign n22134 = ~n22132 & ~n22133 ;
  assign n22135 = n22131 & n22134 ;
  assign n22136 = n22128 & n22135 ;
  assign n22137 = n22121 & n22136 ;
  assign n22138 = \wishbone_bd_ram_mem2_reg[199][19]/P0001  & n13499 ;
  assign n22139 = \wishbone_bd_ram_mem2_reg[71][19]/P0001  & n13636 ;
  assign n22140 = ~n22138 & ~n22139 ;
  assign n22141 = \wishbone_bd_ram_mem2_reg[47][19]/P0001  & n13436 ;
  assign n22142 = \wishbone_bd_ram_mem2_reg[29][19]/P0001  & n13412 ;
  assign n22143 = ~n22141 & ~n22142 ;
  assign n22144 = n22140 & n22143 ;
  assign n22145 = \wishbone_bd_ram_mem2_reg[41][19]/P0001  & n14017 ;
  assign n22146 = \wishbone_bd_ram_mem2_reg[33][19]/P0001  & n13933 ;
  assign n22147 = ~n22145 & ~n22146 ;
  assign n22148 = \wishbone_bd_ram_mem2_reg[198][19]/P0001  & n13592 ;
  assign n22149 = \wishbone_bd_ram_mem2_reg[0][19]/P0001  & n13539 ;
  assign n22150 = ~n22148 & ~n22149 ;
  assign n22151 = n22147 & n22150 ;
  assign n22152 = n22144 & n22151 ;
  assign n22153 = \wishbone_bd_ram_mem2_reg[178][19]/P0001  & n13301 ;
  assign n22154 = \wishbone_bd_ram_mem2_reg[75][19]/P0001  & n13605 ;
  assign n22155 = ~n22153 & ~n22154 ;
  assign n22156 = \wishbone_bd_ram_mem2_reg[53][19]/P0001  & n13875 ;
  assign n22157 = \wishbone_bd_ram_mem2_reg[111][19]/P0001  & n13471 ;
  assign n22158 = ~n22156 & ~n22157 ;
  assign n22159 = n22155 & n22158 ;
  assign n22160 = \wishbone_bd_ram_mem2_reg[110][19]/P0001  & n14030 ;
  assign n22161 = \wishbone_bd_ram_mem2_reg[59][19]/P0001  & n13613 ;
  assign n22162 = ~n22160 & ~n22161 ;
  assign n22163 = \wishbone_bd_ram_mem2_reg[140][19]/P0001  & n13287 ;
  assign n22164 = \wishbone_bd_ram_mem2_reg[9][19]/P0001  & n13580 ;
  assign n22165 = ~n22163 & ~n22164 ;
  assign n22166 = n22162 & n22165 ;
  assign n22167 = n22159 & n22166 ;
  assign n22168 = n22152 & n22167 ;
  assign n22169 = n22137 & n22168 ;
  assign n22170 = n22106 & n22169 ;
  assign n22171 = n22043 & n22170 ;
  assign n22172 = n21916 & n22171 ;
  assign n22173 = n14047 & ~n22172 ;
  assign n22174 = ~n21661 & ~n22173 ;
  assign n22175 = \wishbone_LatchedTxLength_reg[4]/NET0131  & ~n14046 ;
  assign n22176 = ~n17359 & ~n22175 ;
  assign n22177 = \wishbone_LatchedTxLength_reg[5]/NET0131  & ~n14046 ;
  assign n22178 = \wishbone_bd_ram_mem2_reg[68][21]/P0001  & n13379 ;
  assign n22179 = \wishbone_bd_ram_mem2_reg[175][21]/P0001  & n13674 ;
  assign n22180 = ~n22178 & ~n22179 ;
  assign n22181 = \wishbone_bd_ram_mem2_reg[37][21]/P0001  & n13710 ;
  assign n22182 = \wishbone_bd_ram_mem2_reg[169][21]/P0001  & n13541 ;
  assign n22183 = ~n22181 & ~n22182 ;
  assign n22184 = n22180 & n22183 ;
  assign n22185 = \wishbone_bd_ram_mem2_reg[101][21]/P0001  & n13772 ;
  assign n22186 = \wishbone_bd_ram_mem2_reg[99][21]/P0001  & n13996 ;
  assign n22187 = ~n22185 & ~n22186 ;
  assign n22188 = \wishbone_bd_ram_mem2_reg[119][21]/P0001  & n14033 ;
  assign n22189 = \wishbone_bd_ram_mem2_reg[145][21]/P0001  & n13715 ;
  assign n22190 = ~n22188 & ~n22189 ;
  assign n22191 = n22187 & n22190 ;
  assign n22192 = n22184 & n22191 ;
  assign n22193 = \wishbone_bd_ram_mem2_reg[254][21]/P0001  & n13283 ;
  assign n22194 = \wishbone_bd_ram_mem2_reg[183][21]/P0001  & n13645 ;
  assign n22195 = ~n22193 & ~n22194 ;
  assign n22196 = \wishbone_bd_ram_mem2_reg[38][21]/P0001  & n13828 ;
  assign n22197 = \wishbone_bd_ram_mem2_reg[232][21]/P0001  & n13510 ;
  assign n22198 = ~n22196 & ~n22197 ;
  assign n22199 = n22195 & n22198 ;
  assign n22200 = \wishbone_bd_ram_mem2_reg[109][21]/P0001  & n13306 ;
  assign n22201 = \wishbone_bd_ram_mem2_reg[122][21]/P0001  & n13679 ;
  assign n22202 = ~n22200 & ~n22201 ;
  assign n22203 = \wishbone_bd_ram_mem2_reg[28][21]/P0001  & n13810 ;
  assign n22204 = \wishbone_bd_ram_mem2_reg[156][21]/P0001  & n13769 ;
  assign n22205 = ~n22203 & ~n22204 ;
  assign n22206 = n22202 & n22205 ;
  assign n22207 = n22199 & n22206 ;
  assign n22208 = n22192 & n22207 ;
  assign n22209 = \wishbone_bd_ram_mem2_reg[64][21]/P0001  & n13904 ;
  assign n22210 = \wishbone_bd_ram_mem2_reg[157][21]/P0001  & n13445 ;
  assign n22211 = ~n22209 & ~n22210 ;
  assign n22212 = \wishbone_bd_ram_mem2_reg[144][21]/P0001  & n13508 ;
  assign n22213 = \wishbone_bd_ram_mem2_reg[155][21]/P0001  & n13738 ;
  assign n22214 = ~n22212 & ~n22213 ;
  assign n22215 = n22211 & n22214 ;
  assign n22216 = \wishbone_bd_ram_mem2_reg[23][21]/P0001  & n13857 ;
  assign n22217 = \wishbone_bd_ram_mem2_reg[143][21]/P0001  & n13461 ;
  assign n22218 = ~n22216 & ~n22217 ;
  assign n22219 = \wishbone_bd_ram_mem2_reg[48][21]/P0001  & n13917 ;
  assign n22220 = \wishbone_bd_ram_mem2_reg[9][21]/P0001  & n13580 ;
  assign n22221 = ~n22219 & ~n22220 ;
  assign n22222 = n22218 & n22221 ;
  assign n22223 = n22215 & n22222 ;
  assign n22224 = \wishbone_bd_ram_mem2_reg[58][21]/P0001  & n13949 ;
  assign n22225 = \wishbone_bd_ram_mem2_reg[198][21]/P0001  & n13592 ;
  assign n22226 = ~n22224 & ~n22225 ;
  assign n22227 = \wishbone_bd_ram_mem2_reg[246][21]/P0001  & n13981 ;
  assign n22228 = \wishbone_bd_ram_mem2_reg[95][21]/P0001  & n13317 ;
  assign n22229 = ~n22227 & ~n22228 ;
  assign n22230 = n22226 & n22229 ;
  assign n22231 = \wishbone_bd_ram_mem2_reg[24][21]/P0001  & n13970 ;
  assign n22232 = \wishbone_bd_ram_mem2_reg[209][21]/P0001  & n13689 ;
  assign n22233 = ~n22231 & ~n22232 ;
  assign n22234 = \wishbone_bd_ram_mem2_reg[149][21]/P0001  & n13469 ;
  assign n22235 = \wishbone_bd_ram_mem2_reg[207][21]/P0001  & n13826 ;
  assign n22236 = ~n22234 & ~n22235 ;
  assign n22237 = n22233 & n22236 ;
  assign n22238 = n22230 & n22237 ;
  assign n22239 = n22223 & n22238 ;
  assign n22240 = n22208 & n22239 ;
  assign n22241 = \wishbone_bd_ram_mem2_reg[114][21]/P0001  & n13763 ;
  assign n22242 = \wishbone_bd_ram_mem2_reg[129][21]/P0001  & n13629 ;
  assign n22243 = ~n22241 & ~n22242 ;
  assign n22244 = \wishbone_bd_ram_mem2_reg[70][21]/P0001  & n13339 ;
  assign n22245 = \wishbone_bd_ram_mem2_reg[166][21]/P0001  & n13999 ;
  assign n22246 = ~n22244 & ~n22245 ;
  assign n22247 = n22243 & n22246 ;
  assign n22248 = \wishbone_bd_ram_mem2_reg[65][21]/P0001  & n13842 ;
  assign n22249 = \wishbone_bd_ram_mem2_reg[77][21]/P0001  & n13935 ;
  assign n22250 = ~n22248 & ~n22249 ;
  assign n22251 = \wishbone_bd_ram_mem2_reg[195][21]/P0001  & n13700 ;
  assign n22252 = \wishbone_bd_ram_mem2_reg[192][21]/P0001  & n13390 ;
  assign n22253 = ~n22251 & ~n22252 ;
  assign n22254 = n22250 & n22253 ;
  assign n22255 = n22247 & n22254 ;
  assign n22256 = \wishbone_bd_ram_mem2_reg[80][21]/P0001  & n13516 ;
  assign n22257 = \wishbone_bd_ram_mem2_reg[210][21]/P0001  & n13443 ;
  assign n22258 = ~n22256 & ~n22257 ;
  assign n22259 = \wishbone_bd_ram_mem2_reg[208][21]/P0001  & n14010 ;
  assign n22260 = \wishbone_bd_ram_mem2_reg[184][21]/P0001  & n13960 ;
  assign n22261 = ~n22259 & ~n22260 ;
  assign n22262 = n22258 & n22261 ;
  assign n22263 = \wishbone_bd_ram_mem2_reg[14][21]/P0001  & n13972 ;
  assign n22264 = \wishbone_bd_ram_mem2_reg[222][21]/P0001  & n13721 ;
  assign n22265 = ~n22263 & ~n22264 ;
  assign n22266 = \wishbone_bd_ram_mem2_reg[40][21]/P0001  & n13661 ;
  assign n22267 = \wishbone_bd_ram_mem2_reg[181][21]/P0001  & n13587 ;
  assign n22268 = ~n22266 & ~n22267 ;
  assign n22269 = n22265 & n22268 ;
  assign n22270 = n22262 & n22269 ;
  assign n22271 = n22255 & n22270 ;
  assign n22272 = \wishbone_bd_ram_mem2_reg[63][21]/P0001  & n13327 ;
  assign n22273 = \wishbone_bd_ram_mem2_reg[125][21]/P0001  & n13396 ;
  assign n22274 = ~n22272 & ~n22273 ;
  assign n22275 = \wishbone_bd_ram_mem2_reg[104][21]/P0001  & n13684 ;
  assign n22276 = \wishbone_bd_ram_mem2_reg[85][21]/P0001  & n13784 ;
  assign n22277 = ~n22275 & ~n22276 ;
  assign n22278 = n22274 & n22277 ;
  assign n22279 = \wishbone_bd_ram_mem2_reg[81][21]/P0001  & n13409 ;
  assign n22280 = \wishbone_bd_ram_mem2_reg[78][21]/P0001  & n13277 ;
  assign n22281 = ~n22279 & ~n22280 ;
  assign n22282 = \wishbone_bd_ram_mem2_reg[50][21]/P0001  & n13686 ;
  assign n22283 = \wishbone_bd_ram_mem2_reg[127][21]/P0001  & n13803 ;
  assign n22284 = ~n22282 & ~n22283 ;
  assign n22285 = n22281 & n22284 ;
  assign n22286 = n22278 & n22285 ;
  assign n22287 = \wishbone_bd_ram_mem2_reg[196][21]/P0001  & n13977 ;
  assign n22288 = \wishbone_bd_ram_mem2_reg[27][21]/P0001  & n13251 ;
  assign n22289 = ~n22287 & ~n22288 ;
  assign n22290 = \wishbone_bd_ram_mem2_reg[22][21]/P0001  & n13744 ;
  assign n22291 = \wishbone_bd_ram_mem2_reg[1][21]/P0001  & n13888 ;
  assign n22292 = ~n22290 & ~n22291 ;
  assign n22293 = n22289 & n22292 ;
  assign n22294 = \wishbone_bd_ram_mem2_reg[162][21]/P0001  & n13726 ;
  assign n22295 = \wishbone_bd_ram_mem2_reg[7][21]/P0001  & n13546 ;
  assign n22296 = ~n22294 & ~n22295 ;
  assign n22297 = \wishbone_bd_ram_mem2_reg[151][21]/P0001  & n13697 ;
  assign n22298 = \wishbone_bd_ram_mem2_reg[62][21]/P0001  & n13529 ;
  assign n22299 = ~n22297 & ~n22298 ;
  assign n22300 = n22296 & n22299 ;
  assign n22301 = n22293 & n22300 ;
  assign n22302 = n22286 & n22301 ;
  assign n22303 = n22271 & n22302 ;
  assign n22304 = n22240 & n22303 ;
  assign n22305 = \wishbone_bd_ram_mem2_reg[148][21]/P0001  & n13868 ;
  assign n22306 = \wishbone_bd_ram_mem2_reg[193][21]/P0001  & n14022 ;
  assign n22307 = ~n22305 & ~n22306 ;
  assign n22308 = \wishbone_bd_ram_mem2_reg[220][21]/P0001  & n13965 ;
  assign n22309 = \wishbone_bd_ram_mem2_reg[230][21]/P0001  & n13994 ;
  assign n22310 = ~n22308 & ~n22309 ;
  assign n22311 = n22307 & n22310 ;
  assign n22312 = \wishbone_bd_ram_mem2_reg[242][21]/P0001  & n13383 ;
  assign n22313 = \wishbone_bd_ram_mem2_reg[111][21]/P0001  & n13471 ;
  assign n22314 = ~n22312 & ~n22313 ;
  assign n22315 = \wishbone_bd_ram_mem2_reg[2][21]/P0001  & n13975 ;
  assign n22316 = \wishbone_bd_ram_mem2_reg[179][21]/P0001  & n14035 ;
  assign n22317 = ~n22315 & ~n22316 ;
  assign n22318 = n22314 & n22317 ;
  assign n22319 = n22311 & n22318 ;
  assign n22320 = \wishbone_bd_ram_mem2_reg[168][21]/P0001  & n13795 ;
  assign n22321 = \wishbone_bd_ram_mem2_reg[115][21]/P0001  & n13747 ;
  assign n22322 = ~n22320 & ~n22321 ;
  assign n22323 = \wishbone_bd_ram_mem2_reg[82][21]/P0001  & n13374 ;
  assign n22324 = \wishbone_bd_ram_mem2_reg[177][21]/P0001  & n13863 ;
  assign n22325 = ~n22323 & ~n22324 ;
  assign n22326 = n22322 & n22325 ;
  assign n22327 = \wishbone_bd_ram_mem2_reg[87][21]/P0001  & n13691 ;
  assign n22328 = \wishbone_bd_ram_mem2_reg[141][21]/P0001  & n13852 ;
  assign n22329 = ~n22327 & ~n22328 ;
  assign n22330 = \wishbone_bd_ram_mem2_reg[8][21]/P0001  & n13459 ;
  assign n22331 = \wishbone_bd_ram_mem2_reg[186][21]/P0001  & n13616 ;
  assign n22332 = ~n22330 & ~n22331 ;
  assign n22333 = n22329 & n22332 ;
  assign n22334 = n22326 & n22333 ;
  assign n22335 = n22319 & n22334 ;
  assign n22336 = \wishbone_bd_ram_mem2_reg[128][21]/P0001  & n13652 ;
  assign n22337 = \wishbone_bd_ram_mem2_reg[255][21]/P0001  & n13952 ;
  assign n22338 = ~n22336 & ~n22337 ;
  assign n22339 = \wishbone_bd_ram_mem2_reg[90][21]/P0001  & n13906 ;
  assign n22340 = \wishbone_bd_ram_mem2_reg[178][21]/P0001  & n13301 ;
  assign n22341 = ~n22339 & ~n22340 ;
  assign n22342 = n22338 & n22341 ;
  assign n22343 = \wishbone_bd_ram_mem2_reg[44][21]/P0001  & n13291 ;
  assign n22344 = \wishbone_bd_ram_mem2_reg[30][21]/P0001  & n13713 ;
  assign n22345 = ~n22343 & ~n22344 ;
  assign n22346 = \wishbone_bd_ram_mem2_reg[171][21]/P0001  & n13422 ;
  assign n22347 = \wishbone_bd_ram_mem2_reg[17][21]/P0001  & n13324 ;
  assign n22348 = ~n22346 & ~n22347 ;
  assign n22349 = n22345 & n22348 ;
  assign n22350 = n22342 & n22349 ;
  assign n22351 = \wishbone_bd_ram_mem2_reg[212][21]/P0001  & n13634 ;
  assign n22352 = \wishbone_bd_ram_mem2_reg[165][21]/P0001  & n14028 ;
  assign n22353 = ~n22351 & ~n22352 ;
  assign n22354 = \wishbone_bd_ram_mem2_reg[102][21]/P0001  & n13534 ;
  assign n22355 = \wishbone_bd_ram_mem2_reg[213][21]/P0001  & n13870 ;
  assign n22356 = ~n22354 & ~n22355 ;
  assign n22357 = n22353 & n22356 ;
  assign n22358 = \wishbone_bd_ram_mem2_reg[60][21]/P0001  & n13790 ;
  assign n22359 = \wishbone_bd_ram_mem2_reg[238][21]/P0001  & n13819 ;
  assign n22360 = ~n22358 & ~n22359 ;
  assign n22361 = \wishbone_bd_ram_mem2_reg[173][21]/P0001  & n13360 ;
  assign n22362 = \wishbone_bd_ram_mem2_reg[94][21]/P0001  & n13833 ;
  assign n22363 = ~n22361 & ~n22362 ;
  assign n22364 = n22360 & n22363 ;
  assign n22365 = n22357 & n22364 ;
  assign n22366 = n22350 & n22365 ;
  assign n22367 = n22335 & n22366 ;
  assign n22368 = \wishbone_bd_ram_mem2_reg[117][21]/P0001  & n13557 ;
  assign n22369 = \wishbone_bd_ram_mem2_reg[100][21]/P0001  & n13401 ;
  assign n22370 = ~n22368 & ~n22369 ;
  assign n22371 = \wishbone_bd_ram_mem2_reg[182][21]/P0001  & n13598 ;
  assign n22372 = \wishbone_bd_ram_mem2_reg[247][21]/P0001  & n13571 ;
  assign n22373 = ~n22371 & ~n22372 ;
  assign n22374 = n22370 & n22373 ;
  assign n22375 = \wishbone_bd_ram_mem2_reg[191][21]/P0001  & n14012 ;
  assign n22376 = \wishbone_bd_ram_mem2_reg[214][21]/P0001  & n13938 ;
  assign n22377 = ~n22375 & ~n22376 ;
  assign n22378 = \wishbone_bd_ram_mem2_reg[120][21]/P0001  & n13550 ;
  assign n22379 = \wishbone_bd_ram_mem2_reg[5][21]/P0001  & n13243 ;
  assign n22380 = ~n22378 & ~n22379 ;
  assign n22381 = n22377 & n22380 ;
  assign n22382 = n22374 & n22381 ;
  assign n22383 = \wishbone_bd_ram_mem2_reg[237][21]/P0001  & n13924 ;
  assign n22384 = \wishbone_bd_ram_mem2_reg[21][21]/P0001  & n13438 ;
  assign n22385 = ~n22383 & ~n22384 ;
  assign n22386 = \wishbone_bd_ram_mem2_reg[134][21]/P0001  & n13494 ;
  assign n22387 = \wishbone_bd_ram_mem2_reg[211][21]/P0001  & n13805 ;
  assign n22388 = ~n22386 & ~n22387 ;
  assign n22389 = n22385 & n22388 ;
  assign n22390 = \wishbone_bd_ram_mem2_reg[108][21]/P0001  & n13814 ;
  assign n22391 = \wishbone_bd_ram_mem2_reg[190][21]/P0001  & n13365 ;
  assign n22392 = ~n22390 & ~n22391 ;
  assign n22393 = \wishbone_bd_ram_mem2_reg[45][21]/P0001  & n13420 ;
  assign n22394 = \wishbone_bd_ram_mem2_reg[15][21]/P0001  & n13797 ;
  assign n22395 = ~n22393 & ~n22394 ;
  assign n22396 = n22392 & n22395 ;
  assign n22397 = n22389 & n22396 ;
  assign n22398 = n22382 & n22397 ;
  assign n22399 = \wishbone_bd_ram_mem2_reg[203][21]/P0001  & n13816 ;
  assign n22400 = \wishbone_bd_ram_mem2_reg[229][21]/P0001  & n13552 ;
  assign n22401 = ~n22399 & ~n22400 ;
  assign n22402 = \wishbone_bd_ram_mem2_reg[116][21]/P0001  & n13865 ;
  assign n22403 = \wishbone_bd_ram_mem2_reg[234][21]/P0001  & n13781 ;
  assign n22404 = ~n22402 & ~n22403 ;
  assign n22405 = n22401 & n22404 ;
  assign n22406 = \wishbone_bd_ram_mem2_reg[51][21]/P0001  & n13880 ;
  assign n22407 = \wishbone_bd_ram_mem2_reg[93][21]/P0001  & n13891 ;
  assign n22408 = ~n22406 & ~n22407 ;
  assign n22409 = \wishbone_bd_ram_mem2_reg[226][21]/P0001  & n13668 ;
  assign n22410 = \wishbone_bd_ram_mem2_reg[176][21]/P0001  & n13262 ;
  assign n22411 = ~n22409 & ~n22410 ;
  assign n22412 = n22408 & n22411 ;
  assign n22413 = n22405 & n22412 ;
  assign n22414 = \wishbone_bd_ram_mem2_reg[121][21]/P0001  & n13983 ;
  assign n22415 = \wishbone_bd_ram_mem2_reg[10][21]/P0001  & n13837 ;
  assign n22416 = ~n22414 & ~n22415 ;
  assign n22417 = \wishbone_bd_ram_mem2_reg[147][21]/P0001  & n13702 ;
  assign n22418 = \wishbone_bd_ram_mem2_reg[206][21]/P0001  & n13414 ;
  assign n22419 = ~n22417 & ~n22418 ;
  assign n22420 = n22416 & n22419 ;
  assign n22421 = \wishbone_bd_ram_mem2_reg[243][21]/P0001  & n13575 ;
  assign n22422 = \wishbone_bd_ram_mem2_reg[248][21]/P0001  & n13647 ;
  assign n22423 = ~n22421 & ~n22422 ;
  assign n22424 = \wishbone_bd_ram_mem2_reg[189][21]/P0001  & n14001 ;
  assign n22425 = \wishbone_bd_ram_mem2_reg[174][21]/P0001  & n13899 ;
  assign n22426 = ~n22424 & ~n22425 ;
  assign n22427 = n22423 & n22426 ;
  assign n22428 = n22420 & n22427 ;
  assign n22429 = n22413 & n22428 ;
  assign n22430 = n22398 & n22429 ;
  assign n22431 = n22367 & n22430 ;
  assign n22432 = n22304 & n22431 ;
  assign n22433 = \wishbone_bd_ram_mem2_reg[42][21]/P0001  & n13341 ;
  assign n22434 = \wishbone_bd_ram_mem2_reg[26][21]/P0001  & n13521 ;
  assign n22435 = ~n22433 & ~n22434 ;
  assign n22436 = \wishbone_bd_ram_mem2_reg[152][21]/P0001  & n13912 ;
  assign n22437 = \wishbone_bd_ram_mem2_reg[233][21]/P0001  & n13332 ;
  assign n22438 = ~n22436 & ~n22437 ;
  assign n22439 = n22435 & n22438 ;
  assign n22440 = \wishbone_bd_ram_mem2_reg[12][21]/P0001  & n13733 ;
  assign n22441 = \wishbone_bd_ram_mem2_reg[20][21]/P0001  & n13839 ;
  assign n22442 = ~n22440 & ~n22441 ;
  assign n22443 = \wishbone_bd_ram_mem2_reg[221][21]/P0001  & n13641 ;
  assign n22444 = \wishbone_bd_ram_mem2_reg[35][21]/P0001  & n13523 ;
  assign n22445 = ~n22443 & ~n22444 ;
  assign n22446 = n22442 & n22445 ;
  assign n22447 = n22439 & n22446 ;
  assign n22448 = \wishbone_bd_ram_mem2_reg[84][21]/P0001  & n13385 ;
  assign n22449 = \wishbone_bd_ram_mem2_reg[153][21]/P0001  & n13309 ;
  assign n22450 = ~n22448 & ~n22449 ;
  assign n22451 = \wishbone_bd_ram_mem2_reg[106][21]/P0001  & n13555 ;
  assign n22452 = \wishbone_bd_ram_mem2_reg[92][21]/P0001  & n13859 ;
  assign n22453 = ~n22451 & ~n22452 ;
  assign n22454 = n22450 & n22453 ;
  assign n22455 = \wishbone_bd_ram_mem2_reg[160][21]/P0001  & n13271 ;
  assign n22456 = \wishbone_bd_ram_mem2_reg[61][21]/P0001  & n13544 ;
  assign n22457 = ~n22455 & ~n22456 ;
  assign n22458 = \wishbone_bd_ram_mem2_reg[136][21]/P0001  & n13963 ;
  assign n22459 = \wishbone_bd_ram_mem2_reg[41][21]/P0001  & n14017 ;
  assign n22460 = ~n22458 & ~n22459 ;
  assign n22461 = n22457 & n22460 ;
  assign n22462 = n22454 & n22461 ;
  assign n22463 = n22447 & n22462 ;
  assign n22464 = \wishbone_bd_ram_mem2_reg[201][21]/P0001  & n13600 ;
  assign n22465 = \wishbone_bd_ram_mem2_reg[33][21]/P0001  & n13933 ;
  assign n22466 = ~n22464 & ~n22465 ;
  assign n22467 = \wishbone_bd_ram_mem2_reg[223][21]/P0001  & n13335 ;
  assign n22468 = \wishbone_bd_ram_mem2_reg[72][21]/P0001  & n13582 ;
  assign n22469 = ~n22467 & ~n22468 ;
  assign n22470 = n22466 & n22469 ;
  assign n22471 = \wishbone_bd_ram_mem2_reg[76][21]/P0001  & n13831 ;
  assign n22472 = \wishbone_bd_ram_mem2_reg[75][21]/P0001  & n13605 ;
  assign n22473 = ~n22471 & ~n22472 ;
  assign n22474 = \wishbone_bd_ram_mem2_reg[71][21]/P0001  & n13636 ;
  assign n22475 = \wishbone_bd_ram_mem2_reg[105][21]/P0001  & n13503 ;
  assign n22476 = ~n22474 & ~n22475 ;
  assign n22477 = n22473 & n22476 ;
  assign n22478 = n22470 & n22477 ;
  assign n22479 = \wishbone_bd_ram_mem2_reg[236][21]/P0001  & n13480 ;
  assign n22480 = \wishbone_bd_ram_mem2_reg[199][21]/P0001  & n13499 ;
  assign n22481 = ~n22479 & ~n22480 ;
  assign n22482 = \wishbone_bd_ram_mem2_reg[66][21]/P0001  & n13603 ;
  assign n22483 = \wishbone_bd_ram_mem2_reg[31][21]/P0001  & n13758 ;
  assign n22484 = ~n22482 & ~n22483 ;
  assign n22485 = n22481 & n22484 ;
  assign n22486 = \wishbone_bd_ram_mem2_reg[188][21]/P0001  & n13407 ;
  assign n22487 = \wishbone_bd_ram_mem2_reg[158][21]/P0001  & n13294 ;
  assign n22488 = ~n22486 & ~n22487 ;
  assign n22489 = \wishbone_bd_ram_mem2_reg[239][21]/P0001  & n13349 ;
  assign n22490 = \wishbone_bd_ram_mem2_reg[91][21]/P0001  & n13954 ;
  assign n22491 = ~n22489 & ~n22490 ;
  assign n22492 = n22488 & n22491 ;
  assign n22493 = n22485 & n22492 ;
  assign n22494 = n22478 & n22493 ;
  assign n22495 = n22463 & n22494 ;
  assign n22496 = \wishbone_bd_ram_mem2_reg[240][21]/P0001  & n13352 ;
  assign n22497 = \wishbone_bd_ram_mem2_reg[32][21]/P0001  & n13736 ;
  assign n22498 = ~n22496 & ~n22497 ;
  assign n22499 = \wishbone_bd_ram_mem2_reg[88][21]/P0001  & n13347 ;
  assign n22500 = \wishbone_bd_ram_mem2_reg[205][21]/P0001  & n13947 ;
  assign n22501 = ~n22499 & ~n22500 ;
  assign n22502 = n22498 & n22501 ;
  assign n22503 = \wishbone_bd_ram_mem2_reg[219][21]/P0001  & n13577 ;
  assign n22504 = \wishbone_bd_ram_mem2_reg[103][21]/P0001  & n13320 ;
  assign n22505 = ~n22503 & ~n22504 ;
  assign n22506 = \wishbone_bd_ram_mem2_reg[245][21]/P0001  & n13877 ;
  assign n22507 = \wishbone_bd_ram_mem2_reg[251][21]/P0001  & n14019 ;
  assign n22508 = ~n22506 & ~n22507 ;
  assign n22509 = n22505 & n22508 ;
  assign n22510 = n22502 & n22509 ;
  assign n22511 = \wishbone_bd_ram_mem2_reg[96][21]/P0001  & n13425 ;
  assign n22512 = \wishbone_bd_ram_mem2_reg[228][21]/P0001  & n13497 ;
  assign n22513 = ~n22511 & ~n22512 ;
  assign n22514 = \wishbone_bd_ram_mem2_reg[18][21]/P0001  & n13532 ;
  assign n22515 = \wishbone_bd_ram_mem2_reg[126][21]/P0001  & n13786 ;
  assign n22516 = ~n22514 & ~n22515 ;
  assign n22517 = n22513 & n22516 ;
  assign n22518 = \wishbone_bd_ram_mem2_reg[161][21]/P0001  & n13505 ;
  assign n22519 = \wishbone_bd_ram_mem2_reg[36][21]/P0001  & n13639 ;
  assign n22520 = ~n22518 & ~n22519 ;
  assign n22521 = \wishbone_bd_ram_mem2_reg[55][21]/P0001  & n13618 ;
  assign n22522 = \wishbone_bd_ram_mem2_reg[215][21]/P0001  & n13901 ;
  assign n22523 = ~n22521 & ~n22522 ;
  assign n22524 = n22520 & n22523 ;
  assign n22525 = n22517 & n22524 ;
  assign n22526 = n22510 & n22525 ;
  assign n22527 = \wishbone_bd_ram_mem2_reg[118][21]/P0001  & n13589 ;
  assign n22528 = \wishbone_bd_ram_mem2_reg[16][21]/P0001  & n13695 ;
  assign n22529 = ~n22527 & ~n22528 ;
  assign n22530 = \wishbone_bd_ram_mem2_reg[6][21]/P0001  & n13915 ;
  assign n22531 = \wishbone_bd_ram_mem2_reg[139][21]/P0001  & n13566 ;
  assign n22532 = ~n22530 & ~n22531 ;
  assign n22533 = n22529 & n22532 ;
  assign n22534 = \wishbone_bd_ram_mem2_reg[98][21]/P0001  & n13569 ;
  assign n22535 = \wishbone_bd_ram_mem2_reg[200][21]/P0001  & n13922 ;
  assign n22536 = ~n22534 & ~n22535 ;
  assign n22537 = \wishbone_bd_ram_mem2_reg[59][21]/P0001  & n13613 ;
  assign n22538 = \wishbone_bd_ram_mem2_reg[113][21]/P0001  & n13882 ;
  assign n22539 = ~n22537 & ~n22538 ;
  assign n22540 = n22536 & n22539 ;
  assign n22541 = n22533 & n22540 ;
  assign n22542 = \wishbone_bd_ram_mem2_reg[253][21]/P0001  & n13708 ;
  assign n22543 = \wishbone_bd_ram_mem2_reg[39][21]/P0001  & n13893 ;
  assign n22544 = ~n22542 & ~n22543 ;
  assign n22545 = \wishbone_bd_ram_mem2_reg[194][21]/P0001  & n13624 ;
  assign n22546 = \wishbone_bd_ram_mem2_reg[133][21]/P0001  & n13492 ;
  assign n22547 = ~n22545 & ~n22546 ;
  assign n22548 = n22544 & n22547 ;
  assign n22549 = \wishbone_bd_ram_mem2_reg[97][21]/P0001  & n13724 ;
  assign n22550 = \wishbone_bd_ram_mem2_reg[89][21]/P0001  & n13910 ;
  assign n22551 = ~n22549 & ~n22550 ;
  assign n22552 = \wishbone_bd_ram_mem2_reg[0][21]/P0001  & n13539 ;
  assign n22553 = \wishbone_bd_ram_mem2_reg[107][21]/P0001  & n13476 ;
  assign n22554 = ~n22552 & ~n22553 ;
  assign n22555 = n22551 & n22554 ;
  assign n22556 = n22548 & n22555 ;
  assign n22557 = n22541 & n22556 ;
  assign n22558 = n22526 & n22557 ;
  assign n22559 = n22495 & n22558 ;
  assign n22560 = \wishbone_bd_ram_mem2_reg[13][21]/P0001  & n13844 ;
  assign n22561 = \wishbone_bd_ram_mem2_reg[241][21]/P0001  & n13854 ;
  assign n22562 = ~n22560 & ~n22561 ;
  assign n22563 = \wishbone_bd_ram_mem2_reg[167][21]/P0001  & n13940 ;
  assign n22564 = \wishbone_bd_ram_mem2_reg[53][21]/P0001  & n13875 ;
  assign n22565 = ~n22563 & ~n22564 ;
  assign n22566 = n22562 & n22565 ;
  assign n22567 = \wishbone_bd_ram_mem2_reg[135][21]/P0001  & n13672 ;
  assign n22568 = \wishbone_bd_ram_mem2_reg[46][21]/P0001  & n13298 ;
  assign n22569 = ~n22567 & ~n22568 ;
  assign n22570 = \wishbone_bd_ram_mem2_reg[47][21]/P0001  & n13436 ;
  assign n22571 = \wishbone_bd_ram_mem2_reg[132][21]/P0001  & n13927 ;
  assign n22572 = ~n22570 & ~n22571 ;
  assign n22573 = n22569 & n22572 ;
  assign n22574 = n22566 & n22573 ;
  assign n22575 = \wishbone_bd_ram_mem2_reg[83][21]/P0001  & n13454 ;
  assign n22576 = \wishbone_bd_ram_mem2_reg[252][21]/P0001  & n13986 ;
  assign n22577 = ~n22575 & ~n22576 ;
  assign n22578 = \wishbone_bd_ram_mem2_reg[154][21]/P0001  & n13403 ;
  assign n22579 = \wishbone_bd_ram_mem2_reg[231][21]/P0001  & n13363 ;
  assign n22580 = ~n22578 & ~n22579 ;
  assign n22581 = n22577 & n22580 ;
  assign n22582 = \wishbone_bd_ram_mem2_reg[227][21]/P0001  & n13388 ;
  assign n22583 = \wishbone_bd_ram_mem2_reg[34][21]/P0001  & n13450 ;
  assign n22584 = ~n22582 & ~n22583 ;
  assign n22585 = \wishbone_bd_ram_mem2_reg[11][21]/P0001  & n13774 ;
  assign n22586 = \wishbone_bd_ram_mem2_reg[131][21]/P0001  & n13358 ;
  assign n22587 = ~n22585 & ~n22586 ;
  assign n22588 = n22584 & n22587 ;
  assign n22589 = n22581 & n22588 ;
  assign n22590 = n22574 & n22589 ;
  assign n22591 = \wishbone_bd_ram_mem2_reg[57][21]/P0001  & n13731 ;
  assign n22592 = \wishbone_bd_ram_mem2_reg[123][21]/P0001  & n13749 ;
  assign n22593 = ~n22591 & ~n22592 ;
  assign n22594 = \wishbone_bd_ram_mem2_reg[3][21]/P0001  & n13354 ;
  assign n22595 = \wishbone_bd_ram_mem2_reg[130][21]/P0001  & n13427 ;
  assign n22596 = ~n22594 & ~n22595 ;
  assign n22597 = n22593 & n22596 ;
  assign n22598 = \wishbone_bd_ram_mem2_reg[224][21]/P0001  & n13433 ;
  assign n22599 = \wishbone_bd_ram_mem2_reg[54][21]/P0001  & n13622 ;
  assign n22600 = ~n22598 & ~n22599 ;
  assign n22601 = \wishbone_bd_ram_mem2_reg[137][21]/P0001  & n13808 ;
  assign n22602 = \wishbone_bd_ram_mem2_reg[172][21]/P0001  & n13377 ;
  assign n22603 = ~n22601 & ~n22602 ;
  assign n22604 = n22600 & n22603 ;
  assign n22605 = n22597 & n22604 ;
  assign n22606 = \wishbone_bd_ram_mem2_reg[56][21]/P0001  & n13611 ;
  assign n22607 = \wishbone_bd_ram_mem2_reg[150][21]/P0001  & n13666 ;
  assign n22608 = ~n22606 & ~n22607 ;
  assign n22609 = \wishbone_bd_ram_mem2_reg[74][21]/P0001  & n13564 ;
  assign n22610 = \wishbone_bd_ram_mem2_reg[79][21]/P0001  & n13779 ;
  assign n22611 = ~n22609 & ~n22610 ;
  assign n22612 = n22608 & n22611 ;
  assign n22613 = \wishbone_bd_ram_mem2_reg[244][21]/P0001  & n13474 ;
  assign n22614 = \wishbone_bd_ram_mem2_reg[49][21]/P0001  & n13929 ;
  assign n22615 = ~n22613 & ~n22614 ;
  assign n22616 = \wishbone_bd_ram_mem2_reg[217][21]/P0001  & n13767 ;
  assign n22617 = \wishbone_bd_ram_mem2_reg[138][21]/P0001  & n13398 ;
  assign n22618 = ~n22616 & ~n22617 ;
  assign n22619 = n22615 & n22618 ;
  assign n22620 = n22612 & n22619 ;
  assign n22621 = n22605 & n22620 ;
  assign n22622 = n22590 & n22621 ;
  assign n22623 = \wishbone_bd_ram_mem2_reg[185][21]/P0001  & n13372 ;
  assign n22624 = \wishbone_bd_ram_mem2_reg[43][21]/P0001  & n13761 ;
  assign n22625 = ~n22623 & ~n22624 ;
  assign n22626 = \wishbone_bd_ram_mem2_reg[69][21]/P0001  & n13487 ;
  assign n22627 = \wishbone_bd_ram_mem2_reg[249][21]/P0001  & n13431 ;
  assign n22628 = ~n22626 & ~n22627 ;
  assign n22629 = n22625 & n22628 ;
  assign n22630 = \wishbone_bd_ram_mem2_reg[29][21]/P0001  & n13412 ;
  assign n22631 = \wishbone_bd_ram_mem2_reg[110][21]/P0001  & n14030 ;
  assign n22632 = ~n22630 & ~n22631 ;
  assign n22633 = \wishbone_bd_ram_mem2_reg[19][21]/P0001  & n13886 ;
  assign n22634 = \wishbone_bd_ram_mem2_reg[204][21]/P0001  & n13821 ;
  assign n22635 = ~n22633 & ~n22634 ;
  assign n22636 = n22632 & n22635 ;
  assign n22637 = n22629 & n22636 ;
  assign n22638 = \wishbone_bd_ram_mem2_reg[4][21]/P0001  & n13527 ;
  assign n22639 = \wishbone_bd_ram_mem2_reg[202][21]/P0001  & n13268 ;
  assign n22640 = ~n22638 & ~n22639 ;
  assign n22641 = \wishbone_bd_ram_mem2_reg[235][21]/P0001  & n13518 ;
  assign n22642 = \wishbone_bd_ram_mem2_reg[159][21]/P0001  & n13627 ;
  assign n22643 = ~n22641 & ~n22642 ;
  assign n22644 = n22640 & n22643 ;
  assign n22645 = \wishbone_bd_ram_mem2_reg[187][21]/P0001  & n13756 ;
  assign n22646 = \wishbone_bd_ram_mem2_reg[67][21]/P0001  & n13663 ;
  assign n22647 = ~n22645 & ~n22646 ;
  assign n22648 = \wishbone_bd_ram_mem2_reg[73][21]/P0001  & n13456 ;
  assign n22649 = \wishbone_bd_ram_mem2_reg[197][21]/P0001  & n13594 ;
  assign n22650 = ~n22648 & ~n22649 ;
  assign n22651 = n22647 & n22650 ;
  assign n22652 = n22644 & n22651 ;
  assign n22653 = n22637 & n22652 ;
  assign n22654 = \wishbone_bd_ram_mem2_reg[146][21]/P0001  & n13958 ;
  assign n22655 = \wishbone_bd_ram_mem2_reg[124][21]/P0001  & n14024 ;
  assign n22656 = ~n22654 & ~n22655 ;
  assign n22657 = \wishbone_bd_ram_mem2_reg[164][21]/P0001  & n13236 ;
  assign n22658 = \wishbone_bd_ram_mem2_reg[52][21]/P0001  & n13988 ;
  assign n22659 = ~n22657 & ~n22658 ;
  assign n22660 = n22656 & n22659 ;
  assign n22661 = \wishbone_bd_ram_mem2_reg[216][21]/P0001  & n14005 ;
  assign n22662 = \wishbone_bd_ram_mem2_reg[170][21]/P0001  & n14007 ;
  assign n22663 = ~n22661 & ~n22662 ;
  assign n22664 = \wishbone_bd_ram_mem2_reg[142][21]/P0001  & n13448 ;
  assign n22665 = \wishbone_bd_ram_mem2_reg[140][21]/P0001  & n13287 ;
  assign n22666 = ~n22664 & ~n22665 ;
  assign n22667 = n22663 & n22666 ;
  assign n22668 = n22660 & n22667 ;
  assign n22669 = \wishbone_bd_ram_mem2_reg[250][21]/P0001  & n13677 ;
  assign n22670 = \wishbone_bd_ram_mem2_reg[225][21]/P0001  & n13719 ;
  assign n22671 = ~n22669 & ~n22670 ;
  assign n22672 = \wishbone_bd_ram_mem2_reg[112][21]/P0001  & n13482 ;
  assign n22673 = \wishbone_bd_ram_mem2_reg[25][21]/P0001  & n13742 ;
  assign n22674 = ~n22672 & ~n22673 ;
  assign n22675 = n22671 & n22674 ;
  assign n22676 = \wishbone_bd_ram_mem2_reg[163][21]/P0001  & n13255 ;
  assign n22677 = \wishbone_bd_ram_mem2_reg[218][21]/P0001  & n13792 ;
  assign n22678 = ~n22676 & ~n22677 ;
  assign n22679 = \wishbone_bd_ram_mem2_reg[180][21]/P0001  & n13650 ;
  assign n22680 = \wishbone_bd_ram_mem2_reg[86][21]/P0001  & n13485 ;
  assign n22681 = ~n22679 & ~n22680 ;
  assign n22682 = n22678 & n22681 ;
  assign n22683 = n22675 & n22682 ;
  assign n22684 = n22668 & n22683 ;
  assign n22685 = n22653 & n22684 ;
  assign n22686 = n22622 & n22685 ;
  assign n22687 = n22559 & n22686 ;
  assign n22688 = n22432 & n22687 ;
  assign n22689 = n14047 & ~n22688 ;
  assign n22690 = ~n22177 & ~n22689 ;
  assign n22691 = \wishbone_LatchedTxLength_reg[7]/NET0131  & ~n14046 ;
  assign n22692 = \wishbone_bd_ram_mem2_reg[38][23]/P0001  & n13828 ;
  assign n22693 = \wishbone_bd_ram_mem2_reg[85][23]/P0001  & n13784 ;
  assign n22694 = ~n22692 & ~n22693 ;
  assign n22695 = \wishbone_bd_ram_mem2_reg[50][23]/P0001  & n13686 ;
  assign n22696 = \wishbone_bd_ram_mem2_reg[31][23]/P0001  & n13758 ;
  assign n22697 = ~n22695 & ~n22696 ;
  assign n22698 = n22694 & n22697 ;
  assign n22699 = \wishbone_bd_ram_mem2_reg[139][23]/P0001  & n13566 ;
  assign n22700 = \wishbone_bd_ram_mem2_reg[35][23]/P0001  & n13523 ;
  assign n22701 = ~n22699 & ~n22700 ;
  assign n22702 = \wishbone_bd_ram_mem2_reg[5][23]/P0001  & n13243 ;
  assign n22703 = \wishbone_bd_ram_mem2_reg[199][23]/P0001  & n13499 ;
  assign n22704 = ~n22702 & ~n22703 ;
  assign n22705 = n22701 & n22704 ;
  assign n22706 = n22698 & n22705 ;
  assign n22707 = \wishbone_bd_ram_mem2_reg[202][23]/P0001  & n13268 ;
  assign n22708 = \wishbone_bd_ram_mem2_reg[191][23]/P0001  & n14012 ;
  assign n22709 = ~n22707 & ~n22708 ;
  assign n22710 = \wishbone_bd_ram_mem2_reg[68][23]/P0001  & n13379 ;
  assign n22711 = \wishbone_bd_ram_mem2_reg[228][23]/P0001  & n13497 ;
  assign n22712 = ~n22710 & ~n22711 ;
  assign n22713 = n22709 & n22712 ;
  assign n22714 = \wishbone_bd_ram_mem2_reg[11][23]/P0001  & n13774 ;
  assign n22715 = \wishbone_bd_ram_mem2_reg[178][23]/P0001  & n13301 ;
  assign n22716 = ~n22714 & ~n22715 ;
  assign n22717 = \wishbone_bd_ram_mem2_reg[210][23]/P0001  & n13443 ;
  assign n22718 = \wishbone_bd_ram_mem2_reg[231][23]/P0001  & n13363 ;
  assign n22719 = ~n22717 & ~n22718 ;
  assign n22720 = n22716 & n22719 ;
  assign n22721 = n22713 & n22720 ;
  assign n22722 = n22706 & n22721 ;
  assign n22723 = \wishbone_bd_ram_mem2_reg[88][23]/P0001  & n13347 ;
  assign n22724 = \wishbone_bd_ram_mem2_reg[103][23]/P0001  & n13320 ;
  assign n22725 = ~n22723 & ~n22724 ;
  assign n22726 = \wishbone_bd_ram_mem2_reg[61][23]/P0001  & n13544 ;
  assign n22727 = \wishbone_bd_ram_mem2_reg[53][23]/P0001  & n13875 ;
  assign n22728 = ~n22726 & ~n22727 ;
  assign n22729 = n22725 & n22728 ;
  assign n22730 = \wishbone_bd_ram_mem2_reg[249][23]/P0001  & n13431 ;
  assign n22731 = \wishbone_bd_ram_mem2_reg[179][23]/P0001  & n14035 ;
  assign n22732 = ~n22730 & ~n22731 ;
  assign n22733 = \wishbone_bd_ram_mem2_reg[66][23]/P0001  & n13603 ;
  assign n22734 = \wishbone_bd_ram_mem2_reg[180][23]/P0001  & n13650 ;
  assign n22735 = ~n22733 & ~n22734 ;
  assign n22736 = n22732 & n22735 ;
  assign n22737 = n22729 & n22736 ;
  assign n22738 = \wishbone_bd_ram_mem2_reg[3][23]/P0001  & n13354 ;
  assign n22739 = \wishbone_bd_ram_mem2_reg[194][23]/P0001  & n13624 ;
  assign n22740 = ~n22738 & ~n22739 ;
  assign n22741 = \wishbone_bd_ram_mem2_reg[219][23]/P0001  & n13577 ;
  assign n22742 = \wishbone_bd_ram_mem2_reg[79][23]/P0001  & n13779 ;
  assign n22743 = ~n22741 & ~n22742 ;
  assign n22744 = n22740 & n22743 ;
  assign n22745 = \wishbone_bd_ram_mem2_reg[166][23]/P0001  & n13999 ;
  assign n22746 = \wishbone_bd_ram_mem2_reg[126][23]/P0001  & n13786 ;
  assign n22747 = ~n22745 & ~n22746 ;
  assign n22748 = \wishbone_bd_ram_mem2_reg[153][23]/P0001  & n13309 ;
  assign n22749 = \wishbone_bd_ram_mem2_reg[201][23]/P0001  & n13600 ;
  assign n22750 = ~n22748 & ~n22749 ;
  assign n22751 = n22747 & n22750 ;
  assign n22752 = n22744 & n22751 ;
  assign n22753 = n22737 & n22752 ;
  assign n22754 = n22722 & n22753 ;
  assign n22755 = \wishbone_bd_ram_mem2_reg[209][23]/P0001  & n13689 ;
  assign n22756 = \wishbone_bd_ram_mem2_reg[196][23]/P0001  & n13977 ;
  assign n22757 = ~n22755 & ~n22756 ;
  assign n22758 = \wishbone_bd_ram_mem2_reg[10][23]/P0001  & n13837 ;
  assign n22759 = \wishbone_bd_ram_mem2_reg[24][23]/P0001  & n13970 ;
  assign n22760 = ~n22758 & ~n22759 ;
  assign n22761 = n22757 & n22760 ;
  assign n22762 = \wishbone_bd_ram_mem2_reg[175][23]/P0001  & n13674 ;
  assign n22763 = \wishbone_bd_ram_mem2_reg[64][23]/P0001  & n13904 ;
  assign n22764 = ~n22762 & ~n22763 ;
  assign n22765 = \wishbone_bd_ram_mem2_reg[239][23]/P0001  & n13349 ;
  assign n22766 = \wishbone_bd_ram_mem2_reg[118][23]/P0001  & n13589 ;
  assign n22767 = ~n22765 & ~n22766 ;
  assign n22768 = n22764 & n22767 ;
  assign n22769 = n22761 & n22768 ;
  assign n22770 = \wishbone_bd_ram_mem2_reg[78][23]/P0001  & n13277 ;
  assign n22771 = \wishbone_bd_ram_mem2_reg[207][23]/P0001  & n13826 ;
  assign n22772 = ~n22770 & ~n22771 ;
  assign n22773 = \wishbone_bd_ram_mem2_reg[117][23]/P0001  & n13557 ;
  assign n22774 = \wishbone_bd_ram_mem2_reg[237][23]/P0001  & n13924 ;
  assign n22775 = ~n22773 & ~n22774 ;
  assign n22776 = n22772 & n22775 ;
  assign n22777 = \wishbone_bd_ram_mem2_reg[241][23]/P0001  & n13854 ;
  assign n22778 = \wishbone_bd_ram_mem2_reg[227][23]/P0001  & n13388 ;
  assign n22779 = ~n22777 & ~n22778 ;
  assign n22780 = \wishbone_bd_ram_mem2_reg[9][23]/P0001  & n13580 ;
  assign n22781 = \wishbone_bd_ram_mem2_reg[206][23]/P0001  & n13414 ;
  assign n22782 = ~n22780 & ~n22781 ;
  assign n22783 = n22779 & n22782 ;
  assign n22784 = n22776 & n22783 ;
  assign n22785 = n22769 & n22784 ;
  assign n22786 = \wishbone_bd_ram_mem2_reg[92][23]/P0001  & n13859 ;
  assign n22787 = \wishbone_bd_ram_mem2_reg[230][23]/P0001  & n13994 ;
  assign n22788 = ~n22786 & ~n22787 ;
  assign n22789 = \wishbone_bd_ram_mem2_reg[182][23]/P0001  & n13598 ;
  assign n22790 = \wishbone_bd_ram_mem2_reg[80][23]/P0001  & n13516 ;
  assign n22791 = ~n22789 & ~n22790 ;
  assign n22792 = n22788 & n22791 ;
  assign n22793 = \wishbone_bd_ram_mem2_reg[213][23]/P0001  & n13870 ;
  assign n22794 = \wishbone_bd_ram_mem2_reg[212][23]/P0001  & n13634 ;
  assign n22795 = ~n22793 & ~n22794 ;
  assign n22796 = \wishbone_bd_ram_mem2_reg[47][23]/P0001  & n13436 ;
  assign n22797 = \wishbone_bd_ram_mem2_reg[1][23]/P0001  & n13888 ;
  assign n22798 = ~n22796 & ~n22797 ;
  assign n22799 = n22795 & n22798 ;
  assign n22800 = n22792 & n22799 ;
  assign n22801 = \wishbone_bd_ram_mem2_reg[123][23]/P0001  & n13749 ;
  assign n22802 = \wishbone_bd_ram_mem2_reg[149][23]/P0001  & n13469 ;
  assign n22803 = ~n22801 & ~n22802 ;
  assign n22804 = \wishbone_bd_ram_mem2_reg[7][23]/P0001  & n13546 ;
  assign n22805 = \wishbone_bd_ram_mem2_reg[203][23]/P0001  & n13816 ;
  assign n22806 = ~n22804 & ~n22805 ;
  assign n22807 = n22803 & n22806 ;
  assign n22808 = \wishbone_bd_ram_mem2_reg[97][23]/P0001  & n13724 ;
  assign n22809 = \wishbone_bd_ram_mem2_reg[138][23]/P0001  & n13398 ;
  assign n22810 = ~n22808 & ~n22809 ;
  assign n22811 = \wishbone_bd_ram_mem2_reg[8][23]/P0001  & n13459 ;
  assign n22812 = \wishbone_bd_ram_mem2_reg[62][23]/P0001  & n13529 ;
  assign n22813 = ~n22811 & ~n22812 ;
  assign n22814 = n22810 & n22813 ;
  assign n22815 = n22807 & n22814 ;
  assign n22816 = n22800 & n22815 ;
  assign n22817 = n22785 & n22816 ;
  assign n22818 = n22754 & n22817 ;
  assign n22819 = \wishbone_bd_ram_mem2_reg[157][23]/P0001  & n13445 ;
  assign n22820 = \wishbone_bd_ram_mem2_reg[105][23]/P0001  & n13503 ;
  assign n22821 = ~n22819 & ~n22820 ;
  assign n22822 = \wishbone_bd_ram_mem2_reg[220][23]/P0001  & n13965 ;
  assign n22823 = \wishbone_bd_ram_mem2_reg[125][23]/P0001  & n13396 ;
  assign n22824 = ~n22822 & ~n22823 ;
  assign n22825 = n22821 & n22824 ;
  assign n22826 = \wishbone_bd_ram_mem2_reg[243][23]/P0001  & n13575 ;
  assign n22827 = \wishbone_bd_ram_mem2_reg[70][23]/P0001  & n13339 ;
  assign n22828 = ~n22826 & ~n22827 ;
  assign n22829 = \wishbone_bd_ram_mem2_reg[161][23]/P0001  & n13505 ;
  assign n22830 = \wishbone_bd_ram_mem2_reg[29][23]/P0001  & n13412 ;
  assign n22831 = ~n22829 & ~n22830 ;
  assign n22832 = n22828 & n22831 ;
  assign n22833 = n22825 & n22832 ;
  assign n22834 = \wishbone_bd_ram_mem2_reg[82][23]/P0001  & n13374 ;
  assign n22835 = \wishbone_bd_ram_mem2_reg[55][23]/P0001  & n13618 ;
  assign n22836 = ~n22834 & ~n22835 ;
  assign n22837 = \wishbone_bd_ram_mem2_reg[81][23]/P0001  & n13409 ;
  assign n22838 = \wishbone_bd_ram_mem2_reg[223][23]/P0001  & n13335 ;
  assign n22839 = ~n22837 & ~n22838 ;
  assign n22840 = n22836 & n22839 ;
  assign n22841 = \wishbone_bd_ram_mem2_reg[111][23]/P0001  & n13471 ;
  assign n22842 = \wishbone_bd_ram_mem2_reg[160][23]/P0001  & n13271 ;
  assign n22843 = ~n22841 & ~n22842 ;
  assign n22844 = \wishbone_bd_ram_mem2_reg[192][23]/P0001  & n13390 ;
  assign n22845 = \wishbone_bd_ram_mem2_reg[159][23]/P0001  & n13627 ;
  assign n22846 = ~n22844 & ~n22845 ;
  assign n22847 = n22843 & n22846 ;
  assign n22848 = n22840 & n22847 ;
  assign n22849 = n22833 & n22848 ;
  assign n22850 = \wishbone_bd_ram_mem2_reg[189][23]/P0001  & n14001 ;
  assign n22851 = \wishbone_bd_ram_mem2_reg[197][23]/P0001  & n13594 ;
  assign n22852 = ~n22850 & ~n22851 ;
  assign n22853 = \wishbone_bd_ram_mem2_reg[72][23]/P0001  & n13582 ;
  assign n22854 = \wishbone_bd_ram_mem2_reg[6][23]/P0001  & n13915 ;
  assign n22855 = ~n22853 & ~n22854 ;
  assign n22856 = n22852 & n22855 ;
  assign n22857 = \wishbone_bd_ram_mem2_reg[43][23]/P0001  & n13761 ;
  assign n22858 = \wishbone_bd_ram_mem2_reg[18][23]/P0001  & n13532 ;
  assign n22859 = ~n22857 & ~n22858 ;
  assign n22860 = \wishbone_bd_ram_mem2_reg[236][23]/P0001  & n13480 ;
  assign n22861 = \wishbone_bd_ram_mem2_reg[102][23]/P0001  & n13534 ;
  assign n22862 = ~n22860 & ~n22861 ;
  assign n22863 = n22859 & n22862 ;
  assign n22864 = n22856 & n22863 ;
  assign n22865 = \wishbone_bd_ram_mem2_reg[235][23]/P0001  & n13518 ;
  assign n22866 = \wishbone_bd_ram_mem2_reg[112][23]/P0001  & n13482 ;
  assign n22867 = ~n22865 & ~n22866 ;
  assign n22868 = \wishbone_bd_ram_mem2_reg[34][23]/P0001  & n13450 ;
  assign n22869 = \wishbone_bd_ram_mem2_reg[251][23]/P0001  & n14019 ;
  assign n22870 = ~n22868 & ~n22869 ;
  assign n22871 = n22867 & n22870 ;
  assign n22872 = \wishbone_bd_ram_mem2_reg[141][23]/P0001  & n13852 ;
  assign n22873 = \wishbone_bd_ram_mem2_reg[238][23]/P0001  & n13819 ;
  assign n22874 = ~n22872 & ~n22873 ;
  assign n22875 = \wishbone_bd_ram_mem2_reg[114][23]/P0001  & n13763 ;
  assign n22876 = \wishbone_bd_ram_mem2_reg[75][23]/P0001  & n13605 ;
  assign n22877 = ~n22875 & ~n22876 ;
  assign n22878 = n22874 & n22877 ;
  assign n22879 = n22871 & n22878 ;
  assign n22880 = n22864 & n22879 ;
  assign n22881 = n22849 & n22880 ;
  assign n22882 = \wishbone_bd_ram_mem2_reg[109][23]/P0001  & n13306 ;
  assign n22883 = \wishbone_bd_ram_mem2_reg[142][23]/P0001  & n13448 ;
  assign n22884 = ~n22882 & ~n22883 ;
  assign n22885 = \wishbone_bd_ram_mem2_reg[104][23]/P0001  & n13684 ;
  assign n22886 = \wishbone_bd_ram_mem2_reg[151][23]/P0001  & n13697 ;
  assign n22887 = ~n22885 & ~n22886 ;
  assign n22888 = n22884 & n22887 ;
  assign n22889 = \wishbone_bd_ram_mem2_reg[211][23]/P0001  & n13805 ;
  assign n22890 = \wishbone_bd_ram_mem2_reg[240][23]/P0001  & n13352 ;
  assign n22891 = ~n22889 & ~n22890 ;
  assign n22892 = \wishbone_bd_ram_mem2_reg[255][23]/P0001  & n13952 ;
  assign n22893 = \wishbone_bd_ram_mem2_reg[135][23]/P0001  & n13672 ;
  assign n22894 = ~n22892 & ~n22893 ;
  assign n22895 = n22891 & n22894 ;
  assign n22896 = n22888 & n22895 ;
  assign n22897 = \wishbone_bd_ram_mem2_reg[181][23]/P0001  & n13587 ;
  assign n22898 = \wishbone_bd_ram_mem2_reg[144][23]/P0001  & n13508 ;
  assign n22899 = ~n22897 & ~n22898 ;
  assign n22900 = \wishbone_bd_ram_mem2_reg[134][23]/P0001  & n13494 ;
  assign n22901 = \wishbone_bd_ram_mem2_reg[107][23]/P0001  & n13476 ;
  assign n22902 = ~n22900 & ~n22901 ;
  assign n22903 = n22899 & n22902 ;
  assign n22904 = \wishbone_bd_ram_mem2_reg[164][23]/P0001  & n13236 ;
  assign n22905 = \wishbone_bd_ram_mem2_reg[133][23]/P0001  & n13492 ;
  assign n22906 = ~n22904 & ~n22905 ;
  assign n22907 = \wishbone_bd_ram_mem2_reg[163][23]/P0001  & n13255 ;
  assign n22908 = \wishbone_bd_ram_mem2_reg[136][23]/P0001  & n13963 ;
  assign n22909 = ~n22907 & ~n22908 ;
  assign n22910 = n22906 & n22909 ;
  assign n22911 = n22903 & n22910 ;
  assign n22912 = n22896 & n22911 ;
  assign n22913 = \wishbone_bd_ram_mem2_reg[56][23]/P0001  & n13611 ;
  assign n22914 = \wishbone_bd_ram_mem2_reg[59][23]/P0001  & n13613 ;
  assign n22915 = ~n22913 & ~n22914 ;
  assign n22916 = \wishbone_bd_ram_mem2_reg[129][23]/P0001  & n13629 ;
  assign n22917 = \wishbone_bd_ram_mem2_reg[245][23]/P0001  & n13877 ;
  assign n22918 = ~n22916 & ~n22917 ;
  assign n22919 = n22915 & n22918 ;
  assign n22920 = \wishbone_bd_ram_mem2_reg[54][23]/P0001  & n13622 ;
  assign n22921 = \wishbone_bd_ram_mem2_reg[234][23]/P0001  & n13781 ;
  assign n22922 = ~n22920 & ~n22921 ;
  assign n22923 = \wishbone_bd_ram_mem2_reg[222][23]/P0001  & n13721 ;
  assign n22924 = \wishbone_bd_ram_mem2_reg[73][23]/P0001  & n13456 ;
  assign n22925 = ~n22923 & ~n22924 ;
  assign n22926 = n22922 & n22925 ;
  assign n22927 = n22919 & n22926 ;
  assign n22928 = \wishbone_bd_ram_mem2_reg[140][23]/P0001  & n13287 ;
  assign n22929 = \wishbone_bd_ram_mem2_reg[87][23]/P0001  & n13691 ;
  assign n22930 = ~n22928 & ~n22929 ;
  assign n22931 = \wishbone_bd_ram_mem2_reg[51][23]/P0001  & n13880 ;
  assign n22932 = \wishbone_bd_ram_mem2_reg[250][23]/P0001  & n13677 ;
  assign n22933 = ~n22931 & ~n22932 ;
  assign n22934 = n22930 & n22933 ;
  assign n22935 = \wishbone_bd_ram_mem2_reg[242][23]/P0001  & n13383 ;
  assign n22936 = \wishbone_bd_ram_mem2_reg[214][23]/P0001  & n13938 ;
  assign n22937 = ~n22935 & ~n22936 ;
  assign n22938 = \wishbone_bd_ram_mem2_reg[20][23]/P0001  & n13839 ;
  assign n22939 = \wishbone_bd_ram_mem2_reg[65][23]/P0001  & n13842 ;
  assign n22940 = ~n22938 & ~n22939 ;
  assign n22941 = n22937 & n22940 ;
  assign n22942 = n22934 & n22941 ;
  assign n22943 = n22927 & n22942 ;
  assign n22944 = n22912 & n22943 ;
  assign n22945 = n22881 & n22944 ;
  assign n22946 = n22818 & n22945 ;
  assign n22947 = \wishbone_bd_ram_mem2_reg[2][23]/P0001  & n13975 ;
  assign n22948 = \wishbone_bd_ram_mem2_reg[42][23]/P0001  & n13341 ;
  assign n22949 = ~n22947 & ~n22948 ;
  assign n22950 = \wishbone_bd_ram_mem2_reg[218][23]/P0001  & n13792 ;
  assign n22951 = \wishbone_bd_ram_mem2_reg[158][23]/P0001  & n13294 ;
  assign n22952 = ~n22950 & ~n22951 ;
  assign n22953 = n22949 & n22952 ;
  assign n22954 = \wishbone_bd_ram_mem2_reg[12][23]/P0001  & n13733 ;
  assign n22955 = \wishbone_bd_ram_mem2_reg[30][23]/P0001  & n13713 ;
  assign n22956 = ~n22954 & ~n22955 ;
  assign n22957 = \wishbone_bd_ram_mem2_reg[221][23]/P0001  & n13641 ;
  assign n22958 = \wishbone_bd_ram_mem2_reg[188][23]/P0001  & n13407 ;
  assign n22959 = ~n22957 & ~n22958 ;
  assign n22960 = n22956 & n22959 ;
  assign n22961 = n22953 & n22960 ;
  assign n22962 = \wishbone_bd_ram_mem2_reg[98][23]/P0001  & n13569 ;
  assign n22963 = \wishbone_bd_ram_mem2_reg[27][23]/P0001  & n13251 ;
  assign n22964 = ~n22962 & ~n22963 ;
  assign n22965 = \wishbone_bd_ram_mem2_reg[205][23]/P0001  & n13947 ;
  assign n22966 = \wishbone_bd_ram_mem2_reg[71][23]/P0001  & n13636 ;
  assign n22967 = ~n22965 & ~n22966 ;
  assign n22968 = n22964 & n22967 ;
  assign n22969 = \wishbone_bd_ram_mem2_reg[40][23]/P0001  & n13661 ;
  assign n22970 = \wishbone_bd_ram_mem2_reg[21][23]/P0001  & n13438 ;
  assign n22971 = ~n22969 & ~n22970 ;
  assign n22972 = \wishbone_bd_ram_mem2_reg[101][23]/P0001  & n13772 ;
  assign n22973 = \wishbone_bd_ram_mem2_reg[147][23]/P0001  & n13702 ;
  assign n22974 = ~n22972 & ~n22973 ;
  assign n22975 = n22971 & n22974 ;
  assign n22976 = n22968 & n22975 ;
  assign n22977 = n22961 & n22976 ;
  assign n22978 = \wishbone_bd_ram_mem2_reg[233][23]/P0001  & n13332 ;
  assign n22979 = \wishbone_bd_ram_mem2_reg[37][23]/P0001  & n13710 ;
  assign n22980 = ~n22978 & ~n22979 ;
  assign n22981 = \wishbone_bd_ram_mem2_reg[177][23]/P0001  & n13863 ;
  assign n22982 = \wishbone_bd_ram_mem2_reg[174][23]/P0001  & n13899 ;
  assign n22983 = ~n22981 & ~n22982 ;
  assign n22984 = n22980 & n22983 ;
  assign n22985 = \wishbone_bd_ram_mem2_reg[94][23]/P0001  & n13833 ;
  assign n22986 = \wishbone_bd_ram_mem2_reg[176][23]/P0001  & n13262 ;
  assign n22987 = ~n22985 & ~n22986 ;
  assign n22988 = \wishbone_bd_ram_mem2_reg[172][23]/P0001  & n13377 ;
  assign n22989 = \wishbone_bd_ram_mem2_reg[193][23]/P0001  & n14022 ;
  assign n22990 = ~n22988 & ~n22989 ;
  assign n22991 = n22987 & n22990 ;
  assign n22992 = n22984 & n22991 ;
  assign n22993 = \wishbone_bd_ram_mem2_reg[67][23]/P0001  & n13663 ;
  assign n22994 = \wishbone_bd_ram_mem2_reg[121][23]/P0001  & n13983 ;
  assign n22995 = ~n22993 & ~n22994 ;
  assign n22996 = \wishbone_bd_ram_mem2_reg[48][23]/P0001  & n13917 ;
  assign n22997 = \wishbone_bd_ram_mem2_reg[169][23]/P0001  & n13541 ;
  assign n22998 = ~n22996 & ~n22997 ;
  assign n22999 = n22995 & n22998 ;
  assign n23000 = \wishbone_bd_ram_mem2_reg[99][23]/P0001  & n13996 ;
  assign n23001 = \wishbone_bd_ram_mem2_reg[186][23]/P0001  & n13616 ;
  assign n23002 = ~n23000 & ~n23001 ;
  assign n23003 = \wishbone_bd_ram_mem2_reg[195][23]/P0001  & n13700 ;
  assign n23004 = \wishbone_bd_ram_mem2_reg[76][23]/P0001  & n13831 ;
  assign n23005 = ~n23003 & ~n23004 ;
  assign n23006 = n23002 & n23005 ;
  assign n23007 = n22999 & n23006 ;
  assign n23008 = n22992 & n23007 ;
  assign n23009 = n22977 & n23008 ;
  assign n23010 = \wishbone_bd_ram_mem2_reg[217][23]/P0001  & n13767 ;
  assign n23011 = \wishbone_bd_ram_mem2_reg[162][23]/P0001  & n13726 ;
  assign n23012 = ~n23010 & ~n23011 ;
  assign n23013 = \wishbone_bd_ram_mem2_reg[4][23]/P0001  & n13527 ;
  assign n23014 = \wishbone_bd_ram_mem2_reg[106][23]/P0001  & n13555 ;
  assign n23015 = ~n23013 & ~n23014 ;
  assign n23016 = n23012 & n23015 ;
  assign n23017 = \wishbone_bd_ram_mem2_reg[246][23]/P0001  & n13981 ;
  assign n23018 = \wishbone_bd_ram_mem2_reg[156][23]/P0001  & n13769 ;
  assign n23019 = ~n23017 & ~n23018 ;
  assign n23020 = \wishbone_bd_ram_mem2_reg[74][23]/P0001  & n13564 ;
  assign n23021 = \wishbone_bd_ram_mem2_reg[91][23]/P0001  & n13954 ;
  assign n23022 = ~n23020 & ~n23021 ;
  assign n23023 = n23019 & n23022 ;
  assign n23024 = n23016 & n23023 ;
  assign n23025 = \wishbone_bd_ram_mem2_reg[95][23]/P0001  & n13317 ;
  assign n23026 = \wishbone_bd_ram_mem2_reg[232][23]/P0001  & n13510 ;
  assign n23027 = ~n23025 & ~n23026 ;
  assign n23028 = \wishbone_bd_ram_mem2_reg[13][23]/P0001  & n13844 ;
  assign n23029 = \wishbone_bd_ram_mem2_reg[173][23]/P0001  & n13360 ;
  assign n23030 = ~n23028 & ~n23029 ;
  assign n23031 = n23027 & n23030 ;
  assign n23032 = \wishbone_bd_ram_mem2_reg[26][23]/P0001  & n13521 ;
  assign n23033 = \wishbone_bd_ram_mem2_reg[150][23]/P0001  & n13666 ;
  assign n23034 = ~n23032 & ~n23033 ;
  assign n23035 = \wishbone_bd_ram_mem2_reg[22][23]/P0001  & n13744 ;
  assign n23036 = \wishbone_bd_ram_mem2_reg[168][23]/P0001  & n13795 ;
  assign n23037 = ~n23035 & ~n23036 ;
  assign n23038 = n23034 & n23037 ;
  assign n23039 = n23031 & n23038 ;
  assign n23040 = n23024 & n23039 ;
  assign n23041 = \wishbone_bd_ram_mem2_reg[127][23]/P0001  & n13803 ;
  assign n23042 = \wishbone_bd_ram_mem2_reg[224][23]/P0001  & n13433 ;
  assign n23043 = ~n23041 & ~n23042 ;
  assign n23044 = \wishbone_bd_ram_mem2_reg[229][23]/P0001  & n13552 ;
  assign n23045 = \wishbone_bd_ram_mem2_reg[225][23]/P0001  & n13719 ;
  assign n23046 = ~n23044 & ~n23045 ;
  assign n23047 = n23043 & n23046 ;
  assign n23048 = \wishbone_bd_ram_mem2_reg[58][23]/P0001  & n13949 ;
  assign n23049 = \wishbone_bd_ram_mem2_reg[200][23]/P0001  & n13922 ;
  assign n23050 = ~n23048 & ~n23049 ;
  assign n23051 = \wishbone_bd_ram_mem2_reg[254][23]/P0001  & n13283 ;
  assign n23052 = \wishbone_bd_ram_mem2_reg[204][23]/P0001  & n13821 ;
  assign n23053 = ~n23051 & ~n23052 ;
  assign n23054 = n23050 & n23053 ;
  assign n23055 = n23047 & n23054 ;
  assign n23056 = \wishbone_bd_ram_mem2_reg[252][23]/P0001  & n13986 ;
  assign n23057 = \wishbone_bd_ram_mem2_reg[77][23]/P0001  & n13935 ;
  assign n23058 = ~n23056 & ~n23057 ;
  assign n23059 = \wishbone_bd_ram_mem2_reg[116][23]/P0001  & n13865 ;
  assign n23060 = \wishbone_bd_ram_mem2_reg[23][23]/P0001  & n13857 ;
  assign n23061 = ~n23059 & ~n23060 ;
  assign n23062 = n23058 & n23061 ;
  assign n23063 = \wishbone_bd_ram_mem2_reg[83][23]/P0001  & n13454 ;
  assign n23064 = \wishbone_bd_ram_mem2_reg[69][23]/P0001  & n13487 ;
  assign n23065 = ~n23063 & ~n23064 ;
  assign n23066 = \wishbone_bd_ram_mem2_reg[119][23]/P0001  & n14033 ;
  assign n23067 = \wishbone_bd_ram_mem2_reg[146][23]/P0001  & n13958 ;
  assign n23068 = ~n23066 & ~n23067 ;
  assign n23069 = n23065 & n23068 ;
  assign n23070 = n23062 & n23069 ;
  assign n23071 = n23055 & n23070 ;
  assign n23072 = n23040 & n23071 ;
  assign n23073 = n23009 & n23072 ;
  assign n23074 = \wishbone_bd_ram_mem2_reg[0][23]/P0001  & n13539 ;
  assign n23075 = \wishbone_bd_ram_mem2_reg[122][23]/P0001  & n13679 ;
  assign n23076 = ~n23074 & ~n23075 ;
  assign n23077 = \wishbone_bd_ram_mem2_reg[46][23]/P0001  & n13298 ;
  assign n23078 = \wishbone_bd_ram_mem2_reg[155][23]/P0001  & n13738 ;
  assign n23079 = ~n23077 & ~n23078 ;
  assign n23080 = n23076 & n23079 ;
  assign n23081 = \wishbone_bd_ram_mem2_reg[57][23]/P0001  & n13731 ;
  assign n23082 = \wishbone_bd_ram_mem2_reg[28][23]/P0001  & n13810 ;
  assign n23083 = ~n23081 & ~n23082 ;
  assign n23084 = \wishbone_bd_ram_mem2_reg[148][23]/P0001  & n13868 ;
  assign n23085 = \wishbone_bd_ram_mem2_reg[190][23]/P0001  & n13365 ;
  assign n23086 = ~n23084 & ~n23085 ;
  assign n23087 = n23083 & n23086 ;
  assign n23088 = n23080 & n23087 ;
  assign n23089 = \wishbone_bd_ram_mem2_reg[63][23]/P0001  & n13327 ;
  assign n23090 = \wishbone_bd_ram_mem2_reg[253][23]/P0001  & n13708 ;
  assign n23091 = ~n23089 & ~n23090 ;
  assign n23092 = \wishbone_bd_ram_mem2_reg[36][23]/P0001  & n13639 ;
  assign n23093 = \wishbone_bd_ram_mem2_reg[113][23]/P0001  & n13882 ;
  assign n23094 = ~n23092 & ~n23093 ;
  assign n23095 = n23091 & n23094 ;
  assign n23096 = \wishbone_bd_ram_mem2_reg[132][23]/P0001  & n13927 ;
  assign n23097 = \wishbone_bd_ram_mem2_reg[17][23]/P0001  & n13324 ;
  assign n23098 = ~n23096 & ~n23097 ;
  assign n23099 = \wishbone_bd_ram_mem2_reg[208][23]/P0001  & n14010 ;
  assign n23100 = \wishbone_bd_ram_mem2_reg[49][23]/P0001  & n13929 ;
  assign n23101 = ~n23099 & ~n23100 ;
  assign n23102 = n23098 & n23101 ;
  assign n23103 = n23095 & n23102 ;
  assign n23104 = n23088 & n23103 ;
  assign n23105 = \wishbone_bd_ram_mem2_reg[120][23]/P0001  & n13550 ;
  assign n23106 = \wishbone_bd_ram_mem2_reg[115][23]/P0001  & n13747 ;
  assign n23107 = ~n23105 & ~n23106 ;
  assign n23108 = \wishbone_bd_ram_mem2_reg[84][23]/P0001  & n13385 ;
  assign n23109 = \wishbone_bd_ram_mem2_reg[16][23]/P0001  & n13695 ;
  assign n23110 = ~n23108 & ~n23109 ;
  assign n23111 = n23107 & n23110 ;
  assign n23112 = \wishbone_bd_ram_mem2_reg[143][23]/P0001  & n13461 ;
  assign n23113 = \wishbone_bd_ram_mem2_reg[152][23]/P0001  & n13912 ;
  assign n23114 = ~n23112 & ~n23113 ;
  assign n23115 = \wishbone_bd_ram_mem2_reg[25][23]/P0001  & n13742 ;
  assign n23116 = \wishbone_bd_ram_mem2_reg[32][23]/P0001  & n13736 ;
  assign n23117 = ~n23115 & ~n23116 ;
  assign n23118 = n23114 & n23117 ;
  assign n23119 = n23111 & n23118 ;
  assign n23120 = \wishbone_bd_ram_mem2_reg[247][23]/P0001  & n13571 ;
  assign n23121 = \wishbone_bd_ram_mem2_reg[154][23]/P0001  & n13403 ;
  assign n23122 = ~n23120 & ~n23121 ;
  assign n23123 = \wishbone_bd_ram_mem2_reg[93][23]/P0001  & n13891 ;
  assign n23124 = \wishbone_bd_ram_mem2_reg[39][23]/P0001  & n13893 ;
  assign n23125 = ~n23123 & ~n23124 ;
  assign n23126 = n23122 & n23125 ;
  assign n23127 = \wishbone_bd_ram_mem2_reg[33][23]/P0001  & n13933 ;
  assign n23128 = \wishbone_bd_ram_mem2_reg[131][23]/P0001  & n13358 ;
  assign n23129 = ~n23127 & ~n23128 ;
  assign n23130 = \wishbone_bd_ram_mem2_reg[248][23]/P0001  & n13647 ;
  assign n23131 = \wishbone_bd_ram_mem2_reg[15][23]/P0001  & n13797 ;
  assign n23132 = ~n23130 & ~n23131 ;
  assign n23133 = n23129 & n23132 ;
  assign n23134 = n23126 & n23133 ;
  assign n23135 = n23119 & n23134 ;
  assign n23136 = n23104 & n23135 ;
  assign n23137 = \wishbone_bd_ram_mem2_reg[170][23]/P0001  & n14007 ;
  assign n23138 = \wishbone_bd_ram_mem2_reg[44][23]/P0001  & n13291 ;
  assign n23139 = ~n23137 & ~n23138 ;
  assign n23140 = \wishbone_bd_ram_mem2_reg[90][23]/P0001  & n13906 ;
  assign n23141 = \wishbone_bd_ram_mem2_reg[198][23]/P0001  & n13592 ;
  assign n23142 = ~n23140 & ~n23141 ;
  assign n23143 = n23139 & n23142 ;
  assign n23144 = \wishbone_bd_ram_mem2_reg[128][23]/P0001  & n13652 ;
  assign n23145 = \wishbone_bd_ram_mem2_reg[184][23]/P0001  & n13960 ;
  assign n23146 = ~n23144 & ~n23145 ;
  assign n23147 = \wishbone_bd_ram_mem2_reg[19][23]/P0001  & n13886 ;
  assign n23148 = \wishbone_bd_ram_mem2_reg[244][23]/P0001  & n13474 ;
  assign n23149 = ~n23147 & ~n23148 ;
  assign n23150 = n23146 & n23149 ;
  assign n23151 = n23143 & n23150 ;
  assign n23152 = \wishbone_bd_ram_mem2_reg[96][23]/P0001  & n13425 ;
  assign n23153 = \wishbone_bd_ram_mem2_reg[14][23]/P0001  & n13972 ;
  assign n23154 = ~n23152 & ~n23153 ;
  assign n23155 = \wishbone_bd_ram_mem2_reg[89][23]/P0001  & n13910 ;
  assign n23156 = \wishbone_bd_ram_mem2_reg[100][23]/P0001  & n13401 ;
  assign n23157 = ~n23155 & ~n23156 ;
  assign n23158 = n23154 & n23157 ;
  assign n23159 = \wishbone_bd_ram_mem2_reg[216][23]/P0001  & n14005 ;
  assign n23160 = \wishbone_bd_ram_mem2_reg[86][23]/P0001  & n13485 ;
  assign n23161 = ~n23159 & ~n23160 ;
  assign n23162 = \wishbone_bd_ram_mem2_reg[215][23]/P0001  & n13901 ;
  assign n23163 = \wishbone_bd_ram_mem2_reg[145][23]/P0001  & n13715 ;
  assign n23164 = ~n23162 & ~n23163 ;
  assign n23165 = n23161 & n23164 ;
  assign n23166 = n23158 & n23165 ;
  assign n23167 = n23151 & n23166 ;
  assign n23168 = \wishbone_bd_ram_mem2_reg[52][23]/P0001  & n13988 ;
  assign n23169 = \wishbone_bd_ram_mem2_reg[137][23]/P0001  & n13808 ;
  assign n23170 = ~n23168 & ~n23169 ;
  assign n23171 = \wishbone_bd_ram_mem2_reg[108][23]/P0001  & n13814 ;
  assign n23172 = \wishbone_bd_ram_mem2_reg[60][23]/P0001  & n13790 ;
  assign n23173 = ~n23171 & ~n23172 ;
  assign n23174 = n23170 & n23173 ;
  assign n23175 = \wishbone_bd_ram_mem2_reg[187][23]/P0001  & n13756 ;
  assign n23176 = \wishbone_bd_ram_mem2_reg[185][23]/P0001  & n13372 ;
  assign n23177 = ~n23175 & ~n23176 ;
  assign n23178 = \wishbone_bd_ram_mem2_reg[167][23]/P0001  & n13940 ;
  assign n23179 = \wishbone_bd_ram_mem2_reg[130][23]/P0001  & n13427 ;
  assign n23180 = ~n23178 & ~n23179 ;
  assign n23181 = n23177 & n23180 ;
  assign n23182 = n23174 & n23181 ;
  assign n23183 = \wishbone_bd_ram_mem2_reg[41][23]/P0001  & n14017 ;
  assign n23184 = \wishbone_bd_ram_mem2_reg[226][23]/P0001  & n13668 ;
  assign n23185 = ~n23183 & ~n23184 ;
  assign n23186 = \wishbone_bd_ram_mem2_reg[165][23]/P0001  & n14028 ;
  assign n23187 = \wishbone_bd_ram_mem2_reg[124][23]/P0001  & n14024 ;
  assign n23188 = ~n23186 & ~n23187 ;
  assign n23189 = n23185 & n23188 ;
  assign n23190 = \wishbone_bd_ram_mem2_reg[45][23]/P0001  & n13420 ;
  assign n23191 = \wishbone_bd_ram_mem2_reg[110][23]/P0001  & n14030 ;
  assign n23192 = ~n23190 & ~n23191 ;
  assign n23193 = \wishbone_bd_ram_mem2_reg[183][23]/P0001  & n13645 ;
  assign n23194 = \wishbone_bd_ram_mem2_reg[171][23]/P0001  & n13422 ;
  assign n23195 = ~n23193 & ~n23194 ;
  assign n23196 = n23192 & n23195 ;
  assign n23197 = n23189 & n23196 ;
  assign n23198 = n23182 & n23197 ;
  assign n23199 = n23167 & n23198 ;
  assign n23200 = n23136 & n23199 ;
  assign n23201 = n23073 & n23200 ;
  assign n23202 = n22946 & n23201 ;
  assign n23203 = n14047 & ~n23202 ;
  assign n23204 = ~n22691 & ~n23203 ;
  assign n23205 = \wishbone_LatchedTxLength_reg[8]/NET0131  & ~n14046 ;
  assign n23206 = ~n15696 & ~n23205 ;
  assign n23207 = \wishbone_LatchedTxLength_reg[6]/NET0131  & ~n14046 ;
  assign n23208 = \wishbone_bd_ram_mem2_reg[86][22]/P0001  & n13485 ;
  assign n23209 = \wishbone_bd_ram_mem2_reg[79][22]/P0001  & n13779 ;
  assign n23210 = ~n23208 & ~n23209 ;
  assign n23211 = \wishbone_bd_ram_mem2_reg[52][22]/P0001  & n13988 ;
  assign n23212 = \wishbone_bd_ram_mem2_reg[74][22]/P0001  & n13564 ;
  assign n23213 = ~n23211 & ~n23212 ;
  assign n23214 = n23210 & n23213 ;
  assign n23215 = \wishbone_bd_ram_mem2_reg[202][22]/P0001  & n13268 ;
  assign n23216 = \wishbone_bd_ram_mem2_reg[228][22]/P0001  & n13497 ;
  assign n23217 = ~n23215 & ~n23216 ;
  assign n23218 = \wishbone_bd_ram_mem2_reg[64][22]/P0001  & n13904 ;
  assign n23219 = \wishbone_bd_ram_mem2_reg[247][22]/P0001  & n13571 ;
  assign n23220 = ~n23218 & ~n23219 ;
  assign n23221 = n23217 & n23220 ;
  assign n23222 = n23214 & n23221 ;
  assign n23223 = \wishbone_bd_ram_mem2_reg[133][22]/P0001  & n13492 ;
  assign n23224 = \wishbone_bd_ram_mem2_reg[204][22]/P0001  & n13821 ;
  assign n23225 = ~n23223 & ~n23224 ;
  assign n23226 = \wishbone_bd_ram_mem2_reg[135][22]/P0001  & n13672 ;
  assign n23227 = \wishbone_bd_ram_mem2_reg[111][22]/P0001  & n13471 ;
  assign n23228 = ~n23226 & ~n23227 ;
  assign n23229 = n23225 & n23228 ;
  assign n23230 = \wishbone_bd_ram_mem2_reg[32][22]/P0001  & n13736 ;
  assign n23231 = \wishbone_bd_ram_mem2_reg[194][22]/P0001  & n13624 ;
  assign n23232 = ~n23230 & ~n23231 ;
  assign n23233 = \wishbone_bd_ram_mem2_reg[51][22]/P0001  & n13880 ;
  assign n23234 = \wishbone_bd_ram_mem2_reg[180][22]/P0001  & n13650 ;
  assign n23235 = ~n23233 & ~n23234 ;
  assign n23236 = n23232 & n23235 ;
  assign n23237 = n23229 & n23236 ;
  assign n23238 = n23222 & n23237 ;
  assign n23239 = \wishbone_bd_ram_mem2_reg[42][22]/P0001  & n13341 ;
  assign n23240 = \wishbone_bd_ram_mem2_reg[107][22]/P0001  & n13476 ;
  assign n23241 = ~n23239 & ~n23240 ;
  assign n23242 = \wishbone_bd_ram_mem2_reg[2][22]/P0001  & n13975 ;
  assign n23243 = \wishbone_bd_ram_mem2_reg[138][22]/P0001  & n13398 ;
  assign n23244 = ~n23242 & ~n23243 ;
  assign n23245 = n23241 & n23244 ;
  assign n23246 = \wishbone_bd_ram_mem2_reg[248][22]/P0001  & n13647 ;
  assign n23247 = \wishbone_bd_ram_mem2_reg[164][22]/P0001  & n13236 ;
  assign n23248 = ~n23246 & ~n23247 ;
  assign n23249 = \wishbone_bd_ram_mem2_reg[251][22]/P0001  & n14019 ;
  assign n23250 = \wishbone_bd_ram_mem2_reg[50][22]/P0001  & n13686 ;
  assign n23251 = ~n23249 & ~n23250 ;
  assign n23252 = n23248 & n23251 ;
  assign n23253 = n23245 & n23252 ;
  assign n23254 = \wishbone_bd_ram_mem2_reg[174][22]/P0001  & n13899 ;
  assign n23255 = \wishbone_bd_ram_mem2_reg[165][22]/P0001  & n14028 ;
  assign n23256 = ~n23254 & ~n23255 ;
  assign n23257 = \wishbone_bd_ram_mem2_reg[226][22]/P0001  & n13668 ;
  assign n23258 = \wishbone_bd_ram_mem2_reg[243][22]/P0001  & n13575 ;
  assign n23259 = ~n23257 & ~n23258 ;
  assign n23260 = n23256 & n23259 ;
  assign n23261 = \wishbone_bd_ram_mem2_reg[30][22]/P0001  & n13713 ;
  assign n23262 = \wishbone_bd_ram_mem2_reg[212][22]/P0001  & n13634 ;
  assign n23263 = ~n23261 & ~n23262 ;
  assign n23264 = \wishbone_bd_ram_mem2_reg[146][22]/P0001  & n13958 ;
  assign n23265 = \wishbone_bd_ram_mem2_reg[206][22]/P0001  & n13414 ;
  assign n23266 = ~n23264 & ~n23265 ;
  assign n23267 = n23263 & n23266 ;
  assign n23268 = n23260 & n23267 ;
  assign n23269 = n23253 & n23268 ;
  assign n23270 = n23238 & n23269 ;
  assign n23271 = \wishbone_bd_ram_mem2_reg[140][22]/P0001  & n13287 ;
  assign n23272 = \wishbone_bd_ram_mem2_reg[59][22]/P0001  & n13613 ;
  assign n23273 = ~n23271 & ~n23272 ;
  assign n23274 = \wishbone_bd_ram_mem2_reg[176][22]/P0001  & n13262 ;
  assign n23275 = \wishbone_bd_ram_mem2_reg[67][22]/P0001  & n13663 ;
  assign n23276 = ~n23274 & ~n23275 ;
  assign n23277 = n23273 & n23276 ;
  assign n23278 = \wishbone_bd_ram_mem2_reg[106][22]/P0001  & n13555 ;
  assign n23279 = \wishbone_bd_ram_mem2_reg[85][22]/P0001  & n13784 ;
  assign n23280 = ~n23278 & ~n23279 ;
  assign n23281 = \wishbone_bd_ram_mem2_reg[221][22]/P0001  & n13641 ;
  assign n23282 = \wishbone_bd_ram_mem2_reg[128][22]/P0001  & n13652 ;
  assign n23283 = ~n23281 & ~n23282 ;
  assign n23284 = n23280 & n23283 ;
  assign n23285 = n23277 & n23284 ;
  assign n23286 = \wishbone_bd_ram_mem2_reg[104][22]/P0001  & n13684 ;
  assign n23287 = \wishbone_bd_ram_mem2_reg[41][22]/P0001  & n14017 ;
  assign n23288 = ~n23286 & ~n23287 ;
  assign n23289 = \wishbone_bd_ram_mem2_reg[63][22]/P0001  & n13327 ;
  assign n23290 = \wishbone_bd_ram_mem2_reg[210][22]/P0001  & n13443 ;
  assign n23291 = ~n23289 & ~n23290 ;
  assign n23292 = n23288 & n23291 ;
  assign n23293 = \wishbone_bd_ram_mem2_reg[222][22]/P0001  & n13721 ;
  assign n23294 = \wishbone_bd_ram_mem2_reg[254][22]/P0001  & n13283 ;
  assign n23295 = ~n23293 & ~n23294 ;
  assign n23296 = \wishbone_bd_ram_mem2_reg[148][22]/P0001  & n13868 ;
  assign n23297 = \wishbone_bd_ram_mem2_reg[239][22]/P0001  & n13349 ;
  assign n23298 = ~n23296 & ~n23297 ;
  assign n23299 = n23295 & n23298 ;
  assign n23300 = n23292 & n23299 ;
  assign n23301 = n23285 & n23300 ;
  assign n23302 = \wishbone_bd_ram_mem2_reg[116][22]/P0001  & n13865 ;
  assign n23303 = \wishbone_bd_ram_mem2_reg[144][22]/P0001  & n13508 ;
  assign n23304 = ~n23302 & ~n23303 ;
  assign n23305 = \wishbone_bd_ram_mem2_reg[80][22]/P0001  & n13516 ;
  assign n23306 = \wishbone_bd_ram_mem2_reg[108][22]/P0001  & n13814 ;
  assign n23307 = ~n23305 & ~n23306 ;
  assign n23308 = n23304 & n23307 ;
  assign n23309 = \wishbone_bd_ram_mem2_reg[214][22]/P0001  & n13938 ;
  assign n23310 = \wishbone_bd_ram_mem2_reg[173][22]/P0001  & n13360 ;
  assign n23311 = ~n23309 & ~n23310 ;
  assign n23312 = \wishbone_bd_ram_mem2_reg[60][22]/P0001  & n13790 ;
  assign n23313 = \wishbone_bd_ram_mem2_reg[5][22]/P0001  & n13243 ;
  assign n23314 = ~n23312 & ~n23313 ;
  assign n23315 = n23311 & n23314 ;
  assign n23316 = n23308 & n23315 ;
  assign n23317 = \wishbone_bd_ram_mem2_reg[97][22]/P0001  & n13724 ;
  assign n23318 = \wishbone_bd_ram_mem2_reg[141][22]/P0001  & n13852 ;
  assign n23319 = ~n23317 & ~n23318 ;
  assign n23320 = \wishbone_bd_ram_mem2_reg[58][22]/P0001  & n13949 ;
  assign n23321 = \wishbone_bd_ram_mem2_reg[0][22]/P0001  & n13539 ;
  assign n23322 = ~n23320 & ~n23321 ;
  assign n23323 = n23319 & n23322 ;
  assign n23324 = \wishbone_bd_ram_mem2_reg[76][22]/P0001  & n13831 ;
  assign n23325 = \wishbone_bd_ram_mem2_reg[14][22]/P0001  & n13972 ;
  assign n23326 = ~n23324 & ~n23325 ;
  assign n23327 = \wishbone_bd_ram_mem2_reg[57][22]/P0001  & n13731 ;
  assign n23328 = \wishbone_bd_ram_mem2_reg[153][22]/P0001  & n13309 ;
  assign n23329 = ~n23327 & ~n23328 ;
  assign n23330 = n23326 & n23329 ;
  assign n23331 = n23323 & n23330 ;
  assign n23332 = n23316 & n23331 ;
  assign n23333 = n23301 & n23332 ;
  assign n23334 = n23270 & n23333 ;
  assign n23335 = \wishbone_bd_ram_mem2_reg[160][22]/P0001  & n13271 ;
  assign n23336 = \wishbone_bd_ram_mem2_reg[23][22]/P0001  & n13857 ;
  assign n23337 = ~n23335 & ~n23336 ;
  assign n23338 = \wishbone_bd_ram_mem2_reg[191][22]/P0001  & n14012 ;
  assign n23339 = \wishbone_bd_ram_mem2_reg[98][22]/P0001  & n13569 ;
  assign n23340 = ~n23338 & ~n23339 ;
  assign n23341 = n23337 & n23340 ;
  assign n23342 = \wishbone_bd_ram_mem2_reg[200][22]/P0001  & n13922 ;
  assign n23343 = \wishbone_bd_ram_mem2_reg[139][22]/P0001  & n13566 ;
  assign n23344 = ~n23342 & ~n23343 ;
  assign n23345 = \wishbone_bd_ram_mem2_reg[61][22]/P0001  & n13544 ;
  assign n23346 = \wishbone_bd_ram_mem2_reg[17][22]/P0001  & n13324 ;
  assign n23347 = ~n23345 & ~n23346 ;
  assign n23348 = n23344 & n23347 ;
  assign n23349 = n23341 & n23348 ;
  assign n23350 = \wishbone_bd_ram_mem2_reg[112][22]/P0001  & n13482 ;
  assign n23351 = \wishbone_bd_ram_mem2_reg[169][22]/P0001  & n13541 ;
  assign n23352 = ~n23350 & ~n23351 ;
  assign n23353 = \wishbone_bd_ram_mem2_reg[105][22]/P0001  & n13503 ;
  assign n23354 = \wishbone_bd_ram_mem2_reg[220][22]/P0001  & n13965 ;
  assign n23355 = ~n23353 & ~n23354 ;
  assign n23356 = n23352 & n23355 ;
  assign n23357 = \wishbone_bd_ram_mem2_reg[75][22]/P0001  & n13605 ;
  assign n23358 = \wishbone_bd_ram_mem2_reg[157][22]/P0001  & n13445 ;
  assign n23359 = ~n23357 & ~n23358 ;
  assign n23360 = \wishbone_bd_ram_mem2_reg[145][22]/P0001  & n13715 ;
  assign n23361 = \wishbone_bd_ram_mem2_reg[237][22]/P0001  & n13924 ;
  assign n23362 = ~n23360 & ~n23361 ;
  assign n23363 = n23359 & n23362 ;
  assign n23364 = n23356 & n23363 ;
  assign n23365 = n23349 & n23364 ;
  assign n23366 = \wishbone_bd_ram_mem2_reg[56][22]/P0001  & n13611 ;
  assign n23367 = \wishbone_bd_ram_mem2_reg[127][22]/P0001  & n13803 ;
  assign n23368 = ~n23366 & ~n23367 ;
  assign n23369 = \wishbone_bd_ram_mem2_reg[49][22]/P0001  & n13929 ;
  assign n23370 = \wishbone_bd_ram_mem2_reg[15][22]/P0001  & n13797 ;
  assign n23371 = ~n23369 & ~n23370 ;
  assign n23372 = n23368 & n23371 ;
  assign n23373 = \wishbone_bd_ram_mem2_reg[189][22]/P0001  & n14001 ;
  assign n23374 = \wishbone_bd_ram_mem2_reg[166][22]/P0001  & n13999 ;
  assign n23375 = ~n23373 & ~n23374 ;
  assign n23376 = \wishbone_bd_ram_mem2_reg[44][22]/P0001  & n13291 ;
  assign n23377 = \wishbone_bd_ram_mem2_reg[121][22]/P0001  & n13983 ;
  assign n23378 = ~n23376 & ~n23377 ;
  assign n23379 = n23375 & n23378 ;
  assign n23380 = n23372 & n23379 ;
  assign n23381 = \wishbone_bd_ram_mem2_reg[38][22]/P0001  & n13828 ;
  assign n23382 = \wishbone_bd_ram_mem2_reg[234][22]/P0001  & n13781 ;
  assign n23383 = ~n23381 & ~n23382 ;
  assign n23384 = \wishbone_bd_ram_mem2_reg[20][22]/P0001  & n13839 ;
  assign n23385 = \wishbone_bd_ram_mem2_reg[45][22]/P0001  & n13420 ;
  assign n23386 = ~n23384 & ~n23385 ;
  assign n23387 = n23383 & n23386 ;
  assign n23388 = \wishbone_bd_ram_mem2_reg[156][22]/P0001  & n13769 ;
  assign n23389 = \wishbone_bd_ram_mem2_reg[252][22]/P0001  & n13986 ;
  assign n23390 = ~n23388 & ~n23389 ;
  assign n23391 = \wishbone_bd_ram_mem2_reg[175][22]/P0001  & n13674 ;
  assign n23392 = \wishbone_bd_ram_mem2_reg[53][22]/P0001  & n13875 ;
  assign n23393 = ~n23391 & ~n23392 ;
  assign n23394 = n23390 & n23393 ;
  assign n23395 = n23387 & n23394 ;
  assign n23396 = n23380 & n23395 ;
  assign n23397 = n23365 & n23396 ;
  assign n23398 = \wishbone_bd_ram_mem2_reg[35][22]/P0001  & n13523 ;
  assign n23399 = \wishbone_bd_ram_mem2_reg[184][22]/P0001  & n13960 ;
  assign n23400 = ~n23398 & ~n23399 ;
  assign n23401 = \wishbone_bd_ram_mem2_reg[16][22]/P0001  & n13695 ;
  assign n23402 = \wishbone_bd_ram_mem2_reg[130][22]/P0001  & n13427 ;
  assign n23403 = ~n23401 & ~n23402 ;
  assign n23404 = n23400 & n23403 ;
  assign n23405 = \wishbone_bd_ram_mem2_reg[244][22]/P0001  & n13474 ;
  assign n23406 = \wishbone_bd_ram_mem2_reg[215][22]/P0001  & n13901 ;
  assign n23407 = ~n23405 & ~n23406 ;
  assign n23408 = \wishbone_bd_ram_mem2_reg[217][22]/P0001  & n13767 ;
  assign n23409 = \wishbone_bd_ram_mem2_reg[34][22]/P0001  & n13450 ;
  assign n23410 = ~n23408 & ~n23409 ;
  assign n23411 = n23407 & n23410 ;
  assign n23412 = n23404 & n23411 ;
  assign n23413 = \wishbone_bd_ram_mem2_reg[207][22]/P0001  & n13826 ;
  assign n23414 = \wishbone_bd_ram_mem2_reg[26][22]/P0001  & n13521 ;
  assign n23415 = ~n23413 & ~n23414 ;
  assign n23416 = \wishbone_bd_ram_mem2_reg[154][22]/P0001  & n13403 ;
  assign n23417 = \wishbone_bd_ram_mem2_reg[113][22]/P0001  & n13882 ;
  assign n23418 = ~n23416 & ~n23417 ;
  assign n23419 = n23415 & n23418 ;
  assign n23420 = \wishbone_bd_ram_mem2_reg[143][22]/P0001  & n13461 ;
  assign n23421 = \wishbone_bd_ram_mem2_reg[96][22]/P0001  & n13425 ;
  assign n23422 = ~n23420 & ~n23421 ;
  assign n23423 = \wishbone_bd_ram_mem2_reg[136][22]/P0001  & n13963 ;
  assign n23424 = \wishbone_bd_ram_mem2_reg[137][22]/P0001  & n13808 ;
  assign n23425 = ~n23423 & ~n23424 ;
  assign n23426 = n23422 & n23425 ;
  assign n23427 = n23419 & n23426 ;
  assign n23428 = n23412 & n23427 ;
  assign n23429 = \wishbone_bd_ram_mem2_reg[18][22]/P0001  & n13532 ;
  assign n23430 = \wishbone_bd_ram_mem2_reg[55][22]/P0001  & n13618 ;
  assign n23431 = ~n23429 & ~n23430 ;
  assign n23432 = \wishbone_bd_ram_mem2_reg[77][22]/P0001  & n13935 ;
  assign n23433 = \wishbone_bd_ram_mem2_reg[66][22]/P0001  & n13603 ;
  assign n23434 = ~n23432 & ~n23433 ;
  assign n23435 = n23431 & n23434 ;
  assign n23436 = \wishbone_bd_ram_mem2_reg[100][22]/P0001  & n13401 ;
  assign n23437 = \wishbone_bd_ram_mem2_reg[246][22]/P0001  & n13981 ;
  assign n23438 = ~n23436 & ~n23437 ;
  assign n23439 = \wishbone_bd_ram_mem2_reg[10][22]/P0001  & n13837 ;
  assign n23440 = \wishbone_bd_ram_mem2_reg[31][22]/P0001  & n13758 ;
  assign n23441 = ~n23439 & ~n23440 ;
  assign n23442 = n23438 & n23441 ;
  assign n23443 = n23435 & n23442 ;
  assign n23444 = \wishbone_bd_ram_mem2_reg[203][22]/P0001  & n13816 ;
  assign n23445 = \wishbone_bd_ram_mem2_reg[232][22]/P0001  & n13510 ;
  assign n23446 = ~n23444 & ~n23445 ;
  assign n23447 = \wishbone_bd_ram_mem2_reg[159][22]/P0001  & n13627 ;
  assign n23448 = \wishbone_bd_ram_mem2_reg[233][22]/P0001  & n13332 ;
  assign n23449 = ~n23447 & ~n23448 ;
  assign n23450 = n23446 & n23449 ;
  assign n23451 = \wishbone_bd_ram_mem2_reg[114][22]/P0001  & n13763 ;
  assign n23452 = \wishbone_bd_ram_mem2_reg[208][22]/P0001  & n14010 ;
  assign n23453 = ~n23451 & ~n23452 ;
  assign n23454 = \wishbone_bd_ram_mem2_reg[95][22]/P0001  & n13317 ;
  assign n23455 = \wishbone_bd_ram_mem2_reg[24][22]/P0001  & n13970 ;
  assign n23456 = ~n23454 & ~n23455 ;
  assign n23457 = n23453 & n23456 ;
  assign n23458 = n23450 & n23457 ;
  assign n23459 = n23443 & n23458 ;
  assign n23460 = n23428 & n23459 ;
  assign n23461 = n23397 & n23460 ;
  assign n23462 = n23334 & n23461 ;
  assign n23463 = \wishbone_bd_ram_mem2_reg[4][22]/P0001  & n13527 ;
  assign n23464 = \wishbone_bd_ram_mem2_reg[21][22]/P0001  & n13438 ;
  assign n23465 = ~n23463 & ~n23464 ;
  assign n23466 = \wishbone_bd_ram_mem2_reg[167][22]/P0001  & n13940 ;
  assign n23467 = \wishbone_bd_ram_mem2_reg[181][22]/P0001  & n13587 ;
  assign n23468 = ~n23466 & ~n23467 ;
  assign n23469 = n23465 & n23468 ;
  assign n23470 = \wishbone_bd_ram_mem2_reg[149][22]/P0001  & n13469 ;
  assign n23471 = \wishbone_bd_ram_mem2_reg[1][22]/P0001  & n13888 ;
  assign n23472 = ~n23470 & ~n23471 ;
  assign n23473 = \wishbone_bd_ram_mem2_reg[201][22]/P0001  & n13600 ;
  assign n23474 = \wishbone_bd_ram_mem2_reg[117][22]/P0001  & n13557 ;
  assign n23475 = ~n23473 & ~n23474 ;
  assign n23476 = n23472 & n23475 ;
  assign n23477 = n23469 & n23476 ;
  assign n23478 = \wishbone_bd_ram_mem2_reg[72][22]/P0001  & n13582 ;
  assign n23479 = \wishbone_bd_ram_mem2_reg[9][22]/P0001  & n13580 ;
  assign n23480 = ~n23478 & ~n23479 ;
  assign n23481 = \wishbone_bd_ram_mem2_reg[90][22]/P0001  & n13906 ;
  assign n23482 = \wishbone_bd_ram_mem2_reg[168][22]/P0001  & n13795 ;
  assign n23483 = ~n23481 & ~n23482 ;
  assign n23484 = n23480 & n23483 ;
  assign n23485 = \wishbone_bd_ram_mem2_reg[47][22]/P0001  & n13436 ;
  assign n23486 = \wishbone_bd_ram_mem2_reg[125][22]/P0001  & n13396 ;
  assign n23487 = ~n23485 & ~n23486 ;
  assign n23488 = \wishbone_bd_ram_mem2_reg[216][22]/P0001  & n14005 ;
  assign n23489 = \wishbone_bd_ram_mem2_reg[19][22]/P0001  & n13886 ;
  assign n23490 = ~n23488 & ~n23489 ;
  assign n23491 = n23487 & n23490 ;
  assign n23492 = n23484 & n23491 ;
  assign n23493 = n23477 & n23492 ;
  assign n23494 = \wishbone_bd_ram_mem2_reg[250][22]/P0001  & n13677 ;
  assign n23495 = \wishbone_bd_ram_mem2_reg[12][22]/P0001  & n13733 ;
  assign n23496 = ~n23494 & ~n23495 ;
  assign n23497 = \wishbone_bd_ram_mem2_reg[27][22]/P0001  & n13251 ;
  assign n23498 = \wishbone_bd_ram_mem2_reg[88][22]/P0001  & n13347 ;
  assign n23499 = ~n23497 & ~n23498 ;
  assign n23500 = n23496 & n23499 ;
  assign n23501 = \wishbone_bd_ram_mem2_reg[187][22]/P0001  & n13756 ;
  assign n23502 = \wishbone_bd_ram_mem2_reg[172][22]/P0001  & n13377 ;
  assign n23503 = ~n23501 & ~n23502 ;
  assign n23504 = \wishbone_bd_ram_mem2_reg[109][22]/P0001  & n13306 ;
  assign n23505 = \wishbone_bd_ram_mem2_reg[82][22]/P0001  & n13374 ;
  assign n23506 = ~n23504 & ~n23505 ;
  assign n23507 = n23503 & n23506 ;
  assign n23508 = n23500 & n23507 ;
  assign n23509 = \wishbone_bd_ram_mem2_reg[131][22]/P0001  & n13358 ;
  assign n23510 = \wishbone_bd_ram_mem2_reg[68][22]/P0001  & n13379 ;
  assign n23511 = ~n23509 & ~n23510 ;
  assign n23512 = \wishbone_bd_ram_mem2_reg[196][22]/P0001  & n13977 ;
  assign n23513 = \wishbone_bd_ram_mem2_reg[115][22]/P0001  & n13747 ;
  assign n23514 = ~n23512 & ~n23513 ;
  assign n23515 = n23511 & n23514 ;
  assign n23516 = \wishbone_bd_ram_mem2_reg[11][22]/P0001  & n13774 ;
  assign n23517 = \wishbone_bd_ram_mem2_reg[147][22]/P0001  & n13702 ;
  assign n23518 = ~n23516 & ~n23517 ;
  assign n23519 = \wishbone_bd_ram_mem2_reg[36][22]/P0001  & n13639 ;
  assign n23520 = \wishbone_bd_ram_mem2_reg[87][22]/P0001  & n13691 ;
  assign n23521 = ~n23519 & ~n23520 ;
  assign n23522 = n23518 & n23521 ;
  assign n23523 = n23515 & n23522 ;
  assign n23524 = n23508 & n23523 ;
  assign n23525 = n23493 & n23524 ;
  assign n23526 = \wishbone_bd_ram_mem2_reg[190][22]/P0001  & n13365 ;
  assign n23527 = \wishbone_bd_ram_mem2_reg[22][22]/P0001  & n13744 ;
  assign n23528 = ~n23526 & ~n23527 ;
  assign n23529 = \wishbone_bd_ram_mem2_reg[89][22]/P0001  & n13910 ;
  assign n23530 = \wishbone_bd_ram_mem2_reg[197][22]/P0001  & n13594 ;
  assign n23531 = ~n23529 & ~n23530 ;
  assign n23532 = n23528 & n23531 ;
  assign n23533 = \wishbone_bd_ram_mem2_reg[94][22]/P0001  & n13833 ;
  assign n23534 = \wishbone_bd_ram_mem2_reg[177][22]/P0001  & n13863 ;
  assign n23535 = ~n23533 & ~n23534 ;
  assign n23536 = \wishbone_bd_ram_mem2_reg[155][22]/P0001  & n13738 ;
  assign n23537 = \wishbone_bd_ram_mem2_reg[48][22]/P0001  & n13917 ;
  assign n23538 = ~n23536 & ~n23537 ;
  assign n23539 = n23535 & n23538 ;
  assign n23540 = n23532 & n23539 ;
  assign n23541 = \wishbone_bd_ram_mem2_reg[69][22]/P0001  & n13487 ;
  assign n23542 = \wishbone_bd_ram_mem2_reg[188][22]/P0001  & n13407 ;
  assign n23543 = ~n23541 & ~n23542 ;
  assign n23544 = \wishbone_bd_ram_mem2_reg[118][22]/P0001  & n13589 ;
  assign n23545 = \wishbone_bd_ram_mem2_reg[161][22]/P0001  & n13505 ;
  assign n23546 = ~n23544 & ~n23545 ;
  assign n23547 = n23543 & n23546 ;
  assign n23548 = \wishbone_bd_ram_mem2_reg[39][22]/P0001  & n13893 ;
  assign n23549 = \wishbone_bd_ram_mem2_reg[142][22]/P0001  & n13448 ;
  assign n23550 = ~n23548 & ~n23549 ;
  assign n23551 = \wishbone_bd_ram_mem2_reg[122][22]/P0001  & n13679 ;
  assign n23552 = \wishbone_bd_ram_mem2_reg[83][22]/P0001  & n13454 ;
  assign n23553 = ~n23551 & ~n23552 ;
  assign n23554 = n23550 & n23553 ;
  assign n23555 = n23547 & n23554 ;
  assign n23556 = n23540 & n23555 ;
  assign n23557 = \wishbone_bd_ram_mem2_reg[179][22]/P0001  & n14035 ;
  assign n23558 = \wishbone_bd_ram_mem2_reg[126][22]/P0001  & n13786 ;
  assign n23559 = ~n23557 & ~n23558 ;
  assign n23560 = \wishbone_bd_ram_mem2_reg[7][22]/P0001  & n13546 ;
  assign n23561 = \wishbone_bd_ram_mem2_reg[209][22]/P0001  & n13689 ;
  assign n23562 = ~n23560 & ~n23561 ;
  assign n23563 = n23559 & n23562 ;
  assign n23564 = \wishbone_bd_ram_mem2_reg[120][22]/P0001  & n13550 ;
  assign n23565 = \wishbone_bd_ram_mem2_reg[242][22]/P0001  & n13383 ;
  assign n23566 = ~n23564 & ~n23565 ;
  assign n23567 = \wishbone_bd_ram_mem2_reg[249][22]/P0001  & n13431 ;
  assign n23568 = \wishbone_bd_ram_mem2_reg[223][22]/P0001  & n13335 ;
  assign n23569 = ~n23567 & ~n23568 ;
  assign n23570 = n23566 & n23569 ;
  assign n23571 = n23563 & n23570 ;
  assign n23572 = \wishbone_bd_ram_mem2_reg[240][22]/P0001  & n13352 ;
  assign n23573 = \wishbone_bd_ram_mem2_reg[29][22]/P0001  & n13412 ;
  assign n23574 = ~n23572 & ~n23573 ;
  assign n23575 = \wishbone_bd_ram_mem2_reg[25][22]/P0001  & n13742 ;
  assign n23576 = \wishbone_bd_ram_mem2_reg[124][22]/P0001  & n14024 ;
  assign n23577 = ~n23575 & ~n23576 ;
  assign n23578 = n23574 & n23577 ;
  assign n23579 = \wishbone_bd_ram_mem2_reg[253][22]/P0001  & n13708 ;
  assign n23580 = \wishbone_bd_ram_mem2_reg[84][22]/P0001  & n13385 ;
  assign n23581 = ~n23579 & ~n23580 ;
  assign n23582 = \wishbone_bd_ram_mem2_reg[8][22]/P0001  & n13459 ;
  assign n23583 = \wishbone_bd_ram_mem2_reg[37][22]/P0001  & n13710 ;
  assign n23584 = ~n23582 & ~n23583 ;
  assign n23585 = n23581 & n23584 ;
  assign n23586 = n23578 & n23585 ;
  assign n23587 = n23571 & n23586 ;
  assign n23588 = n23556 & n23587 ;
  assign n23589 = n23525 & n23588 ;
  assign n23590 = \wishbone_bd_ram_mem2_reg[70][22]/P0001  & n13339 ;
  assign n23591 = \wishbone_bd_ram_mem2_reg[129][22]/P0001  & n13629 ;
  assign n23592 = ~n23590 & ~n23591 ;
  assign n23593 = \wishbone_bd_ram_mem2_reg[54][22]/P0001  & n13622 ;
  assign n23594 = \wishbone_bd_ram_mem2_reg[73][22]/P0001  & n13456 ;
  assign n23595 = ~n23593 & ~n23594 ;
  assign n23596 = n23592 & n23595 ;
  assign n23597 = \wishbone_bd_ram_mem2_reg[170][22]/P0001  & n14007 ;
  assign n23598 = \wishbone_bd_ram_mem2_reg[152][22]/P0001  & n13912 ;
  assign n23599 = ~n23597 & ~n23598 ;
  assign n23600 = \wishbone_bd_ram_mem2_reg[62][22]/P0001  & n13529 ;
  assign n23601 = \wishbone_bd_ram_mem2_reg[229][22]/P0001  & n13552 ;
  assign n23602 = ~n23600 & ~n23601 ;
  assign n23603 = n23599 & n23602 ;
  assign n23604 = n23596 & n23603 ;
  assign n23605 = \wishbone_bd_ram_mem2_reg[81][22]/P0001  & n13409 ;
  assign n23606 = \wishbone_bd_ram_mem2_reg[238][22]/P0001  & n13819 ;
  assign n23607 = ~n23605 & ~n23606 ;
  assign n23608 = \wishbone_bd_ram_mem2_reg[28][22]/P0001  & n13810 ;
  assign n23609 = \wishbone_bd_ram_mem2_reg[183][22]/P0001  & n13645 ;
  assign n23610 = ~n23608 & ~n23609 ;
  assign n23611 = n23607 & n23610 ;
  assign n23612 = \wishbone_bd_ram_mem2_reg[163][22]/P0001  & n13255 ;
  assign n23613 = \wishbone_bd_ram_mem2_reg[255][22]/P0001  & n13952 ;
  assign n23614 = ~n23612 & ~n23613 ;
  assign n23615 = \wishbone_bd_ram_mem2_reg[99][22]/P0001  & n13996 ;
  assign n23616 = \wishbone_bd_ram_mem2_reg[119][22]/P0001  & n14033 ;
  assign n23617 = ~n23615 & ~n23616 ;
  assign n23618 = n23614 & n23617 ;
  assign n23619 = n23611 & n23618 ;
  assign n23620 = n23604 & n23619 ;
  assign n23621 = \wishbone_bd_ram_mem2_reg[151][22]/P0001  & n13697 ;
  assign n23622 = \wishbone_bd_ram_mem2_reg[6][22]/P0001  & n13915 ;
  assign n23623 = ~n23621 & ~n23622 ;
  assign n23624 = \wishbone_bd_ram_mem2_reg[230][22]/P0001  & n13994 ;
  assign n23625 = \wishbone_bd_ram_mem2_reg[102][22]/P0001  & n13534 ;
  assign n23626 = ~n23624 & ~n23625 ;
  assign n23627 = n23623 & n23626 ;
  assign n23628 = \wishbone_bd_ram_mem2_reg[192][22]/P0001  & n13390 ;
  assign n23629 = \wishbone_bd_ram_mem2_reg[134][22]/P0001  & n13494 ;
  assign n23630 = ~n23628 & ~n23629 ;
  assign n23631 = \wishbone_bd_ram_mem2_reg[225][22]/P0001  & n13719 ;
  assign n23632 = \wishbone_bd_ram_mem2_reg[91][22]/P0001  & n13954 ;
  assign n23633 = ~n23631 & ~n23632 ;
  assign n23634 = n23630 & n23633 ;
  assign n23635 = n23627 & n23634 ;
  assign n23636 = \wishbone_bd_ram_mem2_reg[224][22]/P0001  & n13433 ;
  assign n23637 = \wishbone_bd_ram_mem2_reg[186][22]/P0001  & n13616 ;
  assign n23638 = ~n23636 & ~n23637 ;
  assign n23639 = \wishbone_bd_ram_mem2_reg[193][22]/P0001  & n14022 ;
  assign n23640 = \wishbone_bd_ram_mem2_reg[78][22]/P0001  & n13277 ;
  assign n23641 = ~n23639 & ~n23640 ;
  assign n23642 = n23638 & n23641 ;
  assign n23643 = \wishbone_bd_ram_mem2_reg[40][22]/P0001  & n13661 ;
  assign n23644 = \wishbone_bd_ram_mem2_reg[65][22]/P0001  & n13842 ;
  assign n23645 = ~n23643 & ~n23644 ;
  assign n23646 = \wishbone_bd_ram_mem2_reg[213][22]/P0001  & n13870 ;
  assign n23647 = \wishbone_bd_ram_mem2_reg[71][22]/P0001  & n13636 ;
  assign n23648 = ~n23646 & ~n23647 ;
  assign n23649 = n23645 & n23648 ;
  assign n23650 = n23642 & n23649 ;
  assign n23651 = n23635 & n23650 ;
  assign n23652 = n23620 & n23651 ;
  assign n23653 = \wishbone_bd_ram_mem2_reg[199][22]/P0001  & n13499 ;
  assign n23654 = \wishbone_bd_ram_mem2_reg[235][22]/P0001  & n13518 ;
  assign n23655 = ~n23653 & ~n23654 ;
  assign n23656 = \wishbone_bd_ram_mem2_reg[185][22]/P0001  & n13372 ;
  assign n23657 = \wishbone_bd_ram_mem2_reg[241][22]/P0001  & n13854 ;
  assign n23658 = ~n23656 & ~n23657 ;
  assign n23659 = n23655 & n23658 ;
  assign n23660 = \wishbone_bd_ram_mem2_reg[92][22]/P0001  & n13859 ;
  assign n23661 = \wishbone_bd_ram_mem2_reg[195][22]/P0001  & n13700 ;
  assign n23662 = ~n23660 & ~n23661 ;
  assign n23663 = \wishbone_bd_ram_mem2_reg[150][22]/P0001  & n13666 ;
  assign n23664 = \wishbone_bd_ram_mem2_reg[211][22]/P0001  & n13805 ;
  assign n23665 = ~n23663 & ~n23664 ;
  assign n23666 = n23662 & n23665 ;
  assign n23667 = n23659 & n23666 ;
  assign n23668 = \wishbone_bd_ram_mem2_reg[13][22]/P0001  & n13844 ;
  assign n23669 = \wishbone_bd_ram_mem2_reg[101][22]/P0001  & n13772 ;
  assign n23670 = ~n23668 & ~n23669 ;
  assign n23671 = \wishbone_bd_ram_mem2_reg[43][22]/P0001  & n13761 ;
  assign n23672 = \wishbone_bd_ram_mem2_reg[110][22]/P0001  & n14030 ;
  assign n23673 = ~n23671 & ~n23672 ;
  assign n23674 = n23670 & n23673 ;
  assign n23675 = \wishbone_bd_ram_mem2_reg[227][22]/P0001  & n13388 ;
  assign n23676 = \wishbone_bd_ram_mem2_reg[182][22]/P0001  & n13598 ;
  assign n23677 = ~n23675 & ~n23676 ;
  assign n23678 = \wishbone_bd_ram_mem2_reg[219][22]/P0001  & n13577 ;
  assign n23679 = \wishbone_bd_ram_mem2_reg[3][22]/P0001  & n13354 ;
  assign n23680 = ~n23678 & ~n23679 ;
  assign n23681 = n23677 & n23680 ;
  assign n23682 = n23674 & n23681 ;
  assign n23683 = n23667 & n23682 ;
  assign n23684 = \wishbone_bd_ram_mem2_reg[231][22]/P0001  & n13363 ;
  assign n23685 = \wishbone_bd_ram_mem2_reg[123][22]/P0001  & n13749 ;
  assign n23686 = ~n23684 & ~n23685 ;
  assign n23687 = \wishbone_bd_ram_mem2_reg[171][22]/P0001  & n13422 ;
  assign n23688 = \wishbone_bd_ram_mem2_reg[103][22]/P0001  & n13320 ;
  assign n23689 = ~n23687 & ~n23688 ;
  assign n23690 = n23686 & n23689 ;
  assign n23691 = \wishbone_bd_ram_mem2_reg[245][22]/P0001  & n13877 ;
  assign n23692 = \wishbone_bd_ram_mem2_reg[236][22]/P0001  & n13480 ;
  assign n23693 = ~n23691 & ~n23692 ;
  assign n23694 = \wishbone_bd_ram_mem2_reg[218][22]/P0001  & n13792 ;
  assign n23695 = \wishbone_bd_ram_mem2_reg[162][22]/P0001  & n13726 ;
  assign n23696 = ~n23694 & ~n23695 ;
  assign n23697 = n23693 & n23696 ;
  assign n23698 = n23690 & n23697 ;
  assign n23699 = \wishbone_bd_ram_mem2_reg[46][22]/P0001  & n13298 ;
  assign n23700 = \wishbone_bd_ram_mem2_reg[178][22]/P0001  & n13301 ;
  assign n23701 = ~n23699 & ~n23700 ;
  assign n23702 = \wishbone_bd_ram_mem2_reg[198][22]/P0001  & n13592 ;
  assign n23703 = \wishbone_bd_ram_mem2_reg[132][22]/P0001  & n13927 ;
  assign n23704 = ~n23702 & ~n23703 ;
  assign n23705 = n23701 & n23704 ;
  assign n23706 = \wishbone_bd_ram_mem2_reg[93][22]/P0001  & n13891 ;
  assign n23707 = \wishbone_bd_ram_mem2_reg[158][22]/P0001  & n13294 ;
  assign n23708 = ~n23706 & ~n23707 ;
  assign n23709 = \wishbone_bd_ram_mem2_reg[33][22]/P0001  & n13933 ;
  assign n23710 = \wishbone_bd_ram_mem2_reg[205][22]/P0001  & n13947 ;
  assign n23711 = ~n23709 & ~n23710 ;
  assign n23712 = n23708 & n23711 ;
  assign n23713 = n23705 & n23712 ;
  assign n23714 = n23698 & n23713 ;
  assign n23715 = n23683 & n23714 ;
  assign n23716 = n23652 & n23715 ;
  assign n23717 = n23589 & n23716 ;
  assign n23718 = n23462 & n23717 ;
  assign n23719 = n14047 & ~n23718 ;
  assign n23720 = ~n23207 & ~n23719 ;
  assign n23721 = \wishbone_LatchedTxLength_reg[9]/NET0131  & ~n14046 ;
  assign n23722 = ~n18435 & ~n23721 ;
  assign n23723 = ~\wb_sel_i[0]_pad  & ~\wb_sel_i[1]_pad  ;
  assign n23724 = ~\wb_sel_i[2]_pad  & ~\wb_sel_i[3]_pad  ;
  assign n23725 = n23723 & n23724 ;
  assign n23726 = wb_cyc_i_pad & wb_stb_i_pad ;
  assign n23727 = ~\wb_adr_i[10]_pad  & ~\wb_adr_i[11]_pad  ;
  assign n23728 = n23726 & n23727 ;
  assign n23729 = ~n23725 & n23728 ;
  assign n23730 = ~wb_we_i_pad & n23729 ;
  assign n23731 = ~\wb_adr_i[7]_pad  & ~\wb_adr_i[9]_pad  ;
  assign n23732 = ~\wb_adr_i[6]_pad  & ~\wb_adr_i[8]_pad  ;
  assign n23733 = n23731 & n23732 ;
  assign n23734 = ~\wb_adr_i[2]_pad  & \wb_adr_i[3]_pad  ;
  assign n23735 = \wb_adr_i[4]_pad  & ~\wb_adr_i[5]_pad  ;
  assign n23736 = n23734 & n23735 ;
  assign n23737 = n23733 & n23736 ;
  assign n23738 = \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  & n23737 ;
  assign n23739 = \wb_adr_i[6]_pad  & n23731 ;
  assign n23740 = ~\wb_adr_i[2]_pad  & ~\wb_adr_i[8]_pad  ;
  assign n23741 = n23739 & n23740 ;
  assign n23742 = ~\wb_adr_i[4]_pad  & ~\wb_adr_i[5]_pad  ;
  assign n23743 = \wb_adr_i[3]_pad  & n23742 ;
  assign n23744 = \ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131  & n23743 ;
  assign n23745 = n23741 & n23744 ;
  assign n23746 = \wb_adr_i[2]_pad  & ~\wb_adr_i[8]_pad  ;
  assign n23747 = n23739 & n23746 ;
  assign n23748 = \ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131  & n23743 ;
  assign n23749 = n23747 & n23748 ;
  assign n23750 = ~n23745 & ~n23749 ;
  assign n23751 = ~\wb_adr_i[3]_pad  & n23742 ;
  assign n23752 = \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  & n23751 ;
  assign n23753 = n23741 & n23752 ;
  assign n23754 = n23730 & ~n23753 ;
  assign n23755 = n23750 & n23754 ;
  assign n23756 = ~n23738 & n23755 ;
  assign n23757 = n23730 & ~n23756 ;
  assign n23758 = ~wb_rst_i_pad & ~n23756 ;
  assign n23759 = ~n22688 & n23758 ;
  assign n23760 = ~n23757 & ~n23759 ;
  assign n23761 = \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  & n23737 ;
  assign n23762 = \ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131  & n23743 ;
  assign n23763 = n23741 & n23762 ;
  assign n23764 = \ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131  & n23743 ;
  assign n23765 = n23747 & n23764 ;
  assign n23766 = ~n23763 & ~n23765 ;
  assign n23767 = \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  & n23751 ;
  assign n23768 = n23741 & n23767 ;
  assign n23769 = n23730 & ~n23768 ;
  assign n23770 = n23766 & n23769 ;
  assign n23771 = ~n23761 & n23770 ;
  assign n23772 = n23730 & ~n23771 ;
  assign n23773 = ~wb_rst_i_pad & ~n23771 ;
  assign n23774 = ~n23718 & n23773 ;
  assign n23775 = ~n23772 & ~n23774 ;
  assign n23776 = \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  & n23751 ;
  assign n23777 = n23747 & n23776 ;
  assign n23778 = \wb_adr_i[4]_pad  & ~\wb_adr_i[6]_pad  ;
  assign n23779 = n23740 & n23778 ;
  assign n23780 = \wb_adr_i[3]_pad  & \wb_adr_i[5]_pad  ;
  assign n23781 = n23731 & n23780 ;
  assign n23782 = n23779 & n23781 ;
  assign n23783 = \ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131  & n23782 ;
  assign n23784 = ~n23777 & ~n23783 ;
  assign n23785 = \ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131  & n23743 ;
  assign n23786 = n23741 & n23785 ;
  assign n23787 = \ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131  & n23743 ;
  assign n23788 = n23747 & n23787 ;
  assign n23789 = ~n23786 & ~n23788 ;
  assign n23790 = n23784 & n23789 ;
  assign n23791 = \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  & n23751 ;
  assign n23792 = n23741 & n23791 ;
  assign n23793 = ~\wb_adr_i[3]_pad  & \wb_adr_i[4]_pad  ;
  assign n23794 = ~\wb_adr_i[5]_pad  & n23793 ;
  assign n23795 = \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131  & n23794 ;
  assign n23796 = n23741 & n23795 ;
  assign n23797 = ~n23792 & ~n23796 ;
  assign n23798 = n23730 & n23797 ;
  assign n23799 = n23790 & n23798 ;
  assign n23800 = ~\wb_adr_i[3]_pad  & \wb_adr_i[5]_pad  ;
  assign n23801 = n23731 & n23800 ;
  assign n23802 = n23779 & n23801 ;
  assign n23803 = \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131  & n23802 ;
  assign n23804 = ~\wb_adr_i[3]_pad  & ~\wb_adr_i[5]_pad  ;
  assign n23805 = n23731 & n23804 ;
  assign n23806 = ~\wb_adr_i[4]_pad  & ~\wb_adr_i[6]_pad  ;
  assign n23807 = n23740 & n23806 ;
  assign n23808 = n23805 & n23807 ;
  assign n23809 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & n23808 ;
  assign n23810 = ~n23803 & ~n23809 ;
  assign n23811 = \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  & n23737 ;
  assign n23812 = n23746 & n23778 ;
  assign n23813 = n23801 & n23812 ;
  assign n23814 = \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131  & n23813 ;
  assign n23815 = ~n23811 & ~n23814 ;
  assign n23816 = n23810 & n23815 ;
  assign n23817 = n23799 & n23816 ;
  assign n23818 = n23730 & ~n23817 ;
  assign n23819 = \wishbone_bd_ram_mem1_reg[43][12]/P0001  & n13761 ;
  assign n23820 = \wishbone_bd_ram_mem1_reg[135][12]/P0001  & n13672 ;
  assign n23821 = ~n23819 & ~n23820 ;
  assign n23822 = \wishbone_bd_ram_mem1_reg[103][12]/P0001  & n13320 ;
  assign n23823 = \wishbone_bd_ram_mem1_reg[219][12]/P0001  & n13577 ;
  assign n23824 = ~n23822 & ~n23823 ;
  assign n23825 = n23821 & n23824 ;
  assign n23826 = \wishbone_bd_ram_mem1_reg[82][12]/P0001  & n13374 ;
  assign n23827 = \wishbone_bd_ram_mem1_reg[55][12]/P0001  & n13618 ;
  assign n23828 = ~n23826 & ~n23827 ;
  assign n23829 = \wishbone_bd_ram_mem1_reg[205][12]/P0001  & n13947 ;
  assign n23830 = \wishbone_bd_ram_mem1_reg[175][12]/P0001  & n13674 ;
  assign n23831 = ~n23829 & ~n23830 ;
  assign n23832 = n23828 & n23831 ;
  assign n23833 = n23825 & n23832 ;
  assign n23834 = \wishbone_bd_ram_mem1_reg[252][12]/P0001  & n13986 ;
  assign n23835 = \wishbone_bd_ram_mem1_reg[180][12]/P0001  & n13650 ;
  assign n23836 = ~n23834 & ~n23835 ;
  assign n23837 = \wishbone_bd_ram_mem1_reg[1][12]/P0001  & n13888 ;
  assign n23838 = \wishbone_bd_ram_mem1_reg[31][12]/P0001  & n13758 ;
  assign n23839 = ~n23837 & ~n23838 ;
  assign n23840 = n23836 & n23839 ;
  assign n23841 = \wishbone_bd_ram_mem1_reg[112][12]/P0001  & n13482 ;
  assign n23842 = \wishbone_bd_ram_mem1_reg[249][12]/P0001  & n13431 ;
  assign n23843 = ~n23841 & ~n23842 ;
  assign n23844 = \wishbone_bd_ram_mem1_reg[201][12]/P0001  & n13600 ;
  assign n23845 = \wishbone_bd_ram_mem1_reg[47][12]/P0001  & n13436 ;
  assign n23846 = ~n23844 & ~n23845 ;
  assign n23847 = n23843 & n23846 ;
  assign n23848 = n23840 & n23847 ;
  assign n23849 = n23833 & n23848 ;
  assign n23850 = \wishbone_bd_ram_mem1_reg[118][12]/P0001  & n13589 ;
  assign n23851 = \wishbone_bd_ram_mem1_reg[231][12]/P0001  & n13363 ;
  assign n23852 = ~n23850 & ~n23851 ;
  assign n23853 = \wishbone_bd_ram_mem1_reg[121][12]/P0001  & n13983 ;
  assign n23854 = \wishbone_bd_ram_mem1_reg[229][12]/P0001  & n13552 ;
  assign n23855 = ~n23853 & ~n23854 ;
  assign n23856 = n23852 & n23855 ;
  assign n23857 = \wishbone_bd_ram_mem1_reg[193][12]/P0001  & n14022 ;
  assign n23858 = \wishbone_bd_ram_mem1_reg[126][12]/P0001  & n13786 ;
  assign n23859 = ~n23857 & ~n23858 ;
  assign n23860 = \wishbone_bd_ram_mem1_reg[35][12]/P0001  & n13523 ;
  assign n23861 = \wishbone_bd_ram_mem1_reg[191][12]/P0001  & n14012 ;
  assign n23862 = ~n23860 & ~n23861 ;
  assign n23863 = n23859 & n23862 ;
  assign n23864 = n23856 & n23863 ;
  assign n23865 = \wishbone_bd_ram_mem1_reg[104][12]/P0001  & n13684 ;
  assign n23866 = \wishbone_bd_ram_mem1_reg[248][12]/P0001  & n13647 ;
  assign n23867 = ~n23865 & ~n23866 ;
  assign n23868 = \wishbone_bd_ram_mem1_reg[241][12]/P0001  & n13854 ;
  assign n23869 = \wishbone_bd_ram_mem1_reg[127][12]/P0001  & n13803 ;
  assign n23870 = ~n23868 & ~n23869 ;
  assign n23871 = n23867 & n23870 ;
  assign n23872 = \wishbone_bd_ram_mem1_reg[144][12]/P0001  & n13508 ;
  assign n23873 = \wishbone_bd_ram_mem1_reg[49][12]/P0001  & n13929 ;
  assign n23874 = ~n23872 & ~n23873 ;
  assign n23875 = \wishbone_bd_ram_mem1_reg[220][12]/P0001  & n13965 ;
  assign n23876 = \wishbone_bd_ram_mem1_reg[210][12]/P0001  & n13443 ;
  assign n23877 = ~n23875 & ~n23876 ;
  assign n23878 = n23874 & n23877 ;
  assign n23879 = n23871 & n23878 ;
  assign n23880 = n23864 & n23879 ;
  assign n23881 = n23849 & n23880 ;
  assign n23882 = \wishbone_bd_ram_mem1_reg[8][12]/P0001  & n13459 ;
  assign n23883 = \wishbone_bd_ram_mem1_reg[245][12]/P0001  & n13877 ;
  assign n23884 = ~n23882 & ~n23883 ;
  assign n23885 = \wishbone_bd_ram_mem1_reg[105][12]/P0001  & n13503 ;
  assign n23886 = \wishbone_bd_ram_mem1_reg[106][12]/P0001  & n13555 ;
  assign n23887 = ~n23885 & ~n23886 ;
  assign n23888 = n23884 & n23887 ;
  assign n23889 = \wishbone_bd_ram_mem1_reg[243][12]/P0001  & n13575 ;
  assign n23890 = \wishbone_bd_ram_mem1_reg[96][12]/P0001  & n13425 ;
  assign n23891 = ~n23889 & ~n23890 ;
  assign n23892 = \wishbone_bd_ram_mem1_reg[239][12]/P0001  & n13349 ;
  assign n23893 = \wishbone_bd_ram_mem1_reg[7][12]/P0001  & n13546 ;
  assign n23894 = ~n23892 & ~n23893 ;
  assign n23895 = n23891 & n23894 ;
  assign n23896 = n23888 & n23895 ;
  assign n23897 = \wishbone_bd_ram_mem1_reg[230][12]/P0001  & n13994 ;
  assign n23898 = \wishbone_bd_ram_mem1_reg[158][12]/P0001  & n13294 ;
  assign n23899 = ~n23897 & ~n23898 ;
  assign n23900 = \wishbone_bd_ram_mem1_reg[187][12]/P0001  & n13756 ;
  assign n23901 = \wishbone_bd_ram_mem1_reg[54][12]/P0001  & n13622 ;
  assign n23902 = ~n23900 & ~n23901 ;
  assign n23903 = n23899 & n23902 ;
  assign n23904 = \wishbone_bd_ram_mem1_reg[129][12]/P0001  & n13629 ;
  assign n23905 = \wishbone_bd_ram_mem1_reg[215][12]/P0001  & n13901 ;
  assign n23906 = ~n23904 & ~n23905 ;
  assign n23907 = \wishbone_bd_ram_mem1_reg[52][12]/P0001  & n13988 ;
  assign n23908 = \wishbone_bd_ram_mem1_reg[147][12]/P0001  & n13702 ;
  assign n23909 = ~n23907 & ~n23908 ;
  assign n23910 = n23906 & n23909 ;
  assign n23911 = n23903 & n23910 ;
  assign n23912 = n23896 & n23911 ;
  assign n23913 = \wishbone_bd_ram_mem1_reg[216][12]/P0001  & n14005 ;
  assign n23914 = \wishbone_bd_ram_mem1_reg[174][12]/P0001  & n13899 ;
  assign n23915 = ~n23913 & ~n23914 ;
  assign n23916 = \wishbone_bd_ram_mem1_reg[77][12]/P0001  & n13935 ;
  assign n23917 = \wishbone_bd_ram_mem1_reg[120][12]/P0001  & n13550 ;
  assign n23918 = ~n23916 & ~n23917 ;
  assign n23919 = n23915 & n23918 ;
  assign n23920 = \wishbone_bd_ram_mem1_reg[227][12]/P0001  & n13388 ;
  assign n23921 = \wishbone_bd_ram_mem1_reg[199][12]/P0001  & n13499 ;
  assign n23922 = ~n23920 & ~n23921 ;
  assign n23923 = \wishbone_bd_ram_mem1_reg[244][12]/P0001  & n13474 ;
  assign n23924 = \wishbone_bd_ram_mem1_reg[26][12]/P0001  & n13521 ;
  assign n23925 = ~n23923 & ~n23924 ;
  assign n23926 = n23922 & n23925 ;
  assign n23927 = n23919 & n23926 ;
  assign n23928 = \wishbone_bd_ram_mem1_reg[155][12]/P0001  & n13738 ;
  assign n23929 = \wishbone_bd_ram_mem1_reg[27][12]/P0001  & n13251 ;
  assign n23930 = ~n23928 & ~n23929 ;
  assign n23931 = \wishbone_bd_ram_mem1_reg[111][12]/P0001  & n13471 ;
  assign n23932 = \wishbone_bd_ram_mem1_reg[225][12]/P0001  & n13719 ;
  assign n23933 = ~n23931 & ~n23932 ;
  assign n23934 = n23930 & n23933 ;
  assign n23935 = \wishbone_bd_ram_mem1_reg[217][12]/P0001  & n13767 ;
  assign n23936 = \wishbone_bd_ram_mem1_reg[234][12]/P0001  & n13781 ;
  assign n23937 = ~n23935 & ~n23936 ;
  assign n23938 = \wishbone_bd_ram_mem1_reg[5][12]/P0001  & n13243 ;
  assign n23939 = \wishbone_bd_ram_mem1_reg[62][12]/P0001  & n13529 ;
  assign n23940 = ~n23938 & ~n23939 ;
  assign n23941 = n23937 & n23940 ;
  assign n23942 = n23934 & n23941 ;
  assign n23943 = n23927 & n23942 ;
  assign n23944 = n23912 & n23943 ;
  assign n23945 = n23881 & n23944 ;
  assign n23946 = \wishbone_bd_ram_mem1_reg[33][12]/P0001  & n13933 ;
  assign n23947 = \wishbone_bd_ram_mem1_reg[238][12]/P0001  & n13819 ;
  assign n23948 = ~n23946 & ~n23947 ;
  assign n23949 = \wishbone_bd_ram_mem1_reg[153][12]/P0001  & n13309 ;
  assign n23950 = \wishbone_bd_ram_mem1_reg[24][12]/P0001  & n13970 ;
  assign n23951 = ~n23949 & ~n23950 ;
  assign n23952 = n23948 & n23951 ;
  assign n23953 = \wishbone_bd_ram_mem1_reg[212][12]/P0001  & n13634 ;
  assign n23954 = \wishbone_bd_ram_mem1_reg[59][12]/P0001  & n13613 ;
  assign n23955 = ~n23953 & ~n23954 ;
  assign n23956 = \wishbone_bd_ram_mem1_reg[85][12]/P0001  & n13784 ;
  assign n23957 = \wishbone_bd_ram_mem1_reg[90][12]/P0001  & n13906 ;
  assign n23958 = ~n23956 & ~n23957 ;
  assign n23959 = n23955 & n23958 ;
  assign n23960 = n23952 & n23959 ;
  assign n23961 = \wishbone_bd_ram_mem1_reg[139][12]/P0001  & n13566 ;
  assign n23962 = \wishbone_bd_ram_mem1_reg[97][12]/P0001  & n13724 ;
  assign n23963 = ~n23961 & ~n23962 ;
  assign n23964 = \wishbone_bd_ram_mem1_reg[232][12]/P0001  & n13510 ;
  assign n23965 = \wishbone_bd_ram_mem1_reg[223][12]/P0001  & n13335 ;
  assign n23966 = ~n23964 & ~n23965 ;
  assign n23967 = n23963 & n23966 ;
  assign n23968 = \wishbone_bd_ram_mem1_reg[165][12]/P0001  & n14028 ;
  assign n23969 = \wishbone_bd_ram_mem1_reg[146][12]/P0001  & n13958 ;
  assign n23970 = ~n23968 & ~n23969 ;
  assign n23971 = \wishbone_bd_ram_mem1_reg[128][12]/P0001  & n13652 ;
  assign n23972 = \wishbone_bd_ram_mem1_reg[28][12]/P0001  & n13810 ;
  assign n23973 = ~n23971 & ~n23972 ;
  assign n23974 = n23970 & n23973 ;
  assign n23975 = n23967 & n23974 ;
  assign n23976 = n23960 & n23975 ;
  assign n23977 = \wishbone_bd_ram_mem1_reg[236][12]/P0001  & n13480 ;
  assign n23978 = \wishbone_bd_ram_mem1_reg[86][12]/P0001  & n13485 ;
  assign n23979 = ~n23977 & ~n23978 ;
  assign n23980 = \wishbone_bd_ram_mem1_reg[161][12]/P0001  & n13505 ;
  assign n23981 = \wishbone_bd_ram_mem1_reg[117][12]/P0001  & n13557 ;
  assign n23982 = ~n23980 & ~n23981 ;
  assign n23983 = n23979 & n23982 ;
  assign n23984 = \wishbone_bd_ram_mem1_reg[17][12]/P0001  & n13324 ;
  assign n23985 = \wishbone_bd_ram_mem1_reg[95][12]/P0001  & n13317 ;
  assign n23986 = ~n23984 & ~n23985 ;
  assign n23987 = \wishbone_bd_ram_mem1_reg[189][12]/P0001  & n14001 ;
  assign n23988 = \wishbone_bd_ram_mem1_reg[145][12]/P0001  & n13715 ;
  assign n23989 = ~n23987 & ~n23988 ;
  assign n23990 = n23986 & n23989 ;
  assign n23991 = n23983 & n23990 ;
  assign n23992 = \wishbone_bd_ram_mem1_reg[13][12]/P0001  & n13844 ;
  assign n23993 = \wishbone_bd_ram_mem1_reg[83][12]/P0001  & n13454 ;
  assign n23994 = ~n23992 & ~n23993 ;
  assign n23995 = \wishbone_bd_ram_mem1_reg[125][12]/P0001  & n13396 ;
  assign n23996 = \wishbone_bd_ram_mem1_reg[22][12]/P0001  & n13744 ;
  assign n23997 = ~n23995 & ~n23996 ;
  assign n23998 = n23994 & n23997 ;
  assign n23999 = \wishbone_bd_ram_mem1_reg[211][12]/P0001  & n13805 ;
  assign n24000 = \wishbone_bd_ram_mem1_reg[194][12]/P0001  & n13624 ;
  assign n24001 = ~n23999 & ~n24000 ;
  assign n24002 = \wishbone_bd_ram_mem1_reg[166][12]/P0001  & n13999 ;
  assign n24003 = \wishbone_bd_ram_mem1_reg[208][12]/P0001  & n14010 ;
  assign n24004 = ~n24002 & ~n24003 ;
  assign n24005 = n24001 & n24004 ;
  assign n24006 = n23998 & n24005 ;
  assign n24007 = n23991 & n24006 ;
  assign n24008 = n23976 & n24007 ;
  assign n24009 = \wishbone_bd_ram_mem1_reg[76][12]/P0001  & n13831 ;
  assign n24010 = \wishbone_bd_ram_mem1_reg[233][12]/P0001  & n13332 ;
  assign n24011 = ~n24009 & ~n24010 ;
  assign n24012 = \wishbone_bd_ram_mem1_reg[200][12]/P0001  & n13922 ;
  assign n24013 = \wishbone_bd_ram_mem1_reg[242][12]/P0001  & n13383 ;
  assign n24014 = ~n24012 & ~n24013 ;
  assign n24015 = n24011 & n24014 ;
  assign n24016 = \wishbone_bd_ram_mem1_reg[141][12]/P0001  & n13852 ;
  assign n24017 = \wishbone_bd_ram_mem1_reg[169][12]/P0001  & n13541 ;
  assign n24018 = ~n24016 & ~n24017 ;
  assign n24019 = \wishbone_bd_ram_mem1_reg[4][12]/P0001  & n13527 ;
  assign n24020 = \wishbone_bd_ram_mem1_reg[78][12]/P0001  & n13277 ;
  assign n24021 = ~n24019 & ~n24020 ;
  assign n24022 = n24018 & n24021 ;
  assign n24023 = n24015 & n24022 ;
  assign n24024 = \wishbone_bd_ram_mem1_reg[218][12]/P0001  & n13792 ;
  assign n24025 = \wishbone_bd_ram_mem1_reg[57][12]/P0001  & n13731 ;
  assign n24026 = ~n24024 & ~n24025 ;
  assign n24027 = \wishbone_bd_ram_mem1_reg[134][12]/P0001  & n13494 ;
  assign n24028 = \wishbone_bd_ram_mem1_reg[183][12]/P0001  & n13645 ;
  assign n24029 = ~n24027 & ~n24028 ;
  assign n24030 = n24026 & n24029 ;
  assign n24031 = \wishbone_bd_ram_mem1_reg[247][12]/P0001  & n13571 ;
  assign n24032 = \wishbone_bd_ram_mem1_reg[240][12]/P0001  & n13352 ;
  assign n24033 = ~n24031 & ~n24032 ;
  assign n24034 = \wishbone_bd_ram_mem1_reg[6][12]/P0001  & n13915 ;
  assign n24035 = \wishbone_bd_ram_mem1_reg[81][12]/P0001  & n13409 ;
  assign n24036 = ~n24034 & ~n24035 ;
  assign n24037 = n24033 & n24036 ;
  assign n24038 = n24030 & n24037 ;
  assign n24039 = n24023 & n24038 ;
  assign n24040 = \wishbone_bd_ram_mem1_reg[20][12]/P0001  & n13839 ;
  assign n24041 = \wishbone_bd_ram_mem1_reg[123][12]/P0001  & n13749 ;
  assign n24042 = ~n24040 & ~n24041 ;
  assign n24043 = \wishbone_bd_ram_mem1_reg[63][12]/P0001  & n13327 ;
  assign n24044 = \wishbone_bd_ram_mem1_reg[196][12]/P0001  & n13977 ;
  assign n24045 = ~n24043 & ~n24044 ;
  assign n24046 = n24042 & n24045 ;
  assign n24047 = \wishbone_bd_ram_mem1_reg[250][12]/P0001  & n13677 ;
  assign n24048 = \wishbone_bd_ram_mem1_reg[23][12]/P0001  & n13857 ;
  assign n24049 = ~n24047 & ~n24048 ;
  assign n24050 = \wishbone_bd_ram_mem1_reg[66][12]/P0001  & n13603 ;
  assign n24051 = \wishbone_bd_ram_mem1_reg[116][12]/P0001  & n13865 ;
  assign n24052 = ~n24050 & ~n24051 ;
  assign n24053 = n24049 & n24052 ;
  assign n24054 = n24046 & n24053 ;
  assign n24055 = \wishbone_bd_ram_mem1_reg[235][12]/P0001  & n13518 ;
  assign n24056 = \wishbone_bd_ram_mem1_reg[124][12]/P0001  & n14024 ;
  assign n24057 = ~n24055 & ~n24056 ;
  assign n24058 = \wishbone_bd_ram_mem1_reg[110][12]/P0001  & n14030 ;
  assign n24059 = \wishbone_bd_ram_mem1_reg[181][12]/P0001  & n13587 ;
  assign n24060 = ~n24058 & ~n24059 ;
  assign n24061 = n24057 & n24060 ;
  assign n24062 = \wishbone_bd_ram_mem1_reg[38][12]/P0001  & n13828 ;
  assign n24063 = \wishbone_bd_ram_mem1_reg[202][12]/P0001  & n13268 ;
  assign n24064 = ~n24062 & ~n24063 ;
  assign n24065 = \wishbone_bd_ram_mem1_reg[131][12]/P0001  & n13358 ;
  assign n24066 = \wishbone_bd_ram_mem1_reg[29][12]/P0001  & n13412 ;
  assign n24067 = ~n24065 & ~n24066 ;
  assign n24068 = n24064 & n24067 ;
  assign n24069 = n24061 & n24068 ;
  assign n24070 = n24054 & n24069 ;
  assign n24071 = n24039 & n24070 ;
  assign n24072 = n24008 & n24071 ;
  assign n24073 = n23945 & n24072 ;
  assign n24074 = \wishbone_bd_ram_mem1_reg[108][12]/P0001  & n13814 ;
  assign n24075 = \wishbone_bd_ram_mem1_reg[69][12]/P0001  & n13487 ;
  assign n24076 = ~n24074 & ~n24075 ;
  assign n24077 = \wishbone_bd_ram_mem1_reg[41][12]/P0001  & n14017 ;
  assign n24078 = \wishbone_bd_ram_mem1_reg[207][12]/P0001  & n13826 ;
  assign n24079 = ~n24077 & ~n24078 ;
  assign n24080 = n24076 & n24079 ;
  assign n24081 = \wishbone_bd_ram_mem1_reg[177][12]/P0001  & n13863 ;
  assign n24082 = \wishbone_bd_ram_mem1_reg[89][12]/P0001  & n13910 ;
  assign n24083 = ~n24081 & ~n24082 ;
  assign n24084 = \wishbone_bd_ram_mem1_reg[154][12]/P0001  & n13403 ;
  assign n24085 = \wishbone_bd_ram_mem1_reg[101][12]/P0001  & n13772 ;
  assign n24086 = ~n24084 & ~n24085 ;
  assign n24087 = n24083 & n24086 ;
  assign n24088 = n24080 & n24087 ;
  assign n24089 = \wishbone_bd_ram_mem1_reg[164][12]/P0001  & n13236 ;
  assign n24090 = \wishbone_bd_ram_mem1_reg[149][12]/P0001  & n13469 ;
  assign n24091 = ~n24089 & ~n24090 ;
  assign n24092 = \wishbone_bd_ram_mem1_reg[58][12]/P0001  & n13949 ;
  assign n24093 = \wishbone_bd_ram_mem1_reg[162][12]/P0001  & n13726 ;
  assign n24094 = ~n24092 & ~n24093 ;
  assign n24095 = n24091 & n24094 ;
  assign n24096 = \wishbone_bd_ram_mem1_reg[60][12]/P0001  & n13790 ;
  assign n24097 = \wishbone_bd_ram_mem1_reg[18][12]/P0001  & n13532 ;
  assign n24098 = ~n24096 & ~n24097 ;
  assign n24099 = \wishbone_bd_ram_mem1_reg[10][12]/P0001  & n13837 ;
  assign n24100 = \wishbone_bd_ram_mem1_reg[206][12]/P0001  & n13414 ;
  assign n24101 = ~n24099 & ~n24100 ;
  assign n24102 = n24098 & n24101 ;
  assign n24103 = n24095 & n24102 ;
  assign n24104 = n24088 & n24103 ;
  assign n24105 = \wishbone_bd_ram_mem1_reg[142][12]/P0001  & n13448 ;
  assign n24106 = \wishbone_bd_ram_mem1_reg[204][12]/P0001  & n13821 ;
  assign n24107 = ~n24105 & ~n24106 ;
  assign n24108 = \wishbone_bd_ram_mem1_reg[12][12]/P0001  & n13733 ;
  assign n24109 = \wishbone_bd_ram_mem1_reg[143][12]/P0001  & n13461 ;
  assign n24110 = ~n24108 & ~n24109 ;
  assign n24111 = n24107 & n24110 ;
  assign n24112 = \wishbone_bd_ram_mem1_reg[190][12]/P0001  & n13365 ;
  assign n24113 = \wishbone_bd_ram_mem1_reg[198][12]/P0001  & n13592 ;
  assign n24114 = ~n24112 & ~n24113 ;
  assign n24115 = \wishbone_bd_ram_mem1_reg[122][12]/P0001  & n13679 ;
  assign n24116 = \wishbone_bd_ram_mem1_reg[92][12]/P0001  & n13859 ;
  assign n24117 = ~n24115 & ~n24116 ;
  assign n24118 = n24114 & n24117 ;
  assign n24119 = n24111 & n24118 ;
  assign n24120 = \wishbone_bd_ram_mem1_reg[119][12]/P0001  & n14033 ;
  assign n24121 = \wishbone_bd_ram_mem1_reg[64][12]/P0001  & n13904 ;
  assign n24122 = ~n24120 & ~n24121 ;
  assign n24123 = \wishbone_bd_ram_mem1_reg[25][12]/P0001  & n13742 ;
  assign n24124 = \wishbone_bd_ram_mem1_reg[188][12]/P0001  & n13407 ;
  assign n24125 = ~n24123 & ~n24124 ;
  assign n24126 = n24122 & n24125 ;
  assign n24127 = \wishbone_bd_ram_mem1_reg[132][12]/P0001  & n13927 ;
  assign n24128 = \wishbone_bd_ram_mem1_reg[167][12]/P0001  & n13940 ;
  assign n24129 = ~n24127 & ~n24128 ;
  assign n24130 = \wishbone_bd_ram_mem1_reg[19][12]/P0001  & n13886 ;
  assign n24131 = \wishbone_bd_ram_mem1_reg[115][12]/P0001  & n13747 ;
  assign n24132 = ~n24130 & ~n24131 ;
  assign n24133 = n24129 & n24132 ;
  assign n24134 = n24126 & n24133 ;
  assign n24135 = n24119 & n24134 ;
  assign n24136 = n24104 & n24135 ;
  assign n24137 = \wishbone_bd_ram_mem1_reg[14][12]/P0001  & n13972 ;
  assign n24138 = \wishbone_bd_ram_mem1_reg[163][12]/P0001  & n13255 ;
  assign n24139 = ~n24137 & ~n24138 ;
  assign n24140 = \wishbone_bd_ram_mem1_reg[173][12]/P0001  & n13360 ;
  assign n24141 = \wishbone_bd_ram_mem1_reg[192][12]/P0001  & n13390 ;
  assign n24142 = ~n24140 & ~n24141 ;
  assign n24143 = n24139 & n24142 ;
  assign n24144 = \wishbone_bd_ram_mem1_reg[70][12]/P0001  & n13339 ;
  assign n24145 = \wishbone_bd_ram_mem1_reg[148][12]/P0001  & n13868 ;
  assign n24146 = ~n24144 & ~n24145 ;
  assign n24147 = \wishbone_bd_ram_mem1_reg[138][12]/P0001  & n13398 ;
  assign n24148 = \wishbone_bd_ram_mem1_reg[109][12]/P0001  & n13306 ;
  assign n24149 = ~n24147 & ~n24148 ;
  assign n24150 = n24146 & n24149 ;
  assign n24151 = n24143 & n24150 ;
  assign n24152 = \wishbone_bd_ram_mem1_reg[209][12]/P0001  & n13689 ;
  assign n24153 = \wishbone_bd_ram_mem1_reg[176][12]/P0001  & n13262 ;
  assign n24154 = ~n24152 & ~n24153 ;
  assign n24155 = \wishbone_bd_ram_mem1_reg[65][12]/P0001  & n13842 ;
  assign n24156 = \wishbone_bd_ram_mem1_reg[151][12]/P0001  & n13697 ;
  assign n24157 = ~n24155 & ~n24156 ;
  assign n24158 = n24154 & n24157 ;
  assign n24159 = \wishbone_bd_ram_mem1_reg[185][12]/P0001  & n13372 ;
  assign n24160 = \wishbone_bd_ram_mem1_reg[36][12]/P0001  & n13639 ;
  assign n24161 = ~n24159 & ~n24160 ;
  assign n24162 = \wishbone_bd_ram_mem1_reg[73][12]/P0001  & n13456 ;
  assign n24163 = \wishbone_bd_ram_mem1_reg[136][12]/P0001  & n13963 ;
  assign n24164 = ~n24162 & ~n24163 ;
  assign n24165 = n24161 & n24164 ;
  assign n24166 = n24158 & n24165 ;
  assign n24167 = n24151 & n24166 ;
  assign n24168 = \wishbone_bd_ram_mem1_reg[224][12]/P0001  & n13433 ;
  assign n24169 = \wishbone_bd_ram_mem1_reg[182][12]/P0001  & n13598 ;
  assign n24170 = ~n24168 & ~n24169 ;
  assign n24171 = \wishbone_bd_ram_mem1_reg[0][12]/P0001  & n13539 ;
  assign n24172 = \wishbone_bd_ram_mem1_reg[32][12]/P0001  & n13736 ;
  assign n24173 = ~n24171 & ~n24172 ;
  assign n24174 = n24170 & n24173 ;
  assign n24175 = \wishbone_bd_ram_mem1_reg[56][12]/P0001  & n13611 ;
  assign n24176 = \wishbone_bd_ram_mem1_reg[179][12]/P0001  & n14035 ;
  assign n24177 = ~n24175 & ~n24176 ;
  assign n24178 = \wishbone_bd_ram_mem1_reg[255][12]/P0001  & n13952 ;
  assign n24179 = \wishbone_bd_ram_mem1_reg[37][12]/P0001  & n13710 ;
  assign n24180 = ~n24178 & ~n24179 ;
  assign n24181 = n24177 & n24180 ;
  assign n24182 = n24174 & n24181 ;
  assign n24183 = \wishbone_bd_ram_mem1_reg[45][12]/P0001  & n13420 ;
  assign n24184 = \wishbone_bd_ram_mem1_reg[170][12]/P0001  & n14007 ;
  assign n24185 = ~n24183 & ~n24184 ;
  assign n24186 = \wishbone_bd_ram_mem1_reg[94][12]/P0001  & n13833 ;
  assign n24187 = \wishbone_bd_ram_mem1_reg[74][12]/P0001  & n13564 ;
  assign n24188 = ~n24186 & ~n24187 ;
  assign n24189 = n24185 & n24188 ;
  assign n24190 = \wishbone_bd_ram_mem1_reg[178][12]/P0001  & n13301 ;
  assign n24191 = \wishbone_bd_ram_mem1_reg[30][12]/P0001  & n13713 ;
  assign n24192 = ~n24190 & ~n24191 ;
  assign n24193 = \wishbone_bd_ram_mem1_reg[171][12]/P0001  & n13422 ;
  assign n24194 = \wishbone_bd_ram_mem1_reg[160][12]/P0001  & n13271 ;
  assign n24195 = ~n24193 & ~n24194 ;
  assign n24196 = n24192 & n24195 ;
  assign n24197 = n24189 & n24196 ;
  assign n24198 = n24182 & n24197 ;
  assign n24199 = n24167 & n24198 ;
  assign n24200 = n24136 & n24199 ;
  assign n24201 = \wishbone_bd_ram_mem1_reg[98][12]/P0001  & n13569 ;
  assign n24202 = \wishbone_bd_ram_mem1_reg[130][12]/P0001  & n13427 ;
  assign n24203 = ~n24201 & ~n24202 ;
  assign n24204 = \wishbone_bd_ram_mem1_reg[100][12]/P0001  & n13401 ;
  assign n24205 = \wishbone_bd_ram_mem1_reg[99][12]/P0001  & n13996 ;
  assign n24206 = ~n24204 & ~n24205 ;
  assign n24207 = n24203 & n24206 ;
  assign n24208 = \wishbone_bd_ram_mem1_reg[3][12]/P0001  & n13354 ;
  assign n24209 = \wishbone_bd_ram_mem1_reg[159][12]/P0001  & n13627 ;
  assign n24210 = ~n24208 & ~n24209 ;
  assign n24211 = \wishbone_bd_ram_mem1_reg[156][12]/P0001  & n13769 ;
  assign n24212 = \wishbone_bd_ram_mem1_reg[251][12]/P0001  & n14019 ;
  assign n24213 = ~n24211 & ~n24212 ;
  assign n24214 = n24210 & n24213 ;
  assign n24215 = n24207 & n24214 ;
  assign n24216 = \wishbone_bd_ram_mem1_reg[172][12]/P0001  & n13377 ;
  assign n24217 = \wishbone_bd_ram_mem1_reg[213][12]/P0001  & n13870 ;
  assign n24218 = ~n24216 & ~n24217 ;
  assign n24219 = \wishbone_bd_ram_mem1_reg[150][12]/P0001  & n13666 ;
  assign n24220 = \wishbone_bd_ram_mem1_reg[157][12]/P0001  & n13445 ;
  assign n24221 = ~n24219 & ~n24220 ;
  assign n24222 = n24218 & n24221 ;
  assign n24223 = \wishbone_bd_ram_mem1_reg[71][12]/P0001  & n13636 ;
  assign n24224 = \wishbone_bd_ram_mem1_reg[2][12]/P0001  & n13975 ;
  assign n24225 = ~n24223 & ~n24224 ;
  assign n24226 = \wishbone_bd_ram_mem1_reg[168][12]/P0001  & n13795 ;
  assign n24227 = \wishbone_bd_ram_mem1_reg[203][12]/P0001  & n13816 ;
  assign n24228 = ~n24226 & ~n24227 ;
  assign n24229 = n24225 & n24228 ;
  assign n24230 = n24222 & n24229 ;
  assign n24231 = n24215 & n24230 ;
  assign n24232 = \wishbone_bd_ram_mem1_reg[80][12]/P0001  & n13516 ;
  assign n24233 = \wishbone_bd_ram_mem1_reg[91][12]/P0001  & n13954 ;
  assign n24234 = ~n24232 & ~n24233 ;
  assign n24235 = \wishbone_bd_ram_mem1_reg[102][12]/P0001  & n13534 ;
  assign n24236 = \wishbone_bd_ram_mem1_reg[67][12]/P0001  & n13663 ;
  assign n24237 = ~n24235 & ~n24236 ;
  assign n24238 = n24234 & n24237 ;
  assign n24239 = \wishbone_bd_ram_mem1_reg[72][12]/P0001  & n13582 ;
  assign n24240 = \wishbone_bd_ram_mem1_reg[184][12]/P0001  & n13960 ;
  assign n24241 = ~n24239 & ~n24240 ;
  assign n24242 = \wishbone_bd_ram_mem1_reg[11][12]/P0001  & n13774 ;
  assign n24243 = \wishbone_bd_ram_mem1_reg[214][12]/P0001  & n13938 ;
  assign n24244 = ~n24242 & ~n24243 ;
  assign n24245 = n24241 & n24244 ;
  assign n24246 = n24238 & n24245 ;
  assign n24247 = \wishbone_bd_ram_mem1_reg[133][12]/P0001  & n13492 ;
  assign n24248 = \wishbone_bd_ram_mem1_reg[221][12]/P0001  & n13641 ;
  assign n24249 = ~n24247 & ~n24248 ;
  assign n24250 = \wishbone_bd_ram_mem1_reg[226][12]/P0001  & n13668 ;
  assign n24251 = \wishbone_bd_ram_mem1_reg[88][12]/P0001  & n13347 ;
  assign n24252 = ~n24250 & ~n24251 ;
  assign n24253 = n24249 & n24252 ;
  assign n24254 = \wishbone_bd_ram_mem1_reg[50][12]/P0001  & n13686 ;
  assign n24255 = \wishbone_bd_ram_mem1_reg[61][12]/P0001  & n13544 ;
  assign n24256 = ~n24254 & ~n24255 ;
  assign n24257 = \wishbone_bd_ram_mem1_reg[53][12]/P0001  & n13875 ;
  assign n24258 = \wishbone_bd_ram_mem1_reg[246][12]/P0001  & n13981 ;
  assign n24259 = ~n24257 & ~n24258 ;
  assign n24260 = n24256 & n24259 ;
  assign n24261 = n24253 & n24260 ;
  assign n24262 = n24246 & n24261 ;
  assign n24263 = n24231 & n24262 ;
  assign n24264 = \wishbone_bd_ram_mem1_reg[34][12]/P0001  & n13450 ;
  assign n24265 = \wishbone_bd_ram_mem1_reg[21][12]/P0001  & n13438 ;
  assign n24266 = ~n24264 & ~n24265 ;
  assign n24267 = \wishbone_bd_ram_mem1_reg[140][12]/P0001  & n13287 ;
  assign n24268 = \wishbone_bd_ram_mem1_reg[75][12]/P0001  & n13605 ;
  assign n24269 = ~n24267 & ~n24268 ;
  assign n24270 = n24266 & n24269 ;
  assign n24271 = \wishbone_bd_ram_mem1_reg[39][12]/P0001  & n13893 ;
  assign n24272 = \wishbone_bd_ram_mem1_reg[152][12]/P0001  & n13912 ;
  assign n24273 = ~n24271 & ~n24272 ;
  assign n24274 = \wishbone_bd_ram_mem1_reg[195][12]/P0001  & n13700 ;
  assign n24275 = \wishbone_bd_ram_mem1_reg[113][12]/P0001  & n13882 ;
  assign n24276 = ~n24274 & ~n24275 ;
  assign n24277 = n24273 & n24276 ;
  assign n24278 = n24270 & n24277 ;
  assign n24279 = \wishbone_bd_ram_mem1_reg[68][12]/P0001  & n13379 ;
  assign n24280 = \wishbone_bd_ram_mem1_reg[15][12]/P0001  & n13797 ;
  assign n24281 = ~n24279 & ~n24280 ;
  assign n24282 = \wishbone_bd_ram_mem1_reg[42][12]/P0001  & n13341 ;
  assign n24283 = \wishbone_bd_ram_mem1_reg[46][12]/P0001  & n13298 ;
  assign n24284 = ~n24282 & ~n24283 ;
  assign n24285 = n24281 & n24284 ;
  assign n24286 = \wishbone_bd_ram_mem1_reg[137][12]/P0001  & n13808 ;
  assign n24287 = \wishbone_bd_ram_mem1_reg[197][12]/P0001  & n13594 ;
  assign n24288 = ~n24286 & ~n24287 ;
  assign n24289 = \wishbone_bd_ram_mem1_reg[253][12]/P0001  & n13708 ;
  assign n24290 = \wishbone_bd_ram_mem1_reg[44][12]/P0001  & n13291 ;
  assign n24291 = ~n24289 & ~n24290 ;
  assign n24292 = n24288 & n24291 ;
  assign n24293 = n24285 & n24292 ;
  assign n24294 = n24278 & n24293 ;
  assign n24295 = \wishbone_bd_ram_mem1_reg[9][12]/P0001  & n13580 ;
  assign n24296 = \wishbone_bd_ram_mem1_reg[228][12]/P0001  & n13497 ;
  assign n24297 = ~n24295 & ~n24296 ;
  assign n24298 = \wishbone_bd_ram_mem1_reg[79][12]/P0001  & n13779 ;
  assign n24299 = \wishbone_bd_ram_mem1_reg[40][12]/P0001  & n13661 ;
  assign n24300 = ~n24298 & ~n24299 ;
  assign n24301 = n24297 & n24300 ;
  assign n24302 = \wishbone_bd_ram_mem1_reg[87][12]/P0001  & n13691 ;
  assign n24303 = \wishbone_bd_ram_mem1_reg[84][12]/P0001  & n13385 ;
  assign n24304 = ~n24302 & ~n24303 ;
  assign n24305 = \wishbone_bd_ram_mem1_reg[186][12]/P0001  & n13616 ;
  assign n24306 = \wishbone_bd_ram_mem1_reg[114][12]/P0001  & n13763 ;
  assign n24307 = ~n24305 & ~n24306 ;
  assign n24308 = n24304 & n24307 ;
  assign n24309 = n24301 & n24308 ;
  assign n24310 = \wishbone_bd_ram_mem1_reg[51][12]/P0001  & n13880 ;
  assign n24311 = \wishbone_bd_ram_mem1_reg[93][12]/P0001  & n13891 ;
  assign n24312 = ~n24310 & ~n24311 ;
  assign n24313 = \wishbone_bd_ram_mem1_reg[254][12]/P0001  & n13283 ;
  assign n24314 = \wishbone_bd_ram_mem1_reg[222][12]/P0001  & n13721 ;
  assign n24315 = ~n24313 & ~n24314 ;
  assign n24316 = n24312 & n24315 ;
  assign n24317 = \wishbone_bd_ram_mem1_reg[48][12]/P0001  & n13917 ;
  assign n24318 = \wishbone_bd_ram_mem1_reg[237][12]/P0001  & n13924 ;
  assign n24319 = ~n24317 & ~n24318 ;
  assign n24320 = \wishbone_bd_ram_mem1_reg[107][12]/P0001  & n13476 ;
  assign n24321 = \wishbone_bd_ram_mem1_reg[16][12]/P0001  & n13695 ;
  assign n24322 = ~n24320 & ~n24321 ;
  assign n24323 = n24319 & n24322 ;
  assign n24324 = n24316 & n24323 ;
  assign n24325 = n24309 & n24324 ;
  assign n24326 = n24294 & n24325 ;
  assign n24327 = n24263 & n24326 ;
  assign n24328 = n24200 & n24327 ;
  assign n24329 = n24073 & n24328 ;
  assign n24330 = ~wb_rst_i_pad & ~n23817 ;
  assign n24331 = ~n24329 & n24330 ;
  assign n24332 = ~n23818 & ~n24331 ;
  assign n24333 = \wishbone_TxLength_reg[3]/NET0131  & ~n14049 ;
  assign n24334 = ~n14046 & n24333 ;
  assign n24335 = ~\wishbone_TxLength_reg[2]/NET0131  & n17372 ;
  assign n24336 = \wishbone_TxLength_reg[3]/NET0131  & ~n24335 ;
  assign n24337 = n17371 & ~n17373 ;
  assign n24338 = ~n24336 & n24337 ;
  assign n24339 = n14049 & ~n24338 ;
  assign n24340 = ~n14064 & n24339 ;
  assign n24341 = ~\wishbone_TxLength_reg[1]/NET0131  & ~\wishbone_TxLength_reg[2]/NET0131  ;
  assign n24342 = ~\wishbone_TxLength_reg[2]/NET0131  & ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
  assign n24343 = ~n14068 & n24342 ;
  assign n24344 = ~n24341 & ~n24343 ;
  assign n24345 = ~\wishbone_TxLength_reg[3]/NET0131  & ~n17371 ;
  assign n24346 = n24344 & n24345 ;
  assign n24347 = \wishbone_TxLength_reg[3]/NET0131  & ~n17371 ;
  assign n24348 = ~n24344 & n24347 ;
  assign n24349 = ~n24346 & ~n24348 ;
  assign n24350 = ~n14046 & n24349 ;
  assign n24351 = n24340 & n24350 ;
  assign n24352 = ~n24334 & ~n24351 ;
  assign n24353 = ~n22173 & n24352 ;
  assign n24354 = \wishbone_TxLength_reg[6]/NET0131  & ~n14049 ;
  assign n24355 = ~n17360 & ~n24354 ;
  assign n24356 = ~\wishbone_TxLength_reg[4]/NET0131  & ~\wishbone_TxLength_reg[5]/NET0131  ;
  assign n24357 = n14054 & n24356 ;
  assign n24358 = \wishbone_TxLength_reg[6]/NET0131  & ~n24357 ;
  assign n24359 = ~n14057 & ~n24358 ;
  assign n24360 = n17379 & ~n24359 ;
  assign n24361 = ~n17365 & n24359 ;
  assign n24362 = ~\wishbone_TxLength_reg[6]/NET0131  & n17365 ;
  assign n24363 = n17367 & ~n24362 ;
  assign n24364 = ~n24361 & n24363 ;
  assign n24365 = ~n24360 & ~n24364 ;
  assign n24366 = ~\wishbone_TxLength_reg[0]/NET0131  & \wishbone_TxLength_reg[6]/NET0131  ;
  assign n24367 = ~\wishbone_TxLength_reg[5]/NET0131  & n24366 ;
  assign n24368 = n17383 & n24367 ;
  assign n24369 = \wishbone_TxLength_reg[6]/NET0131  & n17371 ;
  assign n24370 = n17371 & n17372 ;
  assign n24371 = n24357 & n24370 ;
  assign n24372 = ~n24369 & ~n24371 ;
  assign n24373 = ~n24368 & ~n24372 ;
  assign n24374 = ~\wishbone_TxLength_reg[5]/NET0131  & n17383 ;
  assign n24375 = ~\wishbone_TxLength_reg[6]/NET0131  & ~n24374 ;
  assign n24376 = ~\wishbone_TxLength_reg[5]/NET0131  & \wishbone_TxLength_reg[6]/NET0131  ;
  assign n24377 = n17383 & n24376 ;
  assign n24378 = n17381 & ~n24377 ;
  assign n24379 = ~n24375 & n24378 ;
  assign n24380 = ~n24373 & ~n24379 ;
  assign n24381 = ~n24354 & n24380 ;
  assign n24382 = n24365 & n24381 ;
  assign n24383 = ~n24355 & ~n24382 ;
  assign n24384 = ~n14046 & n24383 ;
  assign n24385 = ~n23719 & ~n24384 ;
  assign n24386 = \wishbone_TxPointerLSB_reg[1]/NET0131  & ~n18545 ;
  assign n24387 = ~wb_rst_i_pad & n18545 ;
  assign n24388 = ~n16820 & n24387 ;
  assign n24389 = ~n24386 & ~n24388 ;
  assign n24390 = \wishbone_TxPointerLSB_rst_reg[0]/NET0131  & ~n14049 ;
  assign n24391 = ~n18545 & n24390 ;
  assign n24392 = \wishbone_bd_ram_mem0_reg[153][0]/P0001  & n13309 ;
  assign n24393 = \wishbone_bd_ram_mem0_reg[174][0]/P0001  & n13899 ;
  assign n24394 = ~n24392 & ~n24393 ;
  assign n24395 = \wishbone_bd_ram_mem0_reg[166][0]/P0001  & n13999 ;
  assign n24396 = \wishbone_bd_ram_mem0_reg[150][0]/P0001  & n13666 ;
  assign n24397 = ~n24395 & ~n24396 ;
  assign n24398 = n24394 & n24397 ;
  assign n24399 = \wishbone_bd_ram_mem0_reg[159][0]/P0001  & n13627 ;
  assign n24400 = \wishbone_bd_ram_mem0_reg[25][0]/P0001  & n13742 ;
  assign n24401 = ~n24399 & ~n24400 ;
  assign n24402 = \wishbone_bd_ram_mem0_reg[26][0]/P0001  & n13521 ;
  assign n24403 = \wishbone_bd_ram_mem0_reg[146][0]/P0001  & n13958 ;
  assign n24404 = ~n24402 & ~n24403 ;
  assign n24405 = n24401 & n24404 ;
  assign n24406 = n24398 & n24405 ;
  assign n24407 = \wishbone_bd_ram_mem0_reg[14][0]/P0001  & n13972 ;
  assign n24408 = \wishbone_bd_ram_mem0_reg[189][0]/P0001  & n14001 ;
  assign n24409 = ~n24407 & ~n24408 ;
  assign n24410 = \wishbone_bd_ram_mem0_reg[3][0]/P0001  & n13354 ;
  assign n24411 = \wishbone_bd_ram_mem0_reg[194][0]/P0001  & n13624 ;
  assign n24412 = ~n24410 & ~n24411 ;
  assign n24413 = n24409 & n24412 ;
  assign n24414 = \wishbone_bd_ram_mem0_reg[101][0]/P0001  & n13772 ;
  assign n24415 = \wishbone_bd_ram_mem0_reg[238][0]/P0001  & n13819 ;
  assign n24416 = ~n24414 & ~n24415 ;
  assign n24417 = \wishbone_bd_ram_mem0_reg[115][0]/P0001  & n13747 ;
  assign n24418 = \wishbone_bd_ram_mem0_reg[164][0]/P0001  & n13236 ;
  assign n24419 = ~n24417 & ~n24418 ;
  assign n24420 = n24416 & n24419 ;
  assign n24421 = n24413 & n24420 ;
  assign n24422 = n24406 & n24421 ;
  assign n24423 = \wishbone_bd_ram_mem0_reg[114][0]/P0001  & n13763 ;
  assign n24424 = \wishbone_bd_ram_mem0_reg[79][0]/P0001  & n13779 ;
  assign n24425 = ~n24423 & ~n24424 ;
  assign n24426 = \wishbone_bd_ram_mem0_reg[151][0]/P0001  & n13697 ;
  assign n24427 = \wishbone_bd_ram_mem0_reg[112][0]/P0001  & n13482 ;
  assign n24428 = ~n24426 & ~n24427 ;
  assign n24429 = n24425 & n24428 ;
  assign n24430 = \wishbone_bd_ram_mem0_reg[228][0]/P0001  & n13497 ;
  assign n24431 = \wishbone_bd_ram_mem0_reg[0][0]/P0001  & n13539 ;
  assign n24432 = ~n24430 & ~n24431 ;
  assign n24433 = \wishbone_bd_ram_mem0_reg[184][0]/P0001  & n13960 ;
  assign n24434 = \wishbone_bd_ram_mem0_reg[30][0]/P0001  & n13713 ;
  assign n24435 = ~n24433 & ~n24434 ;
  assign n24436 = n24432 & n24435 ;
  assign n24437 = n24429 & n24436 ;
  assign n24438 = \wishbone_bd_ram_mem0_reg[103][0]/P0001  & n13320 ;
  assign n24439 = \wishbone_bd_ram_mem0_reg[7][0]/P0001  & n13546 ;
  assign n24440 = ~n24438 & ~n24439 ;
  assign n24441 = \wishbone_bd_ram_mem0_reg[45][0]/P0001  & n13420 ;
  assign n24442 = \wishbone_bd_ram_mem0_reg[39][0]/P0001  & n13893 ;
  assign n24443 = ~n24441 & ~n24442 ;
  assign n24444 = n24440 & n24443 ;
  assign n24445 = \wishbone_bd_ram_mem0_reg[126][0]/P0001  & n13786 ;
  assign n24446 = \wishbone_bd_ram_mem0_reg[47][0]/P0001  & n13436 ;
  assign n24447 = ~n24445 & ~n24446 ;
  assign n24448 = \wishbone_bd_ram_mem0_reg[58][0]/P0001  & n13949 ;
  assign n24449 = \wishbone_bd_ram_mem0_reg[196][0]/P0001  & n13977 ;
  assign n24450 = ~n24448 & ~n24449 ;
  assign n24451 = n24447 & n24450 ;
  assign n24452 = n24444 & n24451 ;
  assign n24453 = n24437 & n24452 ;
  assign n24454 = n24422 & n24453 ;
  assign n24455 = \wishbone_bd_ram_mem0_reg[205][0]/P0001  & n13947 ;
  assign n24456 = \wishbone_bd_ram_mem0_reg[207][0]/P0001  & n13826 ;
  assign n24457 = ~n24455 & ~n24456 ;
  assign n24458 = \wishbone_bd_ram_mem0_reg[110][0]/P0001  & n14030 ;
  assign n24459 = \wishbone_bd_ram_mem0_reg[149][0]/P0001  & n13469 ;
  assign n24460 = ~n24458 & ~n24459 ;
  assign n24461 = n24457 & n24460 ;
  assign n24462 = \wishbone_bd_ram_mem0_reg[236][0]/P0001  & n13480 ;
  assign n24463 = \wishbone_bd_ram_mem0_reg[113][0]/P0001  & n13882 ;
  assign n24464 = ~n24462 & ~n24463 ;
  assign n24465 = \wishbone_bd_ram_mem0_reg[109][0]/P0001  & n13306 ;
  assign n24466 = \wishbone_bd_ram_mem0_reg[127][0]/P0001  & n13803 ;
  assign n24467 = ~n24465 & ~n24466 ;
  assign n24468 = n24464 & n24467 ;
  assign n24469 = n24461 & n24468 ;
  assign n24470 = \wishbone_bd_ram_mem0_reg[171][0]/P0001  & n13422 ;
  assign n24471 = \wishbone_bd_ram_mem0_reg[22][0]/P0001  & n13744 ;
  assign n24472 = ~n24470 & ~n24471 ;
  assign n24473 = \wishbone_bd_ram_mem0_reg[132][0]/P0001  & n13927 ;
  assign n24474 = \wishbone_bd_ram_mem0_reg[165][0]/P0001  & n14028 ;
  assign n24475 = ~n24473 & ~n24474 ;
  assign n24476 = n24472 & n24475 ;
  assign n24477 = \wishbone_bd_ram_mem0_reg[241][0]/P0001  & n13854 ;
  assign n24478 = \wishbone_bd_ram_mem0_reg[186][0]/P0001  & n13616 ;
  assign n24479 = ~n24477 & ~n24478 ;
  assign n24480 = \wishbone_bd_ram_mem0_reg[119][0]/P0001  & n14033 ;
  assign n24481 = \wishbone_bd_ram_mem0_reg[48][0]/P0001  & n13917 ;
  assign n24482 = ~n24480 & ~n24481 ;
  assign n24483 = n24479 & n24482 ;
  assign n24484 = n24476 & n24483 ;
  assign n24485 = n24469 & n24484 ;
  assign n24486 = \wishbone_bd_ram_mem0_reg[155][0]/P0001  & n13738 ;
  assign n24487 = \wishbone_bd_ram_mem0_reg[62][0]/P0001  & n13529 ;
  assign n24488 = ~n24486 & ~n24487 ;
  assign n24489 = \wishbone_bd_ram_mem0_reg[148][0]/P0001  & n13868 ;
  assign n24490 = \wishbone_bd_ram_mem0_reg[89][0]/P0001  & n13910 ;
  assign n24491 = ~n24489 & ~n24490 ;
  assign n24492 = n24488 & n24491 ;
  assign n24493 = \wishbone_bd_ram_mem0_reg[213][0]/P0001  & n13870 ;
  assign n24494 = \wishbone_bd_ram_mem0_reg[212][0]/P0001  & n13634 ;
  assign n24495 = ~n24493 & ~n24494 ;
  assign n24496 = \wishbone_bd_ram_mem0_reg[84][0]/P0001  & n13385 ;
  assign n24497 = \wishbone_bd_ram_mem0_reg[1][0]/P0001  & n13888 ;
  assign n24498 = ~n24496 & ~n24497 ;
  assign n24499 = n24495 & n24498 ;
  assign n24500 = n24492 & n24499 ;
  assign n24501 = \wishbone_bd_ram_mem0_reg[252][0]/P0001  & n13986 ;
  assign n24502 = \wishbone_bd_ram_mem0_reg[96][0]/P0001  & n13425 ;
  assign n24503 = ~n24501 & ~n24502 ;
  assign n24504 = \wishbone_bd_ram_mem0_reg[123][0]/P0001  & n13749 ;
  assign n24505 = \wishbone_bd_ram_mem0_reg[102][0]/P0001  & n13534 ;
  assign n24506 = ~n24504 & ~n24505 ;
  assign n24507 = n24503 & n24506 ;
  assign n24508 = \wishbone_bd_ram_mem0_reg[41][0]/P0001  & n14017 ;
  assign n24509 = \wishbone_bd_ram_mem0_reg[46][0]/P0001  & n13298 ;
  assign n24510 = ~n24508 & ~n24509 ;
  assign n24511 = \wishbone_bd_ram_mem0_reg[61][0]/P0001  & n13544 ;
  assign n24512 = \wishbone_bd_ram_mem0_reg[230][0]/P0001  & n13994 ;
  assign n24513 = ~n24511 & ~n24512 ;
  assign n24514 = n24510 & n24513 ;
  assign n24515 = n24507 & n24514 ;
  assign n24516 = n24500 & n24515 ;
  assign n24517 = n24485 & n24516 ;
  assign n24518 = n24454 & n24517 ;
  assign n24519 = \wishbone_bd_ram_mem0_reg[68][0]/P0001  & n13379 ;
  assign n24520 = \wishbone_bd_ram_mem0_reg[31][0]/P0001  & n13758 ;
  assign n24521 = ~n24519 & ~n24520 ;
  assign n24522 = \wishbone_bd_ram_mem0_reg[209][0]/P0001  & n13689 ;
  assign n24523 = \wishbone_bd_ram_mem0_reg[179][0]/P0001  & n14035 ;
  assign n24524 = ~n24522 & ~n24523 ;
  assign n24525 = n24521 & n24524 ;
  assign n24526 = \wishbone_bd_ram_mem0_reg[223][0]/P0001  & n13335 ;
  assign n24527 = \wishbone_bd_ram_mem0_reg[66][0]/P0001  & n13603 ;
  assign n24528 = ~n24526 & ~n24527 ;
  assign n24529 = \wishbone_bd_ram_mem0_reg[12][0]/P0001  & n13733 ;
  assign n24530 = \wishbone_bd_ram_mem0_reg[211][0]/P0001  & n13805 ;
  assign n24531 = ~n24529 & ~n24530 ;
  assign n24532 = n24528 & n24531 ;
  assign n24533 = n24525 & n24532 ;
  assign n24534 = \wishbone_bd_ram_mem0_reg[91][0]/P0001  & n13954 ;
  assign n24535 = \wishbone_bd_ram_mem0_reg[133][0]/P0001  & n13492 ;
  assign n24536 = ~n24534 & ~n24535 ;
  assign n24537 = \wishbone_bd_ram_mem0_reg[234][0]/P0001  & n13781 ;
  assign n24538 = \wishbone_bd_ram_mem0_reg[42][0]/P0001  & n13341 ;
  assign n24539 = ~n24537 & ~n24538 ;
  assign n24540 = n24536 & n24539 ;
  assign n24541 = \wishbone_bd_ram_mem0_reg[237][0]/P0001  & n13924 ;
  assign n24542 = \wishbone_bd_ram_mem0_reg[135][0]/P0001  & n13672 ;
  assign n24543 = ~n24541 & ~n24542 ;
  assign n24544 = \wishbone_bd_ram_mem0_reg[192][0]/P0001  & n13390 ;
  assign n24545 = \wishbone_bd_ram_mem0_reg[198][0]/P0001  & n13592 ;
  assign n24546 = ~n24544 & ~n24545 ;
  assign n24547 = n24543 & n24546 ;
  assign n24548 = n24540 & n24547 ;
  assign n24549 = n24533 & n24548 ;
  assign n24550 = \wishbone_bd_ram_mem0_reg[183][0]/P0001  & n13645 ;
  assign n24551 = \wishbone_bd_ram_mem0_reg[60][0]/P0001  & n13790 ;
  assign n24552 = ~n24550 & ~n24551 ;
  assign n24553 = \wishbone_bd_ram_mem0_reg[86][0]/P0001  & n13485 ;
  assign n24554 = \wishbone_bd_ram_mem0_reg[6][0]/P0001  & n13915 ;
  assign n24555 = ~n24553 & ~n24554 ;
  assign n24556 = n24552 & n24555 ;
  assign n24557 = \wishbone_bd_ram_mem0_reg[185][0]/P0001  & n13372 ;
  assign n24558 = \wishbone_bd_ram_mem0_reg[130][0]/P0001  & n13427 ;
  assign n24559 = ~n24557 & ~n24558 ;
  assign n24560 = \wishbone_bd_ram_mem0_reg[235][0]/P0001  & n13518 ;
  assign n24561 = \wishbone_bd_ram_mem0_reg[21][0]/P0001  & n13438 ;
  assign n24562 = ~n24560 & ~n24561 ;
  assign n24563 = n24559 & n24562 ;
  assign n24564 = n24556 & n24563 ;
  assign n24565 = \wishbone_bd_ram_mem0_reg[175][0]/P0001  & n13674 ;
  assign n24566 = \wishbone_bd_ram_mem0_reg[36][0]/P0001  & n13639 ;
  assign n24567 = ~n24565 & ~n24566 ;
  assign n24568 = \wishbone_bd_ram_mem0_reg[247][0]/P0001  & n13571 ;
  assign n24569 = \wishbone_bd_ram_mem0_reg[215][0]/P0001  & n13901 ;
  assign n24570 = ~n24568 & ~n24569 ;
  assign n24571 = n24567 & n24570 ;
  assign n24572 = \wishbone_bd_ram_mem0_reg[197][0]/P0001  & n13594 ;
  assign n24573 = \wishbone_bd_ram_mem0_reg[122][0]/P0001  & n13679 ;
  assign n24574 = ~n24572 & ~n24573 ;
  assign n24575 = \wishbone_bd_ram_mem0_reg[244][0]/P0001  & n13474 ;
  assign n24576 = \wishbone_bd_ram_mem0_reg[93][0]/P0001  & n13891 ;
  assign n24577 = ~n24575 & ~n24576 ;
  assign n24578 = n24574 & n24577 ;
  assign n24579 = n24571 & n24578 ;
  assign n24580 = n24564 & n24579 ;
  assign n24581 = n24549 & n24580 ;
  assign n24582 = \wishbone_bd_ram_mem0_reg[195][0]/P0001  & n13700 ;
  assign n24583 = \wishbone_bd_ram_mem0_reg[226][0]/P0001  & n13668 ;
  assign n24584 = ~n24582 & ~n24583 ;
  assign n24585 = \wishbone_bd_ram_mem0_reg[24][0]/P0001  & n13970 ;
  assign n24586 = \wishbone_bd_ram_mem0_reg[8][0]/P0001  & n13459 ;
  assign n24587 = ~n24585 & ~n24586 ;
  assign n24588 = n24584 & n24587 ;
  assign n24589 = \wishbone_bd_ram_mem0_reg[199][0]/P0001  & n13499 ;
  assign n24590 = \wishbone_bd_ram_mem0_reg[250][0]/P0001  & n13677 ;
  assign n24591 = ~n24589 & ~n24590 ;
  assign n24592 = \wishbone_bd_ram_mem0_reg[5][0]/P0001  & n13243 ;
  assign n24593 = \wishbone_bd_ram_mem0_reg[9][0]/P0001  & n13580 ;
  assign n24594 = ~n24592 & ~n24593 ;
  assign n24595 = n24591 & n24594 ;
  assign n24596 = n24588 & n24595 ;
  assign n24597 = \wishbone_bd_ram_mem0_reg[214][0]/P0001  & n13938 ;
  assign n24598 = \wishbone_bd_ram_mem0_reg[203][0]/P0001  & n13816 ;
  assign n24599 = ~n24597 & ~n24598 ;
  assign n24600 = \wishbone_bd_ram_mem0_reg[232][0]/P0001  & n13510 ;
  assign n24601 = \wishbone_bd_ram_mem0_reg[140][0]/P0001  & n13287 ;
  assign n24602 = ~n24600 & ~n24601 ;
  assign n24603 = n24599 & n24602 ;
  assign n24604 = \wishbone_bd_ram_mem0_reg[64][0]/P0001  & n13904 ;
  assign n24605 = \wishbone_bd_ram_mem0_reg[222][0]/P0001  & n13721 ;
  assign n24606 = ~n24604 & ~n24605 ;
  assign n24607 = \wishbone_bd_ram_mem0_reg[10][0]/P0001  & n13837 ;
  assign n24608 = \wishbone_bd_ram_mem0_reg[28][0]/P0001  & n13810 ;
  assign n24609 = ~n24607 & ~n24608 ;
  assign n24610 = n24606 & n24609 ;
  assign n24611 = n24603 & n24610 ;
  assign n24612 = n24596 & n24611 ;
  assign n24613 = \wishbone_bd_ram_mem0_reg[144][0]/P0001  & n13508 ;
  assign n24614 = \wishbone_bd_ram_mem0_reg[188][0]/P0001  & n13407 ;
  assign n24615 = ~n24613 & ~n24614 ;
  assign n24616 = \wishbone_bd_ram_mem0_reg[249][0]/P0001  & n13431 ;
  assign n24617 = \wishbone_bd_ram_mem0_reg[251][0]/P0001  & n14019 ;
  assign n24618 = ~n24616 & ~n24617 ;
  assign n24619 = n24615 & n24618 ;
  assign n24620 = \wishbone_bd_ram_mem0_reg[87][0]/P0001  & n13691 ;
  assign n24621 = \wishbone_bd_ram_mem0_reg[82][0]/P0001  & n13374 ;
  assign n24622 = ~n24620 & ~n24621 ;
  assign n24623 = \wishbone_bd_ram_mem0_reg[11][0]/P0001  & n13774 ;
  assign n24624 = \wishbone_bd_ram_mem0_reg[81][0]/P0001  & n13409 ;
  assign n24625 = ~n24623 & ~n24624 ;
  assign n24626 = n24622 & n24625 ;
  assign n24627 = n24619 & n24626 ;
  assign n24628 = \wishbone_bd_ram_mem0_reg[160][0]/P0001  & n13271 ;
  assign n24629 = \wishbone_bd_ram_mem0_reg[32][0]/P0001  & n13736 ;
  assign n24630 = ~n24628 & ~n24629 ;
  assign n24631 = \wishbone_bd_ram_mem0_reg[169][0]/P0001  & n13541 ;
  assign n24632 = \wishbone_bd_ram_mem0_reg[216][0]/P0001  & n14005 ;
  assign n24633 = ~n24631 & ~n24632 ;
  assign n24634 = n24630 & n24633 ;
  assign n24635 = \wishbone_bd_ram_mem0_reg[18][0]/P0001  & n13532 ;
  assign n24636 = \wishbone_bd_ram_mem0_reg[111][0]/P0001  & n13471 ;
  assign n24637 = ~n24635 & ~n24636 ;
  assign n24638 = \wishbone_bd_ram_mem0_reg[242][0]/P0001  & n13383 ;
  assign n24639 = \wishbone_bd_ram_mem0_reg[78][0]/P0001  & n13277 ;
  assign n24640 = ~n24638 & ~n24639 ;
  assign n24641 = n24637 & n24640 ;
  assign n24642 = n24634 & n24641 ;
  assign n24643 = n24627 & n24642 ;
  assign n24644 = n24612 & n24643 ;
  assign n24645 = n24581 & n24644 ;
  assign n24646 = n24518 & n24645 ;
  assign n24647 = \wishbone_bd_ram_mem0_reg[57][0]/P0001  & n13731 ;
  assign n24648 = \wishbone_bd_ram_mem0_reg[177][0]/P0001  & n13863 ;
  assign n24649 = ~n24647 & ~n24648 ;
  assign n24650 = \wishbone_bd_ram_mem0_reg[163][0]/P0001  & n13255 ;
  assign n24651 = \wishbone_bd_ram_mem0_reg[190][0]/P0001  & n13365 ;
  assign n24652 = ~n24650 & ~n24651 ;
  assign n24653 = n24649 & n24652 ;
  assign n24654 = \wishbone_bd_ram_mem0_reg[243][0]/P0001  & n13575 ;
  assign n24655 = \wishbone_bd_ram_mem0_reg[191][0]/P0001  & n14012 ;
  assign n24656 = ~n24654 & ~n24655 ;
  assign n24657 = \wishbone_bd_ram_mem0_reg[217][0]/P0001  & n13767 ;
  assign n24658 = \wishbone_bd_ram_mem0_reg[229][0]/P0001  & n13552 ;
  assign n24659 = ~n24657 & ~n24658 ;
  assign n24660 = n24656 & n24659 ;
  assign n24661 = n24653 & n24660 ;
  assign n24662 = \wishbone_bd_ram_mem0_reg[231][0]/P0001  & n13363 ;
  assign n24663 = \wishbone_bd_ram_mem0_reg[77][0]/P0001  & n13935 ;
  assign n24664 = ~n24662 & ~n24663 ;
  assign n24665 = \wishbone_bd_ram_mem0_reg[37][0]/P0001  & n13710 ;
  assign n24666 = \wishbone_bd_ram_mem0_reg[181][0]/P0001  & n13587 ;
  assign n24667 = ~n24665 & ~n24666 ;
  assign n24668 = n24664 & n24667 ;
  assign n24669 = \wishbone_bd_ram_mem0_reg[120][0]/P0001  & n13550 ;
  assign n24670 = \wishbone_bd_ram_mem0_reg[17][0]/P0001  & n13324 ;
  assign n24671 = ~n24669 & ~n24670 ;
  assign n24672 = \wishbone_bd_ram_mem0_reg[225][0]/P0001  & n13719 ;
  assign n24673 = \wishbone_bd_ram_mem0_reg[219][0]/P0001  & n13577 ;
  assign n24674 = ~n24672 & ~n24673 ;
  assign n24675 = n24671 & n24674 ;
  assign n24676 = n24668 & n24675 ;
  assign n24677 = n24661 & n24676 ;
  assign n24678 = \wishbone_bd_ram_mem0_reg[227][0]/P0001  & n13388 ;
  assign n24679 = \wishbone_bd_ram_mem0_reg[106][0]/P0001  & n13555 ;
  assign n24680 = ~n24678 & ~n24679 ;
  assign n24681 = \wishbone_bd_ram_mem0_reg[161][0]/P0001  & n13505 ;
  assign n24682 = \wishbone_bd_ram_mem0_reg[85][0]/P0001  & n13784 ;
  assign n24683 = ~n24681 & ~n24682 ;
  assign n24684 = n24680 & n24683 ;
  assign n24685 = \wishbone_bd_ram_mem0_reg[75][0]/P0001  & n13605 ;
  assign n24686 = \wishbone_bd_ram_mem0_reg[168][0]/P0001  & n13795 ;
  assign n24687 = ~n24685 & ~n24686 ;
  assign n24688 = \wishbone_bd_ram_mem0_reg[240][0]/P0001  & n13352 ;
  assign n24689 = \wishbone_bd_ram_mem0_reg[152][0]/P0001  & n13912 ;
  assign n24690 = ~n24688 & ~n24689 ;
  assign n24691 = n24687 & n24690 ;
  assign n24692 = n24684 & n24691 ;
  assign n24693 = \wishbone_bd_ram_mem0_reg[90][0]/P0001  & n13906 ;
  assign n24694 = \wishbone_bd_ram_mem0_reg[128][0]/P0001  & n13652 ;
  assign n24695 = ~n24693 & ~n24694 ;
  assign n24696 = \wishbone_bd_ram_mem0_reg[187][0]/P0001  & n13756 ;
  assign n24697 = \wishbone_bd_ram_mem0_reg[248][0]/P0001  & n13647 ;
  assign n24698 = ~n24696 & ~n24697 ;
  assign n24699 = n24695 & n24698 ;
  assign n24700 = \wishbone_bd_ram_mem0_reg[202][0]/P0001  & n13268 ;
  assign n24701 = \wishbone_bd_ram_mem0_reg[23][0]/P0001  & n13857 ;
  assign n24702 = ~n24700 & ~n24701 ;
  assign n24703 = \wishbone_bd_ram_mem0_reg[208][0]/P0001  & n14010 ;
  assign n24704 = \wishbone_bd_ram_mem0_reg[76][0]/P0001  & n13831 ;
  assign n24705 = ~n24703 & ~n24704 ;
  assign n24706 = n24702 & n24705 ;
  assign n24707 = n24699 & n24706 ;
  assign n24708 = n24692 & n24707 ;
  assign n24709 = n24677 & n24708 ;
  assign n24710 = \wishbone_bd_ram_mem0_reg[246][0]/P0001  & n13981 ;
  assign n24711 = \wishbone_bd_ram_mem0_reg[193][0]/P0001  & n14022 ;
  assign n24712 = ~n24710 & ~n24711 ;
  assign n24713 = \wishbone_bd_ram_mem0_reg[50][0]/P0001  & n13686 ;
  assign n24714 = \wishbone_bd_ram_mem0_reg[38][0]/P0001  & n13828 ;
  assign n24715 = ~n24713 & ~n24714 ;
  assign n24716 = n24712 & n24715 ;
  assign n24717 = \wishbone_bd_ram_mem0_reg[147][0]/P0001  & n13702 ;
  assign n24718 = \wishbone_bd_ram_mem0_reg[49][0]/P0001  & n13929 ;
  assign n24719 = ~n24717 & ~n24718 ;
  assign n24720 = \wishbone_bd_ram_mem0_reg[94][0]/P0001  & n13833 ;
  assign n24721 = \wishbone_bd_ram_mem0_reg[74][0]/P0001  & n13564 ;
  assign n24722 = ~n24720 & ~n24721 ;
  assign n24723 = n24719 & n24722 ;
  assign n24724 = n24716 & n24723 ;
  assign n24725 = \wishbone_bd_ram_mem0_reg[33][0]/P0001  & n13933 ;
  assign n24726 = \wishbone_bd_ram_mem0_reg[134][0]/P0001  & n13494 ;
  assign n24727 = ~n24725 & ~n24726 ;
  assign n24728 = \wishbone_bd_ram_mem0_reg[180][0]/P0001  & n13650 ;
  assign n24729 = \wishbone_bd_ram_mem0_reg[98][0]/P0001  & n13569 ;
  assign n24730 = ~n24728 & ~n24729 ;
  assign n24731 = n24727 & n24730 ;
  assign n24732 = \wishbone_bd_ram_mem0_reg[121][0]/P0001  & n13983 ;
  assign n24733 = \wishbone_bd_ram_mem0_reg[162][0]/P0001  & n13726 ;
  assign n24734 = ~n24732 & ~n24733 ;
  assign n24735 = \wishbone_bd_ram_mem0_reg[210][0]/P0001  & n13443 ;
  assign n24736 = \wishbone_bd_ram_mem0_reg[176][0]/P0001  & n13262 ;
  assign n24737 = ~n24735 & ~n24736 ;
  assign n24738 = n24734 & n24737 ;
  assign n24739 = n24731 & n24738 ;
  assign n24740 = n24724 & n24739 ;
  assign n24741 = \wishbone_bd_ram_mem0_reg[200][0]/P0001  & n13922 ;
  assign n24742 = \wishbone_bd_ram_mem0_reg[125][0]/P0001  & n13396 ;
  assign n24743 = ~n24741 & ~n24742 ;
  assign n24744 = \wishbone_bd_ram_mem0_reg[124][0]/P0001  & n14024 ;
  assign n24745 = \wishbone_bd_ram_mem0_reg[15][0]/P0001  & n13797 ;
  assign n24746 = ~n24744 & ~n24745 ;
  assign n24747 = n24743 & n24746 ;
  assign n24748 = \wishbone_bd_ram_mem0_reg[44][0]/P0001  & n13291 ;
  assign n24749 = \wishbone_bd_ram_mem0_reg[118][0]/P0001  & n13589 ;
  assign n24750 = ~n24748 & ~n24749 ;
  assign n24751 = \wishbone_bd_ram_mem0_reg[137][0]/P0001  & n13808 ;
  assign n24752 = \wishbone_bd_ram_mem0_reg[43][0]/P0001  & n13761 ;
  assign n24753 = ~n24751 & ~n24752 ;
  assign n24754 = n24750 & n24753 ;
  assign n24755 = n24747 & n24754 ;
  assign n24756 = \wishbone_bd_ram_mem0_reg[55][0]/P0001  & n13618 ;
  assign n24757 = \wishbone_bd_ram_mem0_reg[131][0]/P0001  & n13358 ;
  assign n24758 = ~n24756 & ~n24757 ;
  assign n24759 = \wishbone_bd_ram_mem0_reg[233][0]/P0001  & n13332 ;
  assign n24760 = \wishbone_bd_ram_mem0_reg[158][0]/P0001  & n13294 ;
  assign n24761 = ~n24759 & ~n24760 ;
  assign n24762 = n24758 & n24761 ;
  assign n24763 = \wishbone_bd_ram_mem0_reg[63][0]/P0001  & n13327 ;
  assign n24764 = \wishbone_bd_ram_mem0_reg[69][0]/P0001  & n13487 ;
  assign n24765 = ~n24763 & ~n24764 ;
  assign n24766 = \wishbone_bd_ram_mem0_reg[40][0]/P0001  & n13661 ;
  assign n24767 = \wishbone_bd_ram_mem0_reg[16][0]/P0001  & n13695 ;
  assign n24768 = ~n24766 & ~n24767 ;
  assign n24769 = n24765 & n24768 ;
  assign n24770 = n24762 & n24769 ;
  assign n24771 = n24755 & n24770 ;
  assign n24772 = n24740 & n24771 ;
  assign n24773 = n24709 & n24772 ;
  assign n24774 = \wishbone_bd_ram_mem0_reg[20][0]/P0001  & n13839 ;
  assign n24775 = \wishbone_bd_ram_mem0_reg[178][0]/P0001  & n13301 ;
  assign n24776 = ~n24774 & ~n24775 ;
  assign n24777 = \wishbone_bd_ram_mem0_reg[139][0]/P0001  & n13566 ;
  assign n24778 = \wishbone_bd_ram_mem0_reg[206][0]/P0001  & n13414 ;
  assign n24779 = ~n24777 & ~n24778 ;
  assign n24780 = n24776 & n24779 ;
  assign n24781 = \wishbone_bd_ram_mem0_reg[255][0]/P0001  & n13952 ;
  assign n24782 = \wishbone_bd_ram_mem0_reg[138][0]/P0001  & n13398 ;
  assign n24783 = ~n24781 & ~n24782 ;
  assign n24784 = \wishbone_bd_ram_mem0_reg[104][0]/P0001  & n13684 ;
  assign n24785 = \wishbone_bd_ram_mem0_reg[167][0]/P0001  & n13940 ;
  assign n24786 = ~n24784 & ~n24785 ;
  assign n24787 = n24783 & n24786 ;
  assign n24788 = n24780 & n24787 ;
  assign n24789 = \wishbone_bd_ram_mem0_reg[218][0]/P0001  & n13792 ;
  assign n24790 = \wishbone_bd_ram_mem0_reg[239][0]/P0001  & n13349 ;
  assign n24791 = ~n24789 & ~n24790 ;
  assign n24792 = \wishbone_bd_ram_mem0_reg[92][0]/P0001  & n13859 ;
  assign n24793 = \wishbone_bd_ram_mem0_reg[173][0]/P0001  & n13360 ;
  assign n24794 = ~n24792 & ~n24793 ;
  assign n24795 = n24791 & n24794 ;
  assign n24796 = \wishbone_bd_ram_mem0_reg[129][0]/P0001  & n13629 ;
  assign n24797 = \wishbone_bd_ram_mem0_reg[56][0]/P0001  & n13611 ;
  assign n24798 = ~n24796 & ~n24797 ;
  assign n24799 = \wishbone_bd_ram_mem0_reg[19][0]/P0001  & n13886 ;
  assign n24800 = \wishbone_bd_ram_mem0_reg[108][0]/P0001  & n13814 ;
  assign n24801 = ~n24799 & ~n24800 ;
  assign n24802 = n24798 & n24801 ;
  assign n24803 = n24795 & n24802 ;
  assign n24804 = n24788 & n24803 ;
  assign n24805 = \wishbone_bd_ram_mem0_reg[52][0]/P0001  & n13988 ;
  assign n24806 = \wishbone_bd_ram_mem0_reg[201][0]/P0001  & n13600 ;
  assign n24807 = ~n24805 & ~n24806 ;
  assign n24808 = \wishbone_bd_ram_mem0_reg[4][0]/P0001  & n13527 ;
  assign n24809 = \wishbone_bd_ram_mem0_reg[107][0]/P0001  & n13476 ;
  assign n24810 = ~n24808 & ~n24809 ;
  assign n24811 = n24807 & n24810 ;
  assign n24812 = \wishbone_bd_ram_mem0_reg[141][0]/P0001  & n13852 ;
  assign n24813 = \wishbone_bd_ram_mem0_reg[105][0]/P0001  & n13503 ;
  assign n24814 = ~n24812 & ~n24813 ;
  assign n24815 = \wishbone_bd_ram_mem0_reg[59][0]/P0001  & n13613 ;
  assign n24816 = \wishbone_bd_ram_mem0_reg[51][0]/P0001  & n13880 ;
  assign n24817 = ~n24815 & ~n24816 ;
  assign n24818 = n24814 & n24817 ;
  assign n24819 = n24811 & n24818 ;
  assign n24820 = \wishbone_bd_ram_mem0_reg[34][0]/P0001  & n13450 ;
  assign n24821 = \wishbone_bd_ram_mem0_reg[70][0]/P0001  & n13339 ;
  assign n24822 = ~n24820 & ~n24821 ;
  assign n24823 = \wishbone_bd_ram_mem0_reg[73][0]/P0001  & n13456 ;
  assign n24824 = \wishbone_bd_ram_mem0_reg[157][0]/P0001  & n13445 ;
  assign n24825 = ~n24823 & ~n24824 ;
  assign n24826 = n24822 & n24825 ;
  assign n24827 = \wishbone_bd_ram_mem0_reg[88][0]/P0001  & n13347 ;
  assign n24828 = \wishbone_bd_ram_mem0_reg[204][0]/P0001  & n13821 ;
  assign n24829 = ~n24827 & ~n24828 ;
  assign n24830 = \wishbone_bd_ram_mem0_reg[54][0]/P0001  & n13622 ;
  assign n24831 = \wishbone_bd_ram_mem0_reg[117][0]/P0001  & n13557 ;
  assign n24832 = ~n24830 & ~n24831 ;
  assign n24833 = n24829 & n24832 ;
  assign n24834 = n24826 & n24833 ;
  assign n24835 = n24819 & n24834 ;
  assign n24836 = n24804 & n24835 ;
  assign n24837 = \wishbone_bd_ram_mem0_reg[95][0]/P0001  & n13317 ;
  assign n24838 = \wishbone_bd_ram_mem0_reg[156][0]/P0001  & n13769 ;
  assign n24839 = ~n24837 & ~n24838 ;
  assign n24840 = \wishbone_bd_ram_mem0_reg[72][0]/P0001  & n13582 ;
  assign n24841 = \wishbone_bd_ram_mem0_reg[142][0]/P0001  & n13448 ;
  assign n24842 = ~n24840 & ~n24841 ;
  assign n24843 = n24839 & n24842 ;
  assign n24844 = \wishbone_bd_ram_mem0_reg[224][0]/P0001  & n13433 ;
  assign n24845 = \wishbone_bd_ram_mem0_reg[53][0]/P0001  & n13875 ;
  assign n24846 = ~n24844 & ~n24845 ;
  assign n24847 = \wishbone_bd_ram_mem0_reg[253][0]/P0001  & n13708 ;
  assign n24848 = \wishbone_bd_ram_mem0_reg[170][0]/P0001  & n14007 ;
  assign n24849 = ~n24847 & ~n24848 ;
  assign n24850 = n24846 & n24849 ;
  assign n24851 = n24843 & n24850 ;
  assign n24852 = \wishbone_bd_ram_mem0_reg[182][0]/P0001  & n13598 ;
  assign n24853 = \wishbone_bd_ram_mem0_reg[99][0]/P0001  & n13996 ;
  assign n24854 = ~n24852 & ~n24853 ;
  assign n24855 = \wishbone_bd_ram_mem0_reg[67][0]/P0001  & n13663 ;
  assign n24856 = \wishbone_bd_ram_mem0_reg[116][0]/P0001  & n13865 ;
  assign n24857 = ~n24855 & ~n24856 ;
  assign n24858 = n24854 & n24857 ;
  assign n24859 = \wishbone_bd_ram_mem0_reg[97][0]/P0001  & n13724 ;
  assign n24860 = \wishbone_bd_ram_mem0_reg[65][0]/P0001  & n13842 ;
  assign n24861 = ~n24859 & ~n24860 ;
  assign n24862 = \wishbone_bd_ram_mem0_reg[245][0]/P0001  & n13877 ;
  assign n24863 = \wishbone_bd_ram_mem0_reg[2][0]/P0001  & n13975 ;
  assign n24864 = ~n24862 & ~n24863 ;
  assign n24865 = n24861 & n24864 ;
  assign n24866 = n24858 & n24865 ;
  assign n24867 = n24851 & n24866 ;
  assign n24868 = \wishbone_bd_ram_mem0_reg[143][0]/P0001  & n13461 ;
  assign n24869 = \wishbone_bd_ram_mem0_reg[254][0]/P0001  & n13283 ;
  assign n24870 = ~n24868 & ~n24869 ;
  assign n24871 = \wishbone_bd_ram_mem0_reg[27][0]/P0001  & n13251 ;
  assign n24872 = \wishbone_bd_ram_mem0_reg[29][0]/P0001  & n13412 ;
  assign n24873 = ~n24871 & ~n24872 ;
  assign n24874 = n24870 & n24873 ;
  assign n24875 = \wishbone_bd_ram_mem0_reg[221][0]/P0001  & n13641 ;
  assign n24876 = \wishbone_bd_ram_mem0_reg[220][0]/P0001  & n13965 ;
  assign n24877 = ~n24875 & ~n24876 ;
  assign n24878 = \wishbone_bd_ram_mem0_reg[136][0]/P0001  & n13963 ;
  assign n24879 = \wishbone_bd_ram_mem0_reg[145][0]/P0001  & n13715 ;
  assign n24880 = ~n24878 & ~n24879 ;
  assign n24881 = n24877 & n24880 ;
  assign n24882 = n24874 & n24881 ;
  assign n24883 = \wishbone_bd_ram_mem0_reg[172][0]/P0001  & n13377 ;
  assign n24884 = \wishbone_bd_ram_mem0_reg[100][0]/P0001  & n13401 ;
  assign n24885 = ~n24883 & ~n24884 ;
  assign n24886 = \wishbone_bd_ram_mem0_reg[71][0]/P0001  & n13636 ;
  assign n24887 = \wishbone_bd_ram_mem0_reg[35][0]/P0001  & n13523 ;
  assign n24888 = ~n24886 & ~n24887 ;
  assign n24889 = n24885 & n24888 ;
  assign n24890 = \wishbone_bd_ram_mem0_reg[154][0]/P0001  & n13403 ;
  assign n24891 = \wishbone_bd_ram_mem0_reg[83][0]/P0001  & n13454 ;
  assign n24892 = ~n24890 & ~n24891 ;
  assign n24893 = \wishbone_bd_ram_mem0_reg[13][0]/P0001  & n13844 ;
  assign n24894 = \wishbone_bd_ram_mem0_reg[80][0]/P0001  & n13516 ;
  assign n24895 = ~n24893 & ~n24894 ;
  assign n24896 = n24892 & n24895 ;
  assign n24897 = n24889 & n24896 ;
  assign n24898 = n24882 & n24897 ;
  assign n24899 = n24867 & n24898 ;
  assign n24900 = n24836 & n24899 ;
  assign n24901 = n24773 & n24900 ;
  assign n24902 = n24646 & n24901 ;
  assign n24903 = n24387 & ~n24902 ;
  assign n24904 = ~n24391 & ~n24903 ;
  assign n24905 = \wishbone_TxPointerLSB_reg[0]/NET0131  & ~n18545 ;
  assign n24906 = ~n24903 & ~n24905 ;
  assign n24907 = \wishbone_TxPointerLSB_rst_reg[1]/NET0131  & ~n14049 ;
  assign n24908 = ~n18545 & n24907 ;
  assign n24909 = ~n24388 & ~n24908 ;
  assign n24910 = \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  & n23737 ;
  assign n24911 = \ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131  & n23743 ;
  assign n24912 = n23741 & n24911 ;
  assign n24913 = \ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131  & n23743 ;
  assign n24914 = n23747 & n24913 ;
  assign n24915 = ~n24912 & ~n24914 ;
  assign n24916 = \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  & n23751 ;
  assign n24917 = n23741 & n24916 ;
  assign n24918 = n23730 & ~n24917 ;
  assign n24919 = n24915 & n24918 ;
  assign n24920 = ~n24910 & n24919 ;
  assign n24921 = n23730 & ~n24920 ;
  assign n24922 = ~wb_rst_i_pad & ~n24920 ;
  assign n24923 = ~n23202 & n24922 ;
  assign n24924 = ~n24921 & ~n24923 ;
  assign n24925 = \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  & n23737 ;
  assign n24926 = \ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131  & n23743 ;
  assign n24927 = n23741 & n24926 ;
  assign n24928 = \ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131  & n23743 ;
  assign n24929 = n23747 & n24928 ;
  assign n24930 = ~n24927 & ~n24929 ;
  assign n24931 = \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  & n23751 ;
  assign n24932 = n23741 & n24931 ;
  assign n24933 = n23730 & ~n24932 ;
  assign n24934 = n24930 & n24933 ;
  assign n24935 = ~n24925 & n24934 ;
  assign n24936 = n23730 & ~n24935 ;
  assign n24937 = ~wb_rst_i_pad & ~n24935 ;
  assign n24938 = ~n15695 & n24937 ;
  assign n24939 = ~n24936 & ~n24938 ;
  assign n24940 = \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  & n23737 ;
  assign n24941 = \ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131  & n23743 ;
  assign n24942 = n23741 & n24941 ;
  assign n24943 = \ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131  & n23743 ;
  assign n24944 = n23747 & n24943 ;
  assign n24945 = ~n24942 & ~n24944 ;
  assign n24946 = \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  & n23751 ;
  assign n24947 = n23741 & n24946 ;
  assign n24948 = n23730 & ~n24947 ;
  assign n24949 = n24945 & n24948 ;
  assign n24950 = ~n24940 & n24949 ;
  assign n24951 = n23730 & ~n24950 ;
  assign n24952 = ~wb_rst_i_pad & ~n24950 ;
  assign n24953 = ~n18434 & n24952 ;
  assign n24954 = ~n24951 & ~n24953 ;
  assign n24955 = \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  & n23737 ;
  assign n24956 = \ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131  & n23743 ;
  assign n24957 = n23741 & n24956 ;
  assign n24958 = \ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131  & n23743 ;
  assign n24959 = n23747 & n24958 ;
  assign n24960 = ~n24957 & ~n24959 ;
  assign n24961 = \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  & n23751 ;
  assign n24962 = n23741 & n24961 ;
  assign n24963 = n23730 & ~n24962 ;
  assign n24964 = n24960 & n24963 ;
  assign n24965 = ~n24955 & n24964 ;
  assign n24966 = n23730 & ~n24965 ;
  assign n24967 = ~wb_rst_i_pad & ~n24965 ;
  assign n24968 = ~n17905 & n24967 ;
  assign n24969 = ~n24966 & ~n24968 ;
  assign n24970 = \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  & n23737 ;
  assign n24971 = \ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131  & n23743 ;
  assign n24972 = n23741 & n24971 ;
  assign n24973 = \ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131  & n23743 ;
  assign n24974 = n23747 & n24973 ;
  assign n24975 = ~n24972 & ~n24974 ;
  assign n24976 = \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  & n23751 ;
  assign n24977 = n23741 & n24976 ;
  assign n24978 = n23730 & ~n24977 ;
  assign n24979 = n24975 & n24978 ;
  assign n24980 = ~n24970 & n24979 ;
  assign n24981 = n23730 & ~n24980 ;
  assign n24982 = ~wb_rst_i_pad & ~n24980 ;
  assign n24983 = ~n21643 & n24982 ;
  assign n24984 = ~n24981 & ~n24983 ;
  assign n24985 = \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  & n23737 ;
  assign n24986 = \ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131  & n23743 ;
  assign n24987 = n23741 & n24986 ;
  assign n24988 = \ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131  & n23743 ;
  assign n24989 = n23747 & n24988 ;
  assign n24990 = ~n24987 & ~n24989 ;
  assign n24991 = \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  & n23751 ;
  assign n24992 = n23741 & n24991 ;
  assign n24993 = n23730 & ~n24992 ;
  assign n24994 = n24990 & n24993 ;
  assign n24995 = ~n24985 & n24994 ;
  assign n24996 = n23730 & ~n24995 ;
  assign n24997 = ~wb_rst_i_pad & ~n24995 ;
  assign n24998 = ~n14044 & n24997 ;
  assign n24999 = ~n24996 & ~n24998 ;
  assign n25000 = \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  & n23737 ;
  assign n25001 = \ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131  & n23743 ;
  assign n25002 = n23741 & n25001 ;
  assign n25003 = \ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131  & n23743 ;
  assign n25004 = n23747 & n25003 ;
  assign n25005 = ~n25002 & ~n25004 ;
  assign n25006 = \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  & n23751 ;
  assign n25007 = n23741 & n25006 ;
  assign n25008 = n23730 & ~n25007 ;
  assign n25009 = n25005 & n25008 ;
  assign n25010 = ~n25000 & n25009 ;
  assign n25011 = n23730 & ~n25010 ;
  assign n25012 = ~wb_rst_i_pad & ~n25010 ;
  assign n25013 = ~n14593 & n25012 ;
  assign n25014 = ~n25011 & ~n25013 ;
  assign n25015 = m_wb_we_o_pad & n13189 ;
  assign n25016 = n13196 & ~n25015 ;
  assign n25017 = \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  & n23737 ;
  assign n25018 = \ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131  & n23743 ;
  assign n25019 = n23741 & n25018 ;
  assign n25020 = \ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131  & n23743 ;
  assign n25021 = n23747 & n25020 ;
  assign n25022 = ~n25019 & ~n25021 ;
  assign n25023 = \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  & n23751 ;
  assign n25024 = n23741 & n25023 ;
  assign n25025 = n23730 & ~n25024 ;
  assign n25026 = n25022 & n25025 ;
  assign n25027 = ~n25017 & n25026 ;
  assign n25028 = n23730 & ~n25027 ;
  assign n25029 = ~wb_rst_i_pad & ~n25027 ;
  assign n25030 = ~n15114 & n25029 ;
  assign n25031 = ~n25028 & ~n25030 ;
  assign n25032 = \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  & n23737 ;
  assign n25033 = \ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131  & n23743 ;
  assign n25034 = n23741 & n25033 ;
  assign n25035 = \ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131  & n23743 ;
  assign n25036 = n23747 & n25035 ;
  assign n25037 = ~n25034 & ~n25036 ;
  assign n25038 = \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  & n23751 ;
  assign n25039 = n23741 & n25038 ;
  assign n25040 = n23730 & ~n25039 ;
  assign n25041 = n25037 & n25040 ;
  assign n25042 = ~n25032 & n25041 ;
  assign n25043 = n23730 & ~n25042 ;
  assign n25044 = ~wb_rst_i_pad & ~n25042 ;
  assign n25045 = ~n20314 & n25044 ;
  assign n25046 = ~n25043 & ~n25045 ;
  assign n25047 = \ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131  & n23743 ;
  assign n25048 = n23747 & n25047 ;
  assign n25049 = \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  & n23751 ;
  assign n25050 = n23741 & n25049 ;
  assign n25051 = ~n25048 & ~n25050 ;
  assign n25052 = \ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131  & n23782 ;
  assign n25053 = \ethreg1_MODER_0_DataOut_reg[3]/NET0131  & n23808 ;
  assign n25054 = ~n25052 & ~n25053 ;
  assign n25055 = n25051 & n25054 ;
  assign n25056 = \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  & n23737 ;
  assign n25057 = \wb_adr_i[2]_pad  & \wb_adr_i[3]_pad  ;
  assign n25058 = n23735 & n25057 ;
  assign n25059 = n23733 & n25058 ;
  assign n25060 = \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  & n25059 ;
  assign n25061 = ~n25056 & ~n25060 ;
  assign n25062 = n25055 & n25061 ;
  assign n25063 = n23746 & n23806 ;
  assign n25064 = n23805 & n25063 ;
  assign n25065 = \ethreg1_irq_rxe_reg/NET0131  & n25064 ;
  assign n25066 = \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131  & n23794 ;
  assign n25067 = n23741 & n25066 ;
  assign n25068 = ~n25065 & ~n25067 ;
  assign n25069 = n23779 & n23805 ;
  assign n25070 = \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131  & n25069 ;
  assign n25071 = \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131  & n23802 ;
  assign n25072 = ~n25070 & ~n25071 ;
  assign n25073 = n25068 & n25072 ;
  assign n25074 = n23730 & n25073 ;
  assign n25075 = \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  & n23751 ;
  assign n25076 = n23747 & n25075 ;
  assign n25077 = \wb_adr_i[3]_pad  & ~\wb_adr_i[5]_pad  ;
  assign n25078 = n23731 & n25077 ;
  assign n25079 = n23807 & n25078 ;
  assign n25080 = \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131  & n25079 ;
  assign n25081 = ~n25076 & ~n25080 ;
  assign n25082 = n23805 & n23812 ;
  assign n25083 = \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131  & n25082 ;
  assign n25084 = n23781 & n23807 ;
  assign n25085 = \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  & n25084 ;
  assign n25086 = ~n25083 & ~n25085 ;
  assign n25087 = n25081 & n25086 ;
  assign n25088 = n23801 & n23807 ;
  assign n25089 = \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131  & n25088 ;
  assign n25090 = n25063 & n25078 ;
  assign n25091 = \ethreg1_IPGT_0_DataOut_reg[3]/NET0131  & n25090 ;
  assign n25092 = ~n25089 & ~n25091 ;
  assign n25093 = \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131  & n23813 ;
  assign n25094 = \ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131  & n23743 ;
  assign n25095 = n23741 & n25094 ;
  assign n25096 = ~n25093 & ~n25095 ;
  assign n25097 = n25092 & n25096 ;
  assign n25098 = n25087 & n25097 ;
  assign n25099 = n25074 & n25098 ;
  assign n25100 = n25062 & n25099 ;
  assign n25101 = n23730 & ~n25100 ;
  assign n25102 = \wishbone_bd_ram_mem0_reg[209][3]/P0001  & n13689 ;
  assign n25103 = \wishbone_bd_ram_mem0_reg[12][3]/P0001  & n13733 ;
  assign n25104 = ~n25102 & ~n25103 ;
  assign n25105 = \wishbone_bd_ram_mem0_reg[37][3]/P0001  & n13710 ;
  assign n25106 = \wishbone_bd_ram_mem0_reg[162][3]/P0001  & n13726 ;
  assign n25107 = ~n25105 & ~n25106 ;
  assign n25108 = n25104 & n25107 ;
  assign n25109 = \wishbone_bd_ram_mem0_reg[94][3]/P0001  & n13833 ;
  assign n25110 = \wishbone_bd_ram_mem0_reg[97][3]/P0001  & n13724 ;
  assign n25111 = ~n25109 & ~n25110 ;
  assign n25112 = \wishbone_bd_ram_mem0_reg[128][3]/P0001  & n13652 ;
  assign n25113 = \wishbone_bd_ram_mem0_reg[175][3]/P0001  & n13674 ;
  assign n25114 = ~n25112 & ~n25113 ;
  assign n25115 = n25111 & n25114 ;
  assign n25116 = n25108 & n25115 ;
  assign n25117 = \wishbone_bd_ram_mem0_reg[187][3]/P0001  & n13756 ;
  assign n25118 = \wishbone_bd_ram_mem0_reg[197][3]/P0001  & n13594 ;
  assign n25119 = ~n25117 & ~n25118 ;
  assign n25120 = \wishbone_bd_ram_mem0_reg[102][3]/P0001  & n13534 ;
  assign n25121 = \wishbone_bd_ram_mem0_reg[228][3]/P0001  & n13497 ;
  assign n25122 = ~n25120 & ~n25121 ;
  assign n25123 = n25119 & n25122 ;
  assign n25124 = \wishbone_bd_ram_mem0_reg[11][3]/P0001  & n13774 ;
  assign n25125 = \wishbone_bd_ram_mem0_reg[246][3]/P0001  & n13981 ;
  assign n25126 = ~n25124 & ~n25125 ;
  assign n25127 = \wishbone_bd_ram_mem0_reg[115][3]/P0001  & n13747 ;
  assign n25128 = \wishbone_bd_ram_mem0_reg[156][3]/P0001  & n13769 ;
  assign n25129 = ~n25127 & ~n25128 ;
  assign n25130 = n25126 & n25129 ;
  assign n25131 = n25123 & n25130 ;
  assign n25132 = n25116 & n25131 ;
  assign n25133 = \wishbone_bd_ram_mem0_reg[144][3]/P0001  & n13508 ;
  assign n25134 = \wishbone_bd_ram_mem0_reg[153][3]/P0001  & n13309 ;
  assign n25135 = ~n25133 & ~n25134 ;
  assign n25136 = \wishbone_bd_ram_mem0_reg[3][3]/P0001  & n13354 ;
  assign n25137 = \wishbone_bd_ram_mem0_reg[122][3]/P0001  & n13679 ;
  assign n25138 = ~n25136 & ~n25137 ;
  assign n25139 = n25135 & n25138 ;
  assign n25140 = \wishbone_bd_ram_mem0_reg[225][3]/P0001  & n13719 ;
  assign n25141 = \wishbone_bd_ram_mem0_reg[179][3]/P0001  & n14035 ;
  assign n25142 = ~n25140 & ~n25141 ;
  assign n25143 = \wishbone_bd_ram_mem0_reg[216][3]/P0001  & n14005 ;
  assign n25144 = \wishbone_bd_ram_mem0_reg[30][3]/P0001  & n13713 ;
  assign n25145 = ~n25143 & ~n25144 ;
  assign n25146 = n25142 & n25145 ;
  assign n25147 = n25139 & n25146 ;
  assign n25148 = \wishbone_bd_ram_mem0_reg[43][3]/P0001  & n13761 ;
  assign n25149 = \wishbone_bd_ram_mem0_reg[194][3]/P0001  & n13624 ;
  assign n25150 = ~n25148 & ~n25149 ;
  assign n25151 = \wishbone_bd_ram_mem0_reg[229][3]/P0001  & n13552 ;
  assign n25152 = \wishbone_bd_ram_mem0_reg[21][3]/P0001  & n13438 ;
  assign n25153 = ~n25151 & ~n25152 ;
  assign n25154 = n25150 & n25153 ;
  assign n25155 = \wishbone_bd_ram_mem0_reg[14][3]/P0001  & n13972 ;
  assign n25156 = \wishbone_bd_ram_mem0_reg[49][3]/P0001  & n13929 ;
  assign n25157 = ~n25155 & ~n25156 ;
  assign n25158 = \wishbone_bd_ram_mem0_reg[231][3]/P0001  & n13363 ;
  assign n25159 = \wishbone_bd_ram_mem0_reg[226][3]/P0001  & n13668 ;
  assign n25160 = ~n25158 & ~n25159 ;
  assign n25161 = n25157 & n25160 ;
  assign n25162 = n25154 & n25161 ;
  assign n25163 = n25147 & n25162 ;
  assign n25164 = n25132 & n25163 ;
  assign n25165 = \wishbone_bd_ram_mem0_reg[247][3]/P0001  & n13571 ;
  assign n25166 = \wishbone_bd_ram_mem0_reg[93][3]/P0001  & n13891 ;
  assign n25167 = ~n25165 & ~n25166 ;
  assign n25168 = \wishbone_bd_ram_mem0_reg[48][3]/P0001  & n13917 ;
  assign n25169 = \wishbone_bd_ram_mem0_reg[96][3]/P0001  & n13425 ;
  assign n25170 = ~n25168 & ~n25169 ;
  assign n25171 = n25167 & n25170 ;
  assign n25172 = \wishbone_bd_ram_mem0_reg[211][3]/P0001  & n13805 ;
  assign n25173 = \wishbone_bd_ram_mem0_reg[106][3]/P0001  & n13555 ;
  assign n25174 = ~n25172 & ~n25173 ;
  assign n25175 = \wishbone_bd_ram_mem0_reg[190][3]/P0001  & n13365 ;
  assign n25176 = \wishbone_bd_ram_mem0_reg[108][3]/P0001  & n13814 ;
  assign n25177 = ~n25175 & ~n25176 ;
  assign n25178 = n25174 & n25177 ;
  assign n25179 = n25171 & n25178 ;
  assign n25180 = \wishbone_bd_ram_mem0_reg[180][3]/P0001  & n13650 ;
  assign n25181 = \wishbone_bd_ram_mem0_reg[109][3]/P0001  & n13306 ;
  assign n25182 = ~n25180 & ~n25181 ;
  assign n25183 = \wishbone_bd_ram_mem0_reg[117][3]/P0001  & n13557 ;
  assign n25184 = \wishbone_bd_ram_mem0_reg[184][3]/P0001  & n13960 ;
  assign n25185 = ~n25183 & ~n25184 ;
  assign n25186 = n25182 & n25185 ;
  assign n25187 = \wishbone_bd_ram_mem0_reg[111][3]/P0001  & n13471 ;
  assign n25188 = \wishbone_bd_ram_mem0_reg[215][3]/P0001  & n13901 ;
  assign n25189 = ~n25187 & ~n25188 ;
  assign n25190 = \wishbone_bd_ram_mem0_reg[119][3]/P0001  & n14033 ;
  assign n25191 = \wishbone_bd_ram_mem0_reg[181][3]/P0001  & n13587 ;
  assign n25192 = ~n25190 & ~n25191 ;
  assign n25193 = n25189 & n25192 ;
  assign n25194 = n25186 & n25193 ;
  assign n25195 = n25179 & n25194 ;
  assign n25196 = \wishbone_bd_ram_mem0_reg[137][3]/P0001  & n13808 ;
  assign n25197 = \wishbone_bd_ram_mem0_reg[174][3]/P0001  & n13899 ;
  assign n25198 = ~n25196 & ~n25197 ;
  assign n25199 = \wishbone_bd_ram_mem0_reg[164][3]/P0001  & n13236 ;
  assign n25200 = \wishbone_bd_ram_mem0_reg[146][3]/P0001  & n13958 ;
  assign n25201 = ~n25199 & ~n25200 ;
  assign n25202 = n25198 & n25201 ;
  assign n25203 = \wishbone_bd_ram_mem0_reg[239][3]/P0001  & n13349 ;
  assign n25204 = \wishbone_bd_ram_mem0_reg[223][3]/P0001  & n13335 ;
  assign n25205 = ~n25203 & ~n25204 ;
  assign n25206 = \wishbone_bd_ram_mem0_reg[149][3]/P0001  & n13469 ;
  assign n25207 = \wishbone_bd_ram_mem0_reg[4][3]/P0001  & n13527 ;
  assign n25208 = ~n25206 & ~n25207 ;
  assign n25209 = n25205 & n25208 ;
  assign n25210 = n25202 & n25209 ;
  assign n25211 = \wishbone_bd_ram_mem0_reg[133][3]/P0001  & n13492 ;
  assign n25212 = \wishbone_bd_ram_mem0_reg[157][3]/P0001  & n13445 ;
  assign n25213 = ~n25211 & ~n25212 ;
  assign n25214 = \wishbone_bd_ram_mem0_reg[123][3]/P0001  & n13749 ;
  assign n25215 = \wishbone_bd_ram_mem0_reg[38][3]/P0001  & n13828 ;
  assign n25216 = ~n25214 & ~n25215 ;
  assign n25217 = n25213 & n25216 ;
  assign n25218 = \wishbone_bd_ram_mem0_reg[105][3]/P0001  & n13503 ;
  assign n25219 = \wishbone_bd_ram_mem0_reg[74][3]/P0001  & n13564 ;
  assign n25220 = ~n25218 & ~n25219 ;
  assign n25221 = \wishbone_bd_ram_mem0_reg[44][3]/P0001  & n13291 ;
  assign n25222 = \wishbone_bd_ram_mem0_reg[120][3]/P0001  & n13550 ;
  assign n25223 = ~n25221 & ~n25222 ;
  assign n25224 = n25220 & n25223 ;
  assign n25225 = n25217 & n25224 ;
  assign n25226 = n25210 & n25225 ;
  assign n25227 = n25195 & n25226 ;
  assign n25228 = n25164 & n25227 ;
  assign n25229 = \wishbone_bd_ram_mem0_reg[148][3]/P0001  & n13868 ;
  assign n25230 = \wishbone_bd_ram_mem0_reg[202][3]/P0001  & n13268 ;
  assign n25231 = ~n25229 & ~n25230 ;
  assign n25232 = \wishbone_bd_ram_mem0_reg[244][3]/P0001  & n13474 ;
  assign n25233 = \wishbone_bd_ram_mem0_reg[125][3]/P0001  & n13396 ;
  assign n25234 = ~n25232 & ~n25233 ;
  assign n25235 = n25231 & n25234 ;
  assign n25236 = \wishbone_bd_ram_mem0_reg[212][3]/P0001  & n13634 ;
  assign n25237 = \wishbone_bd_ram_mem0_reg[241][3]/P0001  & n13854 ;
  assign n25238 = ~n25236 & ~n25237 ;
  assign n25239 = \wishbone_bd_ram_mem0_reg[85][3]/P0001  & n13784 ;
  assign n25240 = \wishbone_bd_ram_mem0_reg[65][3]/P0001  & n13842 ;
  assign n25241 = ~n25239 & ~n25240 ;
  assign n25242 = n25238 & n25241 ;
  assign n25243 = n25235 & n25242 ;
  assign n25244 = \wishbone_bd_ram_mem0_reg[186][3]/P0001  & n13616 ;
  assign n25245 = \wishbone_bd_ram_mem0_reg[101][3]/P0001  & n13772 ;
  assign n25246 = ~n25244 & ~n25245 ;
  assign n25247 = \wishbone_bd_ram_mem0_reg[210][3]/P0001  & n13443 ;
  assign n25248 = \wishbone_bd_ram_mem0_reg[140][3]/P0001  & n13287 ;
  assign n25249 = ~n25247 & ~n25248 ;
  assign n25250 = n25246 & n25249 ;
  assign n25251 = \wishbone_bd_ram_mem0_reg[87][3]/P0001  & n13691 ;
  assign n25252 = \wishbone_bd_ram_mem0_reg[135][3]/P0001  & n13672 ;
  assign n25253 = ~n25251 & ~n25252 ;
  assign n25254 = \wishbone_bd_ram_mem0_reg[98][3]/P0001  & n13569 ;
  assign n25255 = \wishbone_bd_ram_mem0_reg[198][3]/P0001  & n13592 ;
  assign n25256 = ~n25254 & ~n25255 ;
  assign n25257 = n25253 & n25256 ;
  assign n25258 = n25250 & n25257 ;
  assign n25259 = n25243 & n25258 ;
  assign n25260 = \wishbone_bd_ram_mem0_reg[86][3]/P0001  & n13485 ;
  assign n25261 = \wishbone_bd_ram_mem0_reg[236][3]/P0001  & n13480 ;
  assign n25262 = ~n25260 & ~n25261 ;
  assign n25263 = \wishbone_bd_ram_mem0_reg[160][3]/P0001  & n13271 ;
  assign n25264 = \wishbone_bd_ram_mem0_reg[32][3]/P0001  & n13736 ;
  assign n25265 = ~n25263 & ~n25264 ;
  assign n25266 = n25262 & n25265 ;
  assign n25267 = \wishbone_bd_ram_mem0_reg[17][3]/P0001  & n13324 ;
  assign n25268 = \wishbone_bd_ram_mem0_reg[57][3]/P0001  & n13731 ;
  assign n25269 = ~n25267 & ~n25268 ;
  assign n25270 = \wishbone_bd_ram_mem0_reg[40][3]/P0001  & n13661 ;
  assign n25271 = \wishbone_bd_ram_mem0_reg[182][3]/P0001  & n13598 ;
  assign n25272 = ~n25270 & ~n25271 ;
  assign n25273 = n25269 & n25272 ;
  assign n25274 = n25266 & n25273 ;
  assign n25275 = \wishbone_bd_ram_mem0_reg[9][3]/P0001  & n13580 ;
  assign n25276 = \wishbone_bd_ram_mem0_reg[92][3]/P0001  & n13859 ;
  assign n25277 = ~n25275 & ~n25276 ;
  assign n25278 = \wishbone_bd_ram_mem0_reg[39][3]/P0001  & n13893 ;
  assign n25279 = \wishbone_bd_ram_mem0_reg[28][3]/P0001  & n13810 ;
  assign n25280 = ~n25278 & ~n25279 ;
  assign n25281 = n25277 & n25280 ;
  assign n25282 = \wishbone_bd_ram_mem0_reg[189][3]/P0001  & n14001 ;
  assign n25283 = \wishbone_bd_ram_mem0_reg[248][3]/P0001  & n13647 ;
  assign n25284 = ~n25282 & ~n25283 ;
  assign n25285 = \wishbone_bd_ram_mem0_reg[79][3]/P0001  & n13779 ;
  assign n25286 = \wishbone_bd_ram_mem0_reg[167][3]/P0001  & n13940 ;
  assign n25287 = ~n25285 & ~n25286 ;
  assign n25288 = n25284 & n25287 ;
  assign n25289 = n25281 & n25288 ;
  assign n25290 = n25274 & n25289 ;
  assign n25291 = n25259 & n25290 ;
  assign n25292 = \wishbone_bd_ram_mem0_reg[76][3]/P0001  & n13831 ;
  assign n25293 = \wishbone_bd_ram_mem0_reg[196][3]/P0001  & n13977 ;
  assign n25294 = ~n25292 & ~n25293 ;
  assign n25295 = \wishbone_bd_ram_mem0_reg[151][3]/P0001  & n13697 ;
  assign n25296 = \wishbone_bd_ram_mem0_reg[185][3]/P0001  & n13372 ;
  assign n25297 = ~n25295 & ~n25296 ;
  assign n25298 = n25294 & n25297 ;
  assign n25299 = \wishbone_bd_ram_mem0_reg[199][3]/P0001  & n13499 ;
  assign n25300 = \wishbone_bd_ram_mem0_reg[83][3]/P0001  & n13454 ;
  assign n25301 = ~n25299 & ~n25300 ;
  assign n25302 = \wishbone_bd_ram_mem0_reg[5][3]/P0001  & n13243 ;
  assign n25303 = \wishbone_bd_ram_mem0_reg[78][3]/P0001  & n13277 ;
  assign n25304 = ~n25302 & ~n25303 ;
  assign n25305 = n25301 & n25304 ;
  assign n25306 = n25298 & n25305 ;
  assign n25307 = \wishbone_bd_ram_mem0_reg[221][3]/P0001  & n13641 ;
  assign n25308 = \wishbone_bd_ram_mem0_reg[64][3]/P0001  & n13904 ;
  assign n25309 = ~n25307 & ~n25308 ;
  assign n25310 = \wishbone_bd_ram_mem0_reg[139][3]/P0001  & n13566 ;
  assign n25311 = \wishbone_bd_ram_mem0_reg[243][3]/P0001  & n13575 ;
  assign n25312 = ~n25310 & ~n25311 ;
  assign n25313 = n25309 & n25312 ;
  assign n25314 = \wishbone_bd_ram_mem0_reg[59][3]/P0001  & n13613 ;
  assign n25315 = \wishbone_bd_ram_mem0_reg[249][3]/P0001  & n13431 ;
  assign n25316 = ~n25314 & ~n25315 ;
  assign n25317 = \wishbone_bd_ram_mem0_reg[8][3]/P0001  & n13459 ;
  assign n25318 = \wishbone_bd_ram_mem0_reg[81][3]/P0001  & n13409 ;
  assign n25319 = ~n25317 & ~n25318 ;
  assign n25320 = n25316 & n25319 ;
  assign n25321 = n25313 & n25320 ;
  assign n25322 = n25306 & n25321 ;
  assign n25323 = \wishbone_bd_ram_mem0_reg[131][3]/P0001  & n13358 ;
  assign n25324 = \wishbone_bd_ram_mem0_reg[155][3]/P0001  & n13738 ;
  assign n25325 = ~n25323 & ~n25324 ;
  assign n25326 = \wishbone_bd_ram_mem0_reg[222][3]/P0001  & n13721 ;
  assign n25327 = \wishbone_bd_ram_mem0_reg[46][3]/P0001  & n13298 ;
  assign n25328 = ~n25326 & ~n25327 ;
  assign n25329 = n25325 & n25328 ;
  assign n25330 = \wishbone_bd_ram_mem0_reg[150][3]/P0001  & n13666 ;
  assign n25331 = \wishbone_bd_ram_mem0_reg[207][3]/P0001  & n13826 ;
  assign n25332 = ~n25330 & ~n25331 ;
  assign n25333 = \wishbone_bd_ram_mem0_reg[7][3]/P0001  & n13546 ;
  assign n25334 = \wishbone_bd_ram_mem0_reg[142][3]/P0001  & n13448 ;
  assign n25335 = ~n25333 & ~n25334 ;
  assign n25336 = n25332 & n25335 ;
  assign n25337 = n25329 & n25336 ;
  assign n25338 = \wishbone_bd_ram_mem0_reg[235][3]/P0001  & n13518 ;
  assign n25339 = \wishbone_bd_ram_mem0_reg[99][3]/P0001  & n13996 ;
  assign n25340 = ~n25338 & ~n25339 ;
  assign n25341 = \wishbone_bd_ram_mem0_reg[147][3]/P0001  & n13702 ;
  assign n25342 = \wishbone_bd_ram_mem0_reg[206][3]/P0001  & n13414 ;
  assign n25343 = ~n25341 & ~n25342 ;
  assign n25344 = n25340 & n25343 ;
  assign n25345 = \wishbone_bd_ram_mem0_reg[242][3]/P0001  & n13383 ;
  assign n25346 = \wishbone_bd_ram_mem0_reg[238][3]/P0001  & n13819 ;
  assign n25347 = ~n25345 & ~n25346 ;
  assign n25348 = \wishbone_bd_ram_mem0_reg[130][3]/P0001  & n13427 ;
  assign n25349 = \wishbone_bd_ram_mem0_reg[141][3]/P0001  & n13852 ;
  assign n25350 = ~n25348 & ~n25349 ;
  assign n25351 = n25347 & n25350 ;
  assign n25352 = n25344 & n25351 ;
  assign n25353 = n25337 & n25352 ;
  assign n25354 = n25322 & n25353 ;
  assign n25355 = n25291 & n25354 ;
  assign n25356 = n25228 & n25355 ;
  assign n25357 = \wishbone_bd_ram_mem0_reg[2][3]/P0001  & n13975 ;
  assign n25358 = \wishbone_bd_ram_mem0_reg[69][3]/P0001  & n13487 ;
  assign n25359 = ~n25357 & ~n25358 ;
  assign n25360 = \wishbone_bd_ram_mem0_reg[152][3]/P0001  & n13912 ;
  assign n25361 = \wishbone_bd_ram_mem0_reg[253][3]/P0001  & n13708 ;
  assign n25362 = ~n25360 & ~n25361 ;
  assign n25363 = n25359 & n25362 ;
  assign n25364 = \wishbone_bd_ram_mem0_reg[29][3]/P0001  & n13412 ;
  assign n25365 = \wishbone_bd_ram_mem0_reg[72][3]/P0001  & n13582 ;
  assign n25366 = ~n25364 & ~n25365 ;
  assign n25367 = \wishbone_bd_ram_mem0_reg[250][3]/P0001  & n13677 ;
  assign n25368 = \wishbone_bd_ram_mem0_reg[71][3]/P0001  & n13636 ;
  assign n25369 = ~n25367 & ~n25368 ;
  assign n25370 = n25366 & n25369 ;
  assign n25371 = n25363 & n25370 ;
  assign n25372 = \wishbone_bd_ram_mem0_reg[84][3]/P0001  & n13385 ;
  assign n25373 = \wishbone_bd_ram_mem0_reg[50][3]/P0001  & n13686 ;
  assign n25374 = ~n25372 & ~n25373 ;
  assign n25375 = \wishbone_bd_ram_mem0_reg[68][3]/P0001  & n13379 ;
  assign n25376 = \wishbone_bd_ram_mem0_reg[219][3]/P0001  & n13577 ;
  assign n25377 = ~n25375 & ~n25376 ;
  assign n25378 = n25374 & n25377 ;
  assign n25379 = \wishbone_bd_ram_mem0_reg[161][3]/P0001  & n13505 ;
  assign n25380 = \wishbone_bd_ram_mem0_reg[95][3]/P0001  & n13317 ;
  assign n25381 = ~n25379 & ~n25380 ;
  assign n25382 = \wishbone_bd_ram_mem0_reg[132][3]/P0001  & n13927 ;
  assign n25383 = \wishbone_bd_ram_mem0_reg[41][3]/P0001  & n14017 ;
  assign n25384 = ~n25382 & ~n25383 ;
  assign n25385 = n25381 & n25384 ;
  assign n25386 = n25378 & n25385 ;
  assign n25387 = n25371 & n25386 ;
  assign n25388 = \wishbone_bd_ram_mem0_reg[227][3]/P0001  & n13388 ;
  assign n25389 = \wishbone_bd_ram_mem0_reg[33][3]/P0001  & n13933 ;
  assign n25390 = ~n25388 & ~n25389 ;
  assign n25391 = \wishbone_bd_ram_mem0_reg[13][3]/P0001  & n13844 ;
  assign n25392 = \wishbone_bd_ram_mem0_reg[177][3]/P0001  & n13863 ;
  assign n25393 = ~n25391 & ~n25392 ;
  assign n25394 = n25390 & n25393 ;
  assign n25395 = \wishbone_bd_ram_mem0_reg[201][3]/P0001  & n13600 ;
  assign n25396 = \wishbone_bd_ram_mem0_reg[195][3]/P0001  & n13700 ;
  assign n25397 = ~n25395 & ~n25396 ;
  assign n25398 = \wishbone_bd_ram_mem0_reg[188][3]/P0001  & n13407 ;
  assign n25399 = \wishbone_bd_ram_mem0_reg[165][3]/P0001  & n14028 ;
  assign n25400 = ~n25398 & ~n25399 ;
  assign n25401 = n25397 & n25400 ;
  assign n25402 = n25394 & n25401 ;
  assign n25403 = \wishbone_bd_ram_mem0_reg[60][3]/P0001  & n13790 ;
  assign n25404 = \wishbone_bd_ram_mem0_reg[18][3]/P0001  & n13532 ;
  assign n25405 = ~n25403 & ~n25404 ;
  assign n25406 = \wishbone_bd_ram_mem0_reg[25][3]/P0001  & n13742 ;
  assign n25407 = \wishbone_bd_ram_mem0_reg[124][3]/P0001  & n14024 ;
  assign n25408 = ~n25406 & ~n25407 ;
  assign n25409 = n25405 & n25408 ;
  assign n25410 = \wishbone_bd_ram_mem0_reg[10][3]/P0001  & n13837 ;
  assign n25411 = \wishbone_bd_ram_mem0_reg[23][3]/P0001  & n13857 ;
  assign n25412 = ~n25410 & ~n25411 ;
  assign n25413 = \wishbone_bd_ram_mem0_reg[22][3]/P0001  & n13744 ;
  assign n25414 = \wishbone_bd_ram_mem0_reg[134][3]/P0001  & n13494 ;
  assign n25415 = ~n25413 & ~n25414 ;
  assign n25416 = n25412 & n25415 ;
  assign n25417 = n25409 & n25416 ;
  assign n25418 = n25402 & n25417 ;
  assign n25419 = n25387 & n25418 ;
  assign n25420 = \wishbone_bd_ram_mem0_reg[254][3]/P0001  & n13283 ;
  assign n25421 = \wishbone_bd_ram_mem0_reg[6][3]/P0001  & n13915 ;
  assign n25422 = ~n25420 & ~n25421 ;
  assign n25423 = \wishbone_bd_ram_mem0_reg[88][3]/P0001  & n13347 ;
  assign n25424 = \wishbone_bd_ram_mem0_reg[203][3]/P0001  & n13816 ;
  assign n25425 = ~n25423 & ~n25424 ;
  assign n25426 = n25422 & n25425 ;
  assign n25427 = \wishbone_bd_ram_mem0_reg[163][3]/P0001  & n13255 ;
  assign n25428 = \wishbone_bd_ram_mem0_reg[103][3]/P0001  & n13320 ;
  assign n25429 = ~n25427 & ~n25428 ;
  assign n25430 = \wishbone_bd_ram_mem0_reg[100][3]/P0001  & n13401 ;
  assign n25431 = \wishbone_bd_ram_mem0_reg[159][3]/P0001  & n13627 ;
  assign n25432 = ~n25430 & ~n25431 ;
  assign n25433 = n25429 & n25432 ;
  assign n25434 = n25426 & n25433 ;
  assign n25435 = \wishbone_bd_ram_mem0_reg[104][3]/P0001  & n13684 ;
  assign n25436 = \wishbone_bd_ram_mem0_reg[176][3]/P0001  & n13262 ;
  assign n25437 = ~n25435 & ~n25436 ;
  assign n25438 = \wishbone_bd_ram_mem0_reg[80][3]/P0001  & n13516 ;
  assign n25439 = \wishbone_bd_ram_mem0_reg[200][3]/P0001  & n13922 ;
  assign n25440 = ~n25438 & ~n25439 ;
  assign n25441 = n25437 & n25440 ;
  assign n25442 = \wishbone_bd_ram_mem0_reg[26][3]/P0001  & n13521 ;
  assign n25443 = \wishbone_bd_ram_mem0_reg[218][3]/P0001  & n13792 ;
  assign n25444 = ~n25442 & ~n25443 ;
  assign n25445 = \wishbone_bd_ram_mem0_reg[82][3]/P0001  & n13374 ;
  assign n25446 = \wishbone_bd_ram_mem0_reg[19][3]/P0001  & n13886 ;
  assign n25447 = ~n25445 & ~n25446 ;
  assign n25448 = n25444 & n25447 ;
  assign n25449 = n25441 & n25448 ;
  assign n25450 = n25434 & n25449 ;
  assign n25451 = \wishbone_bd_ram_mem0_reg[205][3]/P0001  & n13947 ;
  assign n25452 = \wishbone_bd_ram_mem0_reg[255][3]/P0001  & n13952 ;
  assign n25453 = ~n25451 & ~n25452 ;
  assign n25454 = \wishbone_bd_ram_mem0_reg[45][3]/P0001  & n13420 ;
  assign n25455 = \wishbone_bd_ram_mem0_reg[15][3]/P0001  & n13797 ;
  assign n25456 = ~n25454 & ~n25455 ;
  assign n25457 = n25453 & n25456 ;
  assign n25458 = \wishbone_bd_ram_mem0_reg[192][3]/P0001  & n13390 ;
  assign n25459 = \wishbone_bd_ram_mem0_reg[126][3]/P0001  & n13786 ;
  assign n25460 = ~n25458 & ~n25459 ;
  assign n25461 = \wishbone_bd_ram_mem0_reg[240][3]/P0001  & n13352 ;
  assign n25462 = \wishbone_bd_ram_mem0_reg[113][3]/P0001  & n13882 ;
  assign n25463 = ~n25461 & ~n25462 ;
  assign n25464 = n25460 & n25463 ;
  assign n25465 = n25457 & n25464 ;
  assign n25466 = \wishbone_bd_ram_mem0_reg[252][3]/P0001  & n13986 ;
  assign n25467 = \wishbone_bd_ram_mem0_reg[34][3]/P0001  & n13450 ;
  assign n25468 = ~n25466 & ~n25467 ;
  assign n25469 = \wishbone_bd_ram_mem0_reg[73][3]/P0001  & n13456 ;
  assign n25470 = \wishbone_bd_ram_mem0_reg[234][3]/P0001  & n13781 ;
  assign n25471 = ~n25469 & ~n25470 ;
  assign n25472 = n25468 & n25471 ;
  assign n25473 = \wishbone_bd_ram_mem0_reg[35][3]/P0001  & n13523 ;
  assign n25474 = \wishbone_bd_ram_mem0_reg[62][3]/P0001  & n13529 ;
  assign n25475 = ~n25473 & ~n25474 ;
  assign n25476 = \wishbone_bd_ram_mem0_reg[67][3]/P0001  & n13663 ;
  assign n25477 = \wishbone_bd_ram_mem0_reg[16][3]/P0001  & n13695 ;
  assign n25478 = ~n25476 & ~n25477 ;
  assign n25479 = n25475 & n25478 ;
  assign n25480 = n25472 & n25479 ;
  assign n25481 = n25465 & n25480 ;
  assign n25482 = n25450 & n25481 ;
  assign n25483 = n25419 & n25482 ;
  assign n25484 = \wishbone_bd_ram_mem0_reg[20][3]/P0001  & n13839 ;
  assign n25485 = \wishbone_bd_ram_mem0_reg[112][3]/P0001  & n13482 ;
  assign n25486 = ~n25484 & ~n25485 ;
  assign n25487 = \wishbone_bd_ram_mem0_reg[208][3]/P0001  & n14010 ;
  assign n25488 = \wishbone_bd_ram_mem0_reg[169][3]/P0001  & n13541 ;
  assign n25489 = ~n25487 & ~n25488 ;
  assign n25490 = n25486 & n25489 ;
  assign n25491 = \wishbone_bd_ram_mem0_reg[121][3]/P0001  & n13983 ;
  assign n25492 = \wishbone_bd_ram_mem0_reg[138][3]/P0001  & n13398 ;
  assign n25493 = ~n25491 & ~n25492 ;
  assign n25494 = \wishbone_bd_ram_mem0_reg[47][3]/P0001  & n13436 ;
  assign n25495 = \wishbone_bd_ram_mem0_reg[251][3]/P0001  & n14019 ;
  assign n25496 = ~n25494 & ~n25495 ;
  assign n25497 = n25493 & n25496 ;
  assign n25498 = n25490 & n25497 ;
  assign n25499 = \wishbone_bd_ram_mem0_reg[214][3]/P0001  & n13938 ;
  assign n25500 = \wishbone_bd_ram_mem0_reg[213][3]/P0001  & n13870 ;
  assign n25501 = ~n25499 & ~n25500 ;
  assign n25502 = \wishbone_bd_ram_mem0_reg[51][3]/P0001  & n13880 ;
  assign n25503 = \wishbone_bd_ram_mem0_reg[220][3]/P0001  & n13965 ;
  assign n25504 = ~n25502 & ~n25503 ;
  assign n25505 = n25501 & n25504 ;
  assign n25506 = \wishbone_bd_ram_mem0_reg[55][3]/P0001  & n13618 ;
  assign n25507 = \wishbone_bd_ram_mem0_reg[24][3]/P0001  & n13970 ;
  assign n25508 = ~n25506 & ~n25507 ;
  assign n25509 = \wishbone_bd_ram_mem0_reg[168][3]/P0001  & n13795 ;
  assign n25510 = \wishbone_bd_ram_mem0_reg[118][3]/P0001  & n13589 ;
  assign n25511 = ~n25509 & ~n25510 ;
  assign n25512 = n25508 & n25511 ;
  assign n25513 = n25505 & n25512 ;
  assign n25514 = n25498 & n25513 ;
  assign n25515 = \wishbone_bd_ram_mem0_reg[90][3]/P0001  & n13906 ;
  assign n25516 = \wishbone_bd_ram_mem0_reg[75][3]/P0001  & n13605 ;
  assign n25517 = ~n25515 & ~n25516 ;
  assign n25518 = \wishbone_bd_ram_mem0_reg[61][3]/P0001  & n13544 ;
  assign n25519 = \wishbone_bd_ram_mem0_reg[171][3]/P0001  & n13422 ;
  assign n25520 = ~n25518 & ~n25519 ;
  assign n25521 = n25517 & n25520 ;
  assign n25522 = \wishbone_bd_ram_mem0_reg[89][3]/P0001  & n13910 ;
  assign n25523 = \wishbone_bd_ram_mem0_reg[54][3]/P0001  & n13622 ;
  assign n25524 = ~n25522 & ~n25523 ;
  assign n25525 = \wishbone_bd_ram_mem0_reg[31][3]/P0001  & n13758 ;
  assign n25526 = \wishbone_bd_ram_mem0_reg[172][3]/P0001  & n13377 ;
  assign n25527 = ~n25525 & ~n25526 ;
  assign n25528 = n25524 & n25527 ;
  assign n25529 = n25521 & n25528 ;
  assign n25530 = \wishbone_bd_ram_mem0_reg[114][3]/P0001  & n13763 ;
  assign n25531 = \wishbone_bd_ram_mem0_reg[237][3]/P0001  & n13924 ;
  assign n25532 = ~n25530 & ~n25531 ;
  assign n25533 = \wishbone_bd_ram_mem0_reg[158][3]/P0001  & n13294 ;
  assign n25534 = \wishbone_bd_ram_mem0_reg[173][3]/P0001  & n13360 ;
  assign n25535 = ~n25533 & ~n25534 ;
  assign n25536 = n25532 & n25535 ;
  assign n25537 = \wishbone_bd_ram_mem0_reg[27][3]/P0001  & n13251 ;
  assign n25538 = \wishbone_bd_ram_mem0_reg[166][3]/P0001  & n13999 ;
  assign n25539 = ~n25537 & ~n25538 ;
  assign n25540 = \wishbone_bd_ram_mem0_reg[53][3]/P0001  & n13875 ;
  assign n25541 = \wishbone_bd_ram_mem0_reg[129][3]/P0001  & n13629 ;
  assign n25542 = ~n25540 & ~n25541 ;
  assign n25543 = n25539 & n25542 ;
  assign n25544 = n25536 & n25543 ;
  assign n25545 = n25529 & n25544 ;
  assign n25546 = n25514 & n25545 ;
  assign n25547 = \wishbone_bd_ram_mem0_reg[178][3]/P0001  & n13301 ;
  assign n25548 = \wishbone_bd_ram_mem0_reg[170][3]/P0001  & n14007 ;
  assign n25549 = ~n25547 & ~n25548 ;
  assign n25550 = \wishbone_bd_ram_mem0_reg[191][3]/P0001  & n14012 ;
  assign n25551 = \wishbone_bd_ram_mem0_reg[91][3]/P0001  & n13954 ;
  assign n25552 = ~n25550 & ~n25551 ;
  assign n25553 = n25549 & n25552 ;
  assign n25554 = \wishbone_bd_ram_mem0_reg[145][3]/P0001  & n13715 ;
  assign n25555 = \wishbone_bd_ram_mem0_reg[110][3]/P0001  & n14030 ;
  assign n25556 = ~n25554 & ~n25555 ;
  assign n25557 = \wishbone_bd_ram_mem0_reg[116][3]/P0001  & n13865 ;
  assign n25558 = \wishbone_bd_ram_mem0_reg[204][3]/P0001  & n13821 ;
  assign n25559 = ~n25557 & ~n25558 ;
  assign n25560 = n25556 & n25559 ;
  assign n25561 = n25553 & n25560 ;
  assign n25562 = \wishbone_bd_ram_mem0_reg[1][3]/P0001  & n13888 ;
  assign n25563 = \wishbone_bd_ram_mem0_reg[66][3]/P0001  & n13603 ;
  assign n25564 = ~n25562 & ~n25563 ;
  assign n25565 = \wishbone_bd_ram_mem0_reg[52][3]/P0001  & n13988 ;
  assign n25566 = \wishbone_bd_ram_mem0_reg[232][3]/P0001  & n13510 ;
  assign n25567 = ~n25565 & ~n25566 ;
  assign n25568 = n25564 & n25567 ;
  assign n25569 = \wishbone_bd_ram_mem0_reg[127][3]/P0001  & n13803 ;
  assign n25570 = \wishbone_bd_ram_mem0_reg[107][3]/P0001  & n13476 ;
  assign n25571 = ~n25569 & ~n25570 ;
  assign n25572 = \wishbone_bd_ram_mem0_reg[233][3]/P0001  & n13332 ;
  assign n25573 = \wishbone_bd_ram_mem0_reg[0][3]/P0001  & n13539 ;
  assign n25574 = ~n25572 & ~n25573 ;
  assign n25575 = n25571 & n25574 ;
  assign n25576 = n25568 & n25575 ;
  assign n25577 = n25561 & n25576 ;
  assign n25578 = \wishbone_bd_ram_mem0_reg[143][3]/P0001  & n13461 ;
  assign n25579 = \wishbone_bd_ram_mem0_reg[63][3]/P0001  & n13327 ;
  assign n25580 = ~n25578 & ~n25579 ;
  assign n25581 = \wishbone_bd_ram_mem0_reg[77][3]/P0001  & n13935 ;
  assign n25582 = \wishbone_bd_ram_mem0_reg[230][3]/P0001  & n13994 ;
  assign n25583 = ~n25581 & ~n25582 ;
  assign n25584 = n25580 & n25583 ;
  assign n25585 = \wishbone_bd_ram_mem0_reg[70][3]/P0001  & n13339 ;
  assign n25586 = \wishbone_bd_ram_mem0_reg[58][3]/P0001  & n13949 ;
  assign n25587 = ~n25585 & ~n25586 ;
  assign n25588 = \wishbone_bd_ram_mem0_reg[136][3]/P0001  & n13963 ;
  assign n25589 = \wishbone_bd_ram_mem0_reg[224][3]/P0001  & n13433 ;
  assign n25590 = ~n25588 & ~n25589 ;
  assign n25591 = n25587 & n25590 ;
  assign n25592 = n25584 & n25591 ;
  assign n25593 = \wishbone_bd_ram_mem0_reg[36][3]/P0001  & n13639 ;
  assign n25594 = \wishbone_bd_ram_mem0_reg[245][3]/P0001  & n13877 ;
  assign n25595 = ~n25593 & ~n25594 ;
  assign n25596 = \wishbone_bd_ram_mem0_reg[56][3]/P0001  & n13611 ;
  assign n25597 = \wishbone_bd_ram_mem0_reg[193][3]/P0001  & n14022 ;
  assign n25598 = ~n25596 & ~n25597 ;
  assign n25599 = n25595 & n25598 ;
  assign n25600 = \wishbone_bd_ram_mem0_reg[217][3]/P0001  & n13767 ;
  assign n25601 = \wishbone_bd_ram_mem0_reg[154][3]/P0001  & n13403 ;
  assign n25602 = ~n25600 & ~n25601 ;
  assign n25603 = \wishbone_bd_ram_mem0_reg[42][3]/P0001  & n13341 ;
  assign n25604 = \wishbone_bd_ram_mem0_reg[183][3]/P0001  & n13645 ;
  assign n25605 = ~n25603 & ~n25604 ;
  assign n25606 = n25602 & n25605 ;
  assign n25607 = n25599 & n25606 ;
  assign n25608 = n25592 & n25607 ;
  assign n25609 = n25577 & n25608 ;
  assign n25610 = n25546 & n25609 ;
  assign n25611 = n25483 & n25610 ;
  assign n25612 = n25356 & n25611 ;
  assign n25613 = ~wb_rst_i_pad & ~n25100 ;
  assign n25614 = ~n25612 & n25613 ;
  assign n25615 = ~n25101 & ~n25614 ;
  assign n25616 = \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131  & n25082 ;
  assign n25617 = \ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131  & n23782 ;
  assign n25618 = ~n25616 & ~n25617 ;
  assign n25619 = \ethreg1_MODER_0_DataOut_reg[4]/NET0131  & n23808 ;
  assign n25620 = \ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131  & n23743 ;
  assign n25621 = n23741 & n25620 ;
  assign n25622 = ~n25619 & ~n25621 ;
  assign n25623 = n25618 & n25622 ;
  assign n25624 = \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  & n23737 ;
  assign n25625 = \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  & n25059 ;
  assign n25626 = ~n25624 & ~n25625 ;
  assign n25627 = n25623 & n25626 ;
  assign n25628 = \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131  & n23813 ;
  assign n25629 = \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131  & n25069 ;
  assign n25630 = ~n25628 & ~n25629 ;
  assign n25631 = \ethreg1_IPGT_0_DataOut_reg[4]/NET0131  & n25090 ;
  assign n25632 = \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131  & n25079 ;
  assign n25633 = ~n25631 & ~n25632 ;
  assign n25634 = n25630 & n25633 ;
  assign n25635 = n23730 & n25634 ;
  assign n25636 = \ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131  & n23743 ;
  assign n25637 = n23747 & n25636 ;
  assign n25638 = \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  & n23751 ;
  assign n25639 = n23741 & n25638 ;
  assign n25640 = ~n25637 & ~n25639 ;
  assign n25641 = \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  & n23751 ;
  assign n25642 = n23747 & n25641 ;
  assign n25643 = \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131  & n25088 ;
  assign n25644 = ~n25642 & ~n25643 ;
  assign n25645 = n25640 & n25644 ;
  assign n25646 = \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131  & n23794 ;
  assign n25647 = n23741 & n25646 ;
  assign n25648 = \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  & n25084 ;
  assign n25649 = ~n25647 & ~n25648 ;
  assign n25650 = \ethreg1_irq_busy_reg/NET0131  & n25064 ;
  assign n25651 = \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131  & n23802 ;
  assign n25652 = ~n25650 & ~n25651 ;
  assign n25653 = n25649 & n25652 ;
  assign n25654 = n25645 & n25653 ;
  assign n25655 = n25635 & n25654 ;
  assign n25656 = n25627 & n25655 ;
  assign n25657 = n23730 & ~n25656 ;
  assign n25658 = \wishbone_bd_ram_mem0_reg[61][4]/P0001  & n13544 ;
  assign n25659 = \wishbone_bd_ram_mem0_reg[72][4]/P0001  & n13582 ;
  assign n25660 = ~n25658 & ~n25659 ;
  assign n25661 = \wishbone_bd_ram_mem0_reg[9][4]/P0001  & n13580 ;
  assign n25662 = \wishbone_bd_ram_mem0_reg[35][4]/P0001  & n13523 ;
  assign n25663 = ~n25661 & ~n25662 ;
  assign n25664 = n25660 & n25663 ;
  assign n25665 = \wishbone_bd_ram_mem0_reg[54][4]/P0001  & n13622 ;
  assign n25666 = \wishbone_bd_ram_mem0_reg[87][4]/P0001  & n13691 ;
  assign n25667 = ~n25665 & ~n25666 ;
  assign n25668 = \wishbone_bd_ram_mem0_reg[119][4]/P0001  & n14033 ;
  assign n25669 = \wishbone_bd_ram_mem0_reg[37][4]/P0001  & n13710 ;
  assign n25670 = ~n25668 & ~n25669 ;
  assign n25671 = n25667 & n25670 ;
  assign n25672 = n25664 & n25671 ;
  assign n25673 = \wishbone_bd_ram_mem0_reg[48][4]/P0001  & n13917 ;
  assign n25674 = \wishbone_bd_ram_mem0_reg[95][4]/P0001  & n13317 ;
  assign n25675 = ~n25673 & ~n25674 ;
  assign n25676 = \wishbone_bd_ram_mem0_reg[62][4]/P0001  & n13529 ;
  assign n25677 = \wishbone_bd_ram_mem0_reg[139][4]/P0001  & n13566 ;
  assign n25678 = ~n25676 & ~n25677 ;
  assign n25679 = n25675 & n25678 ;
  assign n25680 = \wishbone_bd_ram_mem0_reg[22][4]/P0001  & n13744 ;
  assign n25681 = \wishbone_bd_ram_mem0_reg[187][4]/P0001  & n13756 ;
  assign n25682 = ~n25680 & ~n25681 ;
  assign n25683 = \wishbone_bd_ram_mem0_reg[25][4]/P0001  & n13742 ;
  assign n25684 = \wishbone_bd_ram_mem0_reg[146][4]/P0001  & n13958 ;
  assign n25685 = ~n25683 & ~n25684 ;
  assign n25686 = n25682 & n25685 ;
  assign n25687 = n25679 & n25686 ;
  assign n25688 = n25672 & n25687 ;
  assign n25689 = \wishbone_bd_ram_mem0_reg[145][4]/P0001  & n13715 ;
  assign n25690 = \wishbone_bd_ram_mem0_reg[107][4]/P0001  & n13476 ;
  assign n25691 = ~n25689 & ~n25690 ;
  assign n25692 = \wishbone_bd_ram_mem0_reg[106][4]/P0001  & n13555 ;
  assign n25693 = \wishbone_bd_ram_mem0_reg[129][4]/P0001  & n13629 ;
  assign n25694 = ~n25692 & ~n25693 ;
  assign n25695 = n25691 & n25694 ;
  assign n25696 = \wishbone_bd_ram_mem0_reg[226][4]/P0001  & n13668 ;
  assign n25697 = \wishbone_bd_ram_mem0_reg[243][4]/P0001  & n13575 ;
  assign n25698 = ~n25696 & ~n25697 ;
  assign n25699 = \wishbone_bd_ram_mem0_reg[36][4]/P0001  & n13639 ;
  assign n25700 = \wishbone_bd_ram_mem0_reg[17][4]/P0001  & n13324 ;
  assign n25701 = ~n25699 & ~n25700 ;
  assign n25702 = n25698 & n25701 ;
  assign n25703 = n25695 & n25702 ;
  assign n25704 = \wishbone_bd_ram_mem0_reg[231][4]/P0001  & n13363 ;
  assign n25705 = \wishbone_bd_ram_mem0_reg[253][4]/P0001  & n13708 ;
  assign n25706 = ~n25704 & ~n25705 ;
  assign n25707 = \wishbone_bd_ram_mem0_reg[225][4]/P0001  & n13719 ;
  assign n25708 = \wishbone_bd_ram_mem0_reg[5][4]/P0001  & n13243 ;
  assign n25709 = ~n25707 & ~n25708 ;
  assign n25710 = n25706 & n25709 ;
  assign n25711 = \wishbone_bd_ram_mem0_reg[12][4]/P0001  & n13733 ;
  assign n25712 = \wishbone_bd_ram_mem0_reg[244][4]/P0001  & n13474 ;
  assign n25713 = ~n25711 & ~n25712 ;
  assign n25714 = \wishbone_bd_ram_mem0_reg[143][4]/P0001  & n13461 ;
  assign n25715 = \wishbone_bd_ram_mem0_reg[97][4]/P0001  & n13724 ;
  assign n25716 = ~n25714 & ~n25715 ;
  assign n25717 = n25713 & n25716 ;
  assign n25718 = n25710 & n25717 ;
  assign n25719 = n25703 & n25718 ;
  assign n25720 = n25688 & n25719 ;
  assign n25721 = \wishbone_bd_ram_mem0_reg[179][4]/P0001  & n14035 ;
  assign n25722 = \wishbone_bd_ram_mem0_reg[184][4]/P0001  & n13960 ;
  assign n25723 = ~n25721 & ~n25722 ;
  assign n25724 = \wishbone_bd_ram_mem0_reg[237][4]/P0001  & n13924 ;
  assign n25725 = \wishbone_bd_ram_mem0_reg[21][4]/P0001  & n13438 ;
  assign n25726 = ~n25724 & ~n25725 ;
  assign n25727 = n25723 & n25726 ;
  assign n25728 = \wishbone_bd_ram_mem0_reg[236][4]/P0001  & n13480 ;
  assign n25729 = \wishbone_bd_ram_mem0_reg[157][4]/P0001  & n13445 ;
  assign n25730 = ~n25728 & ~n25729 ;
  assign n25731 = \wishbone_bd_ram_mem0_reg[111][4]/P0001  & n13471 ;
  assign n25732 = \wishbone_bd_ram_mem0_reg[49][4]/P0001  & n13929 ;
  assign n25733 = ~n25731 & ~n25732 ;
  assign n25734 = n25730 & n25733 ;
  assign n25735 = n25727 & n25734 ;
  assign n25736 = \wishbone_bd_ram_mem0_reg[86][4]/P0001  & n13485 ;
  assign n25737 = \wishbone_bd_ram_mem0_reg[14][4]/P0001  & n13972 ;
  assign n25738 = ~n25736 & ~n25737 ;
  assign n25739 = \wishbone_bd_ram_mem0_reg[116][4]/P0001  & n13865 ;
  assign n25740 = \wishbone_bd_ram_mem0_reg[186][4]/P0001  & n13616 ;
  assign n25741 = ~n25739 & ~n25740 ;
  assign n25742 = n25738 & n25741 ;
  assign n25743 = \wishbone_bd_ram_mem0_reg[165][4]/P0001  & n14028 ;
  assign n25744 = \wishbone_bd_ram_mem0_reg[147][4]/P0001  & n13702 ;
  assign n25745 = ~n25743 & ~n25744 ;
  assign n25746 = \wishbone_bd_ram_mem0_reg[38][4]/P0001  & n13828 ;
  assign n25747 = \wishbone_bd_ram_mem0_reg[233][4]/P0001  & n13332 ;
  assign n25748 = ~n25746 & ~n25747 ;
  assign n25749 = n25745 & n25748 ;
  assign n25750 = n25742 & n25749 ;
  assign n25751 = n25735 & n25750 ;
  assign n25752 = \wishbone_bd_ram_mem0_reg[55][4]/P0001  & n13618 ;
  assign n25753 = \wishbone_bd_ram_mem0_reg[77][4]/P0001  & n13935 ;
  assign n25754 = ~n25752 & ~n25753 ;
  assign n25755 = \wishbone_bd_ram_mem0_reg[153][4]/P0001  & n13309 ;
  assign n25756 = \wishbone_bd_ram_mem0_reg[192][4]/P0001  & n13390 ;
  assign n25757 = ~n25755 & ~n25756 ;
  assign n25758 = n25754 & n25757 ;
  assign n25759 = \wishbone_bd_ram_mem0_reg[215][4]/P0001  & n13901 ;
  assign n25760 = \wishbone_bd_ram_mem0_reg[175][4]/P0001  & n13674 ;
  assign n25761 = ~n25759 & ~n25760 ;
  assign n25762 = \wishbone_bd_ram_mem0_reg[60][4]/P0001  & n13790 ;
  assign n25763 = \wishbone_bd_ram_mem0_reg[193][4]/P0001  & n14022 ;
  assign n25764 = ~n25762 & ~n25763 ;
  assign n25765 = n25761 & n25764 ;
  assign n25766 = n25758 & n25765 ;
  assign n25767 = \wishbone_bd_ram_mem0_reg[196][4]/P0001  & n13977 ;
  assign n25768 = \wishbone_bd_ram_mem0_reg[135][4]/P0001  & n13672 ;
  assign n25769 = ~n25767 & ~n25768 ;
  assign n25770 = \wishbone_bd_ram_mem0_reg[82][4]/P0001  & n13374 ;
  assign n25771 = \wishbone_bd_ram_mem0_reg[166][4]/P0001  & n13999 ;
  assign n25772 = ~n25770 & ~n25771 ;
  assign n25773 = n25769 & n25772 ;
  assign n25774 = \wishbone_bd_ram_mem0_reg[51][4]/P0001  & n13880 ;
  assign n25775 = \wishbone_bd_ram_mem0_reg[206][4]/P0001  & n13414 ;
  assign n25776 = ~n25774 & ~n25775 ;
  assign n25777 = \wishbone_bd_ram_mem0_reg[173][4]/P0001  & n13360 ;
  assign n25778 = \wishbone_bd_ram_mem0_reg[39][4]/P0001  & n13893 ;
  assign n25779 = ~n25777 & ~n25778 ;
  assign n25780 = n25776 & n25779 ;
  assign n25781 = n25773 & n25780 ;
  assign n25782 = n25766 & n25781 ;
  assign n25783 = n25751 & n25782 ;
  assign n25784 = n25720 & n25783 ;
  assign n25785 = \wishbone_bd_ram_mem0_reg[141][4]/P0001  & n13852 ;
  assign n25786 = \wishbone_bd_ram_mem0_reg[133][4]/P0001  & n13492 ;
  assign n25787 = ~n25785 & ~n25786 ;
  assign n25788 = \wishbone_bd_ram_mem0_reg[199][4]/P0001  & n13499 ;
  assign n25789 = \wishbone_bd_ram_mem0_reg[120][4]/P0001  & n13550 ;
  assign n25790 = ~n25788 & ~n25789 ;
  assign n25791 = n25787 & n25790 ;
  assign n25792 = \wishbone_bd_ram_mem0_reg[58][4]/P0001  & n13949 ;
  assign n25793 = \wishbone_bd_ram_mem0_reg[101][4]/P0001  & n13772 ;
  assign n25794 = ~n25792 & ~n25793 ;
  assign n25795 = \wishbone_bd_ram_mem0_reg[4][4]/P0001  & n13527 ;
  assign n25796 = \wishbone_bd_ram_mem0_reg[209][4]/P0001  & n13689 ;
  assign n25797 = ~n25795 & ~n25796 ;
  assign n25798 = n25794 & n25797 ;
  assign n25799 = n25791 & n25798 ;
  assign n25800 = \wishbone_bd_ram_mem0_reg[241][4]/P0001  & n13854 ;
  assign n25801 = \wishbone_bd_ram_mem0_reg[208][4]/P0001  & n14010 ;
  assign n25802 = ~n25800 & ~n25801 ;
  assign n25803 = \wishbone_bd_ram_mem0_reg[93][4]/P0001  & n13891 ;
  assign n25804 = \wishbone_bd_ram_mem0_reg[98][4]/P0001  & n13569 ;
  assign n25805 = ~n25803 & ~n25804 ;
  assign n25806 = n25802 & n25805 ;
  assign n25807 = \wishbone_bd_ram_mem0_reg[228][4]/P0001  & n13497 ;
  assign n25808 = \wishbone_bd_ram_mem0_reg[118][4]/P0001  & n13589 ;
  assign n25809 = ~n25807 & ~n25808 ;
  assign n25810 = \wishbone_bd_ram_mem0_reg[164][4]/P0001  & n13236 ;
  assign n25811 = \wishbone_bd_ram_mem0_reg[202][4]/P0001  & n13268 ;
  assign n25812 = ~n25810 & ~n25811 ;
  assign n25813 = n25809 & n25812 ;
  assign n25814 = n25806 & n25813 ;
  assign n25815 = n25799 & n25814 ;
  assign n25816 = \wishbone_bd_ram_mem0_reg[156][4]/P0001  & n13769 ;
  assign n25817 = \wishbone_bd_ram_mem0_reg[66][4]/P0001  & n13603 ;
  assign n25818 = ~n25816 & ~n25817 ;
  assign n25819 = \wishbone_bd_ram_mem0_reg[171][4]/P0001  & n13422 ;
  assign n25820 = \wishbone_bd_ram_mem0_reg[182][4]/P0001  & n13598 ;
  assign n25821 = ~n25819 & ~n25820 ;
  assign n25822 = n25818 & n25821 ;
  assign n25823 = \wishbone_bd_ram_mem0_reg[0][4]/P0001  & n13539 ;
  assign n25824 = \wishbone_bd_ram_mem0_reg[161][4]/P0001  & n13505 ;
  assign n25825 = ~n25823 & ~n25824 ;
  assign n25826 = \wishbone_bd_ram_mem0_reg[212][4]/P0001  & n13634 ;
  assign n25827 = \wishbone_bd_ram_mem0_reg[108][4]/P0001  & n13814 ;
  assign n25828 = ~n25826 & ~n25827 ;
  assign n25829 = n25825 & n25828 ;
  assign n25830 = n25822 & n25829 ;
  assign n25831 = \wishbone_bd_ram_mem0_reg[1][4]/P0001  & n13888 ;
  assign n25832 = \wishbone_bd_ram_mem0_reg[188][4]/P0001  & n13407 ;
  assign n25833 = ~n25831 & ~n25832 ;
  assign n25834 = \wishbone_bd_ram_mem0_reg[246][4]/P0001  & n13981 ;
  assign n25835 = \wishbone_bd_ram_mem0_reg[6][4]/P0001  & n13915 ;
  assign n25836 = ~n25834 & ~n25835 ;
  assign n25837 = n25833 & n25836 ;
  assign n25838 = \wishbone_bd_ram_mem0_reg[3][4]/P0001  & n13354 ;
  assign n25839 = \wishbone_bd_ram_mem0_reg[83][4]/P0001  & n13454 ;
  assign n25840 = ~n25838 & ~n25839 ;
  assign n25841 = \wishbone_bd_ram_mem0_reg[242][4]/P0001  & n13383 ;
  assign n25842 = \wishbone_bd_ram_mem0_reg[234][4]/P0001  & n13781 ;
  assign n25843 = ~n25841 & ~n25842 ;
  assign n25844 = n25840 & n25843 ;
  assign n25845 = n25837 & n25844 ;
  assign n25846 = n25830 & n25845 ;
  assign n25847 = n25815 & n25846 ;
  assign n25848 = \wishbone_bd_ram_mem0_reg[240][4]/P0001  & n13352 ;
  assign n25849 = \wishbone_bd_ram_mem0_reg[10][4]/P0001  & n13837 ;
  assign n25850 = ~n25848 & ~n25849 ;
  assign n25851 = \wishbone_bd_ram_mem0_reg[130][4]/P0001  & n13427 ;
  assign n25852 = \wishbone_bd_ram_mem0_reg[43][4]/P0001  & n13761 ;
  assign n25853 = ~n25851 & ~n25852 ;
  assign n25854 = n25850 & n25853 ;
  assign n25855 = \wishbone_bd_ram_mem0_reg[203][4]/P0001  & n13816 ;
  assign n25856 = \wishbone_bd_ram_mem0_reg[252][4]/P0001  & n13986 ;
  assign n25857 = ~n25855 & ~n25856 ;
  assign n25858 = \wishbone_bd_ram_mem0_reg[65][4]/P0001  & n13842 ;
  assign n25859 = \wishbone_bd_ram_mem0_reg[103][4]/P0001  & n13320 ;
  assign n25860 = ~n25858 & ~n25859 ;
  assign n25861 = n25857 & n25860 ;
  assign n25862 = n25854 & n25861 ;
  assign n25863 = \wishbone_bd_ram_mem0_reg[207][4]/P0001  & n13826 ;
  assign n25864 = \wishbone_bd_ram_mem0_reg[104][4]/P0001  & n13684 ;
  assign n25865 = ~n25863 & ~n25864 ;
  assign n25866 = \wishbone_bd_ram_mem0_reg[63][4]/P0001  & n13327 ;
  assign n25867 = \wishbone_bd_ram_mem0_reg[127][4]/P0001  & n13803 ;
  assign n25868 = ~n25866 & ~n25867 ;
  assign n25869 = n25865 & n25868 ;
  assign n25870 = \wishbone_bd_ram_mem0_reg[177][4]/P0001  & n13863 ;
  assign n25871 = \wishbone_bd_ram_mem0_reg[251][4]/P0001  & n14019 ;
  assign n25872 = ~n25870 & ~n25871 ;
  assign n25873 = \wishbone_bd_ram_mem0_reg[134][4]/P0001  & n13494 ;
  assign n25874 = \wishbone_bd_ram_mem0_reg[110][4]/P0001  & n14030 ;
  assign n25875 = ~n25873 & ~n25874 ;
  assign n25876 = n25872 & n25875 ;
  assign n25877 = n25869 & n25876 ;
  assign n25878 = n25862 & n25877 ;
  assign n25879 = \wishbone_bd_ram_mem0_reg[88][4]/P0001  & n13347 ;
  assign n25880 = \wishbone_bd_ram_mem0_reg[172][4]/P0001  & n13377 ;
  assign n25881 = ~n25879 & ~n25880 ;
  assign n25882 = \wishbone_bd_ram_mem0_reg[94][4]/P0001  & n13833 ;
  assign n25883 = \wishbone_bd_ram_mem0_reg[213][4]/P0001  & n13870 ;
  assign n25884 = ~n25882 & ~n25883 ;
  assign n25885 = n25881 & n25884 ;
  assign n25886 = \wishbone_bd_ram_mem0_reg[100][4]/P0001  & n13401 ;
  assign n25887 = \wishbone_bd_ram_mem0_reg[168][4]/P0001  & n13795 ;
  assign n25888 = ~n25886 & ~n25887 ;
  assign n25889 = \wishbone_bd_ram_mem0_reg[23][4]/P0001  & n13857 ;
  assign n25890 = \wishbone_bd_ram_mem0_reg[137][4]/P0001  & n13808 ;
  assign n25891 = ~n25889 & ~n25890 ;
  assign n25892 = n25888 & n25891 ;
  assign n25893 = n25885 & n25892 ;
  assign n25894 = \wishbone_bd_ram_mem0_reg[33][4]/P0001  & n13933 ;
  assign n25895 = \wishbone_bd_ram_mem0_reg[123][4]/P0001  & n13749 ;
  assign n25896 = ~n25894 & ~n25895 ;
  assign n25897 = \wishbone_bd_ram_mem0_reg[28][4]/P0001  & n13810 ;
  assign n25898 = \wishbone_bd_ram_mem0_reg[201][4]/P0001  & n13600 ;
  assign n25899 = ~n25897 & ~n25898 ;
  assign n25900 = n25896 & n25899 ;
  assign n25901 = \wishbone_bd_ram_mem0_reg[140][4]/P0001  & n13287 ;
  assign n25902 = \wishbone_bd_ram_mem0_reg[249][4]/P0001  & n13431 ;
  assign n25903 = ~n25901 & ~n25902 ;
  assign n25904 = \wishbone_bd_ram_mem0_reg[189][4]/P0001  & n14001 ;
  assign n25905 = \wishbone_bd_ram_mem0_reg[34][4]/P0001  & n13450 ;
  assign n25906 = ~n25904 & ~n25905 ;
  assign n25907 = n25903 & n25906 ;
  assign n25908 = n25900 & n25907 ;
  assign n25909 = n25893 & n25908 ;
  assign n25910 = n25878 & n25909 ;
  assign n25911 = n25847 & n25910 ;
  assign n25912 = n25784 & n25911 ;
  assign n25913 = \wishbone_bd_ram_mem0_reg[13][4]/P0001  & n13844 ;
  assign n25914 = \wishbone_bd_ram_mem0_reg[114][4]/P0001  & n13763 ;
  assign n25915 = ~n25913 & ~n25914 ;
  assign n25916 = \wishbone_bd_ram_mem0_reg[142][4]/P0001  & n13448 ;
  assign n25917 = \wishbone_bd_ram_mem0_reg[178][4]/P0001  & n13301 ;
  assign n25918 = ~n25916 & ~n25917 ;
  assign n25919 = n25915 & n25918 ;
  assign n25920 = \wishbone_bd_ram_mem0_reg[64][4]/P0001  & n13904 ;
  assign n25921 = \wishbone_bd_ram_mem0_reg[113][4]/P0001  & n13882 ;
  assign n25922 = ~n25920 & ~n25921 ;
  assign n25923 = \wishbone_bd_ram_mem0_reg[227][4]/P0001  & n13388 ;
  assign n25924 = \wishbone_bd_ram_mem0_reg[105][4]/P0001  & n13503 ;
  assign n25925 = ~n25923 & ~n25924 ;
  assign n25926 = n25922 & n25925 ;
  assign n25927 = n25919 & n25926 ;
  assign n25928 = \wishbone_bd_ram_mem0_reg[125][4]/P0001  & n13396 ;
  assign n25929 = \wishbone_bd_ram_mem0_reg[30][4]/P0001  & n13713 ;
  assign n25930 = ~n25928 & ~n25929 ;
  assign n25931 = \wishbone_bd_ram_mem0_reg[220][4]/P0001  & n13965 ;
  assign n25932 = \wishbone_bd_ram_mem0_reg[218][4]/P0001  & n13792 ;
  assign n25933 = ~n25931 & ~n25932 ;
  assign n25934 = n25930 & n25933 ;
  assign n25935 = \wishbone_bd_ram_mem0_reg[56][4]/P0001  & n13611 ;
  assign n25936 = \wishbone_bd_ram_mem0_reg[84][4]/P0001  & n13385 ;
  assign n25937 = ~n25935 & ~n25936 ;
  assign n25938 = \wishbone_bd_ram_mem0_reg[232][4]/P0001  & n13510 ;
  assign n25939 = \wishbone_bd_ram_mem0_reg[159][4]/P0001  & n13627 ;
  assign n25940 = ~n25938 & ~n25939 ;
  assign n25941 = n25937 & n25940 ;
  assign n25942 = n25934 & n25941 ;
  assign n25943 = n25927 & n25942 ;
  assign n25944 = \wishbone_bd_ram_mem0_reg[229][4]/P0001  & n13552 ;
  assign n25945 = \wishbone_bd_ram_mem0_reg[52][4]/P0001  & n13988 ;
  assign n25946 = ~n25944 & ~n25945 ;
  assign n25947 = \wishbone_bd_ram_mem0_reg[126][4]/P0001  & n13786 ;
  assign n25948 = \wishbone_bd_ram_mem0_reg[89][4]/P0001  & n13910 ;
  assign n25949 = ~n25947 & ~n25948 ;
  assign n25950 = n25946 & n25949 ;
  assign n25951 = \wishbone_bd_ram_mem0_reg[254][4]/P0001  & n13283 ;
  assign n25952 = \wishbone_bd_ram_mem0_reg[91][4]/P0001  & n13954 ;
  assign n25953 = ~n25951 & ~n25952 ;
  assign n25954 = \wishbone_bd_ram_mem0_reg[222][4]/P0001  & n13721 ;
  assign n25955 = \wishbone_bd_ram_mem0_reg[154][4]/P0001  & n13403 ;
  assign n25956 = ~n25954 & ~n25955 ;
  assign n25957 = n25953 & n25956 ;
  assign n25958 = n25950 & n25957 ;
  assign n25959 = \wishbone_bd_ram_mem0_reg[69][4]/P0001  & n13487 ;
  assign n25960 = \wishbone_bd_ram_mem0_reg[42][4]/P0001  & n13341 ;
  assign n25961 = ~n25959 & ~n25960 ;
  assign n25962 = \wishbone_bd_ram_mem0_reg[7][4]/P0001  & n13546 ;
  assign n25963 = \wishbone_bd_ram_mem0_reg[19][4]/P0001  & n13886 ;
  assign n25964 = ~n25962 & ~n25963 ;
  assign n25965 = n25961 & n25964 ;
  assign n25966 = \wishbone_bd_ram_mem0_reg[219][4]/P0001  & n13577 ;
  assign n25967 = \wishbone_bd_ram_mem0_reg[31][4]/P0001  & n13758 ;
  assign n25968 = ~n25966 & ~n25967 ;
  assign n25969 = \wishbone_bd_ram_mem0_reg[248][4]/P0001  & n13647 ;
  assign n25970 = \wishbone_bd_ram_mem0_reg[81][4]/P0001  & n13409 ;
  assign n25971 = ~n25969 & ~n25970 ;
  assign n25972 = n25968 & n25971 ;
  assign n25973 = n25965 & n25972 ;
  assign n25974 = n25958 & n25973 ;
  assign n25975 = n25943 & n25974 ;
  assign n25976 = \wishbone_bd_ram_mem0_reg[194][4]/P0001  & n13624 ;
  assign n25977 = \wishbone_bd_ram_mem0_reg[132][4]/P0001  & n13927 ;
  assign n25978 = ~n25976 & ~n25977 ;
  assign n25979 = \wishbone_bd_ram_mem0_reg[2][4]/P0001  & n13975 ;
  assign n25980 = \wishbone_bd_ram_mem0_reg[255][4]/P0001  & n13952 ;
  assign n25981 = ~n25979 & ~n25980 ;
  assign n25982 = n25978 & n25981 ;
  assign n25983 = \wishbone_bd_ram_mem0_reg[221][4]/P0001  & n13641 ;
  assign n25984 = \wishbone_bd_ram_mem0_reg[180][4]/P0001  & n13650 ;
  assign n25985 = ~n25983 & ~n25984 ;
  assign n25986 = \wishbone_bd_ram_mem0_reg[76][4]/P0001  & n13831 ;
  assign n25987 = \wishbone_bd_ram_mem0_reg[74][4]/P0001  & n13564 ;
  assign n25988 = ~n25986 & ~n25987 ;
  assign n25989 = n25985 & n25988 ;
  assign n25990 = n25982 & n25989 ;
  assign n25991 = \wishbone_bd_ram_mem0_reg[50][4]/P0001  & n13686 ;
  assign n25992 = \wishbone_bd_ram_mem0_reg[92][4]/P0001  & n13859 ;
  assign n25993 = ~n25991 & ~n25992 ;
  assign n25994 = \wishbone_bd_ram_mem0_reg[96][4]/P0001  & n13425 ;
  assign n25995 = \wishbone_bd_ram_mem0_reg[224][4]/P0001  & n13433 ;
  assign n25996 = ~n25994 & ~n25995 ;
  assign n25997 = n25993 & n25996 ;
  assign n25998 = \wishbone_bd_ram_mem0_reg[29][4]/P0001  & n13412 ;
  assign n25999 = \wishbone_bd_ram_mem0_reg[136][4]/P0001  & n13963 ;
  assign n26000 = ~n25998 & ~n25999 ;
  assign n26001 = \wishbone_bd_ram_mem0_reg[162][4]/P0001  & n13726 ;
  assign n26002 = \wishbone_bd_ram_mem0_reg[75][4]/P0001  & n13605 ;
  assign n26003 = ~n26001 & ~n26002 ;
  assign n26004 = n26000 & n26003 ;
  assign n26005 = n25997 & n26004 ;
  assign n26006 = n25990 & n26005 ;
  assign n26007 = \wishbone_bd_ram_mem0_reg[185][4]/P0001  & n13372 ;
  assign n26008 = \wishbone_bd_ram_mem0_reg[197][4]/P0001  & n13594 ;
  assign n26009 = ~n26007 & ~n26008 ;
  assign n26010 = \wishbone_bd_ram_mem0_reg[169][4]/P0001  & n13541 ;
  assign n26011 = \wishbone_bd_ram_mem0_reg[73][4]/P0001  & n13456 ;
  assign n26012 = ~n26010 & ~n26011 ;
  assign n26013 = n26009 & n26012 ;
  assign n26014 = \wishbone_bd_ram_mem0_reg[57][4]/P0001  & n13731 ;
  assign n26015 = \wishbone_bd_ram_mem0_reg[79][4]/P0001  & n13779 ;
  assign n26016 = ~n26014 & ~n26015 ;
  assign n26017 = \wishbone_bd_ram_mem0_reg[163][4]/P0001  & n13255 ;
  assign n26018 = \wishbone_bd_ram_mem0_reg[211][4]/P0001  & n13805 ;
  assign n26019 = ~n26017 & ~n26018 ;
  assign n26020 = n26016 & n26019 ;
  assign n26021 = n26013 & n26020 ;
  assign n26022 = \wishbone_bd_ram_mem0_reg[190][4]/P0001  & n13365 ;
  assign n26023 = \wishbone_bd_ram_mem0_reg[18][4]/P0001  & n13532 ;
  assign n26024 = ~n26022 & ~n26023 ;
  assign n26025 = \wishbone_bd_ram_mem0_reg[217][4]/P0001  & n13767 ;
  assign n26026 = \wishbone_bd_ram_mem0_reg[205][4]/P0001  & n13947 ;
  assign n26027 = ~n26025 & ~n26026 ;
  assign n26028 = n26024 & n26027 ;
  assign n26029 = \wishbone_bd_ram_mem0_reg[15][4]/P0001  & n13797 ;
  assign n26030 = \wishbone_bd_ram_mem0_reg[78][4]/P0001  & n13277 ;
  assign n26031 = ~n26029 & ~n26030 ;
  assign n26032 = \wishbone_bd_ram_mem0_reg[204][4]/P0001  & n13821 ;
  assign n26033 = \wishbone_bd_ram_mem0_reg[24][4]/P0001  & n13970 ;
  assign n26034 = ~n26032 & ~n26033 ;
  assign n26035 = n26031 & n26034 ;
  assign n26036 = n26028 & n26035 ;
  assign n26037 = n26021 & n26036 ;
  assign n26038 = n26006 & n26037 ;
  assign n26039 = n25975 & n26038 ;
  assign n26040 = \wishbone_bd_ram_mem0_reg[80][4]/P0001  & n13516 ;
  assign n26041 = \wishbone_bd_ram_mem0_reg[53][4]/P0001  & n13875 ;
  assign n26042 = ~n26040 & ~n26041 ;
  assign n26043 = \wishbone_bd_ram_mem0_reg[59][4]/P0001  & n13613 ;
  assign n26044 = \wishbone_bd_ram_mem0_reg[150][4]/P0001  & n13666 ;
  assign n26045 = ~n26043 & ~n26044 ;
  assign n26046 = n26042 & n26045 ;
  assign n26047 = \wishbone_bd_ram_mem0_reg[230][4]/P0001  & n13994 ;
  assign n26048 = \wishbone_bd_ram_mem0_reg[45][4]/P0001  & n13420 ;
  assign n26049 = ~n26047 & ~n26048 ;
  assign n26050 = \wishbone_bd_ram_mem0_reg[160][4]/P0001  & n13271 ;
  assign n26051 = \wishbone_bd_ram_mem0_reg[41][4]/P0001  & n14017 ;
  assign n26052 = ~n26050 & ~n26051 ;
  assign n26053 = n26049 & n26052 ;
  assign n26054 = n26046 & n26053 ;
  assign n26055 = \wishbone_bd_ram_mem0_reg[117][4]/P0001  & n13557 ;
  assign n26056 = \wishbone_bd_ram_mem0_reg[70][4]/P0001  & n13339 ;
  assign n26057 = ~n26055 & ~n26056 ;
  assign n26058 = \wishbone_bd_ram_mem0_reg[115][4]/P0001  & n13747 ;
  assign n26059 = \wishbone_bd_ram_mem0_reg[183][4]/P0001  & n13645 ;
  assign n26060 = ~n26058 & ~n26059 ;
  assign n26061 = n26057 & n26060 ;
  assign n26062 = \wishbone_bd_ram_mem0_reg[109][4]/P0001  & n13306 ;
  assign n26063 = \wishbone_bd_ram_mem0_reg[170][4]/P0001  & n14007 ;
  assign n26064 = ~n26062 & ~n26063 ;
  assign n26065 = \wishbone_bd_ram_mem0_reg[32][4]/P0001  & n13736 ;
  assign n26066 = \wishbone_bd_ram_mem0_reg[128][4]/P0001  & n13652 ;
  assign n26067 = ~n26065 & ~n26066 ;
  assign n26068 = n26064 & n26067 ;
  assign n26069 = n26061 & n26068 ;
  assign n26070 = n26054 & n26069 ;
  assign n26071 = \wishbone_bd_ram_mem0_reg[47][4]/P0001  & n13436 ;
  assign n26072 = \wishbone_bd_ram_mem0_reg[181][4]/P0001  & n13587 ;
  assign n26073 = ~n26071 & ~n26072 ;
  assign n26074 = \wishbone_bd_ram_mem0_reg[20][4]/P0001  & n13839 ;
  assign n26075 = \wishbone_bd_ram_mem0_reg[155][4]/P0001  & n13738 ;
  assign n26076 = ~n26074 & ~n26075 ;
  assign n26077 = n26073 & n26076 ;
  assign n26078 = \wishbone_bd_ram_mem0_reg[148][4]/P0001  & n13868 ;
  assign n26079 = \wishbone_bd_ram_mem0_reg[167][4]/P0001  & n13940 ;
  assign n26080 = ~n26078 & ~n26079 ;
  assign n26081 = \wishbone_bd_ram_mem0_reg[216][4]/P0001  & n14005 ;
  assign n26082 = \wishbone_bd_ram_mem0_reg[11][4]/P0001  & n13774 ;
  assign n26083 = ~n26081 & ~n26082 ;
  assign n26084 = n26080 & n26083 ;
  assign n26085 = n26077 & n26084 ;
  assign n26086 = \wishbone_bd_ram_mem0_reg[68][4]/P0001  & n13379 ;
  assign n26087 = \wishbone_bd_ram_mem0_reg[198][4]/P0001  & n13592 ;
  assign n26088 = ~n26086 & ~n26087 ;
  assign n26089 = \wishbone_bd_ram_mem0_reg[176][4]/P0001  & n13262 ;
  assign n26090 = \wishbone_bd_ram_mem0_reg[26][4]/P0001  & n13521 ;
  assign n26091 = ~n26089 & ~n26090 ;
  assign n26092 = n26088 & n26091 ;
  assign n26093 = \wishbone_bd_ram_mem0_reg[40][4]/P0001  & n13661 ;
  assign n26094 = \wishbone_bd_ram_mem0_reg[149][4]/P0001  & n13469 ;
  assign n26095 = ~n26093 & ~n26094 ;
  assign n26096 = \wishbone_bd_ram_mem0_reg[250][4]/P0001  & n13677 ;
  assign n26097 = \wishbone_bd_ram_mem0_reg[138][4]/P0001  & n13398 ;
  assign n26098 = ~n26096 & ~n26097 ;
  assign n26099 = n26095 & n26098 ;
  assign n26100 = n26092 & n26099 ;
  assign n26101 = n26085 & n26100 ;
  assign n26102 = n26070 & n26101 ;
  assign n26103 = \wishbone_bd_ram_mem0_reg[223][4]/P0001  & n13335 ;
  assign n26104 = \wishbone_bd_ram_mem0_reg[27][4]/P0001  & n13251 ;
  assign n26105 = ~n26103 & ~n26104 ;
  assign n26106 = \wishbone_bd_ram_mem0_reg[247][4]/P0001  & n13571 ;
  assign n26107 = \wishbone_bd_ram_mem0_reg[152][4]/P0001  & n13912 ;
  assign n26108 = ~n26106 & ~n26107 ;
  assign n26109 = n26105 & n26108 ;
  assign n26110 = \wishbone_bd_ram_mem0_reg[90][4]/P0001  & n13906 ;
  assign n26111 = \wishbone_bd_ram_mem0_reg[210][4]/P0001  & n13443 ;
  assign n26112 = ~n26110 & ~n26111 ;
  assign n26113 = \wishbone_bd_ram_mem0_reg[71][4]/P0001  & n13636 ;
  assign n26114 = \wishbone_bd_ram_mem0_reg[191][4]/P0001  & n14012 ;
  assign n26115 = ~n26113 & ~n26114 ;
  assign n26116 = n26112 & n26115 ;
  assign n26117 = n26109 & n26116 ;
  assign n26118 = \wishbone_bd_ram_mem0_reg[121][4]/P0001  & n13983 ;
  assign n26119 = \wishbone_bd_ram_mem0_reg[214][4]/P0001  & n13938 ;
  assign n26120 = ~n26118 & ~n26119 ;
  assign n26121 = \wishbone_bd_ram_mem0_reg[67][4]/P0001  & n13663 ;
  assign n26122 = \wishbone_bd_ram_mem0_reg[124][4]/P0001  & n14024 ;
  assign n26123 = ~n26121 & ~n26122 ;
  assign n26124 = n26120 & n26123 ;
  assign n26125 = \wishbone_bd_ram_mem0_reg[239][4]/P0001  & n13349 ;
  assign n26126 = \wishbone_bd_ram_mem0_reg[174][4]/P0001  & n13899 ;
  assign n26127 = ~n26125 & ~n26126 ;
  assign n26128 = \wishbone_bd_ram_mem0_reg[245][4]/P0001  & n13877 ;
  assign n26129 = \wishbone_bd_ram_mem0_reg[16][4]/P0001  & n13695 ;
  assign n26130 = ~n26128 & ~n26129 ;
  assign n26131 = n26127 & n26130 ;
  assign n26132 = n26124 & n26131 ;
  assign n26133 = n26117 & n26132 ;
  assign n26134 = \wishbone_bd_ram_mem0_reg[151][4]/P0001  & n13697 ;
  assign n26135 = \wishbone_bd_ram_mem0_reg[131][4]/P0001  & n13358 ;
  assign n26136 = ~n26134 & ~n26135 ;
  assign n26137 = \wishbone_bd_ram_mem0_reg[144][4]/P0001  & n13508 ;
  assign n26138 = \wishbone_bd_ram_mem0_reg[102][4]/P0001  & n13534 ;
  assign n26139 = ~n26137 & ~n26138 ;
  assign n26140 = n26136 & n26139 ;
  assign n26141 = \wishbone_bd_ram_mem0_reg[238][4]/P0001  & n13819 ;
  assign n26142 = \wishbone_bd_ram_mem0_reg[200][4]/P0001  & n13922 ;
  assign n26143 = ~n26141 & ~n26142 ;
  assign n26144 = \wishbone_bd_ram_mem0_reg[122][4]/P0001  & n13679 ;
  assign n26145 = \wishbone_bd_ram_mem0_reg[235][4]/P0001  & n13518 ;
  assign n26146 = ~n26144 & ~n26145 ;
  assign n26147 = n26143 & n26146 ;
  assign n26148 = n26140 & n26147 ;
  assign n26149 = \wishbone_bd_ram_mem0_reg[46][4]/P0001  & n13298 ;
  assign n26150 = \wishbone_bd_ram_mem0_reg[44][4]/P0001  & n13291 ;
  assign n26151 = ~n26149 & ~n26150 ;
  assign n26152 = \wishbone_bd_ram_mem0_reg[195][4]/P0001  & n13700 ;
  assign n26153 = \wishbone_bd_ram_mem0_reg[112][4]/P0001  & n13482 ;
  assign n26154 = ~n26152 & ~n26153 ;
  assign n26155 = n26151 & n26154 ;
  assign n26156 = \wishbone_bd_ram_mem0_reg[99][4]/P0001  & n13996 ;
  assign n26157 = \wishbone_bd_ram_mem0_reg[158][4]/P0001  & n13294 ;
  assign n26158 = ~n26156 & ~n26157 ;
  assign n26159 = \wishbone_bd_ram_mem0_reg[8][4]/P0001  & n13459 ;
  assign n26160 = \wishbone_bd_ram_mem0_reg[85][4]/P0001  & n13784 ;
  assign n26161 = ~n26159 & ~n26160 ;
  assign n26162 = n26158 & n26161 ;
  assign n26163 = n26155 & n26162 ;
  assign n26164 = n26148 & n26163 ;
  assign n26165 = n26133 & n26164 ;
  assign n26166 = n26102 & n26165 ;
  assign n26167 = n26039 & n26166 ;
  assign n26168 = n25912 & n26167 ;
  assign n26169 = ~wb_rst_i_pad & ~n25656 ;
  assign n26170 = ~n26168 & n26169 ;
  assign n26171 = ~n25657 & ~n26170 ;
  assign n26172 = \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  & n25059 ;
  assign n26173 = \ethreg1_irq_txc_reg/NET0131  & n25064 ;
  assign n26174 = \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  & n25084 ;
  assign n26175 = ~n26173 & ~n26174 ;
  assign n26176 = \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  & n23737 ;
  assign n26177 = \ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131  & n23782 ;
  assign n26178 = ~n26176 & ~n26177 ;
  assign n26179 = n26175 & n26178 ;
  assign n26180 = ~n26172 & n26179 ;
  assign n26181 = \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131  & n23813 ;
  assign n26182 = \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  & n23751 ;
  assign n26183 = n23747 & n26182 ;
  assign n26184 = ~n26181 & ~n26183 ;
  assign n26185 = \ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131  & n23743 ;
  assign n26186 = n23747 & n26185 ;
  assign n26187 = \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131  & n25069 ;
  assign n26188 = ~n26186 & ~n26187 ;
  assign n26189 = n26184 & n26188 ;
  assign n26190 = n23730 & n26189 ;
  assign n26191 = \ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131  & n23743 ;
  assign n26192 = n23741 & n26191 ;
  assign n26193 = \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131  & n25079 ;
  assign n26194 = ~n26192 & ~n26193 ;
  assign n26195 = \ethreg1_IPGT_0_DataOut_reg[5]/NET0131  & n25090 ;
  assign n26196 = \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131  & n25088 ;
  assign n26197 = ~n26195 & ~n26196 ;
  assign n26198 = n26194 & n26197 ;
  assign n26199 = \ethreg1_MODER_0_DataOut_reg[5]/NET0131  & n23808 ;
  assign n26200 = \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  & n23751 ;
  assign n26201 = n23741 & n26200 ;
  assign n26202 = ~n26199 & ~n26201 ;
  assign n26203 = \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131  & n23794 ;
  assign n26204 = n23741 & n26203 ;
  assign n26205 = \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131  & n25082 ;
  assign n26206 = ~n26204 & ~n26205 ;
  assign n26207 = n26202 & n26206 ;
  assign n26208 = n26198 & n26207 ;
  assign n26209 = n26190 & n26208 ;
  assign n26210 = n26180 & n26209 ;
  assign n26211 = n23730 & ~n26210 ;
  assign n26212 = \wishbone_bd_ram_mem0_reg[80][5]/P0001  & n13516 ;
  assign n26213 = \wishbone_bd_ram_mem0_reg[37][5]/P0001  & n13710 ;
  assign n26214 = ~n26212 & ~n26213 ;
  assign n26215 = \wishbone_bd_ram_mem0_reg[18][5]/P0001  & n13532 ;
  assign n26216 = \wishbone_bd_ram_mem0_reg[73][5]/P0001  & n13456 ;
  assign n26217 = ~n26215 & ~n26216 ;
  assign n26218 = n26214 & n26217 ;
  assign n26219 = \wishbone_bd_ram_mem0_reg[241][5]/P0001  & n13854 ;
  assign n26220 = \wishbone_bd_ram_mem0_reg[193][5]/P0001  & n14022 ;
  assign n26221 = ~n26219 & ~n26220 ;
  assign n26222 = \wishbone_bd_ram_mem0_reg[141][5]/P0001  & n13852 ;
  assign n26223 = \wishbone_bd_ram_mem0_reg[203][5]/P0001  & n13816 ;
  assign n26224 = ~n26222 & ~n26223 ;
  assign n26225 = n26221 & n26224 ;
  assign n26226 = n26218 & n26225 ;
  assign n26227 = \wishbone_bd_ram_mem0_reg[187][5]/P0001  & n13756 ;
  assign n26228 = \wishbone_bd_ram_mem0_reg[170][5]/P0001  & n14007 ;
  assign n26229 = ~n26227 & ~n26228 ;
  assign n26230 = \wishbone_bd_ram_mem0_reg[29][5]/P0001  & n13412 ;
  assign n26231 = \wishbone_bd_ram_mem0_reg[210][5]/P0001  & n13443 ;
  assign n26232 = ~n26230 & ~n26231 ;
  assign n26233 = n26229 & n26232 ;
  assign n26234 = \wishbone_bd_ram_mem0_reg[159][5]/P0001  & n13627 ;
  assign n26235 = \wishbone_bd_ram_mem0_reg[248][5]/P0001  & n13647 ;
  assign n26236 = ~n26234 & ~n26235 ;
  assign n26237 = \wishbone_bd_ram_mem0_reg[48][5]/P0001  & n13917 ;
  assign n26238 = \wishbone_bd_ram_mem0_reg[121][5]/P0001  & n13983 ;
  assign n26239 = ~n26237 & ~n26238 ;
  assign n26240 = n26236 & n26239 ;
  assign n26241 = n26233 & n26240 ;
  assign n26242 = n26226 & n26241 ;
  assign n26243 = \wishbone_bd_ram_mem0_reg[23][5]/P0001  & n13857 ;
  assign n26244 = \wishbone_bd_ram_mem0_reg[145][5]/P0001  & n13715 ;
  assign n26245 = ~n26243 & ~n26244 ;
  assign n26246 = \wishbone_bd_ram_mem0_reg[44][5]/P0001  & n13291 ;
  assign n26247 = \wishbone_bd_ram_mem0_reg[136][5]/P0001  & n13963 ;
  assign n26248 = ~n26246 & ~n26247 ;
  assign n26249 = n26245 & n26248 ;
  assign n26250 = \wishbone_bd_ram_mem0_reg[201][5]/P0001  & n13600 ;
  assign n26251 = \wishbone_bd_ram_mem0_reg[183][5]/P0001  & n13645 ;
  assign n26252 = ~n26250 & ~n26251 ;
  assign n26253 = \wishbone_bd_ram_mem0_reg[76][5]/P0001  & n13831 ;
  assign n26254 = \wishbone_bd_ram_mem0_reg[43][5]/P0001  & n13761 ;
  assign n26255 = ~n26253 & ~n26254 ;
  assign n26256 = n26252 & n26255 ;
  assign n26257 = n26249 & n26256 ;
  assign n26258 = \wishbone_bd_ram_mem0_reg[236][5]/P0001  & n13480 ;
  assign n26259 = \wishbone_bd_ram_mem0_reg[207][5]/P0001  & n13826 ;
  assign n26260 = ~n26258 & ~n26259 ;
  assign n26261 = \wishbone_bd_ram_mem0_reg[227][5]/P0001  & n13388 ;
  assign n26262 = \wishbone_bd_ram_mem0_reg[138][5]/P0001  & n13398 ;
  assign n26263 = ~n26261 & ~n26262 ;
  assign n26264 = n26260 & n26263 ;
  assign n26265 = \wishbone_bd_ram_mem0_reg[13][5]/P0001  & n13844 ;
  assign n26266 = \wishbone_bd_ram_mem0_reg[74][5]/P0001  & n13564 ;
  assign n26267 = ~n26265 & ~n26266 ;
  assign n26268 = \wishbone_bd_ram_mem0_reg[125][5]/P0001  & n13396 ;
  assign n26269 = \wishbone_bd_ram_mem0_reg[216][5]/P0001  & n14005 ;
  assign n26270 = ~n26268 & ~n26269 ;
  assign n26271 = n26267 & n26270 ;
  assign n26272 = n26264 & n26271 ;
  assign n26273 = n26257 & n26272 ;
  assign n26274 = n26242 & n26273 ;
  assign n26275 = \wishbone_bd_ram_mem0_reg[243][5]/P0001  & n13575 ;
  assign n26276 = \wishbone_bd_ram_mem0_reg[99][5]/P0001  & n13996 ;
  assign n26277 = ~n26275 & ~n26276 ;
  assign n26278 = \wishbone_bd_ram_mem0_reg[93][5]/P0001  & n13891 ;
  assign n26279 = \wishbone_bd_ram_mem0_reg[65][5]/P0001  & n13842 ;
  assign n26280 = ~n26278 & ~n26279 ;
  assign n26281 = n26277 & n26280 ;
  assign n26282 = \wishbone_bd_ram_mem0_reg[220][5]/P0001  & n13965 ;
  assign n26283 = \wishbone_bd_ram_mem0_reg[245][5]/P0001  & n13877 ;
  assign n26284 = ~n26282 & ~n26283 ;
  assign n26285 = \wishbone_bd_ram_mem0_reg[214][5]/P0001  & n13938 ;
  assign n26286 = \wishbone_bd_ram_mem0_reg[108][5]/P0001  & n13814 ;
  assign n26287 = ~n26285 & ~n26286 ;
  assign n26288 = n26284 & n26287 ;
  assign n26289 = n26281 & n26288 ;
  assign n26290 = \wishbone_bd_ram_mem0_reg[153][5]/P0001  & n13309 ;
  assign n26291 = \wishbone_bd_ram_mem0_reg[70][5]/P0001  & n13339 ;
  assign n26292 = ~n26290 & ~n26291 ;
  assign n26293 = \wishbone_bd_ram_mem0_reg[167][5]/P0001  & n13940 ;
  assign n26294 = \wishbone_bd_ram_mem0_reg[132][5]/P0001  & n13927 ;
  assign n26295 = ~n26293 & ~n26294 ;
  assign n26296 = n26292 & n26295 ;
  assign n26297 = \wishbone_bd_ram_mem0_reg[111][5]/P0001  & n13471 ;
  assign n26298 = \wishbone_bd_ram_mem0_reg[229][5]/P0001  & n13552 ;
  assign n26299 = ~n26297 & ~n26298 ;
  assign n26300 = \wishbone_bd_ram_mem0_reg[164][5]/P0001  & n13236 ;
  assign n26301 = \wishbone_bd_ram_mem0_reg[225][5]/P0001  & n13719 ;
  assign n26302 = ~n26300 & ~n26301 ;
  assign n26303 = n26299 & n26302 ;
  assign n26304 = n26296 & n26303 ;
  assign n26305 = n26289 & n26304 ;
  assign n26306 = \wishbone_bd_ram_mem0_reg[208][5]/P0001  & n14010 ;
  assign n26307 = \wishbone_bd_ram_mem0_reg[102][5]/P0001  & n13534 ;
  assign n26308 = ~n26306 & ~n26307 ;
  assign n26309 = \wishbone_bd_ram_mem0_reg[174][5]/P0001  & n13899 ;
  assign n26310 = \wishbone_bd_ram_mem0_reg[231][5]/P0001  & n13363 ;
  assign n26311 = ~n26309 & ~n26310 ;
  assign n26312 = n26308 & n26311 ;
  assign n26313 = \wishbone_bd_ram_mem0_reg[206][5]/P0001  & n13414 ;
  assign n26314 = \wishbone_bd_ram_mem0_reg[204][5]/P0001  & n13821 ;
  assign n26315 = ~n26313 & ~n26314 ;
  assign n26316 = \wishbone_bd_ram_mem0_reg[20][5]/P0001  & n13839 ;
  assign n26317 = \wishbone_bd_ram_mem0_reg[4][5]/P0001  & n13527 ;
  assign n26318 = ~n26316 & ~n26317 ;
  assign n26319 = n26315 & n26318 ;
  assign n26320 = n26312 & n26319 ;
  assign n26321 = \wishbone_bd_ram_mem0_reg[186][5]/P0001  & n13616 ;
  assign n26322 = \wishbone_bd_ram_mem0_reg[26][5]/P0001  & n13521 ;
  assign n26323 = ~n26321 & ~n26322 ;
  assign n26324 = \wishbone_bd_ram_mem0_reg[134][5]/P0001  & n13494 ;
  assign n26325 = \wishbone_bd_ram_mem0_reg[38][5]/P0001  & n13828 ;
  assign n26326 = ~n26324 & ~n26325 ;
  assign n26327 = n26323 & n26326 ;
  assign n26328 = \wishbone_bd_ram_mem0_reg[171][5]/P0001  & n13422 ;
  assign n26329 = \wishbone_bd_ram_mem0_reg[35][5]/P0001  & n13523 ;
  assign n26330 = ~n26328 & ~n26329 ;
  assign n26331 = \wishbone_bd_ram_mem0_reg[3][5]/P0001  & n13354 ;
  assign n26332 = \wishbone_bd_ram_mem0_reg[88][5]/P0001  & n13347 ;
  assign n26333 = ~n26331 & ~n26332 ;
  assign n26334 = n26330 & n26333 ;
  assign n26335 = n26327 & n26334 ;
  assign n26336 = n26320 & n26335 ;
  assign n26337 = n26305 & n26336 ;
  assign n26338 = n26274 & n26337 ;
  assign n26339 = \wishbone_bd_ram_mem0_reg[57][5]/P0001  & n13731 ;
  assign n26340 = \wishbone_bd_ram_mem0_reg[198][5]/P0001  & n13592 ;
  assign n26341 = ~n26339 & ~n26340 ;
  assign n26342 = \wishbone_bd_ram_mem0_reg[242][5]/P0001  & n13383 ;
  assign n26343 = \wishbone_bd_ram_mem0_reg[180][5]/P0001  & n13650 ;
  assign n26344 = ~n26342 & ~n26343 ;
  assign n26345 = n26341 & n26344 ;
  assign n26346 = \wishbone_bd_ram_mem0_reg[127][5]/P0001  & n13803 ;
  assign n26347 = \wishbone_bd_ram_mem0_reg[232][5]/P0001  & n13510 ;
  assign n26348 = ~n26346 & ~n26347 ;
  assign n26349 = \wishbone_bd_ram_mem0_reg[56][5]/P0001  & n13611 ;
  assign n26350 = \wishbone_bd_ram_mem0_reg[1][5]/P0001  & n13888 ;
  assign n26351 = ~n26349 & ~n26350 ;
  assign n26352 = n26348 & n26351 ;
  assign n26353 = n26345 & n26352 ;
  assign n26354 = \wishbone_bd_ram_mem0_reg[237][5]/P0001  & n13924 ;
  assign n26355 = \wishbone_bd_ram_mem0_reg[100][5]/P0001  & n13401 ;
  assign n26356 = ~n26354 & ~n26355 ;
  assign n26357 = \wishbone_bd_ram_mem0_reg[154][5]/P0001  & n13403 ;
  assign n26358 = \wishbone_bd_ram_mem0_reg[173][5]/P0001  & n13360 ;
  assign n26359 = ~n26357 & ~n26358 ;
  assign n26360 = n26356 & n26359 ;
  assign n26361 = \wishbone_bd_ram_mem0_reg[91][5]/P0001  & n13954 ;
  assign n26362 = \wishbone_bd_ram_mem0_reg[49][5]/P0001  & n13929 ;
  assign n26363 = ~n26361 & ~n26362 ;
  assign n26364 = \wishbone_bd_ram_mem0_reg[98][5]/P0001  & n13569 ;
  assign n26365 = \wishbone_bd_ram_mem0_reg[105][5]/P0001  & n13503 ;
  assign n26366 = ~n26364 & ~n26365 ;
  assign n26367 = n26363 & n26366 ;
  assign n26368 = n26360 & n26367 ;
  assign n26369 = n26353 & n26368 ;
  assign n26370 = \wishbone_bd_ram_mem0_reg[61][5]/P0001  & n13544 ;
  assign n26371 = \wishbone_bd_ram_mem0_reg[200][5]/P0001  & n13922 ;
  assign n26372 = ~n26370 & ~n26371 ;
  assign n26373 = \wishbone_bd_ram_mem0_reg[149][5]/P0001  & n13469 ;
  assign n26374 = \wishbone_bd_ram_mem0_reg[32][5]/P0001  & n13736 ;
  assign n26375 = ~n26373 & ~n26374 ;
  assign n26376 = n26372 & n26375 ;
  assign n26377 = \wishbone_bd_ram_mem0_reg[30][5]/P0001  & n13713 ;
  assign n26378 = \wishbone_bd_ram_mem0_reg[60][5]/P0001  & n13790 ;
  assign n26379 = ~n26377 & ~n26378 ;
  assign n26380 = \wishbone_bd_ram_mem0_reg[33][5]/P0001  & n13933 ;
  assign n26381 = \wishbone_bd_ram_mem0_reg[95][5]/P0001  & n13317 ;
  assign n26382 = ~n26380 & ~n26381 ;
  assign n26383 = n26379 & n26382 ;
  assign n26384 = n26376 & n26383 ;
  assign n26385 = \wishbone_bd_ram_mem0_reg[50][5]/P0001  & n13686 ;
  assign n26386 = \wishbone_bd_ram_mem0_reg[94][5]/P0001  & n13833 ;
  assign n26387 = ~n26385 & ~n26386 ;
  assign n26388 = \wishbone_bd_ram_mem0_reg[39][5]/P0001  & n13893 ;
  assign n26389 = \wishbone_bd_ram_mem0_reg[51][5]/P0001  & n13880 ;
  assign n26390 = ~n26388 & ~n26389 ;
  assign n26391 = n26387 & n26390 ;
  assign n26392 = \wishbone_bd_ram_mem0_reg[166][5]/P0001  & n13999 ;
  assign n26393 = \wishbone_bd_ram_mem0_reg[246][5]/P0001  & n13981 ;
  assign n26394 = ~n26392 & ~n26393 ;
  assign n26395 = \wishbone_bd_ram_mem0_reg[175][5]/P0001  & n13674 ;
  assign n26396 = \wishbone_bd_ram_mem0_reg[150][5]/P0001  & n13666 ;
  assign n26397 = ~n26395 & ~n26396 ;
  assign n26398 = n26394 & n26397 ;
  assign n26399 = n26391 & n26398 ;
  assign n26400 = n26384 & n26399 ;
  assign n26401 = n26369 & n26400 ;
  assign n26402 = \wishbone_bd_ram_mem0_reg[14][5]/P0001  & n13972 ;
  assign n26403 = \wishbone_bd_ram_mem0_reg[169][5]/P0001  & n13541 ;
  assign n26404 = ~n26402 & ~n26403 ;
  assign n26405 = \wishbone_bd_ram_mem0_reg[143][5]/P0001  & n13461 ;
  assign n26406 = \wishbone_bd_ram_mem0_reg[185][5]/P0001  & n13372 ;
  assign n26407 = ~n26405 & ~n26406 ;
  assign n26408 = n26404 & n26407 ;
  assign n26409 = \wishbone_bd_ram_mem0_reg[106][5]/P0001  & n13555 ;
  assign n26410 = \wishbone_bd_ram_mem0_reg[215][5]/P0001  & n13901 ;
  assign n26411 = ~n26409 & ~n26410 ;
  assign n26412 = \wishbone_bd_ram_mem0_reg[12][5]/P0001  & n13733 ;
  assign n26413 = \wishbone_bd_ram_mem0_reg[118][5]/P0001  & n13589 ;
  assign n26414 = ~n26412 & ~n26413 ;
  assign n26415 = n26411 & n26414 ;
  assign n26416 = n26408 & n26415 ;
  assign n26417 = \wishbone_bd_ram_mem0_reg[15][5]/P0001  & n13797 ;
  assign n26418 = \wishbone_bd_ram_mem0_reg[131][5]/P0001  & n13358 ;
  assign n26419 = ~n26417 & ~n26418 ;
  assign n26420 = \wishbone_bd_ram_mem0_reg[172][5]/P0001  & n13377 ;
  assign n26421 = \wishbone_bd_ram_mem0_reg[209][5]/P0001  & n13689 ;
  assign n26422 = ~n26420 & ~n26421 ;
  assign n26423 = n26419 & n26422 ;
  assign n26424 = \wishbone_bd_ram_mem0_reg[120][5]/P0001  & n13550 ;
  assign n26425 = \wishbone_bd_ram_mem0_reg[239][5]/P0001  & n13349 ;
  assign n26426 = ~n26424 & ~n26425 ;
  assign n26427 = \wishbone_bd_ram_mem0_reg[116][5]/P0001  & n13865 ;
  assign n26428 = \wishbone_bd_ram_mem0_reg[122][5]/P0001  & n13679 ;
  assign n26429 = ~n26427 & ~n26428 ;
  assign n26430 = n26426 & n26429 ;
  assign n26431 = n26423 & n26430 ;
  assign n26432 = n26416 & n26431 ;
  assign n26433 = \wishbone_bd_ram_mem0_reg[64][5]/P0001  & n13904 ;
  assign n26434 = \wishbone_bd_ram_mem0_reg[71][5]/P0001  & n13636 ;
  assign n26435 = ~n26433 & ~n26434 ;
  assign n26436 = \wishbone_bd_ram_mem0_reg[195][5]/P0001  & n13700 ;
  assign n26437 = \wishbone_bd_ram_mem0_reg[41][5]/P0001  & n14017 ;
  assign n26438 = ~n26436 & ~n26437 ;
  assign n26439 = n26435 & n26438 ;
  assign n26440 = \wishbone_bd_ram_mem0_reg[123][5]/P0001  & n13749 ;
  assign n26441 = \wishbone_bd_ram_mem0_reg[181][5]/P0001  & n13587 ;
  assign n26442 = ~n26440 & ~n26441 ;
  assign n26443 = \wishbone_bd_ram_mem0_reg[28][5]/P0001  & n13810 ;
  assign n26444 = \wishbone_bd_ram_mem0_reg[218][5]/P0001  & n13792 ;
  assign n26445 = ~n26443 & ~n26444 ;
  assign n26446 = n26442 & n26445 ;
  assign n26447 = n26439 & n26446 ;
  assign n26448 = \wishbone_bd_ram_mem0_reg[247][5]/P0001  & n13571 ;
  assign n26449 = \wishbone_bd_ram_mem0_reg[197][5]/P0001  & n13594 ;
  assign n26450 = ~n26448 & ~n26449 ;
  assign n26451 = \wishbone_bd_ram_mem0_reg[55][5]/P0001  & n13618 ;
  assign n26452 = \wishbone_bd_ram_mem0_reg[194][5]/P0001  & n13624 ;
  assign n26453 = ~n26451 & ~n26452 ;
  assign n26454 = n26450 & n26453 ;
  assign n26455 = \wishbone_bd_ram_mem0_reg[211][5]/P0001  & n13805 ;
  assign n26456 = \wishbone_bd_ram_mem0_reg[189][5]/P0001  & n14001 ;
  assign n26457 = ~n26455 & ~n26456 ;
  assign n26458 = \wishbone_bd_ram_mem0_reg[146][5]/P0001  & n13958 ;
  assign n26459 = \wishbone_bd_ram_mem0_reg[157][5]/P0001  & n13445 ;
  assign n26460 = ~n26458 & ~n26459 ;
  assign n26461 = n26457 & n26460 ;
  assign n26462 = n26454 & n26461 ;
  assign n26463 = n26447 & n26462 ;
  assign n26464 = n26432 & n26463 ;
  assign n26465 = n26401 & n26464 ;
  assign n26466 = n26338 & n26465 ;
  assign n26467 = \wishbone_bd_ram_mem0_reg[52][5]/P0001  & n13988 ;
  assign n26468 = \wishbone_bd_ram_mem0_reg[8][5]/P0001  & n13459 ;
  assign n26469 = ~n26467 & ~n26468 ;
  assign n26470 = \wishbone_bd_ram_mem0_reg[101][5]/P0001  & n13772 ;
  assign n26471 = \wishbone_bd_ram_mem0_reg[217][5]/P0001  & n13767 ;
  assign n26472 = ~n26470 & ~n26471 ;
  assign n26473 = n26469 & n26472 ;
  assign n26474 = \wishbone_bd_ram_mem0_reg[84][5]/P0001  & n13385 ;
  assign n26475 = \wishbone_bd_ram_mem0_reg[17][5]/P0001  & n13324 ;
  assign n26476 = ~n26474 & ~n26475 ;
  assign n26477 = \wishbone_bd_ram_mem0_reg[252][5]/P0001  & n13986 ;
  assign n26478 = \wishbone_bd_ram_mem0_reg[155][5]/P0001  & n13738 ;
  assign n26479 = ~n26477 & ~n26478 ;
  assign n26480 = n26476 & n26479 ;
  assign n26481 = n26473 & n26480 ;
  assign n26482 = \wishbone_bd_ram_mem0_reg[89][5]/P0001  & n13910 ;
  assign n26483 = \wishbone_bd_ram_mem0_reg[2][5]/P0001  & n13975 ;
  assign n26484 = ~n26482 & ~n26483 ;
  assign n26485 = \wishbone_bd_ram_mem0_reg[212][5]/P0001  & n13634 ;
  assign n26486 = \wishbone_bd_ram_mem0_reg[86][5]/P0001  & n13485 ;
  assign n26487 = ~n26485 & ~n26486 ;
  assign n26488 = n26484 & n26487 ;
  assign n26489 = \wishbone_bd_ram_mem0_reg[77][5]/P0001  & n13935 ;
  assign n26490 = \wishbone_bd_ram_mem0_reg[182][5]/P0001  & n13598 ;
  assign n26491 = ~n26489 & ~n26490 ;
  assign n26492 = \wishbone_bd_ram_mem0_reg[158][5]/P0001  & n13294 ;
  assign n26493 = \wishbone_bd_ram_mem0_reg[7][5]/P0001  & n13546 ;
  assign n26494 = ~n26492 & ~n26493 ;
  assign n26495 = n26491 & n26494 ;
  assign n26496 = n26488 & n26495 ;
  assign n26497 = n26481 & n26496 ;
  assign n26498 = \wishbone_bd_ram_mem0_reg[219][5]/P0001  & n13577 ;
  assign n26499 = \wishbone_bd_ram_mem0_reg[0][5]/P0001  & n13539 ;
  assign n26500 = ~n26498 & ~n26499 ;
  assign n26501 = \wishbone_bd_ram_mem0_reg[79][5]/P0001  & n13779 ;
  assign n26502 = \wishbone_bd_ram_mem0_reg[156][5]/P0001  & n13769 ;
  assign n26503 = ~n26501 & ~n26502 ;
  assign n26504 = n26500 & n26503 ;
  assign n26505 = \wishbone_bd_ram_mem0_reg[250][5]/P0001  & n13677 ;
  assign n26506 = \wishbone_bd_ram_mem0_reg[184][5]/P0001  & n13960 ;
  assign n26507 = ~n26505 & ~n26506 ;
  assign n26508 = \wishbone_bd_ram_mem0_reg[16][5]/P0001  & n13695 ;
  assign n26509 = \wishbone_bd_ram_mem0_reg[176][5]/P0001  & n13262 ;
  assign n26510 = ~n26508 & ~n26509 ;
  assign n26511 = n26507 & n26510 ;
  assign n26512 = n26504 & n26511 ;
  assign n26513 = \wishbone_bd_ram_mem0_reg[47][5]/P0001  & n13436 ;
  assign n26514 = \wishbone_bd_ram_mem0_reg[40][5]/P0001  & n13661 ;
  assign n26515 = ~n26513 & ~n26514 ;
  assign n26516 = \wishbone_bd_ram_mem0_reg[115][5]/P0001  & n13747 ;
  assign n26517 = \wishbone_bd_ram_mem0_reg[22][5]/P0001  & n13744 ;
  assign n26518 = ~n26516 & ~n26517 ;
  assign n26519 = n26515 & n26518 ;
  assign n26520 = \wishbone_bd_ram_mem0_reg[66][5]/P0001  & n13603 ;
  assign n26521 = \wishbone_bd_ram_mem0_reg[163][5]/P0001  & n13255 ;
  assign n26522 = ~n26520 & ~n26521 ;
  assign n26523 = \wishbone_bd_ram_mem0_reg[83][5]/P0001  & n13454 ;
  assign n26524 = \wishbone_bd_ram_mem0_reg[152][5]/P0001  & n13912 ;
  assign n26525 = ~n26523 & ~n26524 ;
  assign n26526 = n26522 & n26525 ;
  assign n26527 = n26519 & n26526 ;
  assign n26528 = n26512 & n26527 ;
  assign n26529 = n26497 & n26528 ;
  assign n26530 = \wishbone_bd_ram_mem0_reg[253][5]/P0001  & n13708 ;
  assign n26531 = \wishbone_bd_ram_mem0_reg[109][5]/P0001  & n13306 ;
  assign n26532 = ~n26530 & ~n26531 ;
  assign n26533 = \wishbone_bd_ram_mem0_reg[72][5]/P0001  & n13582 ;
  assign n26534 = \wishbone_bd_ram_mem0_reg[199][5]/P0001  & n13499 ;
  assign n26535 = ~n26533 & ~n26534 ;
  assign n26536 = n26532 & n26535 ;
  assign n26537 = \wishbone_bd_ram_mem0_reg[213][5]/P0001  & n13870 ;
  assign n26538 = \wishbone_bd_ram_mem0_reg[130][5]/P0001  & n13427 ;
  assign n26539 = ~n26537 & ~n26538 ;
  assign n26540 = \wishbone_bd_ram_mem0_reg[54][5]/P0001  & n13622 ;
  assign n26541 = \wishbone_bd_ram_mem0_reg[36][5]/P0001  & n13639 ;
  assign n26542 = ~n26540 & ~n26541 ;
  assign n26543 = n26539 & n26542 ;
  assign n26544 = n26536 & n26543 ;
  assign n26545 = \wishbone_bd_ram_mem0_reg[234][5]/P0001  & n13781 ;
  assign n26546 = \wishbone_bd_ram_mem0_reg[124][5]/P0001  & n14024 ;
  assign n26547 = ~n26545 & ~n26546 ;
  assign n26548 = \wishbone_bd_ram_mem0_reg[34][5]/P0001  & n13450 ;
  assign n26549 = \wishbone_bd_ram_mem0_reg[196][5]/P0001  & n13977 ;
  assign n26550 = ~n26548 & ~n26549 ;
  assign n26551 = n26547 & n26550 ;
  assign n26552 = \wishbone_bd_ram_mem0_reg[160][5]/P0001  & n13271 ;
  assign n26553 = \wishbone_bd_ram_mem0_reg[117][5]/P0001  & n13557 ;
  assign n26554 = ~n26552 & ~n26553 ;
  assign n26555 = \wishbone_bd_ram_mem0_reg[137][5]/P0001  & n13808 ;
  assign n26556 = \wishbone_bd_ram_mem0_reg[147][5]/P0001  & n13702 ;
  assign n26557 = ~n26555 & ~n26556 ;
  assign n26558 = n26554 & n26557 ;
  assign n26559 = n26551 & n26558 ;
  assign n26560 = n26544 & n26559 ;
  assign n26561 = \wishbone_bd_ram_mem0_reg[126][5]/P0001  & n13786 ;
  assign n26562 = \wishbone_bd_ram_mem0_reg[191][5]/P0001  & n14012 ;
  assign n26563 = ~n26561 & ~n26562 ;
  assign n26564 = \wishbone_bd_ram_mem0_reg[45][5]/P0001  & n13420 ;
  assign n26565 = \wishbone_bd_ram_mem0_reg[19][5]/P0001  & n13886 ;
  assign n26566 = ~n26564 & ~n26565 ;
  assign n26567 = n26563 & n26566 ;
  assign n26568 = \wishbone_bd_ram_mem0_reg[230][5]/P0001  & n13994 ;
  assign n26569 = \wishbone_bd_ram_mem0_reg[205][5]/P0001  & n13947 ;
  assign n26570 = ~n26568 & ~n26569 ;
  assign n26571 = \wishbone_bd_ram_mem0_reg[240][5]/P0001  & n13352 ;
  assign n26572 = \wishbone_bd_ram_mem0_reg[255][5]/P0001  & n13952 ;
  assign n26573 = ~n26571 & ~n26572 ;
  assign n26574 = n26570 & n26573 ;
  assign n26575 = n26567 & n26574 ;
  assign n26576 = \wishbone_bd_ram_mem0_reg[233][5]/P0001  & n13332 ;
  assign n26577 = \wishbone_bd_ram_mem0_reg[161][5]/P0001  & n13505 ;
  assign n26578 = ~n26576 & ~n26577 ;
  assign n26579 = \wishbone_bd_ram_mem0_reg[6][5]/P0001  & n13915 ;
  assign n26580 = \wishbone_bd_ram_mem0_reg[188][5]/P0001  & n13407 ;
  assign n26581 = ~n26579 & ~n26580 ;
  assign n26582 = n26578 & n26581 ;
  assign n26583 = \wishbone_bd_ram_mem0_reg[119][5]/P0001  & n14033 ;
  assign n26584 = \wishbone_bd_ram_mem0_reg[148][5]/P0001  & n13868 ;
  assign n26585 = ~n26583 & ~n26584 ;
  assign n26586 = \wishbone_bd_ram_mem0_reg[21][5]/P0001  & n13438 ;
  assign n26587 = \wishbone_bd_ram_mem0_reg[68][5]/P0001  & n13379 ;
  assign n26588 = ~n26586 & ~n26587 ;
  assign n26589 = n26585 & n26588 ;
  assign n26590 = n26582 & n26589 ;
  assign n26591 = n26575 & n26590 ;
  assign n26592 = n26560 & n26591 ;
  assign n26593 = n26529 & n26592 ;
  assign n26594 = \wishbone_bd_ram_mem0_reg[62][5]/P0001  & n13529 ;
  assign n26595 = \wishbone_bd_ram_mem0_reg[112][5]/P0001  & n13482 ;
  assign n26596 = ~n26594 & ~n26595 ;
  assign n26597 = \wishbone_bd_ram_mem0_reg[92][5]/P0001  & n13859 ;
  assign n26598 = \wishbone_bd_ram_mem0_reg[168][5]/P0001  & n13795 ;
  assign n26599 = ~n26597 & ~n26598 ;
  assign n26600 = n26596 & n26599 ;
  assign n26601 = \wishbone_bd_ram_mem0_reg[107][5]/P0001  & n13476 ;
  assign n26602 = \wishbone_bd_ram_mem0_reg[165][5]/P0001  & n14028 ;
  assign n26603 = ~n26601 & ~n26602 ;
  assign n26604 = \wishbone_bd_ram_mem0_reg[128][5]/P0001  & n13652 ;
  assign n26605 = \wishbone_bd_ram_mem0_reg[254][5]/P0001  & n13283 ;
  assign n26606 = ~n26604 & ~n26605 ;
  assign n26607 = n26603 & n26606 ;
  assign n26608 = n26600 & n26607 ;
  assign n26609 = \wishbone_bd_ram_mem0_reg[81][5]/P0001  & n13409 ;
  assign n26610 = \wishbone_bd_ram_mem0_reg[178][5]/P0001  & n13301 ;
  assign n26611 = ~n26609 & ~n26610 ;
  assign n26612 = \wishbone_bd_ram_mem0_reg[11][5]/P0001  & n13774 ;
  assign n26613 = \wishbone_bd_ram_mem0_reg[5][5]/P0001  & n13243 ;
  assign n26614 = ~n26612 & ~n26613 ;
  assign n26615 = n26611 & n26614 ;
  assign n26616 = \wishbone_bd_ram_mem0_reg[46][5]/P0001  & n13298 ;
  assign n26617 = \wishbone_bd_ram_mem0_reg[24][5]/P0001  & n13970 ;
  assign n26618 = ~n26616 & ~n26617 ;
  assign n26619 = \wishbone_bd_ram_mem0_reg[59][5]/P0001  & n13613 ;
  assign n26620 = \wishbone_bd_ram_mem0_reg[135][5]/P0001  & n13672 ;
  assign n26621 = ~n26619 & ~n26620 ;
  assign n26622 = n26618 & n26621 ;
  assign n26623 = n26615 & n26622 ;
  assign n26624 = n26608 & n26623 ;
  assign n26625 = \wishbone_bd_ram_mem0_reg[192][5]/P0001  & n13390 ;
  assign n26626 = \wishbone_bd_ram_mem0_reg[25][5]/P0001  & n13742 ;
  assign n26627 = ~n26625 & ~n26626 ;
  assign n26628 = \wishbone_bd_ram_mem0_reg[226][5]/P0001  & n13668 ;
  assign n26629 = \wishbone_bd_ram_mem0_reg[144][5]/P0001  & n13508 ;
  assign n26630 = ~n26628 & ~n26629 ;
  assign n26631 = n26627 & n26630 ;
  assign n26632 = \wishbone_bd_ram_mem0_reg[151][5]/P0001  & n13697 ;
  assign n26633 = \wishbone_bd_ram_mem0_reg[129][5]/P0001  & n13629 ;
  assign n26634 = ~n26632 & ~n26633 ;
  assign n26635 = \wishbone_bd_ram_mem0_reg[31][5]/P0001  & n13758 ;
  assign n26636 = \wishbone_bd_ram_mem0_reg[75][5]/P0001  & n13605 ;
  assign n26637 = ~n26635 & ~n26636 ;
  assign n26638 = n26634 & n26637 ;
  assign n26639 = n26631 & n26638 ;
  assign n26640 = \wishbone_bd_ram_mem0_reg[114][5]/P0001  & n13763 ;
  assign n26641 = \wishbone_bd_ram_mem0_reg[228][5]/P0001  & n13497 ;
  assign n26642 = ~n26640 & ~n26641 ;
  assign n26643 = \wishbone_bd_ram_mem0_reg[110][5]/P0001  & n14030 ;
  assign n26644 = \wishbone_bd_ram_mem0_reg[78][5]/P0001  & n13277 ;
  assign n26645 = ~n26643 & ~n26644 ;
  assign n26646 = n26642 & n26645 ;
  assign n26647 = \wishbone_bd_ram_mem0_reg[224][5]/P0001  & n13433 ;
  assign n26648 = \wishbone_bd_ram_mem0_reg[85][5]/P0001  & n13784 ;
  assign n26649 = ~n26647 & ~n26648 ;
  assign n26650 = \wishbone_bd_ram_mem0_reg[67][5]/P0001  & n13663 ;
  assign n26651 = \wishbone_bd_ram_mem0_reg[142][5]/P0001  & n13448 ;
  assign n26652 = ~n26650 & ~n26651 ;
  assign n26653 = n26649 & n26652 ;
  assign n26654 = n26646 & n26653 ;
  assign n26655 = n26639 & n26654 ;
  assign n26656 = n26624 & n26655 ;
  assign n26657 = \wishbone_bd_ram_mem0_reg[140][5]/P0001  & n13287 ;
  assign n26658 = \wishbone_bd_ram_mem0_reg[69][5]/P0001  & n13487 ;
  assign n26659 = ~n26657 & ~n26658 ;
  assign n26660 = \wishbone_bd_ram_mem0_reg[244][5]/P0001  & n13474 ;
  assign n26661 = \wishbone_bd_ram_mem0_reg[202][5]/P0001  & n13268 ;
  assign n26662 = ~n26660 & ~n26661 ;
  assign n26663 = n26659 & n26662 ;
  assign n26664 = \wishbone_bd_ram_mem0_reg[177][5]/P0001  & n13863 ;
  assign n26665 = \wishbone_bd_ram_mem0_reg[133][5]/P0001  & n13492 ;
  assign n26666 = ~n26664 & ~n26665 ;
  assign n26667 = \wishbone_bd_ram_mem0_reg[87][5]/P0001  & n13691 ;
  assign n26668 = \wishbone_bd_ram_mem0_reg[179][5]/P0001  & n14035 ;
  assign n26669 = ~n26667 & ~n26668 ;
  assign n26670 = n26666 & n26669 ;
  assign n26671 = n26663 & n26670 ;
  assign n26672 = \wishbone_bd_ram_mem0_reg[42][5]/P0001  & n13341 ;
  assign n26673 = \wishbone_bd_ram_mem0_reg[10][5]/P0001  & n13837 ;
  assign n26674 = ~n26672 & ~n26673 ;
  assign n26675 = \wishbone_bd_ram_mem0_reg[27][5]/P0001  & n13251 ;
  assign n26676 = \wishbone_bd_ram_mem0_reg[162][5]/P0001  & n13726 ;
  assign n26677 = ~n26675 & ~n26676 ;
  assign n26678 = n26674 & n26677 ;
  assign n26679 = \wishbone_bd_ram_mem0_reg[190][5]/P0001  & n13365 ;
  assign n26680 = \wishbone_bd_ram_mem0_reg[103][5]/P0001  & n13320 ;
  assign n26681 = ~n26679 & ~n26680 ;
  assign n26682 = \wishbone_bd_ram_mem0_reg[221][5]/P0001  & n13641 ;
  assign n26683 = \wishbone_bd_ram_mem0_reg[9][5]/P0001  & n13580 ;
  assign n26684 = ~n26682 & ~n26683 ;
  assign n26685 = n26681 & n26684 ;
  assign n26686 = n26678 & n26685 ;
  assign n26687 = n26671 & n26686 ;
  assign n26688 = \wishbone_bd_ram_mem0_reg[104][5]/P0001  & n13684 ;
  assign n26689 = \wishbone_bd_ram_mem0_reg[63][5]/P0001  & n13327 ;
  assign n26690 = ~n26688 & ~n26689 ;
  assign n26691 = \wishbone_bd_ram_mem0_reg[90][5]/P0001  & n13906 ;
  assign n26692 = \wishbone_bd_ram_mem0_reg[96][5]/P0001  & n13425 ;
  assign n26693 = ~n26691 & ~n26692 ;
  assign n26694 = n26690 & n26693 ;
  assign n26695 = \wishbone_bd_ram_mem0_reg[251][5]/P0001  & n14019 ;
  assign n26696 = \wishbone_bd_ram_mem0_reg[235][5]/P0001  & n13518 ;
  assign n26697 = ~n26695 & ~n26696 ;
  assign n26698 = \wishbone_bd_ram_mem0_reg[53][5]/P0001  & n13875 ;
  assign n26699 = \wishbone_bd_ram_mem0_reg[223][5]/P0001  & n13335 ;
  assign n26700 = ~n26698 & ~n26699 ;
  assign n26701 = n26697 & n26700 ;
  assign n26702 = n26694 & n26701 ;
  assign n26703 = \wishbone_bd_ram_mem0_reg[249][5]/P0001  & n13431 ;
  assign n26704 = \wishbone_bd_ram_mem0_reg[238][5]/P0001  & n13819 ;
  assign n26705 = ~n26703 & ~n26704 ;
  assign n26706 = \wishbone_bd_ram_mem0_reg[139][5]/P0001  & n13566 ;
  assign n26707 = \wishbone_bd_ram_mem0_reg[97][5]/P0001  & n13724 ;
  assign n26708 = ~n26706 & ~n26707 ;
  assign n26709 = n26705 & n26708 ;
  assign n26710 = \wishbone_bd_ram_mem0_reg[82][5]/P0001  & n13374 ;
  assign n26711 = \wishbone_bd_ram_mem0_reg[222][5]/P0001  & n13721 ;
  assign n26712 = ~n26710 & ~n26711 ;
  assign n26713 = \wishbone_bd_ram_mem0_reg[58][5]/P0001  & n13949 ;
  assign n26714 = \wishbone_bd_ram_mem0_reg[113][5]/P0001  & n13882 ;
  assign n26715 = ~n26713 & ~n26714 ;
  assign n26716 = n26712 & n26715 ;
  assign n26717 = n26709 & n26716 ;
  assign n26718 = n26702 & n26717 ;
  assign n26719 = n26687 & n26718 ;
  assign n26720 = n26656 & n26719 ;
  assign n26721 = n26593 & n26720 ;
  assign n26722 = n26466 & n26721 ;
  assign n26723 = ~wb_rst_i_pad & ~n26210 ;
  assign n26724 = ~n26722 & n26723 ;
  assign n26725 = ~n26211 & ~n26724 ;
  assign n26726 = \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  & n23751 ;
  assign n26727 = n23741 & n26726 ;
  assign n26728 = \ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131  & n25088 ;
  assign n26729 = ~n26727 & ~n26728 ;
  assign n26730 = \ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131  & n23782 ;
  assign n26731 = \ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131  & n23743 ;
  assign n26732 = n23741 & n26731 ;
  assign n26733 = ~n26730 & ~n26732 ;
  assign n26734 = n26729 & n26733 ;
  assign n26735 = \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  & n25084 ;
  assign n26736 = \ethreg1_MODER_0_DataOut_reg[7]/NET0131  & n23808 ;
  assign n26737 = ~n26735 & ~n26736 ;
  assign n26738 = n23730 & n26737 ;
  assign n26739 = n26734 & n26738 ;
  assign n26740 = \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  & n23737 ;
  assign n26741 = \ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131  & n23743 ;
  assign n26742 = n23747 & n26741 ;
  assign n26743 = \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  & n23751 ;
  assign n26744 = n23747 & n26743 ;
  assign n26745 = ~n26742 & ~n26744 ;
  assign n26746 = \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131  & n23794 ;
  assign n26747 = n23741 & n26746 ;
  assign n26748 = \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131  & n23813 ;
  assign n26749 = ~n26747 & ~n26748 ;
  assign n26750 = n26745 & n26749 ;
  assign n26751 = ~n26740 & n26750 ;
  assign n26752 = n26739 & n26751 ;
  assign n26753 = n23730 & ~n26752 ;
  assign n26754 = \wishbone_bd_ram_mem0_reg[49][7]/P0001  & n13929 ;
  assign n26755 = \wishbone_bd_ram_mem0_reg[69][7]/P0001  & n13487 ;
  assign n26756 = ~n26754 & ~n26755 ;
  assign n26757 = \wishbone_bd_ram_mem0_reg[21][7]/P0001  & n13438 ;
  assign n26758 = \wishbone_bd_ram_mem0_reg[105][7]/P0001  & n13503 ;
  assign n26759 = ~n26757 & ~n26758 ;
  assign n26760 = n26756 & n26759 ;
  assign n26761 = \wishbone_bd_ram_mem0_reg[222][7]/P0001  & n13721 ;
  assign n26762 = \wishbone_bd_ram_mem0_reg[193][7]/P0001  & n14022 ;
  assign n26763 = ~n26761 & ~n26762 ;
  assign n26764 = \wishbone_bd_ram_mem0_reg[85][7]/P0001  & n13784 ;
  assign n26765 = \wishbone_bd_ram_mem0_reg[242][7]/P0001  & n13383 ;
  assign n26766 = ~n26764 & ~n26765 ;
  assign n26767 = n26763 & n26766 ;
  assign n26768 = n26760 & n26767 ;
  assign n26769 = \wishbone_bd_ram_mem0_reg[240][7]/P0001  & n13352 ;
  assign n26770 = \wishbone_bd_ram_mem0_reg[183][7]/P0001  & n13645 ;
  assign n26771 = ~n26769 & ~n26770 ;
  assign n26772 = \wishbone_bd_ram_mem0_reg[118][7]/P0001  & n13589 ;
  assign n26773 = \wishbone_bd_ram_mem0_reg[213][7]/P0001  & n13870 ;
  assign n26774 = ~n26772 & ~n26773 ;
  assign n26775 = n26771 & n26774 ;
  assign n26776 = \wishbone_bd_ram_mem0_reg[116][7]/P0001  & n13865 ;
  assign n26777 = \wishbone_bd_ram_mem0_reg[248][7]/P0001  & n13647 ;
  assign n26778 = ~n26776 & ~n26777 ;
  assign n26779 = \wishbone_bd_ram_mem0_reg[28][7]/P0001  & n13810 ;
  assign n26780 = \wishbone_bd_ram_mem0_reg[144][7]/P0001  & n13508 ;
  assign n26781 = ~n26779 & ~n26780 ;
  assign n26782 = n26778 & n26781 ;
  assign n26783 = n26775 & n26782 ;
  assign n26784 = n26768 & n26783 ;
  assign n26785 = \wishbone_bd_ram_mem0_reg[156][7]/P0001  & n13769 ;
  assign n26786 = \wishbone_bd_ram_mem0_reg[153][7]/P0001  & n13309 ;
  assign n26787 = ~n26785 & ~n26786 ;
  assign n26788 = \wishbone_bd_ram_mem0_reg[44][7]/P0001  & n13291 ;
  assign n26789 = \wishbone_bd_ram_mem0_reg[59][7]/P0001  & n13613 ;
  assign n26790 = ~n26788 & ~n26789 ;
  assign n26791 = n26787 & n26790 ;
  assign n26792 = \wishbone_bd_ram_mem0_reg[176][7]/P0001  & n13262 ;
  assign n26793 = \wishbone_bd_ram_mem0_reg[235][7]/P0001  & n13518 ;
  assign n26794 = ~n26792 & ~n26793 ;
  assign n26795 = \wishbone_bd_ram_mem0_reg[163][7]/P0001  & n13255 ;
  assign n26796 = \wishbone_bd_ram_mem0_reg[9][7]/P0001  & n13580 ;
  assign n26797 = ~n26795 & ~n26796 ;
  assign n26798 = n26794 & n26797 ;
  assign n26799 = n26791 & n26798 ;
  assign n26800 = \wishbone_bd_ram_mem0_reg[166][7]/P0001  & n13999 ;
  assign n26801 = \wishbone_bd_ram_mem0_reg[251][7]/P0001  & n14019 ;
  assign n26802 = ~n26800 & ~n26801 ;
  assign n26803 = \wishbone_bd_ram_mem0_reg[178][7]/P0001  & n13301 ;
  assign n26804 = \wishbone_bd_ram_mem0_reg[37][7]/P0001  & n13710 ;
  assign n26805 = ~n26803 & ~n26804 ;
  assign n26806 = n26802 & n26805 ;
  assign n26807 = \wishbone_bd_ram_mem0_reg[17][7]/P0001  & n13324 ;
  assign n26808 = \wishbone_bd_ram_mem0_reg[170][7]/P0001  & n14007 ;
  assign n26809 = ~n26807 & ~n26808 ;
  assign n26810 = \wishbone_bd_ram_mem0_reg[192][7]/P0001  & n13390 ;
  assign n26811 = \wishbone_bd_ram_mem0_reg[207][7]/P0001  & n13826 ;
  assign n26812 = ~n26810 & ~n26811 ;
  assign n26813 = n26809 & n26812 ;
  assign n26814 = n26806 & n26813 ;
  assign n26815 = n26799 & n26814 ;
  assign n26816 = n26784 & n26815 ;
  assign n26817 = \wishbone_bd_ram_mem0_reg[244][7]/P0001  & n13474 ;
  assign n26818 = \wishbone_bd_ram_mem0_reg[101][7]/P0001  & n13772 ;
  assign n26819 = ~n26817 & ~n26818 ;
  assign n26820 = \wishbone_bd_ram_mem0_reg[169][7]/P0001  & n13541 ;
  assign n26821 = \wishbone_bd_ram_mem0_reg[104][7]/P0001  & n13684 ;
  assign n26822 = ~n26820 & ~n26821 ;
  assign n26823 = n26819 & n26822 ;
  assign n26824 = \wishbone_bd_ram_mem0_reg[161][7]/P0001  & n13505 ;
  assign n26825 = \wishbone_bd_ram_mem0_reg[173][7]/P0001  & n13360 ;
  assign n26826 = ~n26824 & ~n26825 ;
  assign n26827 = \wishbone_bd_ram_mem0_reg[233][7]/P0001  & n13332 ;
  assign n26828 = \wishbone_bd_ram_mem0_reg[98][7]/P0001  & n13569 ;
  assign n26829 = ~n26827 & ~n26828 ;
  assign n26830 = n26826 & n26829 ;
  assign n26831 = n26823 & n26830 ;
  assign n26832 = \wishbone_bd_ram_mem0_reg[243][7]/P0001  & n13575 ;
  assign n26833 = \wishbone_bd_ram_mem0_reg[19][7]/P0001  & n13886 ;
  assign n26834 = ~n26832 & ~n26833 ;
  assign n26835 = \wishbone_bd_ram_mem0_reg[190][7]/P0001  & n13365 ;
  assign n26836 = \wishbone_bd_ram_mem0_reg[188][7]/P0001  & n13407 ;
  assign n26837 = ~n26835 & ~n26836 ;
  assign n26838 = n26834 & n26837 ;
  assign n26839 = \wishbone_bd_ram_mem0_reg[112][7]/P0001  & n13482 ;
  assign n26840 = \wishbone_bd_ram_mem0_reg[252][7]/P0001  & n13986 ;
  assign n26841 = ~n26839 & ~n26840 ;
  assign n26842 = \wishbone_bd_ram_mem0_reg[60][7]/P0001  & n13790 ;
  assign n26843 = \wishbone_bd_ram_mem0_reg[181][7]/P0001  & n13587 ;
  assign n26844 = ~n26842 & ~n26843 ;
  assign n26845 = n26841 & n26844 ;
  assign n26846 = n26838 & n26845 ;
  assign n26847 = n26831 & n26846 ;
  assign n26848 = \wishbone_bd_ram_mem0_reg[218][7]/P0001  & n13792 ;
  assign n26849 = \wishbone_bd_ram_mem0_reg[130][7]/P0001  & n13427 ;
  assign n26850 = ~n26848 & ~n26849 ;
  assign n26851 = \wishbone_bd_ram_mem0_reg[79][7]/P0001  & n13779 ;
  assign n26852 = \wishbone_bd_ram_mem0_reg[189][7]/P0001  & n14001 ;
  assign n26853 = ~n26851 & ~n26852 ;
  assign n26854 = n26850 & n26853 ;
  assign n26855 = \wishbone_bd_ram_mem0_reg[91][7]/P0001  & n13954 ;
  assign n26856 = \wishbone_bd_ram_mem0_reg[72][7]/P0001  & n13582 ;
  assign n26857 = ~n26855 & ~n26856 ;
  assign n26858 = \wishbone_bd_ram_mem0_reg[149][7]/P0001  & n13469 ;
  assign n26859 = \wishbone_bd_ram_mem0_reg[24][7]/P0001  & n13970 ;
  assign n26860 = ~n26858 & ~n26859 ;
  assign n26861 = n26857 & n26860 ;
  assign n26862 = n26854 & n26861 ;
  assign n26863 = \wishbone_bd_ram_mem0_reg[22][7]/P0001  & n13744 ;
  assign n26864 = \wishbone_bd_ram_mem0_reg[34][7]/P0001  & n13450 ;
  assign n26865 = ~n26863 & ~n26864 ;
  assign n26866 = \wishbone_bd_ram_mem0_reg[136][7]/P0001  & n13963 ;
  assign n26867 = \wishbone_bd_ram_mem0_reg[39][7]/P0001  & n13893 ;
  assign n26868 = ~n26866 & ~n26867 ;
  assign n26869 = n26865 & n26868 ;
  assign n26870 = \wishbone_bd_ram_mem0_reg[172][7]/P0001  & n13377 ;
  assign n26871 = \wishbone_bd_ram_mem0_reg[55][7]/P0001  & n13618 ;
  assign n26872 = ~n26870 & ~n26871 ;
  assign n26873 = \wishbone_bd_ram_mem0_reg[95][7]/P0001  & n13317 ;
  assign n26874 = \wishbone_bd_ram_mem0_reg[180][7]/P0001  & n13650 ;
  assign n26875 = ~n26873 & ~n26874 ;
  assign n26876 = n26872 & n26875 ;
  assign n26877 = n26869 & n26876 ;
  assign n26878 = n26862 & n26877 ;
  assign n26879 = n26847 & n26878 ;
  assign n26880 = n26816 & n26879 ;
  assign n26881 = \wishbone_bd_ram_mem0_reg[61][7]/P0001  & n13544 ;
  assign n26882 = \wishbone_bd_ram_mem0_reg[124][7]/P0001  & n14024 ;
  assign n26883 = ~n26881 & ~n26882 ;
  assign n26884 = \wishbone_bd_ram_mem0_reg[247][7]/P0001  & n13571 ;
  assign n26885 = \wishbone_bd_ram_mem0_reg[212][7]/P0001  & n13634 ;
  assign n26886 = ~n26884 & ~n26885 ;
  assign n26887 = n26883 & n26886 ;
  assign n26888 = \wishbone_bd_ram_mem0_reg[255][7]/P0001  & n13952 ;
  assign n26889 = \wishbone_bd_ram_mem0_reg[237][7]/P0001  & n13924 ;
  assign n26890 = ~n26888 & ~n26889 ;
  assign n26891 = \wishbone_bd_ram_mem0_reg[128][7]/P0001  & n13652 ;
  assign n26892 = \wishbone_bd_ram_mem0_reg[5][7]/P0001  & n13243 ;
  assign n26893 = ~n26891 & ~n26892 ;
  assign n26894 = n26890 & n26893 ;
  assign n26895 = n26887 & n26894 ;
  assign n26896 = \wishbone_bd_ram_mem0_reg[196][7]/P0001  & n13977 ;
  assign n26897 = \wishbone_bd_ram_mem0_reg[82][7]/P0001  & n13374 ;
  assign n26898 = ~n26896 & ~n26897 ;
  assign n26899 = \wishbone_bd_ram_mem0_reg[253][7]/P0001  & n13708 ;
  assign n26900 = \wishbone_bd_ram_mem0_reg[211][7]/P0001  & n13805 ;
  assign n26901 = ~n26899 & ~n26900 ;
  assign n26902 = n26898 & n26901 ;
  assign n26903 = \wishbone_bd_ram_mem0_reg[70][7]/P0001  & n13339 ;
  assign n26904 = \wishbone_bd_ram_mem0_reg[141][7]/P0001  & n13852 ;
  assign n26905 = ~n26903 & ~n26904 ;
  assign n26906 = \wishbone_bd_ram_mem0_reg[108][7]/P0001  & n13814 ;
  assign n26907 = \wishbone_bd_ram_mem0_reg[186][7]/P0001  & n13616 ;
  assign n26908 = ~n26906 & ~n26907 ;
  assign n26909 = n26905 & n26908 ;
  assign n26910 = n26902 & n26909 ;
  assign n26911 = n26895 & n26910 ;
  assign n26912 = \wishbone_bd_ram_mem0_reg[57][7]/P0001  & n13731 ;
  assign n26913 = \wishbone_bd_ram_mem0_reg[179][7]/P0001  & n14035 ;
  assign n26914 = ~n26912 & ~n26913 ;
  assign n26915 = \wishbone_bd_ram_mem0_reg[42][7]/P0001  & n13341 ;
  assign n26916 = \wishbone_bd_ram_mem0_reg[31][7]/P0001  & n13758 ;
  assign n26917 = ~n26915 & ~n26916 ;
  assign n26918 = n26914 & n26917 ;
  assign n26919 = \wishbone_bd_ram_mem0_reg[8][7]/P0001  & n13459 ;
  assign n26920 = \wishbone_bd_ram_mem0_reg[80][7]/P0001  & n13516 ;
  assign n26921 = ~n26919 & ~n26920 ;
  assign n26922 = \wishbone_bd_ram_mem0_reg[230][7]/P0001  & n13994 ;
  assign n26923 = \wishbone_bd_ram_mem0_reg[64][7]/P0001  & n13904 ;
  assign n26924 = ~n26922 & ~n26923 ;
  assign n26925 = n26921 & n26924 ;
  assign n26926 = n26918 & n26925 ;
  assign n26927 = \wishbone_bd_ram_mem0_reg[16][7]/P0001  & n13695 ;
  assign n26928 = \wishbone_bd_ram_mem0_reg[219][7]/P0001  & n13577 ;
  assign n26929 = ~n26927 & ~n26928 ;
  assign n26930 = \wishbone_bd_ram_mem0_reg[38][7]/P0001  & n13828 ;
  assign n26931 = \wishbone_bd_ram_mem0_reg[23][7]/P0001  & n13857 ;
  assign n26932 = ~n26930 & ~n26931 ;
  assign n26933 = n26929 & n26932 ;
  assign n26934 = \wishbone_bd_ram_mem0_reg[107][7]/P0001  & n13476 ;
  assign n26935 = \wishbone_bd_ram_mem0_reg[246][7]/P0001  & n13981 ;
  assign n26936 = ~n26934 & ~n26935 ;
  assign n26937 = \wishbone_bd_ram_mem0_reg[77][7]/P0001  & n13935 ;
  assign n26938 = \wishbone_bd_ram_mem0_reg[109][7]/P0001  & n13306 ;
  assign n26939 = ~n26937 & ~n26938 ;
  assign n26940 = n26936 & n26939 ;
  assign n26941 = n26933 & n26940 ;
  assign n26942 = n26926 & n26941 ;
  assign n26943 = n26911 & n26942 ;
  assign n26944 = \wishbone_bd_ram_mem0_reg[7][7]/P0001  & n13546 ;
  assign n26945 = \wishbone_bd_ram_mem0_reg[158][7]/P0001  & n13294 ;
  assign n26946 = ~n26944 & ~n26945 ;
  assign n26947 = \wishbone_bd_ram_mem0_reg[102][7]/P0001  & n13534 ;
  assign n26948 = \wishbone_bd_ram_mem0_reg[114][7]/P0001  & n13763 ;
  assign n26949 = ~n26947 & ~n26948 ;
  assign n26950 = n26946 & n26949 ;
  assign n26951 = \wishbone_bd_ram_mem0_reg[191][7]/P0001  & n14012 ;
  assign n26952 = \wishbone_bd_ram_mem0_reg[92][7]/P0001  & n13859 ;
  assign n26953 = ~n26951 & ~n26952 ;
  assign n26954 = \wishbone_bd_ram_mem0_reg[30][7]/P0001  & n13713 ;
  assign n26955 = \wishbone_bd_ram_mem0_reg[26][7]/P0001  & n13521 ;
  assign n26956 = ~n26954 & ~n26955 ;
  assign n26957 = n26953 & n26956 ;
  assign n26958 = n26950 & n26957 ;
  assign n26959 = \wishbone_bd_ram_mem0_reg[221][7]/P0001  & n13641 ;
  assign n26960 = \wishbone_bd_ram_mem0_reg[131][7]/P0001  & n13358 ;
  assign n26961 = ~n26959 & ~n26960 ;
  assign n26962 = \wishbone_bd_ram_mem0_reg[210][7]/P0001  & n13443 ;
  assign n26963 = \wishbone_bd_ram_mem0_reg[223][7]/P0001  & n13335 ;
  assign n26964 = ~n26962 & ~n26963 ;
  assign n26965 = n26961 & n26964 ;
  assign n26966 = \wishbone_bd_ram_mem0_reg[151][7]/P0001  & n13697 ;
  assign n26967 = \wishbone_bd_ram_mem0_reg[227][7]/P0001  & n13388 ;
  assign n26968 = ~n26966 & ~n26967 ;
  assign n26969 = \wishbone_bd_ram_mem0_reg[122][7]/P0001  & n13679 ;
  assign n26970 = \wishbone_bd_ram_mem0_reg[117][7]/P0001  & n13557 ;
  assign n26971 = ~n26969 & ~n26970 ;
  assign n26972 = n26968 & n26971 ;
  assign n26973 = n26965 & n26972 ;
  assign n26974 = n26958 & n26973 ;
  assign n26975 = \wishbone_bd_ram_mem0_reg[3][7]/P0001  & n13354 ;
  assign n26976 = \wishbone_bd_ram_mem0_reg[10][7]/P0001  & n13837 ;
  assign n26977 = ~n26975 & ~n26976 ;
  assign n26978 = \wishbone_bd_ram_mem0_reg[198][7]/P0001  & n13592 ;
  assign n26979 = \wishbone_bd_ram_mem0_reg[232][7]/P0001  & n13510 ;
  assign n26980 = ~n26978 & ~n26979 ;
  assign n26981 = n26977 & n26980 ;
  assign n26982 = \wishbone_bd_ram_mem0_reg[150][7]/P0001  & n13666 ;
  assign n26983 = \wishbone_bd_ram_mem0_reg[245][7]/P0001  & n13877 ;
  assign n26984 = ~n26982 & ~n26983 ;
  assign n26985 = \wishbone_bd_ram_mem0_reg[74][7]/P0001  & n13564 ;
  assign n26986 = \wishbone_bd_ram_mem0_reg[138][7]/P0001  & n13398 ;
  assign n26987 = ~n26985 & ~n26986 ;
  assign n26988 = n26984 & n26987 ;
  assign n26989 = n26981 & n26988 ;
  assign n26990 = \wishbone_bd_ram_mem0_reg[224][7]/P0001  & n13433 ;
  assign n26991 = \wishbone_bd_ram_mem0_reg[152][7]/P0001  & n13912 ;
  assign n26992 = ~n26990 & ~n26991 ;
  assign n26993 = \wishbone_bd_ram_mem0_reg[35][7]/P0001  & n13523 ;
  assign n26994 = \wishbone_bd_ram_mem0_reg[238][7]/P0001  & n13819 ;
  assign n26995 = ~n26993 & ~n26994 ;
  assign n26996 = n26992 & n26995 ;
  assign n26997 = \wishbone_bd_ram_mem0_reg[120][7]/P0001  & n13550 ;
  assign n26998 = \wishbone_bd_ram_mem0_reg[206][7]/P0001  & n13414 ;
  assign n26999 = ~n26997 & ~n26998 ;
  assign n27000 = \wishbone_bd_ram_mem0_reg[13][7]/P0001  & n13844 ;
  assign n27001 = \wishbone_bd_ram_mem0_reg[119][7]/P0001  & n14033 ;
  assign n27002 = ~n27000 & ~n27001 ;
  assign n27003 = n26999 & n27002 ;
  assign n27004 = n26996 & n27003 ;
  assign n27005 = n26989 & n27004 ;
  assign n27006 = n26974 & n27005 ;
  assign n27007 = n26943 & n27006 ;
  assign n27008 = n26880 & n27007 ;
  assign n27009 = \wishbone_bd_ram_mem0_reg[29][7]/P0001  & n13412 ;
  assign n27010 = \wishbone_bd_ram_mem0_reg[0][7]/P0001  & n13539 ;
  assign n27011 = ~n27009 & ~n27010 ;
  assign n27012 = \wishbone_bd_ram_mem0_reg[99][7]/P0001  & n13996 ;
  assign n27013 = \wishbone_bd_ram_mem0_reg[239][7]/P0001  & n13349 ;
  assign n27014 = ~n27012 & ~n27013 ;
  assign n27015 = n27011 & n27014 ;
  assign n27016 = \wishbone_bd_ram_mem0_reg[160][7]/P0001  & n13271 ;
  assign n27017 = \wishbone_bd_ram_mem0_reg[2][7]/P0001  & n13975 ;
  assign n27018 = ~n27016 & ~n27017 ;
  assign n27019 = \wishbone_bd_ram_mem0_reg[254][7]/P0001  & n13283 ;
  assign n27020 = \wishbone_bd_ram_mem0_reg[155][7]/P0001  & n13738 ;
  assign n27021 = ~n27019 & ~n27020 ;
  assign n27022 = n27018 & n27021 ;
  assign n27023 = n27015 & n27022 ;
  assign n27024 = \wishbone_bd_ram_mem0_reg[217][7]/P0001  & n13767 ;
  assign n27025 = \wishbone_bd_ram_mem0_reg[1][7]/P0001  & n13888 ;
  assign n27026 = ~n27024 & ~n27025 ;
  assign n27027 = \wishbone_bd_ram_mem0_reg[84][7]/P0001  & n13385 ;
  assign n27028 = \wishbone_bd_ram_mem0_reg[214][7]/P0001  & n13938 ;
  assign n27029 = ~n27027 & ~n27028 ;
  assign n27030 = n27026 & n27029 ;
  assign n27031 = \wishbone_bd_ram_mem0_reg[62][7]/P0001  & n13529 ;
  assign n27032 = \wishbone_bd_ram_mem0_reg[182][7]/P0001  & n13598 ;
  assign n27033 = ~n27031 & ~n27032 ;
  assign n27034 = \wishbone_bd_ram_mem0_reg[94][7]/P0001  & n13833 ;
  assign n27035 = \wishbone_bd_ram_mem0_reg[41][7]/P0001  & n14017 ;
  assign n27036 = ~n27034 & ~n27035 ;
  assign n27037 = n27033 & n27036 ;
  assign n27038 = n27030 & n27037 ;
  assign n27039 = n27023 & n27038 ;
  assign n27040 = \wishbone_bd_ram_mem0_reg[201][7]/P0001  & n13600 ;
  assign n27041 = \wishbone_bd_ram_mem0_reg[33][7]/P0001  & n13933 ;
  assign n27042 = ~n27040 & ~n27041 ;
  assign n27043 = \wishbone_bd_ram_mem0_reg[52][7]/P0001  & n13988 ;
  assign n27044 = \wishbone_bd_ram_mem0_reg[78][7]/P0001  & n13277 ;
  assign n27045 = ~n27043 & ~n27044 ;
  assign n27046 = n27042 & n27045 ;
  assign n27047 = \wishbone_bd_ram_mem0_reg[226][7]/P0001  & n13668 ;
  assign n27048 = \wishbone_bd_ram_mem0_reg[215][7]/P0001  & n13901 ;
  assign n27049 = ~n27047 & ~n27048 ;
  assign n27050 = \wishbone_bd_ram_mem0_reg[184][7]/P0001  & n13960 ;
  assign n27051 = \wishbone_bd_ram_mem0_reg[83][7]/P0001  & n13454 ;
  assign n27052 = ~n27050 & ~n27051 ;
  assign n27053 = n27049 & n27052 ;
  assign n27054 = n27046 & n27053 ;
  assign n27055 = \wishbone_bd_ram_mem0_reg[171][7]/P0001  & n13422 ;
  assign n27056 = \wishbone_bd_ram_mem0_reg[65][7]/P0001  & n13842 ;
  assign n27057 = ~n27055 & ~n27056 ;
  assign n27058 = \wishbone_bd_ram_mem0_reg[14][7]/P0001  & n13972 ;
  assign n27059 = \wishbone_bd_ram_mem0_reg[25][7]/P0001  & n13742 ;
  assign n27060 = ~n27058 & ~n27059 ;
  assign n27061 = n27057 & n27060 ;
  assign n27062 = \wishbone_bd_ram_mem0_reg[66][7]/P0001  & n13603 ;
  assign n27063 = \wishbone_bd_ram_mem0_reg[46][7]/P0001  & n13298 ;
  assign n27064 = ~n27062 & ~n27063 ;
  assign n27065 = \wishbone_bd_ram_mem0_reg[159][7]/P0001  & n13627 ;
  assign n27066 = \wishbone_bd_ram_mem0_reg[89][7]/P0001  & n13910 ;
  assign n27067 = ~n27065 & ~n27066 ;
  assign n27068 = n27064 & n27067 ;
  assign n27069 = n27061 & n27068 ;
  assign n27070 = n27054 & n27069 ;
  assign n27071 = n27039 & n27070 ;
  assign n27072 = \wishbone_bd_ram_mem0_reg[250][7]/P0001  & n13677 ;
  assign n27073 = \wishbone_bd_ram_mem0_reg[51][7]/P0001  & n13880 ;
  assign n27074 = ~n27072 & ~n27073 ;
  assign n27075 = \wishbone_bd_ram_mem0_reg[209][7]/P0001  & n13689 ;
  assign n27076 = \wishbone_bd_ram_mem0_reg[127][7]/P0001  & n13803 ;
  assign n27077 = ~n27075 & ~n27076 ;
  assign n27078 = n27074 & n27077 ;
  assign n27079 = \wishbone_bd_ram_mem0_reg[87][7]/P0001  & n13691 ;
  assign n27080 = \wishbone_bd_ram_mem0_reg[103][7]/P0001  & n13320 ;
  assign n27081 = ~n27079 & ~n27080 ;
  assign n27082 = \wishbone_bd_ram_mem0_reg[234][7]/P0001  & n13781 ;
  assign n27083 = \wishbone_bd_ram_mem0_reg[81][7]/P0001  & n13409 ;
  assign n27084 = ~n27082 & ~n27083 ;
  assign n27085 = n27081 & n27084 ;
  assign n27086 = n27078 & n27085 ;
  assign n27087 = \wishbone_bd_ram_mem0_reg[88][7]/P0001  & n13347 ;
  assign n27088 = \wishbone_bd_ram_mem0_reg[133][7]/P0001  & n13492 ;
  assign n27089 = ~n27087 & ~n27088 ;
  assign n27090 = \wishbone_bd_ram_mem0_reg[20][7]/P0001  & n13839 ;
  assign n27091 = \wishbone_bd_ram_mem0_reg[204][7]/P0001  & n13821 ;
  assign n27092 = ~n27090 & ~n27091 ;
  assign n27093 = n27089 & n27092 ;
  assign n27094 = \wishbone_bd_ram_mem0_reg[140][7]/P0001  & n13287 ;
  assign n27095 = \wishbone_bd_ram_mem0_reg[137][7]/P0001  & n13808 ;
  assign n27096 = ~n27094 & ~n27095 ;
  assign n27097 = \wishbone_bd_ram_mem0_reg[123][7]/P0001  & n13749 ;
  assign n27098 = \wishbone_bd_ram_mem0_reg[76][7]/P0001  & n13831 ;
  assign n27099 = ~n27097 & ~n27098 ;
  assign n27100 = n27096 & n27099 ;
  assign n27101 = n27093 & n27100 ;
  assign n27102 = n27086 & n27101 ;
  assign n27103 = \wishbone_bd_ram_mem0_reg[126][7]/P0001  & n13786 ;
  assign n27104 = \wishbone_bd_ram_mem0_reg[174][7]/P0001  & n13899 ;
  assign n27105 = ~n27103 & ~n27104 ;
  assign n27106 = \wishbone_bd_ram_mem0_reg[63][7]/P0001  & n13327 ;
  assign n27107 = \wishbone_bd_ram_mem0_reg[115][7]/P0001  & n13747 ;
  assign n27108 = ~n27106 & ~n27107 ;
  assign n27109 = n27105 & n27108 ;
  assign n27110 = \wishbone_bd_ram_mem0_reg[231][7]/P0001  & n13363 ;
  assign n27111 = \wishbone_bd_ram_mem0_reg[205][7]/P0001  & n13947 ;
  assign n27112 = ~n27110 & ~n27111 ;
  assign n27113 = \wishbone_bd_ram_mem0_reg[187][7]/P0001  & n13756 ;
  assign n27114 = \wishbone_bd_ram_mem0_reg[113][7]/P0001  & n13882 ;
  assign n27115 = ~n27113 & ~n27114 ;
  assign n27116 = n27112 & n27115 ;
  assign n27117 = n27109 & n27116 ;
  assign n27118 = \wishbone_bd_ram_mem0_reg[139][7]/P0001  & n13566 ;
  assign n27119 = \wishbone_bd_ram_mem0_reg[157][7]/P0001  & n13445 ;
  assign n27120 = ~n27118 & ~n27119 ;
  assign n27121 = \wishbone_bd_ram_mem0_reg[15][7]/P0001  & n13797 ;
  assign n27122 = \wishbone_bd_ram_mem0_reg[132][7]/P0001  & n13927 ;
  assign n27123 = ~n27121 & ~n27122 ;
  assign n27124 = n27120 & n27123 ;
  assign n27125 = \wishbone_bd_ram_mem0_reg[147][7]/P0001  & n13702 ;
  assign n27126 = \wishbone_bd_ram_mem0_reg[75][7]/P0001  & n13605 ;
  assign n27127 = ~n27125 & ~n27126 ;
  assign n27128 = \wishbone_bd_ram_mem0_reg[18][7]/P0001  & n13532 ;
  assign n27129 = \wishbone_bd_ram_mem0_reg[40][7]/P0001  & n13661 ;
  assign n27130 = ~n27128 & ~n27129 ;
  assign n27131 = n27127 & n27130 ;
  assign n27132 = n27124 & n27131 ;
  assign n27133 = n27117 & n27132 ;
  assign n27134 = n27102 & n27133 ;
  assign n27135 = n27071 & n27134 ;
  assign n27136 = \wishbone_bd_ram_mem0_reg[135][7]/P0001  & n13672 ;
  assign n27137 = \wishbone_bd_ram_mem0_reg[111][7]/P0001  & n13471 ;
  assign n27138 = ~n27136 & ~n27137 ;
  assign n27139 = \wishbone_bd_ram_mem0_reg[134][7]/P0001  & n13494 ;
  assign n27140 = \wishbone_bd_ram_mem0_reg[165][7]/P0001  & n14028 ;
  assign n27141 = ~n27139 & ~n27140 ;
  assign n27142 = n27138 & n27141 ;
  assign n27143 = \wishbone_bd_ram_mem0_reg[90][7]/P0001  & n13906 ;
  assign n27144 = \wishbone_bd_ram_mem0_reg[100][7]/P0001  & n13401 ;
  assign n27145 = ~n27143 & ~n27144 ;
  assign n27146 = \wishbone_bd_ram_mem0_reg[47][7]/P0001  & n13436 ;
  assign n27147 = \wishbone_bd_ram_mem0_reg[249][7]/P0001  & n13431 ;
  assign n27148 = ~n27146 & ~n27147 ;
  assign n27149 = n27145 & n27148 ;
  assign n27150 = n27142 & n27149 ;
  assign n27151 = \wishbone_bd_ram_mem0_reg[162][7]/P0001  & n13726 ;
  assign n27152 = \wishbone_bd_ram_mem0_reg[225][7]/P0001  & n13719 ;
  assign n27153 = ~n27151 & ~n27152 ;
  assign n27154 = \wishbone_bd_ram_mem0_reg[6][7]/P0001  & n13915 ;
  assign n27155 = \wishbone_bd_ram_mem0_reg[220][7]/P0001  & n13965 ;
  assign n27156 = ~n27154 & ~n27155 ;
  assign n27157 = n27153 & n27156 ;
  assign n27158 = \wishbone_bd_ram_mem0_reg[73][7]/P0001  & n13456 ;
  assign n27159 = \wishbone_bd_ram_mem0_reg[4][7]/P0001  & n13527 ;
  assign n27160 = ~n27158 & ~n27159 ;
  assign n27161 = \wishbone_bd_ram_mem0_reg[129][7]/P0001  & n13629 ;
  assign n27162 = \wishbone_bd_ram_mem0_reg[56][7]/P0001  & n13611 ;
  assign n27163 = ~n27161 & ~n27162 ;
  assign n27164 = n27160 & n27163 ;
  assign n27165 = n27157 & n27164 ;
  assign n27166 = n27150 & n27165 ;
  assign n27167 = \wishbone_bd_ram_mem0_reg[145][7]/P0001  & n13715 ;
  assign n27168 = \wishbone_bd_ram_mem0_reg[11][7]/P0001  & n13774 ;
  assign n27169 = ~n27167 & ~n27168 ;
  assign n27170 = \wishbone_bd_ram_mem0_reg[148][7]/P0001  & n13868 ;
  assign n27171 = \wishbone_bd_ram_mem0_reg[121][7]/P0001  & n13983 ;
  assign n27172 = ~n27170 & ~n27171 ;
  assign n27173 = n27169 & n27172 ;
  assign n27174 = \wishbone_bd_ram_mem0_reg[125][7]/P0001  & n13396 ;
  assign n27175 = \wishbone_bd_ram_mem0_reg[54][7]/P0001  & n13622 ;
  assign n27176 = ~n27174 & ~n27175 ;
  assign n27177 = \wishbone_bd_ram_mem0_reg[32][7]/P0001  & n13736 ;
  assign n27178 = \wishbone_bd_ram_mem0_reg[96][7]/P0001  & n13425 ;
  assign n27179 = ~n27177 & ~n27178 ;
  assign n27180 = n27176 & n27179 ;
  assign n27181 = n27173 & n27180 ;
  assign n27182 = \wishbone_bd_ram_mem0_reg[185][7]/P0001  & n13372 ;
  assign n27183 = \wishbone_bd_ram_mem0_reg[241][7]/P0001  & n13854 ;
  assign n27184 = ~n27182 & ~n27183 ;
  assign n27185 = \wishbone_bd_ram_mem0_reg[93][7]/P0001  & n13891 ;
  assign n27186 = \wishbone_bd_ram_mem0_reg[58][7]/P0001  & n13949 ;
  assign n27187 = ~n27185 & ~n27186 ;
  assign n27188 = n27184 & n27187 ;
  assign n27189 = \wishbone_bd_ram_mem0_reg[27][7]/P0001  & n13251 ;
  assign n27190 = \wishbone_bd_ram_mem0_reg[164][7]/P0001  & n13236 ;
  assign n27191 = ~n27189 & ~n27190 ;
  assign n27192 = \wishbone_bd_ram_mem0_reg[216][7]/P0001  & n14005 ;
  assign n27193 = \wishbone_bd_ram_mem0_reg[168][7]/P0001  & n13795 ;
  assign n27194 = ~n27192 & ~n27193 ;
  assign n27195 = n27191 & n27194 ;
  assign n27196 = n27188 & n27195 ;
  assign n27197 = n27181 & n27196 ;
  assign n27198 = n27166 & n27197 ;
  assign n27199 = \wishbone_bd_ram_mem0_reg[203][7]/P0001  & n13816 ;
  assign n27200 = \wishbone_bd_ram_mem0_reg[68][7]/P0001  & n13379 ;
  assign n27201 = ~n27199 & ~n27200 ;
  assign n27202 = \wishbone_bd_ram_mem0_reg[197][7]/P0001  & n13594 ;
  assign n27203 = \wishbone_bd_ram_mem0_reg[228][7]/P0001  & n13497 ;
  assign n27204 = ~n27202 & ~n27203 ;
  assign n27205 = n27201 & n27204 ;
  assign n27206 = \wishbone_bd_ram_mem0_reg[143][7]/P0001  & n13461 ;
  assign n27207 = \wishbone_bd_ram_mem0_reg[110][7]/P0001  & n14030 ;
  assign n27208 = ~n27206 & ~n27207 ;
  assign n27209 = \wishbone_bd_ram_mem0_reg[167][7]/P0001  & n13940 ;
  assign n27210 = \wishbone_bd_ram_mem0_reg[200][7]/P0001  & n13922 ;
  assign n27211 = ~n27209 & ~n27210 ;
  assign n27212 = n27208 & n27211 ;
  assign n27213 = n27205 & n27212 ;
  assign n27214 = \wishbone_bd_ram_mem0_reg[50][7]/P0001  & n13686 ;
  assign n27215 = \wishbone_bd_ram_mem0_reg[97][7]/P0001  & n13724 ;
  assign n27216 = ~n27214 & ~n27215 ;
  assign n27217 = \wishbone_bd_ram_mem0_reg[175][7]/P0001  & n13674 ;
  assign n27218 = \wishbone_bd_ram_mem0_reg[195][7]/P0001  & n13700 ;
  assign n27219 = ~n27217 & ~n27218 ;
  assign n27220 = n27216 & n27219 ;
  assign n27221 = \wishbone_bd_ram_mem0_reg[229][7]/P0001  & n13552 ;
  assign n27222 = \wishbone_bd_ram_mem0_reg[86][7]/P0001  & n13485 ;
  assign n27223 = ~n27221 & ~n27222 ;
  assign n27224 = \wishbone_bd_ram_mem0_reg[208][7]/P0001  & n14010 ;
  assign n27225 = \wishbone_bd_ram_mem0_reg[67][7]/P0001  & n13663 ;
  assign n27226 = ~n27224 & ~n27225 ;
  assign n27227 = n27223 & n27226 ;
  assign n27228 = n27220 & n27227 ;
  assign n27229 = n27213 & n27228 ;
  assign n27230 = \wishbone_bd_ram_mem0_reg[146][7]/P0001  & n13958 ;
  assign n27231 = \wishbone_bd_ram_mem0_reg[45][7]/P0001  & n13420 ;
  assign n27232 = ~n27230 & ~n27231 ;
  assign n27233 = \wishbone_bd_ram_mem0_reg[106][7]/P0001  & n13555 ;
  assign n27234 = \wishbone_bd_ram_mem0_reg[177][7]/P0001  & n13863 ;
  assign n27235 = ~n27233 & ~n27234 ;
  assign n27236 = n27232 & n27235 ;
  assign n27237 = \wishbone_bd_ram_mem0_reg[48][7]/P0001  & n13917 ;
  assign n27238 = \wishbone_bd_ram_mem0_reg[43][7]/P0001  & n13761 ;
  assign n27239 = ~n27237 & ~n27238 ;
  assign n27240 = \wishbone_bd_ram_mem0_reg[142][7]/P0001  & n13448 ;
  assign n27241 = \wishbone_bd_ram_mem0_reg[199][7]/P0001  & n13499 ;
  assign n27242 = ~n27240 & ~n27241 ;
  assign n27243 = n27239 & n27242 ;
  assign n27244 = n27236 & n27243 ;
  assign n27245 = \wishbone_bd_ram_mem0_reg[36][7]/P0001  & n13639 ;
  assign n27246 = \wishbone_bd_ram_mem0_reg[194][7]/P0001  & n13624 ;
  assign n27247 = ~n27245 & ~n27246 ;
  assign n27248 = \wishbone_bd_ram_mem0_reg[202][7]/P0001  & n13268 ;
  assign n27249 = \wishbone_bd_ram_mem0_reg[71][7]/P0001  & n13636 ;
  assign n27250 = ~n27248 & ~n27249 ;
  assign n27251 = n27247 & n27250 ;
  assign n27252 = \wishbone_bd_ram_mem0_reg[53][7]/P0001  & n13875 ;
  assign n27253 = \wishbone_bd_ram_mem0_reg[154][7]/P0001  & n13403 ;
  assign n27254 = ~n27252 & ~n27253 ;
  assign n27255 = \wishbone_bd_ram_mem0_reg[12][7]/P0001  & n13733 ;
  assign n27256 = \wishbone_bd_ram_mem0_reg[236][7]/P0001  & n13480 ;
  assign n27257 = ~n27255 & ~n27256 ;
  assign n27258 = n27254 & n27257 ;
  assign n27259 = n27251 & n27258 ;
  assign n27260 = n27244 & n27259 ;
  assign n27261 = n27229 & n27260 ;
  assign n27262 = n27198 & n27261 ;
  assign n27263 = n27135 & n27262 ;
  assign n27264 = n27008 & n27263 ;
  assign n27265 = ~wb_rst_i_pad & ~n26752 ;
  assign n27266 = ~n27264 & n27265 ;
  assign n27267 = ~n26753 & ~n27266 ;
  assign n27268 = \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  & n23751 ;
  assign n27269 = n23741 & n27268 ;
  assign n27270 = \ethreg1_MODER_1_DataOut_reg[0]/NET0131  & n23808 ;
  assign n27271 = ~n27269 & ~n27270 ;
  assign n27272 = \ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131  & n23782 ;
  assign n27273 = \ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131  & n23743 ;
  assign n27274 = n23741 & n27273 ;
  assign n27275 = ~n27272 & ~n27274 ;
  assign n27276 = n27271 & n27275 ;
  assign n27277 = \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131  & n23813 ;
  assign n27278 = \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131  & n25084 ;
  assign n27279 = ~n27277 & ~n27278 ;
  assign n27280 = n23730 & n27279 ;
  assign n27281 = n27276 & n27280 ;
  assign n27282 = \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  & n23737 ;
  assign n27283 = \ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131  & n23743 ;
  assign n27284 = n23747 & n27283 ;
  assign n27285 = \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  & n23751 ;
  assign n27286 = n23747 & n27285 ;
  assign n27287 = ~n27284 & ~n27286 ;
  assign n27288 = \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131  & n23794 ;
  assign n27289 = n23741 & n27288 ;
  assign n27290 = \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131  & n23802 ;
  assign n27291 = ~n27289 & ~n27290 ;
  assign n27292 = n27287 & n27291 ;
  assign n27293 = ~n27282 & n27292 ;
  assign n27294 = n27281 & n27293 ;
  assign n27295 = n23730 & ~n27294 ;
  assign n27296 = \wishbone_bd_ram_mem1_reg[239][8]/P0001  & n13349 ;
  assign n27297 = \wishbone_bd_ram_mem1_reg[33][8]/P0001  & n13933 ;
  assign n27298 = ~n27296 & ~n27297 ;
  assign n27299 = \wishbone_bd_ram_mem1_reg[72][8]/P0001  & n13582 ;
  assign n27300 = \wishbone_bd_ram_mem1_reg[223][8]/P0001  & n13335 ;
  assign n27301 = ~n27299 & ~n27300 ;
  assign n27302 = n27298 & n27301 ;
  assign n27303 = \wishbone_bd_ram_mem1_reg[92][8]/P0001  & n13859 ;
  assign n27304 = \wishbone_bd_ram_mem1_reg[232][8]/P0001  & n13510 ;
  assign n27305 = ~n27303 & ~n27304 ;
  assign n27306 = \wishbone_bd_ram_mem1_reg[118][8]/P0001  & n13589 ;
  assign n27307 = \wishbone_bd_ram_mem1_reg[4][8]/P0001  & n13527 ;
  assign n27308 = ~n27306 & ~n27307 ;
  assign n27309 = n27305 & n27308 ;
  assign n27310 = n27302 & n27309 ;
  assign n27311 = \wishbone_bd_ram_mem1_reg[190][8]/P0001  & n13365 ;
  assign n27312 = \wishbone_bd_ram_mem1_reg[43][8]/P0001  & n13761 ;
  assign n27313 = ~n27311 & ~n27312 ;
  assign n27314 = \wishbone_bd_ram_mem1_reg[57][8]/P0001  & n13731 ;
  assign n27315 = \wishbone_bd_ram_mem1_reg[188][8]/P0001  & n13407 ;
  assign n27316 = ~n27314 & ~n27315 ;
  assign n27317 = n27313 & n27316 ;
  assign n27318 = \wishbone_bd_ram_mem1_reg[35][8]/P0001  & n13523 ;
  assign n27319 = \wishbone_bd_ram_mem1_reg[226][8]/P0001  & n13668 ;
  assign n27320 = ~n27318 & ~n27319 ;
  assign n27321 = \wishbone_bd_ram_mem1_reg[66][8]/P0001  & n13603 ;
  assign n27322 = \wishbone_bd_ram_mem1_reg[89][8]/P0001  & n13910 ;
  assign n27323 = ~n27321 & ~n27322 ;
  assign n27324 = n27320 & n27323 ;
  assign n27325 = n27317 & n27324 ;
  assign n27326 = n27310 & n27325 ;
  assign n27327 = \wishbone_bd_ram_mem1_reg[145][8]/P0001  & n13715 ;
  assign n27328 = \wishbone_bd_ram_mem1_reg[174][8]/P0001  & n13899 ;
  assign n27329 = ~n27327 & ~n27328 ;
  assign n27330 = \wishbone_bd_ram_mem1_reg[42][8]/P0001  & n13341 ;
  assign n27331 = \wishbone_bd_ram_mem1_reg[117][8]/P0001  & n13557 ;
  assign n27332 = ~n27330 & ~n27331 ;
  assign n27333 = n27329 & n27332 ;
  assign n27334 = \wishbone_bd_ram_mem1_reg[229][8]/P0001  & n13552 ;
  assign n27335 = \wishbone_bd_ram_mem1_reg[127][8]/P0001  & n13803 ;
  assign n27336 = ~n27334 & ~n27335 ;
  assign n27337 = \wishbone_bd_ram_mem1_reg[46][8]/P0001  & n13298 ;
  assign n27338 = \wishbone_bd_ram_mem1_reg[44][8]/P0001  & n13291 ;
  assign n27339 = ~n27337 & ~n27338 ;
  assign n27340 = n27336 & n27339 ;
  assign n27341 = n27333 & n27340 ;
  assign n27342 = \wishbone_bd_ram_mem1_reg[180][8]/P0001  & n13650 ;
  assign n27343 = \wishbone_bd_ram_mem1_reg[178][8]/P0001  & n13301 ;
  assign n27344 = ~n27342 & ~n27343 ;
  assign n27345 = \wishbone_bd_ram_mem1_reg[252][8]/P0001  & n13986 ;
  assign n27346 = \wishbone_bd_ram_mem1_reg[5][8]/P0001  & n13243 ;
  assign n27347 = ~n27345 & ~n27346 ;
  assign n27348 = n27344 & n27347 ;
  assign n27349 = \wishbone_bd_ram_mem1_reg[18][8]/P0001  & n13532 ;
  assign n27350 = \wishbone_bd_ram_mem1_reg[211][8]/P0001  & n13805 ;
  assign n27351 = ~n27349 & ~n27350 ;
  assign n27352 = \wishbone_bd_ram_mem1_reg[171][8]/P0001  & n13422 ;
  assign n27353 = \wishbone_bd_ram_mem1_reg[48][8]/P0001  & n13917 ;
  assign n27354 = ~n27352 & ~n27353 ;
  assign n27355 = n27351 & n27354 ;
  assign n27356 = n27348 & n27355 ;
  assign n27357 = n27341 & n27356 ;
  assign n27358 = n27326 & n27357 ;
  assign n27359 = \wishbone_bd_ram_mem1_reg[255][8]/P0001  & n13952 ;
  assign n27360 = \wishbone_bd_ram_mem1_reg[111][8]/P0001  & n13471 ;
  assign n27361 = ~n27359 & ~n27360 ;
  assign n27362 = \wishbone_bd_ram_mem1_reg[210][8]/P0001  & n13443 ;
  assign n27363 = \wishbone_bd_ram_mem1_reg[19][8]/P0001  & n13886 ;
  assign n27364 = ~n27362 & ~n27363 ;
  assign n27365 = n27361 & n27364 ;
  assign n27366 = \wishbone_bd_ram_mem1_reg[204][8]/P0001  & n13821 ;
  assign n27367 = \wishbone_bd_ram_mem1_reg[160][8]/P0001  & n13271 ;
  assign n27368 = ~n27366 & ~n27367 ;
  assign n27369 = \wishbone_bd_ram_mem1_reg[97][8]/P0001  & n13724 ;
  assign n27370 = \wishbone_bd_ram_mem1_reg[120][8]/P0001  & n13550 ;
  assign n27371 = ~n27369 & ~n27370 ;
  assign n27372 = n27368 & n27371 ;
  assign n27373 = n27365 & n27372 ;
  assign n27374 = \wishbone_bd_ram_mem1_reg[156][8]/P0001  & n13769 ;
  assign n27375 = \wishbone_bd_ram_mem1_reg[31][8]/P0001  & n13758 ;
  assign n27376 = ~n27374 & ~n27375 ;
  assign n27377 = \wishbone_bd_ram_mem1_reg[99][8]/P0001  & n13996 ;
  assign n27378 = \wishbone_bd_ram_mem1_reg[91][8]/P0001  & n13954 ;
  assign n27379 = ~n27377 & ~n27378 ;
  assign n27380 = n27376 & n27379 ;
  assign n27381 = \wishbone_bd_ram_mem1_reg[198][8]/P0001  & n13592 ;
  assign n27382 = \wishbone_bd_ram_mem1_reg[32][8]/P0001  & n13736 ;
  assign n27383 = ~n27381 & ~n27382 ;
  assign n27384 = \wishbone_bd_ram_mem1_reg[49][8]/P0001  & n13929 ;
  assign n27385 = \wishbone_bd_ram_mem1_reg[251][8]/P0001  & n14019 ;
  assign n27386 = ~n27384 & ~n27385 ;
  assign n27387 = n27383 & n27386 ;
  assign n27388 = n27380 & n27387 ;
  assign n27389 = n27373 & n27388 ;
  assign n27390 = \wishbone_bd_ram_mem1_reg[129][8]/P0001  & n13629 ;
  assign n27391 = \wishbone_bd_ram_mem1_reg[104][8]/P0001  & n13684 ;
  assign n27392 = ~n27390 & ~n27391 ;
  assign n27393 = \wishbone_bd_ram_mem1_reg[107][8]/P0001  & n13476 ;
  assign n27394 = \wishbone_bd_ram_mem1_reg[231][8]/P0001  & n13363 ;
  assign n27395 = ~n27393 & ~n27394 ;
  assign n27396 = n27392 & n27395 ;
  assign n27397 = \wishbone_bd_ram_mem1_reg[181][8]/P0001  & n13587 ;
  assign n27398 = \wishbone_bd_ram_mem1_reg[113][8]/P0001  & n13882 ;
  assign n27399 = ~n27397 & ~n27398 ;
  assign n27400 = \wishbone_bd_ram_mem1_reg[85][8]/P0001  & n13784 ;
  assign n27401 = \wishbone_bd_ram_mem1_reg[30][8]/P0001  & n13713 ;
  assign n27402 = ~n27400 & ~n27401 ;
  assign n27403 = n27399 & n27402 ;
  assign n27404 = n27396 & n27403 ;
  assign n27405 = \wishbone_bd_ram_mem1_reg[202][8]/P0001  & n13268 ;
  assign n27406 = \wishbone_bd_ram_mem1_reg[86][8]/P0001  & n13485 ;
  assign n27407 = ~n27405 & ~n27406 ;
  assign n27408 = \wishbone_bd_ram_mem1_reg[137][8]/P0001  & n13808 ;
  assign n27409 = \wishbone_bd_ram_mem1_reg[29][8]/P0001  & n13412 ;
  assign n27410 = ~n27408 & ~n27409 ;
  assign n27411 = n27407 & n27410 ;
  assign n27412 = \wishbone_bd_ram_mem1_reg[159][8]/P0001  & n13627 ;
  assign n27413 = \wishbone_bd_ram_mem1_reg[240][8]/P0001  & n13352 ;
  assign n27414 = ~n27412 & ~n27413 ;
  assign n27415 = \wishbone_bd_ram_mem1_reg[16][8]/P0001  & n13695 ;
  assign n27416 = \wishbone_bd_ram_mem1_reg[68][8]/P0001  & n13379 ;
  assign n27417 = ~n27415 & ~n27416 ;
  assign n27418 = n27414 & n27417 ;
  assign n27419 = n27411 & n27418 ;
  assign n27420 = n27404 & n27419 ;
  assign n27421 = n27389 & n27420 ;
  assign n27422 = n27358 & n27421 ;
  assign n27423 = \wishbone_bd_ram_mem1_reg[78][8]/P0001  & n13277 ;
  assign n27424 = \wishbone_bd_ram_mem1_reg[228][8]/P0001  & n13497 ;
  assign n27425 = ~n27423 & ~n27424 ;
  assign n27426 = \wishbone_bd_ram_mem1_reg[236][8]/P0001  & n13480 ;
  assign n27427 = \wishbone_bd_ram_mem1_reg[144][8]/P0001  & n13508 ;
  assign n27428 = ~n27426 & ~n27427 ;
  assign n27429 = n27425 & n27428 ;
  assign n27430 = \wishbone_bd_ram_mem1_reg[166][8]/P0001  & n13999 ;
  assign n27431 = \wishbone_bd_ram_mem1_reg[133][8]/P0001  & n13492 ;
  assign n27432 = ~n27430 & ~n27431 ;
  assign n27433 = \wishbone_bd_ram_mem1_reg[170][8]/P0001  & n14007 ;
  assign n27434 = \wishbone_bd_ram_mem1_reg[173][8]/P0001  & n13360 ;
  assign n27435 = ~n27433 & ~n27434 ;
  assign n27436 = n27432 & n27435 ;
  assign n27437 = n27429 & n27436 ;
  assign n27438 = \wishbone_bd_ram_mem1_reg[237][8]/P0001  & n13924 ;
  assign n27439 = \wishbone_bd_ram_mem1_reg[59][8]/P0001  & n13613 ;
  assign n27440 = ~n27438 & ~n27439 ;
  assign n27441 = \wishbone_bd_ram_mem1_reg[184][8]/P0001  & n13960 ;
  assign n27442 = \wishbone_bd_ram_mem1_reg[95][8]/P0001  & n13317 ;
  assign n27443 = ~n27441 & ~n27442 ;
  assign n27444 = n27440 & n27443 ;
  assign n27445 = \wishbone_bd_ram_mem1_reg[186][8]/P0001  & n13616 ;
  assign n27446 = \wishbone_bd_ram_mem1_reg[131][8]/P0001  & n13358 ;
  assign n27447 = ~n27445 & ~n27446 ;
  assign n27448 = \wishbone_bd_ram_mem1_reg[143][8]/P0001  & n13461 ;
  assign n27449 = \wishbone_bd_ram_mem1_reg[193][8]/P0001  & n14022 ;
  assign n27450 = ~n27448 & ~n27449 ;
  assign n27451 = n27447 & n27450 ;
  assign n27452 = n27444 & n27451 ;
  assign n27453 = n27437 & n27452 ;
  assign n27454 = \wishbone_bd_ram_mem1_reg[98][8]/P0001  & n13569 ;
  assign n27455 = \wishbone_bd_ram_mem1_reg[84][8]/P0001  & n13385 ;
  assign n27456 = ~n27454 & ~n27455 ;
  assign n27457 = \wishbone_bd_ram_mem1_reg[148][8]/P0001  & n13868 ;
  assign n27458 = \wishbone_bd_ram_mem1_reg[115][8]/P0001  & n13747 ;
  assign n27459 = ~n27457 & ~n27458 ;
  assign n27460 = n27456 & n27459 ;
  assign n27461 = \wishbone_bd_ram_mem1_reg[2][8]/P0001  & n13975 ;
  assign n27462 = \wishbone_bd_ram_mem1_reg[56][8]/P0001  & n13611 ;
  assign n27463 = ~n27461 & ~n27462 ;
  assign n27464 = \wishbone_bd_ram_mem1_reg[27][8]/P0001  & n13251 ;
  assign n27465 = \wishbone_bd_ram_mem1_reg[189][8]/P0001  & n14001 ;
  assign n27466 = ~n27464 & ~n27465 ;
  assign n27467 = n27463 & n27466 ;
  assign n27468 = n27460 & n27467 ;
  assign n27469 = \wishbone_bd_ram_mem1_reg[50][8]/P0001  & n13686 ;
  assign n27470 = \wishbone_bd_ram_mem1_reg[177][8]/P0001  & n13863 ;
  assign n27471 = ~n27469 & ~n27470 ;
  assign n27472 = \wishbone_bd_ram_mem1_reg[135][8]/P0001  & n13672 ;
  assign n27473 = \wishbone_bd_ram_mem1_reg[51][8]/P0001  & n13880 ;
  assign n27474 = ~n27472 & ~n27473 ;
  assign n27475 = n27471 & n27474 ;
  assign n27476 = \wishbone_bd_ram_mem1_reg[3][8]/P0001  & n13354 ;
  assign n27477 = \wishbone_bd_ram_mem1_reg[253][8]/P0001  & n13708 ;
  assign n27478 = ~n27476 & ~n27477 ;
  assign n27479 = \wishbone_bd_ram_mem1_reg[191][8]/P0001  & n14012 ;
  assign n27480 = \wishbone_bd_ram_mem1_reg[152][8]/P0001  & n13912 ;
  assign n27481 = ~n27479 & ~n27480 ;
  assign n27482 = n27478 & n27481 ;
  assign n27483 = n27475 & n27482 ;
  assign n27484 = n27468 & n27483 ;
  assign n27485 = n27453 & n27484 ;
  assign n27486 = \wishbone_bd_ram_mem1_reg[165][8]/P0001  & n14028 ;
  assign n27487 = \wishbone_bd_ram_mem1_reg[10][8]/P0001  & n13837 ;
  assign n27488 = ~n27486 & ~n27487 ;
  assign n27489 = \wishbone_bd_ram_mem1_reg[125][8]/P0001  & n13396 ;
  assign n27490 = \wishbone_bd_ram_mem1_reg[140][8]/P0001  & n13287 ;
  assign n27491 = ~n27489 & ~n27490 ;
  assign n27492 = n27488 & n27491 ;
  assign n27493 = \wishbone_bd_ram_mem1_reg[205][8]/P0001  & n13947 ;
  assign n27494 = \wishbone_bd_ram_mem1_reg[201][8]/P0001  & n13600 ;
  assign n27495 = ~n27493 & ~n27494 ;
  assign n27496 = \wishbone_bd_ram_mem1_reg[1][8]/P0001  & n13888 ;
  assign n27497 = \wishbone_bd_ram_mem1_reg[96][8]/P0001  & n13425 ;
  assign n27498 = ~n27496 & ~n27497 ;
  assign n27499 = n27495 & n27498 ;
  assign n27500 = n27492 & n27499 ;
  assign n27501 = \wishbone_bd_ram_mem1_reg[213][8]/P0001  & n13870 ;
  assign n27502 = \wishbone_bd_ram_mem1_reg[161][8]/P0001  & n13505 ;
  assign n27503 = ~n27501 & ~n27502 ;
  assign n27504 = \wishbone_bd_ram_mem1_reg[163][8]/P0001  & n13255 ;
  assign n27505 = \wishbone_bd_ram_mem1_reg[185][8]/P0001  & n13372 ;
  assign n27506 = ~n27504 & ~n27505 ;
  assign n27507 = n27503 & n27506 ;
  assign n27508 = \wishbone_bd_ram_mem1_reg[121][8]/P0001  & n13983 ;
  assign n27509 = \wishbone_bd_ram_mem1_reg[254][8]/P0001  & n13283 ;
  assign n27510 = ~n27508 & ~n27509 ;
  assign n27511 = \wishbone_bd_ram_mem1_reg[101][8]/P0001  & n13772 ;
  assign n27512 = \wishbone_bd_ram_mem1_reg[162][8]/P0001  & n13726 ;
  assign n27513 = ~n27511 & ~n27512 ;
  assign n27514 = n27510 & n27513 ;
  assign n27515 = n27507 & n27514 ;
  assign n27516 = n27500 & n27515 ;
  assign n27517 = \wishbone_bd_ram_mem1_reg[119][8]/P0001  & n14033 ;
  assign n27518 = \wishbone_bd_ram_mem1_reg[138][8]/P0001  & n13398 ;
  assign n27519 = ~n27517 & ~n27518 ;
  assign n27520 = \wishbone_bd_ram_mem1_reg[241][8]/P0001  & n13854 ;
  assign n27521 = \wishbone_bd_ram_mem1_reg[36][8]/P0001  & n13639 ;
  assign n27522 = ~n27520 & ~n27521 ;
  assign n27523 = n27519 & n27522 ;
  assign n27524 = \wishbone_bd_ram_mem1_reg[168][8]/P0001  & n13795 ;
  assign n27525 = \wishbone_bd_ram_mem1_reg[221][8]/P0001  & n13641 ;
  assign n27526 = ~n27524 & ~n27525 ;
  assign n27527 = \wishbone_bd_ram_mem1_reg[25][8]/P0001  & n13742 ;
  assign n27528 = \wishbone_bd_ram_mem1_reg[218][8]/P0001  & n13792 ;
  assign n27529 = ~n27527 & ~n27528 ;
  assign n27530 = n27526 & n27529 ;
  assign n27531 = n27523 & n27530 ;
  assign n27532 = \wishbone_bd_ram_mem1_reg[58][8]/P0001  & n13949 ;
  assign n27533 = \wishbone_bd_ram_mem1_reg[123][8]/P0001  & n13749 ;
  assign n27534 = ~n27532 & ~n27533 ;
  assign n27535 = \wishbone_bd_ram_mem1_reg[75][8]/P0001  & n13605 ;
  assign n27536 = \wishbone_bd_ram_mem1_reg[215][8]/P0001  & n13901 ;
  assign n27537 = ~n27535 & ~n27536 ;
  assign n27538 = n27534 & n27537 ;
  assign n27539 = \wishbone_bd_ram_mem1_reg[200][8]/P0001  & n13922 ;
  assign n27540 = \wishbone_bd_ram_mem1_reg[249][8]/P0001  & n13431 ;
  assign n27541 = ~n27539 & ~n27540 ;
  assign n27542 = \wishbone_bd_ram_mem1_reg[151][8]/P0001  & n13697 ;
  assign n27543 = \wishbone_bd_ram_mem1_reg[157][8]/P0001  & n13445 ;
  assign n27544 = ~n27542 & ~n27543 ;
  assign n27545 = n27541 & n27544 ;
  assign n27546 = n27538 & n27545 ;
  assign n27547 = n27531 & n27546 ;
  assign n27548 = n27516 & n27547 ;
  assign n27549 = n27485 & n27548 ;
  assign n27550 = n27422 & n27549 ;
  assign n27551 = \wishbone_bd_ram_mem1_reg[21][8]/P0001  & n13438 ;
  assign n27552 = \wishbone_bd_ram_mem1_reg[164][8]/P0001  & n13236 ;
  assign n27553 = ~n27551 & ~n27552 ;
  assign n27554 = \wishbone_bd_ram_mem1_reg[81][8]/P0001  & n13409 ;
  assign n27555 = \wishbone_bd_ram_mem1_reg[187][8]/P0001  & n13756 ;
  assign n27556 = ~n27554 & ~n27555 ;
  assign n27557 = n27553 & n27556 ;
  assign n27558 = \wishbone_bd_ram_mem1_reg[126][8]/P0001  & n13786 ;
  assign n27559 = \wishbone_bd_ram_mem1_reg[209][8]/P0001  & n13689 ;
  assign n27560 = ~n27558 & ~n27559 ;
  assign n27561 = \wishbone_bd_ram_mem1_reg[245][8]/P0001  & n13877 ;
  assign n27562 = \wishbone_bd_ram_mem1_reg[208][8]/P0001  & n14010 ;
  assign n27563 = ~n27561 & ~n27562 ;
  assign n27564 = n27560 & n27563 ;
  assign n27565 = n27557 & n27564 ;
  assign n27566 = \wishbone_bd_ram_mem1_reg[146][8]/P0001  & n13958 ;
  assign n27567 = \wishbone_bd_ram_mem1_reg[67][8]/P0001  & n13663 ;
  assign n27568 = ~n27566 & ~n27567 ;
  assign n27569 = \wishbone_bd_ram_mem1_reg[183][8]/P0001  & n13645 ;
  assign n27570 = \wishbone_bd_ram_mem1_reg[167][8]/P0001  & n13940 ;
  assign n27571 = ~n27569 & ~n27570 ;
  assign n27572 = n27568 & n27571 ;
  assign n27573 = \wishbone_bd_ram_mem1_reg[38][8]/P0001  & n13828 ;
  assign n27574 = \wishbone_bd_ram_mem1_reg[230][8]/P0001  & n13994 ;
  assign n27575 = ~n27573 & ~n27574 ;
  assign n27576 = \wishbone_bd_ram_mem1_reg[124][8]/P0001  & n14024 ;
  assign n27577 = \wishbone_bd_ram_mem1_reg[73][8]/P0001  & n13456 ;
  assign n27578 = ~n27576 & ~n27577 ;
  assign n27579 = n27575 & n27578 ;
  assign n27580 = n27572 & n27579 ;
  assign n27581 = n27565 & n27580 ;
  assign n27582 = \wishbone_bd_ram_mem1_reg[246][8]/P0001  & n13981 ;
  assign n27583 = \wishbone_bd_ram_mem1_reg[65][8]/P0001  & n13842 ;
  assign n27584 = ~n27582 & ~n27583 ;
  assign n27585 = \wishbone_bd_ram_mem1_reg[64][8]/P0001  & n13904 ;
  assign n27586 = \wishbone_bd_ram_mem1_reg[103][8]/P0001  & n13320 ;
  assign n27587 = ~n27585 & ~n27586 ;
  assign n27588 = n27584 & n27587 ;
  assign n27589 = \wishbone_bd_ram_mem1_reg[250][8]/P0001  & n13677 ;
  assign n27590 = \wishbone_bd_ram_mem1_reg[110][8]/P0001  & n14030 ;
  assign n27591 = ~n27589 & ~n27590 ;
  assign n27592 = \wishbone_bd_ram_mem1_reg[222][8]/P0001  & n13721 ;
  assign n27593 = \wishbone_bd_ram_mem1_reg[158][8]/P0001  & n13294 ;
  assign n27594 = ~n27592 & ~n27593 ;
  assign n27595 = n27591 & n27594 ;
  assign n27596 = n27588 & n27595 ;
  assign n27597 = \wishbone_bd_ram_mem1_reg[149][8]/P0001  & n13469 ;
  assign n27598 = \wishbone_bd_ram_mem1_reg[8][8]/P0001  & n13459 ;
  assign n27599 = ~n27597 & ~n27598 ;
  assign n27600 = \wishbone_bd_ram_mem1_reg[11][8]/P0001  & n13774 ;
  assign n27601 = \wishbone_bd_ram_mem1_reg[55][8]/P0001  & n13618 ;
  assign n27602 = ~n27600 & ~n27601 ;
  assign n27603 = n27599 & n27602 ;
  assign n27604 = \wishbone_bd_ram_mem1_reg[109][8]/P0001  & n13306 ;
  assign n27605 = \wishbone_bd_ram_mem1_reg[219][8]/P0001  & n13577 ;
  assign n27606 = ~n27604 & ~n27605 ;
  assign n27607 = \wishbone_bd_ram_mem1_reg[71][8]/P0001  & n13636 ;
  assign n27608 = \wishbone_bd_ram_mem1_reg[54][8]/P0001  & n13622 ;
  assign n27609 = ~n27607 & ~n27608 ;
  assign n27610 = n27606 & n27609 ;
  assign n27611 = n27603 & n27610 ;
  assign n27612 = n27596 & n27611 ;
  assign n27613 = n27581 & n27612 ;
  assign n27614 = \wishbone_bd_ram_mem1_reg[225][8]/P0001  & n13719 ;
  assign n27615 = \wishbone_bd_ram_mem1_reg[7][8]/P0001  & n13546 ;
  assign n27616 = ~n27614 & ~n27615 ;
  assign n27617 = \wishbone_bd_ram_mem1_reg[9][8]/P0001  & n13580 ;
  assign n27618 = \wishbone_bd_ram_mem1_reg[242][8]/P0001  & n13383 ;
  assign n27619 = ~n27617 & ~n27618 ;
  assign n27620 = n27616 & n27619 ;
  assign n27621 = \wishbone_bd_ram_mem1_reg[207][8]/P0001  & n13826 ;
  assign n27622 = \wishbone_bd_ram_mem1_reg[90][8]/P0001  & n13906 ;
  assign n27623 = ~n27621 & ~n27622 ;
  assign n27624 = \wishbone_bd_ram_mem1_reg[150][8]/P0001  & n13666 ;
  assign n27625 = \wishbone_bd_ram_mem1_reg[147][8]/P0001  & n13702 ;
  assign n27626 = ~n27624 & ~n27625 ;
  assign n27627 = n27623 & n27626 ;
  assign n27628 = n27620 & n27627 ;
  assign n27629 = \wishbone_bd_ram_mem1_reg[52][8]/P0001  & n13988 ;
  assign n27630 = \wishbone_bd_ram_mem1_reg[105][8]/P0001  & n13503 ;
  assign n27631 = ~n27629 & ~n27630 ;
  assign n27632 = \wishbone_bd_ram_mem1_reg[79][8]/P0001  & n13779 ;
  assign n27633 = \wishbone_bd_ram_mem1_reg[224][8]/P0001  & n13433 ;
  assign n27634 = ~n27632 & ~n27633 ;
  assign n27635 = n27631 & n27634 ;
  assign n27636 = \wishbone_bd_ram_mem1_reg[61][8]/P0001  & n13544 ;
  assign n27637 = \wishbone_bd_ram_mem1_reg[93][8]/P0001  & n13891 ;
  assign n27638 = ~n27636 & ~n27637 ;
  assign n27639 = \wishbone_bd_ram_mem1_reg[83][8]/P0001  & n13454 ;
  assign n27640 = \wishbone_bd_ram_mem1_reg[41][8]/P0001  & n14017 ;
  assign n27641 = ~n27639 & ~n27640 ;
  assign n27642 = n27638 & n27641 ;
  assign n27643 = n27635 & n27642 ;
  assign n27644 = n27628 & n27643 ;
  assign n27645 = \wishbone_bd_ram_mem1_reg[197][8]/P0001  & n13594 ;
  assign n27646 = \wishbone_bd_ram_mem1_reg[203][8]/P0001  & n13816 ;
  assign n27647 = ~n27645 & ~n27646 ;
  assign n27648 = \wishbone_bd_ram_mem1_reg[116][8]/P0001  & n13865 ;
  assign n27649 = \wishbone_bd_ram_mem1_reg[6][8]/P0001  & n13915 ;
  assign n27650 = ~n27648 & ~n27649 ;
  assign n27651 = n27647 & n27650 ;
  assign n27652 = \wishbone_bd_ram_mem1_reg[130][8]/P0001  & n13427 ;
  assign n27653 = \wishbone_bd_ram_mem1_reg[243][8]/P0001  & n13575 ;
  assign n27654 = ~n27652 & ~n27653 ;
  assign n27655 = \wishbone_bd_ram_mem1_reg[227][8]/P0001  & n13388 ;
  assign n27656 = \wishbone_bd_ram_mem1_reg[235][8]/P0001  & n13518 ;
  assign n27657 = ~n27655 & ~n27656 ;
  assign n27658 = n27654 & n27657 ;
  assign n27659 = n27651 & n27658 ;
  assign n27660 = \wishbone_bd_ram_mem1_reg[238][8]/P0001  & n13819 ;
  assign n27661 = \wishbone_bd_ram_mem1_reg[128][8]/P0001  & n13652 ;
  assign n27662 = ~n27660 & ~n27661 ;
  assign n27663 = \wishbone_bd_ram_mem1_reg[214][8]/P0001  & n13938 ;
  assign n27664 = \wishbone_bd_ram_mem1_reg[172][8]/P0001  & n13377 ;
  assign n27665 = ~n27663 & ~n27664 ;
  assign n27666 = n27662 & n27665 ;
  assign n27667 = \wishbone_bd_ram_mem1_reg[15][8]/P0001  & n13797 ;
  assign n27668 = \wishbone_bd_ram_mem1_reg[47][8]/P0001  & n13436 ;
  assign n27669 = ~n27667 & ~n27668 ;
  assign n27670 = \wishbone_bd_ram_mem1_reg[114][8]/P0001  & n13763 ;
  assign n27671 = \wishbone_bd_ram_mem1_reg[106][8]/P0001  & n13555 ;
  assign n27672 = ~n27670 & ~n27671 ;
  assign n27673 = n27669 & n27672 ;
  assign n27674 = n27666 & n27673 ;
  assign n27675 = n27659 & n27674 ;
  assign n27676 = n27644 & n27675 ;
  assign n27677 = n27613 & n27676 ;
  assign n27678 = \wishbone_bd_ram_mem1_reg[34][8]/P0001  & n13450 ;
  assign n27679 = \wishbone_bd_ram_mem1_reg[139][8]/P0001  & n13566 ;
  assign n27680 = ~n27678 & ~n27679 ;
  assign n27681 = \wishbone_bd_ram_mem1_reg[45][8]/P0001  & n13420 ;
  assign n27682 = \wishbone_bd_ram_mem1_reg[100][8]/P0001  & n13401 ;
  assign n27683 = ~n27681 & ~n27682 ;
  assign n27684 = n27680 & n27683 ;
  assign n27685 = \wishbone_bd_ram_mem1_reg[102][8]/P0001  & n13534 ;
  assign n27686 = \wishbone_bd_ram_mem1_reg[53][8]/P0001  & n13875 ;
  assign n27687 = ~n27685 & ~n27686 ;
  assign n27688 = \wishbone_bd_ram_mem1_reg[80][8]/P0001  & n13516 ;
  assign n27689 = \wishbone_bd_ram_mem1_reg[70][8]/P0001  & n13339 ;
  assign n27690 = ~n27688 & ~n27689 ;
  assign n27691 = n27687 & n27690 ;
  assign n27692 = n27684 & n27691 ;
  assign n27693 = \wishbone_bd_ram_mem1_reg[142][8]/P0001  & n13448 ;
  assign n27694 = \wishbone_bd_ram_mem1_reg[169][8]/P0001  & n13541 ;
  assign n27695 = ~n27693 & ~n27694 ;
  assign n27696 = \wishbone_bd_ram_mem1_reg[74][8]/P0001  & n13564 ;
  assign n27697 = \wishbone_bd_ram_mem1_reg[212][8]/P0001  & n13634 ;
  assign n27698 = ~n27696 & ~n27697 ;
  assign n27699 = n27695 & n27698 ;
  assign n27700 = \wishbone_bd_ram_mem1_reg[14][8]/P0001  & n13972 ;
  assign n27701 = \wishbone_bd_ram_mem1_reg[13][8]/P0001  & n13844 ;
  assign n27702 = ~n27700 & ~n27701 ;
  assign n27703 = \wishbone_bd_ram_mem1_reg[216][8]/P0001  & n14005 ;
  assign n27704 = \wishbone_bd_ram_mem1_reg[26][8]/P0001  & n13521 ;
  assign n27705 = ~n27703 & ~n27704 ;
  assign n27706 = n27702 & n27705 ;
  assign n27707 = n27699 & n27706 ;
  assign n27708 = n27692 & n27707 ;
  assign n27709 = \wishbone_bd_ram_mem1_reg[77][8]/P0001  & n13935 ;
  assign n27710 = \wishbone_bd_ram_mem1_reg[217][8]/P0001  & n13767 ;
  assign n27711 = ~n27709 & ~n27710 ;
  assign n27712 = \wishbone_bd_ram_mem1_reg[20][8]/P0001  & n13839 ;
  assign n27713 = \wishbone_bd_ram_mem1_reg[88][8]/P0001  & n13347 ;
  assign n27714 = ~n27712 & ~n27713 ;
  assign n27715 = n27711 & n27714 ;
  assign n27716 = \wishbone_bd_ram_mem1_reg[39][8]/P0001  & n13893 ;
  assign n27717 = \wishbone_bd_ram_mem1_reg[82][8]/P0001  & n13374 ;
  assign n27718 = ~n27716 & ~n27717 ;
  assign n27719 = \wishbone_bd_ram_mem1_reg[22][8]/P0001  & n13744 ;
  assign n27720 = \wishbone_bd_ram_mem1_reg[28][8]/P0001  & n13810 ;
  assign n27721 = ~n27719 & ~n27720 ;
  assign n27722 = n27718 & n27721 ;
  assign n27723 = n27715 & n27722 ;
  assign n27724 = \wishbone_bd_ram_mem1_reg[199][8]/P0001  & n13499 ;
  assign n27725 = \wishbone_bd_ram_mem1_reg[234][8]/P0001  & n13781 ;
  assign n27726 = ~n27724 & ~n27725 ;
  assign n27727 = \wishbone_bd_ram_mem1_reg[154][8]/P0001  & n13403 ;
  assign n27728 = \wishbone_bd_ram_mem1_reg[141][8]/P0001  & n13852 ;
  assign n27729 = ~n27727 & ~n27728 ;
  assign n27730 = n27726 & n27729 ;
  assign n27731 = \wishbone_bd_ram_mem1_reg[69][8]/P0001  & n13487 ;
  assign n27732 = \wishbone_bd_ram_mem1_reg[60][8]/P0001  & n13790 ;
  assign n27733 = ~n27731 & ~n27732 ;
  assign n27734 = \wishbone_bd_ram_mem1_reg[233][8]/P0001  & n13332 ;
  assign n27735 = \wishbone_bd_ram_mem1_reg[122][8]/P0001  & n13679 ;
  assign n27736 = ~n27734 & ~n27735 ;
  assign n27737 = n27733 & n27736 ;
  assign n27738 = n27730 & n27737 ;
  assign n27739 = n27723 & n27738 ;
  assign n27740 = n27708 & n27739 ;
  assign n27741 = \wishbone_bd_ram_mem1_reg[179][8]/P0001  & n14035 ;
  assign n27742 = \wishbone_bd_ram_mem1_reg[40][8]/P0001  & n13661 ;
  assign n27743 = ~n27741 & ~n27742 ;
  assign n27744 = \wishbone_bd_ram_mem1_reg[244][8]/P0001  & n13474 ;
  assign n27745 = \wishbone_bd_ram_mem1_reg[63][8]/P0001  & n13327 ;
  assign n27746 = ~n27744 & ~n27745 ;
  assign n27747 = n27743 & n27746 ;
  assign n27748 = \wishbone_bd_ram_mem1_reg[192][8]/P0001  & n13390 ;
  assign n27749 = \wishbone_bd_ram_mem1_reg[94][8]/P0001  & n13833 ;
  assign n27750 = ~n27748 & ~n27749 ;
  assign n27751 = \wishbone_bd_ram_mem1_reg[248][8]/P0001  & n13647 ;
  assign n27752 = \wishbone_bd_ram_mem1_reg[175][8]/P0001  & n13674 ;
  assign n27753 = ~n27751 & ~n27752 ;
  assign n27754 = n27750 & n27753 ;
  assign n27755 = n27747 & n27754 ;
  assign n27756 = \wishbone_bd_ram_mem1_reg[0][8]/P0001  & n13539 ;
  assign n27757 = \wishbone_bd_ram_mem1_reg[23][8]/P0001  & n13857 ;
  assign n27758 = ~n27756 & ~n27757 ;
  assign n27759 = \wishbone_bd_ram_mem1_reg[37][8]/P0001  & n13710 ;
  assign n27760 = \wishbone_bd_ram_mem1_reg[112][8]/P0001  & n13482 ;
  assign n27761 = ~n27759 & ~n27760 ;
  assign n27762 = n27758 & n27761 ;
  assign n27763 = \wishbone_bd_ram_mem1_reg[194][8]/P0001  & n13624 ;
  assign n27764 = \wishbone_bd_ram_mem1_reg[153][8]/P0001  & n13309 ;
  assign n27765 = ~n27763 & ~n27764 ;
  assign n27766 = \wishbone_bd_ram_mem1_reg[206][8]/P0001  & n13414 ;
  assign n27767 = \wishbone_bd_ram_mem1_reg[17][8]/P0001  & n13324 ;
  assign n27768 = ~n27766 & ~n27767 ;
  assign n27769 = n27765 & n27768 ;
  assign n27770 = n27762 & n27769 ;
  assign n27771 = n27755 & n27770 ;
  assign n27772 = \wishbone_bd_ram_mem1_reg[182][8]/P0001  & n13598 ;
  assign n27773 = \wishbone_bd_ram_mem1_reg[136][8]/P0001  & n13963 ;
  assign n27774 = ~n27772 & ~n27773 ;
  assign n27775 = \wishbone_bd_ram_mem1_reg[195][8]/P0001  & n13700 ;
  assign n27776 = \wishbone_bd_ram_mem1_reg[108][8]/P0001  & n13814 ;
  assign n27777 = ~n27775 & ~n27776 ;
  assign n27778 = n27774 & n27777 ;
  assign n27779 = \wishbone_bd_ram_mem1_reg[12][8]/P0001  & n13733 ;
  assign n27780 = \wishbone_bd_ram_mem1_reg[62][8]/P0001  & n13529 ;
  assign n27781 = ~n27779 & ~n27780 ;
  assign n27782 = \wishbone_bd_ram_mem1_reg[155][8]/P0001  & n13738 ;
  assign n27783 = \wishbone_bd_ram_mem1_reg[247][8]/P0001  & n13571 ;
  assign n27784 = ~n27782 & ~n27783 ;
  assign n27785 = n27781 & n27784 ;
  assign n27786 = n27778 & n27785 ;
  assign n27787 = \wishbone_bd_ram_mem1_reg[76][8]/P0001  & n13831 ;
  assign n27788 = \wishbone_bd_ram_mem1_reg[87][8]/P0001  & n13691 ;
  assign n27789 = ~n27787 & ~n27788 ;
  assign n27790 = \wishbone_bd_ram_mem1_reg[132][8]/P0001  & n13927 ;
  assign n27791 = \wishbone_bd_ram_mem1_reg[196][8]/P0001  & n13977 ;
  assign n27792 = ~n27790 & ~n27791 ;
  assign n27793 = n27789 & n27792 ;
  assign n27794 = \wishbone_bd_ram_mem1_reg[134][8]/P0001  & n13494 ;
  assign n27795 = \wishbone_bd_ram_mem1_reg[176][8]/P0001  & n13262 ;
  assign n27796 = ~n27794 & ~n27795 ;
  assign n27797 = \wishbone_bd_ram_mem1_reg[24][8]/P0001  & n13970 ;
  assign n27798 = \wishbone_bd_ram_mem1_reg[220][8]/P0001  & n13965 ;
  assign n27799 = ~n27797 & ~n27798 ;
  assign n27800 = n27796 & n27799 ;
  assign n27801 = n27793 & n27800 ;
  assign n27802 = n27786 & n27801 ;
  assign n27803 = n27771 & n27802 ;
  assign n27804 = n27740 & n27803 ;
  assign n27805 = n27677 & n27804 ;
  assign n27806 = n27550 & n27805 ;
  assign n27807 = ~wb_rst_i_pad & ~n27294 ;
  assign n27808 = ~n27806 & n27807 ;
  assign n27809 = ~n27295 & ~n27808 ;
  assign n27810 = \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  & n23751 ;
  assign n27811 = n23747 & n27810 ;
  assign n27812 = \ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131  & n23782 ;
  assign n27813 = ~n27811 & ~n27812 ;
  assign n27814 = \ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131  & n23743 ;
  assign n27815 = n23741 & n27814 ;
  assign n27816 = \ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131  & n23743 ;
  assign n27817 = n23747 & n27816 ;
  assign n27818 = ~n27815 & ~n27817 ;
  assign n27819 = n27813 & n27818 ;
  assign n27820 = \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  & n23751 ;
  assign n27821 = n23741 & n27820 ;
  assign n27822 = \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131  & n23794 ;
  assign n27823 = n23741 & n27822 ;
  assign n27824 = ~n27821 & ~n27823 ;
  assign n27825 = n23730 & n27824 ;
  assign n27826 = n27819 & n27825 ;
  assign n27827 = \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131  & n23802 ;
  assign n27828 = \ethreg1_MODER_1_DataOut_reg[1]/NET0131  & n23808 ;
  assign n27829 = ~n27827 & ~n27828 ;
  assign n27830 = \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  & n23737 ;
  assign n27831 = \ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131  & n23813 ;
  assign n27832 = ~n27830 & ~n27831 ;
  assign n27833 = n27829 & n27832 ;
  assign n27834 = n27826 & n27833 ;
  assign n27835 = n23730 & ~n27834 ;
  assign n27836 = \wishbone_bd_ram_mem1_reg[39][9]/P0001  & n13893 ;
  assign n27837 = \wishbone_bd_ram_mem1_reg[109][9]/P0001  & n13306 ;
  assign n27838 = ~n27836 & ~n27837 ;
  assign n27839 = \wishbone_bd_ram_mem1_reg[82][9]/P0001  & n13374 ;
  assign n27840 = \wishbone_bd_ram_mem1_reg[32][9]/P0001  & n13736 ;
  assign n27841 = ~n27839 & ~n27840 ;
  assign n27842 = n27838 & n27841 ;
  assign n27843 = \wishbone_bd_ram_mem1_reg[48][9]/P0001  & n13917 ;
  assign n27844 = \wishbone_bd_ram_mem1_reg[241][9]/P0001  & n13854 ;
  assign n27845 = ~n27843 & ~n27844 ;
  assign n27846 = \wishbone_bd_ram_mem1_reg[57][9]/P0001  & n13731 ;
  assign n27847 = \wishbone_bd_ram_mem1_reg[209][9]/P0001  & n13689 ;
  assign n27848 = ~n27846 & ~n27847 ;
  assign n27849 = n27845 & n27848 ;
  assign n27850 = n27842 & n27849 ;
  assign n27851 = \wishbone_bd_ram_mem1_reg[178][9]/P0001  & n13301 ;
  assign n27852 = \wishbone_bd_ram_mem1_reg[244][9]/P0001  & n13474 ;
  assign n27853 = ~n27851 & ~n27852 ;
  assign n27854 = \wishbone_bd_ram_mem1_reg[160][9]/P0001  & n13271 ;
  assign n27855 = \wishbone_bd_ram_mem1_reg[133][9]/P0001  & n13492 ;
  assign n27856 = ~n27854 & ~n27855 ;
  assign n27857 = n27853 & n27856 ;
  assign n27858 = \wishbone_bd_ram_mem1_reg[7][9]/P0001  & n13546 ;
  assign n27859 = \wishbone_bd_ram_mem1_reg[238][9]/P0001  & n13819 ;
  assign n27860 = ~n27858 & ~n27859 ;
  assign n27861 = \wishbone_bd_ram_mem1_reg[36][9]/P0001  & n13639 ;
  assign n27862 = \wishbone_bd_ram_mem1_reg[251][9]/P0001  & n14019 ;
  assign n27863 = ~n27861 & ~n27862 ;
  assign n27864 = n27860 & n27863 ;
  assign n27865 = n27857 & n27864 ;
  assign n27866 = n27850 & n27865 ;
  assign n27867 = \wishbone_bd_ram_mem1_reg[107][9]/P0001  & n13476 ;
  assign n27868 = \wishbone_bd_ram_mem1_reg[174][9]/P0001  & n13899 ;
  assign n27869 = ~n27867 & ~n27868 ;
  assign n27870 = \wishbone_bd_ram_mem1_reg[1][9]/P0001  & n13888 ;
  assign n27871 = \wishbone_bd_ram_mem1_reg[142][9]/P0001  & n13448 ;
  assign n27872 = ~n27870 & ~n27871 ;
  assign n27873 = n27869 & n27872 ;
  assign n27874 = \wishbone_bd_ram_mem1_reg[194][9]/P0001  & n13624 ;
  assign n27875 = \wishbone_bd_ram_mem1_reg[224][9]/P0001  & n13433 ;
  assign n27876 = ~n27874 & ~n27875 ;
  assign n27877 = \wishbone_bd_ram_mem1_reg[185][9]/P0001  & n13372 ;
  assign n27878 = \wishbone_bd_ram_mem1_reg[27][9]/P0001  & n13251 ;
  assign n27879 = ~n27877 & ~n27878 ;
  assign n27880 = n27876 & n27879 ;
  assign n27881 = n27873 & n27880 ;
  assign n27882 = \wishbone_bd_ram_mem1_reg[95][9]/P0001  & n13317 ;
  assign n27883 = \wishbone_bd_ram_mem1_reg[249][9]/P0001  & n13431 ;
  assign n27884 = ~n27882 & ~n27883 ;
  assign n27885 = \wishbone_bd_ram_mem1_reg[201][9]/P0001  & n13600 ;
  assign n27886 = \wishbone_bd_ram_mem1_reg[40][9]/P0001  & n13661 ;
  assign n27887 = ~n27885 & ~n27886 ;
  assign n27888 = n27884 & n27887 ;
  assign n27889 = \wishbone_bd_ram_mem1_reg[52][9]/P0001  & n13988 ;
  assign n27890 = \wishbone_bd_ram_mem1_reg[126][9]/P0001  & n13786 ;
  assign n27891 = ~n27889 & ~n27890 ;
  assign n27892 = \wishbone_bd_ram_mem1_reg[171][9]/P0001  & n13422 ;
  assign n27893 = \wishbone_bd_ram_mem1_reg[250][9]/P0001  & n13677 ;
  assign n27894 = ~n27892 & ~n27893 ;
  assign n27895 = n27891 & n27894 ;
  assign n27896 = n27888 & n27895 ;
  assign n27897 = n27881 & n27896 ;
  assign n27898 = n27866 & n27897 ;
  assign n27899 = \wishbone_bd_ram_mem1_reg[223][9]/P0001  & n13335 ;
  assign n27900 = \wishbone_bd_ram_mem1_reg[87][9]/P0001  & n13691 ;
  assign n27901 = ~n27899 & ~n27900 ;
  assign n27902 = \wishbone_bd_ram_mem1_reg[97][9]/P0001  & n13724 ;
  assign n27903 = \wishbone_bd_ram_mem1_reg[4][9]/P0001  & n13527 ;
  assign n27904 = ~n27902 & ~n27903 ;
  assign n27905 = n27901 & n27904 ;
  assign n27906 = \wishbone_bd_ram_mem1_reg[197][9]/P0001  & n13594 ;
  assign n27907 = \wishbone_bd_ram_mem1_reg[64][9]/P0001  & n13904 ;
  assign n27908 = ~n27906 & ~n27907 ;
  assign n27909 = \wishbone_bd_ram_mem1_reg[206][9]/P0001  & n13414 ;
  assign n27910 = \wishbone_bd_ram_mem1_reg[102][9]/P0001  & n13534 ;
  assign n27911 = ~n27909 & ~n27910 ;
  assign n27912 = n27908 & n27911 ;
  assign n27913 = n27905 & n27912 ;
  assign n27914 = \wishbone_bd_ram_mem1_reg[189][9]/P0001  & n14001 ;
  assign n27915 = \wishbone_bd_ram_mem1_reg[181][9]/P0001  & n13587 ;
  assign n27916 = ~n27914 & ~n27915 ;
  assign n27917 = \wishbone_bd_ram_mem1_reg[129][9]/P0001  & n13629 ;
  assign n27918 = \wishbone_bd_ram_mem1_reg[235][9]/P0001  & n13518 ;
  assign n27919 = ~n27917 & ~n27918 ;
  assign n27920 = n27916 & n27919 ;
  assign n27921 = \wishbone_bd_ram_mem1_reg[202][9]/P0001  & n13268 ;
  assign n27922 = \wishbone_bd_ram_mem1_reg[217][9]/P0001  & n13767 ;
  assign n27923 = ~n27921 & ~n27922 ;
  assign n27924 = \wishbone_bd_ram_mem1_reg[157][9]/P0001  & n13445 ;
  assign n27925 = \wishbone_bd_ram_mem1_reg[215][9]/P0001  & n13901 ;
  assign n27926 = ~n27924 & ~n27925 ;
  assign n27927 = n27923 & n27926 ;
  assign n27928 = n27920 & n27927 ;
  assign n27929 = n27913 & n27928 ;
  assign n27930 = \wishbone_bd_ram_mem1_reg[134][9]/P0001  & n13494 ;
  assign n27931 = \wishbone_bd_ram_mem1_reg[170][9]/P0001  & n14007 ;
  assign n27932 = ~n27930 & ~n27931 ;
  assign n27933 = \wishbone_bd_ram_mem1_reg[45][9]/P0001  & n13420 ;
  assign n27934 = \wishbone_bd_ram_mem1_reg[120][9]/P0001  & n13550 ;
  assign n27935 = ~n27933 & ~n27934 ;
  assign n27936 = n27932 & n27935 ;
  assign n27937 = \wishbone_bd_ram_mem1_reg[42][9]/P0001  & n13341 ;
  assign n27938 = \wishbone_bd_ram_mem1_reg[208][9]/P0001  & n14010 ;
  assign n27939 = ~n27937 & ~n27938 ;
  assign n27940 = \wishbone_bd_ram_mem1_reg[85][9]/P0001  & n13784 ;
  assign n27941 = \wishbone_bd_ram_mem1_reg[17][9]/P0001  & n13324 ;
  assign n27942 = ~n27940 & ~n27941 ;
  assign n27943 = n27939 & n27942 ;
  assign n27944 = n27936 & n27943 ;
  assign n27945 = \wishbone_bd_ram_mem1_reg[132][9]/P0001  & n13927 ;
  assign n27946 = \wishbone_bd_ram_mem1_reg[86][9]/P0001  & n13485 ;
  assign n27947 = ~n27945 & ~n27946 ;
  assign n27948 = \wishbone_bd_ram_mem1_reg[117][9]/P0001  & n13557 ;
  assign n27949 = \wishbone_bd_ram_mem1_reg[56][9]/P0001  & n13611 ;
  assign n27950 = ~n27948 & ~n27949 ;
  assign n27951 = n27947 & n27950 ;
  assign n27952 = \wishbone_bd_ram_mem1_reg[10][9]/P0001  & n13837 ;
  assign n27953 = \wishbone_bd_ram_mem1_reg[83][9]/P0001  & n13454 ;
  assign n27954 = ~n27952 & ~n27953 ;
  assign n27955 = \wishbone_bd_ram_mem1_reg[21][9]/P0001  & n13438 ;
  assign n27956 = \wishbone_bd_ram_mem1_reg[156][9]/P0001  & n13769 ;
  assign n27957 = ~n27955 & ~n27956 ;
  assign n27958 = n27954 & n27957 ;
  assign n27959 = n27951 & n27958 ;
  assign n27960 = n27944 & n27959 ;
  assign n27961 = n27929 & n27960 ;
  assign n27962 = n27898 & n27961 ;
  assign n27963 = \wishbone_bd_ram_mem1_reg[73][9]/P0001  & n13456 ;
  assign n27964 = \wishbone_bd_ram_mem1_reg[186][9]/P0001  & n13616 ;
  assign n27965 = ~n27963 & ~n27964 ;
  assign n27966 = \wishbone_bd_ram_mem1_reg[236][9]/P0001  & n13480 ;
  assign n27967 = \wishbone_bd_ram_mem1_reg[130][9]/P0001  & n13427 ;
  assign n27968 = ~n27966 & ~n27967 ;
  assign n27969 = n27965 & n27968 ;
  assign n27970 = \wishbone_bd_ram_mem1_reg[68][9]/P0001  & n13379 ;
  assign n27971 = \wishbone_bd_ram_mem1_reg[195][9]/P0001  & n13700 ;
  assign n27972 = ~n27970 & ~n27971 ;
  assign n27973 = \wishbone_bd_ram_mem1_reg[166][9]/P0001  & n13999 ;
  assign n27974 = \wishbone_bd_ram_mem1_reg[106][9]/P0001  & n13555 ;
  assign n27975 = ~n27973 & ~n27974 ;
  assign n27976 = n27972 & n27975 ;
  assign n27977 = n27969 & n27976 ;
  assign n27978 = \wishbone_bd_ram_mem1_reg[139][9]/P0001  & n13566 ;
  assign n27979 = \wishbone_bd_ram_mem1_reg[123][9]/P0001  & n13749 ;
  assign n27980 = ~n27978 & ~n27979 ;
  assign n27981 = \wishbone_bd_ram_mem1_reg[196][9]/P0001  & n13977 ;
  assign n27982 = \wishbone_bd_ram_mem1_reg[204][9]/P0001  & n13821 ;
  assign n27983 = ~n27981 & ~n27982 ;
  assign n27984 = n27980 & n27983 ;
  assign n27985 = \wishbone_bd_ram_mem1_reg[193][9]/P0001  & n14022 ;
  assign n27986 = \wishbone_bd_ram_mem1_reg[149][9]/P0001  & n13469 ;
  assign n27987 = ~n27985 & ~n27986 ;
  assign n27988 = \wishbone_bd_ram_mem1_reg[151][9]/P0001  & n13697 ;
  assign n27989 = \wishbone_bd_ram_mem1_reg[154][9]/P0001  & n13403 ;
  assign n27990 = ~n27988 & ~n27989 ;
  assign n27991 = n27987 & n27990 ;
  assign n27992 = n27984 & n27991 ;
  assign n27993 = n27977 & n27992 ;
  assign n27994 = \wishbone_bd_ram_mem1_reg[84][9]/P0001  & n13385 ;
  assign n27995 = \wishbone_bd_ram_mem1_reg[173][9]/P0001  & n13360 ;
  assign n27996 = ~n27994 & ~n27995 ;
  assign n27997 = \wishbone_bd_ram_mem1_reg[119][9]/P0001  & n14033 ;
  assign n27998 = \wishbone_bd_ram_mem1_reg[25][9]/P0001  & n13742 ;
  assign n27999 = ~n27997 & ~n27998 ;
  assign n28000 = n27996 & n27999 ;
  assign n28001 = \wishbone_bd_ram_mem1_reg[9][9]/P0001  & n13580 ;
  assign n28002 = \wishbone_bd_ram_mem1_reg[20][9]/P0001  & n13839 ;
  assign n28003 = ~n28001 & ~n28002 ;
  assign n28004 = \wishbone_bd_ram_mem1_reg[30][9]/P0001  & n13713 ;
  assign n28005 = \wishbone_bd_ram_mem1_reg[144][9]/P0001  & n13508 ;
  assign n28006 = ~n28004 & ~n28005 ;
  assign n28007 = n28003 & n28006 ;
  assign n28008 = n28000 & n28007 ;
  assign n28009 = \wishbone_bd_ram_mem1_reg[13][9]/P0001  & n13844 ;
  assign n28010 = \wishbone_bd_ram_mem1_reg[111][9]/P0001  & n13471 ;
  assign n28011 = ~n28009 & ~n28010 ;
  assign n28012 = \wishbone_bd_ram_mem1_reg[118][9]/P0001  & n13589 ;
  assign n28013 = \wishbone_bd_ram_mem1_reg[22][9]/P0001  & n13744 ;
  assign n28014 = ~n28012 & ~n28013 ;
  assign n28015 = n28011 & n28014 ;
  assign n28016 = \wishbone_bd_ram_mem1_reg[231][9]/P0001  & n13363 ;
  assign n28017 = \wishbone_bd_ram_mem1_reg[254][9]/P0001  & n13283 ;
  assign n28018 = ~n28016 & ~n28017 ;
  assign n28019 = \wishbone_bd_ram_mem1_reg[205][9]/P0001  & n13947 ;
  assign n28020 = \wishbone_bd_ram_mem1_reg[138][9]/P0001  & n13398 ;
  assign n28021 = ~n28019 & ~n28020 ;
  assign n28022 = n28018 & n28021 ;
  assign n28023 = n28015 & n28022 ;
  assign n28024 = n28008 & n28023 ;
  assign n28025 = n27993 & n28024 ;
  assign n28026 = \wishbone_bd_ram_mem1_reg[165][9]/P0001  & n14028 ;
  assign n28027 = \wishbone_bd_ram_mem1_reg[237][9]/P0001  & n13924 ;
  assign n28028 = ~n28026 & ~n28027 ;
  assign n28029 = \wishbone_bd_ram_mem1_reg[146][9]/P0001  & n13958 ;
  assign n28030 = \wishbone_bd_ram_mem1_reg[127][9]/P0001  & n13803 ;
  assign n28031 = ~n28029 & ~n28030 ;
  assign n28032 = n28028 & n28031 ;
  assign n28033 = \wishbone_bd_ram_mem1_reg[220][9]/P0001  & n13965 ;
  assign n28034 = \wishbone_bd_ram_mem1_reg[246][9]/P0001  & n13981 ;
  assign n28035 = ~n28033 & ~n28034 ;
  assign n28036 = \wishbone_bd_ram_mem1_reg[2][9]/P0001  & n13975 ;
  assign n28037 = \wishbone_bd_ram_mem1_reg[77][9]/P0001  & n13935 ;
  assign n28038 = ~n28036 & ~n28037 ;
  assign n28039 = n28035 & n28038 ;
  assign n28040 = n28032 & n28039 ;
  assign n28041 = \wishbone_bd_ram_mem1_reg[213][9]/P0001  & n13870 ;
  assign n28042 = \wishbone_bd_ram_mem1_reg[34][9]/P0001  & n13450 ;
  assign n28043 = ~n28041 & ~n28042 ;
  assign n28044 = \wishbone_bd_ram_mem1_reg[184][9]/P0001  & n13960 ;
  assign n28045 = \wishbone_bd_ram_mem1_reg[54][9]/P0001  & n13622 ;
  assign n28046 = ~n28044 & ~n28045 ;
  assign n28047 = n28043 & n28046 ;
  assign n28048 = \wishbone_bd_ram_mem1_reg[180][9]/P0001  & n13650 ;
  assign n28049 = \wishbone_bd_ram_mem1_reg[252][9]/P0001  & n13986 ;
  assign n28050 = ~n28048 & ~n28049 ;
  assign n28051 = \wishbone_bd_ram_mem1_reg[167][9]/P0001  & n13940 ;
  assign n28052 = \wishbone_bd_ram_mem1_reg[92][9]/P0001  & n13859 ;
  assign n28053 = ~n28051 & ~n28052 ;
  assign n28054 = n28050 & n28053 ;
  assign n28055 = n28047 & n28054 ;
  assign n28056 = n28040 & n28055 ;
  assign n28057 = \wishbone_bd_ram_mem1_reg[61][9]/P0001  & n13544 ;
  assign n28058 = \wishbone_bd_ram_mem1_reg[99][9]/P0001  & n13996 ;
  assign n28059 = ~n28057 & ~n28058 ;
  assign n28060 = \wishbone_bd_ram_mem1_reg[228][9]/P0001  & n13497 ;
  assign n28061 = \wishbone_bd_ram_mem1_reg[115][9]/P0001  & n13747 ;
  assign n28062 = ~n28060 & ~n28061 ;
  assign n28063 = n28059 & n28062 ;
  assign n28064 = \wishbone_bd_ram_mem1_reg[168][9]/P0001  & n13795 ;
  assign n28065 = \wishbone_bd_ram_mem1_reg[227][9]/P0001  & n13388 ;
  assign n28066 = ~n28064 & ~n28065 ;
  assign n28067 = \wishbone_bd_ram_mem1_reg[55][9]/P0001  & n13618 ;
  assign n28068 = \wishbone_bd_ram_mem1_reg[116][9]/P0001  & n13865 ;
  assign n28069 = ~n28067 & ~n28068 ;
  assign n28070 = n28066 & n28069 ;
  assign n28071 = n28063 & n28070 ;
  assign n28072 = \wishbone_bd_ram_mem1_reg[49][9]/P0001  & n13929 ;
  assign n28073 = \wishbone_bd_ram_mem1_reg[100][9]/P0001  & n13401 ;
  assign n28074 = ~n28072 & ~n28073 ;
  assign n28075 = \wishbone_bd_ram_mem1_reg[80][9]/P0001  & n13516 ;
  assign n28076 = \wishbone_bd_ram_mem1_reg[90][9]/P0001  & n13906 ;
  assign n28077 = ~n28075 & ~n28076 ;
  assign n28078 = n28074 & n28077 ;
  assign n28079 = \wishbone_bd_ram_mem1_reg[255][9]/P0001  & n13952 ;
  assign n28080 = \wishbone_bd_ram_mem1_reg[207][9]/P0001  & n13826 ;
  assign n28081 = ~n28079 & ~n28080 ;
  assign n28082 = \wishbone_bd_ram_mem1_reg[121][9]/P0001  & n13983 ;
  assign n28083 = \wishbone_bd_ram_mem1_reg[29][9]/P0001  & n13412 ;
  assign n28084 = ~n28082 & ~n28083 ;
  assign n28085 = n28081 & n28084 ;
  assign n28086 = n28078 & n28085 ;
  assign n28087 = n28071 & n28086 ;
  assign n28088 = n28056 & n28087 ;
  assign n28089 = n28025 & n28088 ;
  assign n28090 = n27962 & n28089 ;
  assign n28091 = \wishbone_bd_ram_mem1_reg[0][9]/P0001  & n13539 ;
  assign n28092 = \wishbone_bd_ram_mem1_reg[164][9]/P0001  & n13236 ;
  assign n28093 = ~n28091 & ~n28092 ;
  assign n28094 = \wishbone_bd_ram_mem1_reg[65][9]/P0001  & n13842 ;
  assign n28095 = \wishbone_bd_ram_mem1_reg[47][9]/P0001  & n13436 ;
  assign n28096 = ~n28094 & ~n28095 ;
  assign n28097 = n28093 & n28096 ;
  assign n28098 = \wishbone_bd_ram_mem1_reg[148][9]/P0001  & n13868 ;
  assign n28099 = \wishbone_bd_ram_mem1_reg[58][9]/P0001  & n13949 ;
  assign n28100 = ~n28098 & ~n28099 ;
  assign n28101 = \wishbone_bd_ram_mem1_reg[245][9]/P0001  & n13877 ;
  assign n28102 = \wishbone_bd_ram_mem1_reg[137][9]/P0001  & n13808 ;
  assign n28103 = ~n28101 & ~n28102 ;
  assign n28104 = n28100 & n28103 ;
  assign n28105 = n28097 & n28104 ;
  assign n28106 = \wishbone_bd_ram_mem1_reg[182][9]/P0001  & n13598 ;
  assign n28107 = \wishbone_bd_ram_mem1_reg[67][9]/P0001  & n13663 ;
  assign n28108 = ~n28106 & ~n28107 ;
  assign n28109 = \wishbone_bd_ram_mem1_reg[24][9]/P0001  & n13970 ;
  assign n28110 = \wishbone_bd_ram_mem1_reg[71][9]/P0001  & n13636 ;
  assign n28111 = ~n28109 & ~n28110 ;
  assign n28112 = n28108 & n28111 ;
  assign n28113 = \wishbone_bd_ram_mem1_reg[113][9]/P0001  & n13882 ;
  assign n28114 = \wishbone_bd_ram_mem1_reg[192][9]/P0001  & n13390 ;
  assign n28115 = ~n28113 & ~n28114 ;
  assign n28116 = \wishbone_bd_ram_mem1_reg[222][9]/P0001  & n13721 ;
  assign n28117 = \wishbone_bd_ram_mem1_reg[75][9]/P0001  & n13605 ;
  assign n28118 = ~n28116 & ~n28117 ;
  assign n28119 = n28115 & n28118 ;
  assign n28120 = n28112 & n28119 ;
  assign n28121 = n28105 & n28120 ;
  assign n28122 = \wishbone_bd_ram_mem1_reg[221][9]/P0001  & n13641 ;
  assign n28123 = \wishbone_bd_ram_mem1_reg[72][9]/P0001  & n13582 ;
  assign n28124 = ~n28122 & ~n28123 ;
  assign n28125 = \wishbone_bd_ram_mem1_reg[37][9]/P0001  & n13710 ;
  assign n28126 = \wishbone_bd_ram_mem1_reg[161][9]/P0001  & n13505 ;
  assign n28127 = ~n28125 & ~n28126 ;
  assign n28128 = n28124 & n28127 ;
  assign n28129 = \wishbone_bd_ram_mem1_reg[190][9]/P0001  & n13365 ;
  assign n28130 = \wishbone_bd_ram_mem1_reg[253][9]/P0001  & n13708 ;
  assign n28131 = ~n28129 & ~n28130 ;
  assign n28132 = \wishbone_bd_ram_mem1_reg[158][9]/P0001  & n13294 ;
  assign n28133 = \wishbone_bd_ram_mem1_reg[38][9]/P0001  & n13828 ;
  assign n28134 = ~n28132 & ~n28133 ;
  assign n28135 = n28131 & n28134 ;
  assign n28136 = n28128 & n28135 ;
  assign n28137 = \wishbone_bd_ram_mem1_reg[135][9]/P0001  & n13672 ;
  assign n28138 = \wishbone_bd_ram_mem1_reg[5][9]/P0001  & n13243 ;
  assign n28139 = ~n28137 & ~n28138 ;
  assign n28140 = \wishbone_bd_ram_mem1_reg[28][9]/P0001  & n13810 ;
  assign n28141 = \wishbone_bd_ram_mem1_reg[159][9]/P0001  & n13627 ;
  assign n28142 = ~n28140 & ~n28141 ;
  assign n28143 = n28139 & n28142 ;
  assign n28144 = \wishbone_bd_ram_mem1_reg[6][9]/P0001  & n13915 ;
  assign n28145 = \wishbone_bd_ram_mem1_reg[51][9]/P0001  & n13880 ;
  assign n28146 = ~n28144 & ~n28145 ;
  assign n28147 = \wishbone_bd_ram_mem1_reg[147][9]/P0001  & n13702 ;
  assign n28148 = \wishbone_bd_ram_mem1_reg[230][9]/P0001  & n13994 ;
  assign n28149 = ~n28147 & ~n28148 ;
  assign n28150 = n28146 & n28149 ;
  assign n28151 = n28143 & n28150 ;
  assign n28152 = n28136 & n28151 ;
  assign n28153 = n28121 & n28152 ;
  assign n28154 = \wishbone_bd_ram_mem1_reg[239][9]/P0001  & n13349 ;
  assign n28155 = \wishbone_bd_ram_mem1_reg[19][9]/P0001  & n13886 ;
  assign n28156 = ~n28154 & ~n28155 ;
  assign n28157 = \wishbone_bd_ram_mem1_reg[44][9]/P0001  & n13291 ;
  assign n28158 = \wishbone_bd_ram_mem1_reg[191][9]/P0001  & n14012 ;
  assign n28159 = ~n28157 & ~n28158 ;
  assign n28160 = n28156 & n28159 ;
  assign n28161 = \wishbone_bd_ram_mem1_reg[31][9]/P0001  & n13758 ;
  assign n28162 = \wishbone_bd_ram_mem1_reg[89][9]/P0001  & n13910 ;
  assign n28163 = ~n28161 & ~n28162 ;
  assign n28164 = \wishbone_bd_ram_mem1_reg[136][9]/P0001  & n13963 ;
  assign n28165 = \wishbone_bd_ram_mem1_reg[23][9]/P0001  & n13857 ;
  assign n28166 = ~n28164 & ~n28165 ;
  assign n28167 = n28163 & n28166 ;
  assign n28168 = n28160 & n28167 ;
  assign n28169 = \wishbone_bd_ram_mem1_reg[3][9]/P0001  & n13354 ;
  assign n28170 = \wishbone_bd_ram_mem1_reg[216][9]/P0001  & n14005 ;
  assign n28171 = ~n28169 & ~n28170 ;
  assign n28172 = \wishbone_bd_ram_mem1_reg[104][9]/P0001  & n13684 ;
  assign n28173 = \wishbone_bd_ram_mem1_reg[183][9]/P0001  & n13645 ;
  assign n28174 = ~n28172 & ~n28173 ;
  assign n28175 = n28171 & n28174 ;
  assign n28176 = \wishbone_bd_ram_mem1_reg[128][9]/P0001  & n13652 ;
  assign n28177 = \wishbone_bd_ram_mem1_reg[93][9]/P0001  & n13891 ;
  assign n28178 = ~n28176 & ~n28177 ;
  assign n28179 = \wishbone_bd_ram_mem1_reg[105][9]/P0001  & n13503 ;
  assign n28180 = \wishbone_bd_ram_mem1_reg[243][9]/P0001  & n13575 ;
  assign n28181 = ~n28179 & ~n28180 ;
  assign n28182 = n28178 & n28181 ;
  assign n28183 = n28175 & n28182 ;
  assign n28184 = n28168 & n28183 ;
  assign n28185 = \wishbone_bd_ram_mem1_reg[200][9]/P0001  & n13922 ;
  assign n28186 = \wishbone_bd_ram_mem1_reg[179][9]/P0001  & n14035 ;
  assign n28187 = ~n28185 & ~n28186 ;
  assign n28188 = \wishbone_bd_ram_mem1_reg[59][9]/P0001  & n13613 ;
  assign n28189 = \wishbone_bd_ram_mem1_reg[11][9]/P0001  & n13774 ;
  assign n28190 = ~n28188 & ~n28189 ;
  assign n28191 = n28187 & n28190 ;
  assign n28192 = \wishbone_bd_ram_mem1_reg[177][9]/P0001  & n13863 ;
  assign n28193 = \wishbone_bd_ram_mem1_reg[247][9]/P0001  & n13571 ;
  assign n28194 = ~n28192 & ~n28193 ;
  assign n28195 = \wishbone_bd_ram_mem1_reg[229][9]/P0001  & n13552 ;
  assign n28196 = \wishbone_bd_ram_mem1_reg[175][9]/P0001  & n13674 ;
  assign n28197 = ~n28195 & ~n28196 ;
  assign n28198 = n28194 & n28197 ;
  assign n28199 = n28191 & n28198 ;
  assign n28200 = \wishbone_bd_ram_mem1_reg[225][9]/P0001  & n13719 ;
  assign n28201 = \wishbone_bd_ram_mem1_reg[62][9]/P0001  & n13529 ;
  assign n28202 = ~n28200 & ~n28201 ;
  assign n28203 = \wishbone_bd_ram_mem1_reg[219][9]/P0001  & n13577 ;
  assign n28204 = \wishbone_bd_ram_mem1_reg[172][9]/P0001  & n13377 ;
  assign n28205 = ~n28203 & ~n28204 ;
  assign n28206 = n28202 & n28205 ;
  assign n28207 = \wishbone_bd_ram_mem1_reg[46][9]/P0001  & n13298 ;
  assign n28208 = \wishbone_bd_ram_mem1_reg[232][9]/P0001  & n13510 ;
  assign n28209 = ~n28207 & ~n28208 ;
  assign n28210 = \wishbone_bd_ram_mem1_reg[79][9]/P0001  & n13779 ;
  assign n28211 = \wishbone_bd_ram_mem1_reg[50][9]/P0001  & n13686 ;
  assign n28212 = ~n28210 & ~n28211 ;
  assign n28213 = n28209 & n28212 ;
  assign n28214 = n28206 & n28213 ;
  assign n28215 = n28199 & n28214 ;
  assign n28216 = n28184 & n28215 ;
  assign n28217 = n28153 & n28216 ;
  assign n28218 = \wishbone_bd_ram_mem1_reg[26][9]/P0001  & n13521 ;
  assign n28219 = \wishbone_bd_ram_mem1_reg[124][9]/P0001  & n14024 ;
  assign n28220 = ~n28218 & ~n28219 ;
  assign n28221 = \wishbone_bd_ram_mem1_reg[33][9]/P0001  & n13933 ;
  assign n28222 = \wishbone_bd_ram_mem1_reg[112][9]/P0001  & n13482 ;
  assign n28223 = ~n28221 & ~n28222 ;
  assign n28224 = n28220 & n28223 ;
  assign n28225 = \wishbone_bd_ram_mem1_reg[145][9]/P0001  & n13715 ;
  assign n28226 = \wishbone_bd_ram_mem1_reg[218][9]/P0001  & n13792 ;
  assign n28227 = ~n28225 & ~n28226 ;
  assign n28228 = \wishbone_bd_ram_mem1_reg[78][9]/P0001  & n13277 ;
  assign n28229 = \wishbone_bd_ram_mem1_reg[53][9]/P0001  & n13875 ;
  assign n28230 = ~n28228 & ~n28229 ;
  assign n28231 = n28227 & n28230 ;
  assign n28232 = n28224 & n28231 ;
  assign n28233 = \wishbone_bd_ram_mem1_reg[155][9]/P0001  & n13738 ;
  assign n28234 = \wishbone_bd_ram_mem1_reg[163][9]/P0001  & n13255 ;
  assign n28235 = ~n28233 & ~n28234 ;
  assign n28236 = \wishbone_bd_ram_mem1_reg[74][9]/P0001  & n13564 ;
  assign n28237 = \wishbone_bd_ram_mem1_reg[212][9]/P0001  & n13634 ;
  assign n28238 = ~n28236 & ~n28237 ;
  assign n28239 = n28235 & n28238 ;
  assign n28240 = \wishbone_bd_ram_mem1_reg[15][9]/P0001  & n13797 ;
  assign n28241 = \wishbone_bd_ram_mem1_reg[8][9]/P0001  & n13459 ;
  assign n28242 = ~n28240 & ~n28241 ;
  assign n28243 = \wishbone_bd_ram_mem1_reg[169][9]/P0001  & n13541 ;
  assign n28244 = \wishbone_bd_ram_mem1_reg[141][9]/P0001  & n13852 ;
  assign n28245 = ~n28243 & ~n28244 ;
  assign n28246 = n28242 & n28245 ;
  assign n28247 = n28239 & n28246 ;
  assign n28248 = n28232 & n28247 ;
  assign n28249 = \wishbone_bd_ram_mem1_reg[43][9]/P0001  & n13761 ;
  assign n28250 = \wishbone_bd_ram_mem1_reg[70][9]/P0001  & n13339 ;
  assign n28251 = ~n28249 & ~n28250 ;
  assign n28252 = \wishbone_bd_ram_mem1_reg[60][9]/P0001  & n13790 ;
  assign n28253 = \wishbone_bd_ram_mem1_reg[88][9]/P0001  & n13347 ;
  assign n28254 = ~n28252 & ~n28253 ;
  assign n28255 = n28251 & n28254 ;
  assign n28256 = \wishbone_bd_ram_mem1_reg[96][9]/P0001  & n13425 ;
  assign n28257 = \wishbone_bd_ram_mem1_reg[81][9]/P0001  & n13409 ;
  assign n28258 = ~n28256 & ~n28257 ;
  assign n28259 = \wishbone_bd_ram_mem1_reg[14][9]/P0001  & n13972 ;
  assign n28260 = \wishbone_bd_ram_mem1_reg[66][9]/P0001  & n13603 ;
  assign n28261 = ~n28259 & ~n28260 ;
  assign n28262 = n28258 & n28261 ;
  assign n28263 = n28255 & n28262 ;
  assign n28264 = \wishbone_bd_ram_mem1_reg[203][9]/P0001  & n13816 ;
  assign n28265 = \wishbone_bd_ram_mem1_reg[234][9]/P0001  & n13781 ;
  assign n28266 = ~n28264 & ~n28265 ;
  assign n28267 = \wishbone_bd_ram_mem1_reg[198][9]/P0001  & n13592 ;
  assign n28268 = \wishbone_bd_ram_mem1_reg[131][9]/P0001  & n13358 ;
  assign n28269 = ~n28267 & ~n28268 ;
  assign n28270 = n28266 & n28269 ;
  assign n28271 = \wishbone_bd_ram_mem1_reg[69][9]/P0001  & n13487 ;
  assign n28272 = \wishbone_bd_ram_mem1_reg[108][9]/P0001  & n13814 ;
  assign n28273 = ~n28271 & ~n28272 ;
  assign n28274 = \wishbone_bd_ram_mem1_reg[248][9]/P0001  & n13647 ;
  assign n28275 = \wishbone_bd_ram_mem1_reg[101][9]/P0001  & n13772 ;
  assign n28276 = ~n28274 & ~n28275 ;
  assign n28277 = n28273 & n28276 ;
  assign n28278 = n28270 & n28277 ;
  assign n28279 = n28263 & n28278 ;
  assign n28280 = n28248 & n28279 ;
  assign n28281 = \wishbone_bd_ram_mem1_reg[211][9]/P0001  & n13805 ;
  assign n28282 = \wishbone_bd_ram_mem1_reg[187][9]/P0001  & n13756 ;
  assign n28283 = ~n28281 & ~n28282 ;
  assign n28284 = \wishbone_bd_ram_mem1_reg[140][9]/P0001  & n13287 ;
  assign n28285 = \wishbone_bd_ram_mem1_reg[162][9]/P0001  & n13726 ;
  assign n28286 = ~n28284 & ~n28285 ;
  assign n28287 = n28283 & n28286 ;
  assign n28288 = \wishbone_bd_ram_mem1_reg[125][9]/P0001  & n13396 ;
  assign n28289 = \wishbone_bd_ram_mem1_reg[91][9]/P0001  & n13954 ;
  assign n28290 = ~n28288 & ~n28289 ;
  assign n28291 = \wishbone_bd_ram_mem1_reg[152][9]/P0001  & n13912 ;
  assign n28292 = \wishbone_bd_ram_mem1_reg[94][9]/P0001  & n13833 ;
  assign n28293 = ~n28291 & ~n28292 ;
  assign n28294 = n28290 & n28293 ;
  assign n28295 = n28287 & n28294 ;
  assign n28296 = \wishbone_bd_ram_mem1_reg[12][9]/P0001  & n13733 ;
  assign n28297 = \wishbone_bd_ram_mem1_reg[35][9]/P0001  & n13523 ;
  assign n28298 = ~n28296 & ~n28297 ;
  assign n28299 = \wishbone_bd_ram_mem1_reg[16][9]/P0001  & n13695 ;
  assign n28300 = \wishbone_bd_ram_mem1_reg[103][9]/P0001  & n13320 ;
  assign n28301 = ~n28299 & ~n28300 ;
  assign n28302 = n28298 & n28301 ;
  assign n28303 = \wishbone_bd_ram_mem1_reg[233][9]/P0001  & n13332 ;
  assign n28304 = \wishbone_bd_ram_mem1_reg[143][9]/P0001  & n13461 ;
  assign n28305 = ~n28303 & ~n28304 ;
  assign n28306 = \wishbone_bd_ram_mem1_reg[226][9]/P0001  & n13668 ;
  assign n28307 = \wishbone_bd_ram_mem1_reg[18][9]/P0001  & n13532 ;
  assign n28308 = ~n28306 & ~n28307 ;
  assign n28309 = n28305 & n28308 ;
  assign n28310 = n28302 & n28309 ;
  assign n28311 = n28295 & n28310 ;
  assign n28312 = \wishbone_bd_ram_mem1_reg[153][9]/P0001  & n13309 ;
  assign n28313 = \wishbone_bd_ram_mem1_reg[122][9]/P0001  & n13679 ;
  assign n28314 = ~n28312 & ~n28313 ;
  assign n28315 = \wishbone_bd_ram_mem1_reg[98][9]/P0001  & n13569 ;
  assign n28316 = \wishbone_bd_ram_mem1_reg[110][9]/P0001  & n14030 ;
  assign n28317 = ~n28315 & ~n28316 ;
  assign n28318 = n28314 & n28317 ;
  assign n28319 = \wishbone_bd_ram_mem1_reg[240][9]/P0001  & n13352 ;
  assign n28320 = \wishbone_bd_ram_mem1_reg[114][9]/P0001  & n13763 ;
  assign n28321 = ~n28319 & ~n28320 ;
  assign n28322 = \wishbone_bd_ram_mem1_reg[150][9]/P0001  & n13666 ;
  assign n28323 = \wishbone_bd_ram_mem1_reg[242][9]/P0001  & n13383 ;
  assign n28324 = ~n28322 & ~n28323 ;
  assign n28325 = n28321 & n28324 ;
  assign n28326 = n28318 & n28325 ;
  assign n28327 = \wishbone_bd_ram_mem1_reg[76][9]/P0001  & n13831 ;
  assign n28328 = \wishbone_bd_ram_mem1_reg[214][9]/P0001  & n13938 ;
  assign n28329 = ~n28327 & ~n28328 ;
  assign n28330 = \wishbone_bd_ram_mem1_reg[210][9]/P0001  & n13443 ;
  assign n28331 = \wishbone_bd_ram_mem1_reg[188][9]/P0001  & n13407 ;
  assign n28332 = ~n28330 & ~n28331 ;
  assign n28333 = n28329 & n28332 ;
  assign n28334 = \wishbone_bd_ram_mem1_reg[63][9]/P0001  & n13327 ;
  assign n28335 = \wishbone_bd_ram_mem1_reg[176][9]/P0001  & n13262 ;
  assign n28336 = ~n28334 & ~n28335 ;
  assign n28337 = \wishbone_bd_ram_mem1_reg[41][9]/P0001  & n14017 ;
  assign n28338 = \wishbone_bd_ram_mem1_reg[199][9]/P0001  & n13499 ;
  assign n28339 = ~n28337 & ~n28338 ;
  assign n28340 = n28336 & n28339 ;
  assign n28341 = n28333 & n28340 ;
  assign n28342 = n28326 & n28341 ;
  assign n28343 = n28311 & n28342 ;
  assign n28344 = n28280 & n28343 ;
  assign n28345 = n28217 & n28344 ;
  assign n28346 = n28090 & n28345 ;
  assign n28347 = ~wb_rst_i_pad & ~n27834 ;
  assign n28348 = ~n28346 & n28347 ;
  assign n28349 = ~n27835 & ~n28348 ;
  assign n28350 = \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  & n23737 ;
  assign n28351 = \ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131  & n23743 ;
  assign n28352 = n23741 & n28351 ;
  assign n28353 = \ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131  & n23743 ;
  assign n28354 = n23747 & n28353 ;
  assign n28355 = ~n28352 & ~n28354 ;
  assign n28356 = \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  & n23751 ;
  assign n28357 = n23741 & n28356 ;
  assign n28358 = n23730 & ~n28357 ;
  assign n28359 = n28355 & n28358 ;
  assign n28360 = ~n28350 & n28359 ;
  assign n28361 = n23730 & ~n28360 ;
  assign n28362 = ~wb_rst_i_pad & ~n28360 ;
  assign n28363 = ~n17358 & n28362 ;
  assign n28364 = ~n28361 & ~n28363 ;
  assign n28365 = \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  & n23751 ;
  assign n28366 = n23747 & n28365 ;
  assign n28367 = \ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131  & n23782 ;
  assign n28368 = ~n28366 & ~n28367 ;
  assign n28369 = \ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131  & n23743 ;
  assign n28370 = n23741 & n28369 ;
  assign n28371 = \ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131  & n23743 ;
  assign n28372 = n23747 & n28371 ;
  assign n28373 = ~n28370 & ~n28372 ;
  assign n28374 = n28368 & n28373 ;
  assign n28375 = \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  & n23751 ;
  assign n28376 = n23741 & n28375 ;
  assign n28377 = \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131  & n23794 ;
  assign n28378 = n23741 & n28377 ;
  assign n28379 = ~n28376 & ~n28378 ;
  assign n28380 = n23730 & n28379 ;
  assign n28381 = n28374 & n28380 ;
  assign n28382 = \ethreg1_MODER_1_DataOut_reg[3]/NET0131  & n23808 ;
  assign n28383 = \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131  & n23802 ;
  assign n28384 = ~n28382 & ~n28383 ;
  assign n28385 = \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  & n23737 ;
  assign n28386 = \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131  & n23813 ;
  assign n28387 = ~n28385 & ~n28386 ;
  assign n28388 = n28384 & n28387 ;
  assign n28389 = n28381 & n28388 ;
  assign n28390 = n23730 & ~n28389 ;
  assign n28391 = \wishbone_bd_ram_mem1_reg[16][11]/P0001  & n13695 ;
  assign n28392 = \wishbone_bd_ram_mem1_reg[84][11]/P0001  & n13385 ;
  assign n28393 = ~n28391 & ~n28392 ;
  assign n28394 = \wishbone_bd_ram_mem1_reg[18][11]/P0001  & n13532 ;
  assign n28395 = \wishbone_bd_ram_mem1_reg[138][11]/P0001  & n13398 ;
  assign n28396 = ~n28394 & ~n28395 ;
  assign n28397 = n28393 & n28396 ;
  assign n28398 = \wishbone_bd_ram_mem1_reg[31][11]/P0001  & n13758 ;
  assign n28399 = \wishbone_bd_ram_mem1_reg[142][11]/P0001  & n13448 ;
  assign n28400 = ~n28398 & ~n28399 ;
  assign n28401 = \wishbone_bd_ram_mem1_reg[58][11]/P0001  & n13949 ;
  assign n28402 = \wishbone_bd_ram_mem1_reg[4][11]/P0001  & n13527 ;
  assign n28403 = ~n28401 & ~n28402 ;
  assign n28404 = n28400 & n28403 ;
  assign n28405 = n28397 & n28404 ;
  assign n28406 = \wishbone_bd_ram_mem1_reg[210][11]/P0001  & n13443 ;
  assign n28407 = \wishbone_bd_ram_mem1_reg[151][11]/P0001  & n13697 ;
  assign n28408 = ~n28406 & ~n28407 ;
  assign n28409 = \wishbone_bd_ram_mem1_reg[80][11]/P0001  & n13516 ;
  assign n28410 = \wishbone_bd_ram_mem1_reg[83][11]/P0001  & n13454 ;
  assign n28411 = ~n28409 & ~n28410 ;
  assign n28412 = n28408 & n28411 ;
  assign n28413 = \wishbone_bd_ram_mem1_reg[110][11]/P0001  & n14030 ;
  assign n28414 = \wishbone_bd_ram_mem1_reg[239][11]/P0001  & n13349 ;
  assign n28415 = ~n28413 & ~n28414 ;
  assign n28416 = \wishbone_bd_ram_mem1_reg[178][11]/P0001  & n13301 ;
  assign n28417 = \wishbone_bd_ram_mem1_reg[179][11]/P0001  & n14035 ;
  assign n28418 = ~n28416 & ~n28417 ;
  assign n28419 = n28415 & n28418 ;
  assign n28420 = n28412 & n28419 ;
  assign n28421 = n28405 & n28420 ;
  assign n28422 = \wishbone_bd_ram_mem1_reg[161][11]/P0001  & n13505 ;
  assign n28423 = \wishbone_bd_ram_mem1_reg[224][11]/P0001  & n13433 ;
  assign n28424 = ~n28422 & ~n28423 ;
  assign n28425 = \wishbone_bd_ram_mem1_reg[146][11]/P0001  & n13958 ;
  assign n28426 = \wishbone_bd_ram_mem1_reg[168][11]/P0001  & n13795 ;
  assign n28427 = ~n28425 & ~n28426 ;
  assign n28428 = n28424 & n28427 ;
  assign n28429 = \wishbone_bd_ram_mem1_reg[48][11]/P0001  & n13917 ;
  assign n28430 = \wishbone_bd_ram_mem1_reg[231][11]/P0001  & n13363 ;
  assign n28431 = ~n28429 & ~n28430 ;
  assign n28432 = \wishbone_bd_ram_mem1_reg[136][11]/P0001  & n13963 ;
  assign n28433 = \wishbone_bd_ram_mem1_reg[127][11]/P0001  & n13803 ;
  assign n28434 = ~n28432 & ~n28433 ;
  assign n28435 = n28431 & n28434 ;
  assign n28436 = n28428 & n28435 ;
  assign n28437 = \wishbone_bd_ram_mem1_reg[189][11]/P0001  & n14001 ;
  assign n28438 = \wishbone_bd_ram_mem1_reg[237][11]/P0001  & n13924 ;
  assign n28439 = ~n28437 & ~n28438 ;
  assign n28440 = \wishbone_bd_ram_mem1_reg[213][11]/P0001  & n13870 ;
  assign n28441 = \wishbone_bd_ram_mem1_reg[42][11]/P0001  & n13341 ;
  assign n28442 = ~n28440 & ~n28441 ;
  assign n28443 = n28439 & n28442 ;
  assign n28444 = \wishbone_bd_ram_mem1_reg[65][11]/P0001  & n13842 ;
  assign n28445 = \wishbone_bd_ram_mem1_reg[197][11]/P0001  & n13594 ;
  assign n28446 = ~n28444 & ~n28445 ;
  assign n28447 = \wishbone_bd_ram_mem1_reg[125][11]/P0001  & n13396 ;
  assign n28448 = \wishbone_bd_ram_mem1_reg[202][11]/P0001  & n13268 ;
  assign n28449 = ~n28447 & ~n28448 ;
  assign n28450 = n28446 & n28449 ;
  assign n28451 = n28443 & n28450 ;
  assign n28452 = n28436 & n28451 ;
  assign n28453 = n28421 & n28452 ;
  assign n28454 = \wishbone_bd_ram_mem1_reg[175][11]/P0001  & n13674 ;
  assign n28455 = \wishbone_bd_ram_mem1_reg[71][11]/P0001  & n13636 ;
  assign n28456 = ~n28454 & ~n28455 ;
  assign n28457 = \wishbone_bd_ram_mem1_reg[196][11]/P0001  & n13977 ;
  assign n28458 = \wishbone_bd_ram_mem1_reg[119][11]/P0001  & n14033 ;
  assign n28459 = ~n28457 & ~n28458 ;
  assign n28460 = n28456 & n28459 ;
  assign n28461 = \wishbone_bd_ram_mem1_reg[164][11]/P0001  & n13236 ;
  assign n28462 = \wishbone_bd_ram_mem1_reg[78][11]/P0001  & n13277 ;
  assign n28463 = ~n28461 & ~n28462 ;
  assign n28464 = \wishbone_bd_ram_mem1_reg[35][11]/P0001  & n13523 ;
  assign n28465 = \wishbone_bd_ram_mem1_reg[160][11]/P0001  & n13271 ;
  assign n28466 = ~n28464 & ~n28465 ;
  assign n28467 = n28463 & n28466 ;
  assign n28468 = n28460 & n28467 ;
  assign n28469 = \wishbone_bd_ram_mem1_reg[96][11]/P0001  & n13425 ;
  assign n28470 = \wishbone_bd_ram_mem1_reg[6][11]/P0001  & n13915 ;
  assign n28471 = ~n28469 & ~n28470 ;
  assign n28472 = \wishbone_bd_ram_mem1_reg[54][11]/P0001  & n13622 ;
  assign n28473 = \wishbone_bd_ram_mem1_reg[194][11]/P0001  & n13624 ;
  assign n28474 = ~n28472 & ~n28473 ;
  assign n28475 = n28471 & n28474 ;
  assign n28476 = \wishbone_bd_ram_mem1_reg[207][11]/P0001  & n13826 ;
  assign n28477 = \wishbone_bd_ram_mem1_reg[32][11]/P0001  & n13736 ;
  assign n28478 = ~n28476 & ~n28477 ;
  assign n28479 = \wishbone_bd_ram_mem1_reg[203][11]/P0001  & n13816 ;
  assign n28480 = \wishbone_bd_ram_mem1_reg[7][11]/P0001  & n13546 ;
  assign n28481 = ~n28479 & ~n28480 ;
  assign n28482 = n28478 & n28481 ;
  assign n28483 = n28475 & n28482 ;
  assign n28484 = n28468 & n28483 ;
  assign n28485 = \wishbone_bd_ram_mem1_reg[91][11]/P0001  & n13954 ;
  assign n28486 = \wishbone_bd_ram_mem1_reg[44][11]/P0001  & n13291 ;
  assign n28487 = ~n28485 & ~n28486 ;
  assign n28488 = \wishbone_bd_ram_mem1_reg[30][11]/P0001  & n13713 ;
  assign n28489 = \wishbone_bd_ram_mem1_reg[220][11]/P0001  & n13965 ;
  assign n28490 = ~n28488 & ~n28489 ;
  assign n28491 = n28487 & n28490 ;
  assign n28492 = \wishbone_bd_ram_mem1_reg[214][11]/P0001  & n13938 ;
  assign n28493 = \wishbone_bd_ram_mem1_reg[173][11]/P0001  & n13360 ;
  assign n28494 = ~n28492 & ~n28493 ;
  assign n28495 = \wishbone_bd_ram_mem1_reg[20][11]/P0001  & n13839 ;
  assign n28496 = \wishbone_bd_ram_mem1_reg[40][11]/P0001  & n13661 ;
  assign n28497 = ~n28495 & ~n28496 ;
  assign n28498 = n28494 & n28497 ;
  assign n28499 = n28491 & n28498 ;
  assign n28500 = \wishbone_bd_ram_mem1_reg[181][11]/P0001  & n13587 ;
  assign n28501 = \wishbone_bd_ram_mem1_reg[26][11]/P0001  & n13521 ;
  assign n28502 = ~n28500 & ~n28501 ;
  assign n28503 = \wishbone_bd_ram_mem1_reg[147][11]/P0001  & n13702 ;
  assign n28504 = \wishbone_bd_ram_mem1_reg[211][11]/P0001  & n13805 ;
  assign n28505 = ~n28503 & ~n28504 ;
  assign n28506 = n28502 & n28505 ;
  assign n28507 = \wishbone_bd_ram_mem1_reg[75][11]/P0001  & n13605 ;
  assign n28508 = \wishbone_bd_ram_mem1_reg[10][11]/P0001  & n13837 ;
  assign n28509 = ~n28507 & ~n28508 ;
  assign n28510 = \wishbone_bd_ram_mem1_reg[12][11]/P0001  & n13733 ;
  assign n28511 = \wishbone_bd_ram_mem1_reg[61][11]/P0001  & n13544 ;
  assign n28512 = ~n28510 & ~n28511 ;
  assign n28513 = n28509 & n28512 ;
  assign n28514 = n28506 & n28513 ;
  assign n28515 = n28499 & n28514 ;
  assign n28516 = n28484 & n28515 ;
  assign n28517 = n28453 & n28516 ;
  assign n28518 = \wishbone_bd_ram_mem1_reg[121][11]/P0001  & n13983 ;
  assign n28519 = \wishbone_bd_ram_mem1_reg[176][11]/P0001  & n13262 ;
  assign n28520 = ~n28518 & ~n28519 ;
  assign n28521 = \wishbone_bd_ram_mem1_reg[242][11]/P0001  & n13383 ;
  assign n28522 = \wishbone_bd_ram_mem1_reg[79][11]/P0001  & n13779 ;
  assign n28523 = ~n28521 & ~n28522 ;
  assign n28524 = n28520 & n28523 ;
  assign n28525 = \wishbone_bd_ram_mem1_reg[182][11]/P0001  & n13598 ;
  assign n28526 = \wishbone_bd_ram_mem1_reg[74][11]/P0001  & n13564 ;
  assign n28527 = ~n28525 & ~n28526 ;
  assign n28528 = \wishbone_bd_ram_mem1_reg[131][11]/P0001  & n13358 ;
  assign n28529 = \wishbone_bd_ram_mem1_reg[38][11]/P0001  & n13828 ;
  assign n28530 = ~n28528 & ~n28529 ;
  assign n28531 = n28527 & n28530 ;
  assign n28532 = n28524 & n28531 ;
  assign n28533 = \wishbone_bd_ram_mem1_reg[221][11]/P0001  & n13641 ;
  assign n28534 = \wishbone_bd_ram_mem1_reg[218][11]/P0001  & n13792 ;
  assign n28535 = ~n28533 & ~n28534 ;
  assign n28536 = \wishbone_bd_ram_mem1_reg[162][11]/P0001  & n13726 ;
  assign n28537 = \wishbone_bd_ram_mem1_reg[21][11]/P0001  & n13438 ;
  assign n28538 = ~n28536 & ~n28537 ;
  assign n28539 = n28535 & n28538 ;
  assign n28540 = \wishbone_bd_ram_mem1_reg[245][11]/P0001  & n13877 ;
  assign n28541 = \wishbone_bd_ram_mem1_reg[56][11]/P0001  & n13611 ;
  assign n28542 = ~n28540 & ~n28541 ;
  assign n28543 = \wishbone_bd_ram_mem1_reg[183][11]/P0001  & n13645 ;
  assign n28544 = \wishbone_bd_ram_mem1_reg[124][11]/P0001  & n14024 ;
  assign n28545 = ~n28543 & ~n28544 ;
  assign n28546 = n28542 & n28545 ;
  assign n28547 = n28539 & n28546 ;
  assign n28548 = n28532 & n28547 ;
  assign n28549 = \wishbone_bd_ram_mem1_reg[64][11]/P0001  & n13904 ;
  assign n28550 = \wishbone_bd_ram_mem1_reg[95][11]/P0001  & n13317 ;
  assign n28551 = ~n28549 & ~n28550 ;
  assign n28552 = \wishbone_bd_ram_mem1_reg[68][11]/P0001  & n13379 ;
  assign n28553 = \wishbone_bd_ram_mem1_reg[46][11]/P0001  & n13298 ;
  assign n28554 = ~n28552 & ~n28553 ;
  assign n28555 = n28551 & n28554 ;
  assign n28556 = \wishbone_bd_ram_mem1_reg[69][11]/P0001  & n13487 ;
  assign n28557 = \wishbone_bd_ram_mem1_reg[157][11]/P0001  & n13445 ;
  assign n28558 = ~n28556 & ~n28557 ;
  assign n28559 = \wishbone_bd_ram_mem1_reg[106][11]/P0001  & n13555 ;
  assign n28560 = \wishbone_bd_ram_mem1_reg[177][11]/P0001  & n13863 ;
  assign n28561 = ~n28559 & ~n28560 ;
  assign n28562 = n28558 & n28561 ;
  assign n28563 = n28555 & n28562 ;
  assign n28564 = \wishbone_bd_ram_mem1_reg[27][11]/P0001  & n13251 ;
  assign n28565 = \wishbone_bd_ram_mem1_reg[190][11]/P0001  & n13365 ;
  assign n28566 = ~n28564 & ~n28565 ;
  assign n28567 = \wishbone_bd_ram_mem1_reg[107][11]/P0001  & n13476 ;
  assign n28568 = \wishbone_bd_ram_mem1_reg[36][11]/P0001  & n13639 ;
  assign n28569 = ~n28567 & ~n28568 ;
  assign n28570 = n28566 & n28569 ;
  assign n28571 = \wishbone_bd_ram_mem1_reg[118][11]/P0001  & n13589 ;
  assign n28572 = \wishbone_bd_ram_mem1_reg[28][11]/P0001  & n13810 ;
  assign n28573 = ~n28571 & ~n28572 ;
  assign n28574 = \wishbone_bd_ram_mem1_reg[171][11]/P0001  & n13422 ;
  assign n28575 = \wishbone_bd_ram_mem1_reg[163][11]/P0001  & n13255 ;
  assign n28576 = ~n28574 & ~n28575 ;
  assign n28577 = n28573 & n28576 ;
  assign n28578 = n28570 & n28577 ;
  assign n28579 = n28563 & n28578 ;
  assign n28580 = n28548 & n28579 ;
  assign n28581 = \wishbone_bd_ram_mem1_reg[246][11]/P0001  & n13981 ;
  assign n28582 = \wishbone_bd_ram_mem1_reg[122][11]/P0001  & n13679 ;
  assign n28583 = ~n28581 & ~n28582 ;
  assign n28584 = \wishbone_bd_ram_mem1_reg[174][11]/P0001  & n13899 ;
  assign n28585 = \wishbone_bd_ram_mem1_reg[180][11]/P0001  & n13650 ;
  assign n28586 = ~n28584 & ~n28585 ;
  assign n28587 = n28583 & n28586 ;
  assign n28588 = \wishbone_bd_ram_mem1_reg[8][11]/P0001  & n13459 ;
  assign n28589 = \wishbone_bd_ram_mem1_reg[234][11]/P0001  & n13781 ;
  assign n28590 = ~n28588 & ~n28589 ;
  assign n28591 = \wishbone_bd_ram_mem1_reg[148][11]/P0001  & n13868 ;
  assign n28592 = \wishbone_bd_ram_mem1_reg[98][11]/P0001  & n13569 ;
  assign n28593 = ~n28591 & ~n28592 ;
  assign n28594 = n28590 & n28593 ;
  assign n28595 = n28587 & n28594 ;
  assign n28596 = \wishbone_bd_ram_mem1_reg[222][11]/P0001  & n13721 ;
  assign n28597 = \wishbone_bd_ram_mem1_reg[191][11]/P0001  & n14012 ;
  assign n28598 = ~n28596 & ~n28597 ;
  assign n28599 = \wishbone_bd_ram_mem1_reg[99][11]/P0001  & n13996 ;
  assign n28600 = \wishbone_bd_ram_mem1_reg[192][11]/P0001  & n13390 ;
  assign n28601 = ~n28599 & ~n28600 ;
  assign n28602 = n28598 & n28601 ;
  assign n28603 = \wishbone_bd_ram_mem1_reg[90][11]/P0001  & n13906 ;
  assign n28604 = \wishbone_bd_ram_mem1_reg[206][11]/P0001  & n13414 ;
  assign n28605 = ~n28603 & ~n28604 ;
  assign n28606 = \wishbone_bd_ram_mem1_reg[82][11]/P0001  & n13374 ;
  assign n28607 = \wishbone_bd_ram_mem1_reg[111][11]/P0001  & n13471 ;
  assign n28608 = ~n28606 & ~n28607 ;
  assign n28609 = n28605 & n28608 ;
  assign n28610 = n28602 & n28609 ;
  assign n28611 = n28595 & n28610 ;
  assign n28612 = \wishbone_bd_ram_mem1_reg[62][11]/P0001  & n13529 ;
  assign n28613 = \wishbone_bd_ram_mem1_reg[134][11]/P0001  & n13494 ;
  assign n28614 = ~n28612 & ~n28613 ;
  assign n28615 = \wishbone_bd_ram_mem1_reg[184][11]/P0001  & n13960 ;
  assign n28616 = \wishbone_bd_ram_mem1_reg[219][11]/P0001  & n13577 ;
  assign n28617 = ~n28615 & ~n28616 ;
  assign n28618 = n28614 & n28617 ;
  assign n28619 = \wishbone_bd_ram_mem1_reg[123][11]/P0001  & n13749 ;
  assign n28620 = \wishbone_bd_ram_mem1_reg[217][11]/P0001  & n13767 ;
  assign n28621 = ~n28619 & ~n28620 ;
  assign n28622 = \wishbone_bd_ram_mem1_reg[250][11]/P0001  & n13677 ;
  assign n28623 = \wishbone_bd_ram_mem1_reg[154][11]/P0001  & n13403 ;
  assign n28624 = ~n28622 & ~n28623 ;
  assign n28625 = n28621 & n28624 ;
  assign n28626 = n28618 & n28625 ;
  assign n28627 = \wishbone_bd_ram_mem1_reg[185][11]/P0001  & n13372 ;
  assign n28628 = \wishbone_bd_ram_mem1_reg[232][11]/P0001  & n13510 ;
  assign n28629 = ~n28627 & ~n28628 ;
  assign n28630 = \wishbone_bd_ram_mem1_reg[55][11]/P0001  & n13618 ;
  assign n28631 = \wishbone_bd_ram_mem1_reg[101][11]/P0001  & n13772 ;
  assign n28632 = ~n28630 & ~n28631 ;
  assign n28633 = n28629 & n28632 ;
  assign n28634 = \wishbone_bd_ram_mem1_reg[33][11]/P0001  & n13933 ;
  assign n28635 = \wishbone_bd_ram_mem1_reg[253][11]/P0001  & n13708 ;
  assign n28636 = ~n28634 & ~n28635 ;
  assign n28637 = \wishbone_bd_ram_mem1_reg[113][11]/P0001  & n13882 ;
  assign n28638 = \wishbone_bd_ram_mem1_reg[153][11]/P0001  & n13309 ;
  assign n28639 = ~n28637 & ~n28638 ;
  assign n28640 = n28636 & n28639 ;
  assign n28641 = n28633 & n28640 ;
  assign n28642 = n28626 & n28641 ;
  assign n28643 = n28611 & n28642 ;
  assign n28644 = n28580 & n28643 ;
  assign n28645 = n28517 & n28644 ;
  assign n28646 = \wishbone_bd_ram_mem1_reg[103][11]/P0001  & n13320 ;
  assign n28647 = \wishbone_bd_ram_mem1_reg[205][11]/P0001  & n13947 ;
  assign n28648 = ~n28646 & ~n28647 ;
  assign n28649 = \wishbone_bd_ram_mem1_reg[132][11]/P0001  & n13927 ;
  assign n28650 = \wishbone_bd_ram_mem1_reg[247][11]/P0001  & n13571 ;
  assign n28651 = ~n28649 & ~n28650 ;
  assign n28652 = n28648 & n28651 ;
  assign n28653 = \wishbone_bd_ram_mem1_reg[200][11]/P0001  & n13922 ;
  assign n28654 = \wishbone_bd_ram_mem1_reg[114][11]/P0001  & n13763 ;
  assign n28655 = ~n28653 & ~n28654 ;
  assign n28656 = \wishbone_bd_ram_mem1_reg[252][11]/P0001  & n13986 ;
  assign n28657 = \wishbone_bd_ram_mem1_reg[201][11]/P0001  & n13600 ;
  assign n28658 = ~n28656 & ~n28657 ;
  assign n28659 = n28655 & n28658 ;
  assign n28660 = n28652 & n28659 ;
  assign n28661 = \wishbone_bd_ram_mem1_reg[236][11]/P0001  & n13480 ;
  assign n28662 = \wishbone_bd_ram_mem1_reg[2][11]/P0001  & n13975 ;
  assign n28663 = ~n28661 & ~n28662 ;
  assign n28664 = \wishbone_bd_ram_mem1_reg[199][11]/P0001  & n13499 ;
  assign n28665 = \wishbone_bd_ram_mem1_reg[81][11]/P0001  & n13409 ;
  assign n28666 = ~n28664 & ~n28665 ;
  assign n28667 = n28663 & n28666 ;
  assign n28668 = \wishbone_bd_ram_mem1_reg[241][11]/P0001  & n13854 ;
  assign n28669 = \wishbone_bd_ram_mem1_reg[141][11]/P0001  & n13852 ;
  assign n28670 = ~n28668 & ~n28669 ;
  assign n28671 = \wishbone_bd_ram_mem1_reg[51][11]/P0001  & n13880 ;
  assign n28672 = \wishbone_bd_ram_mem1_reg[129][11]/P0001  & n13629 ;
  assign n28673 = ~n28671 & ~n28672 ;
  assign n28674 = n28670 & n28673 ;
  assign n28675 = n28667 & n28674 ;
  assign n28676 = n28660 & n28675 ;
  assign n28677 = \wishbone_bd_ram_mem1_reg[14][11]/P0001  & n13972 ;
  assign n28678 = \wishbone_bd_ram_mem1_reg[128][11]/P0001  & n13652 ;
  assign n28679 = ~n28677 & ~n28678 ;
  assign n28680 = \wishbone_bd_ram_mem1_reg[144][11]/P0001  & n13508 ;
  assign n28681 = \wishbone_bd_ram_mem1_reg[170][11]/P0001  & n14007 ;
  assign n28682 = ~n28680 & ~n28681 ;
  assign n28683 = n28679 & n28682 ;
  assign n28684 = \wishbone_bd_ram_mem1_reg[150][11]/P0001  & n13666 ;
  assign n28685 = \wishbone_bd_ram_mem1_reg[216][11]/P0001  & n14005 ;
  assign n28686 = ~n28684 & ~n28685 ;
  assign n28687 = \wishbone_bd_ram_mem1_reg[208][11]/P0001  & n14010 ;
  assign n28688 = \wishbone_bd_ram_mem1_reg[115][11]/P0001  & n13747 ;
  assign n28689 = ~n28687 & ~n28688 ;
  assign n28690 = n28686 & n28689 ;
  assign n28691 = n28683 & n28690 ;
  assign n28692 = \wishbone_bd_ram_mem1_reg[49][11]/P0001  & n13929 ;
  assign n28693 = \wishbone_bd_ram_mem1_reg[104][11]/P0001  & n13684 ;
  assign n28694 = ~n28692 & ~n28693 ;
  assign n28695 = \wishbone_bd_ram_mem1_reg[76][11]/P0001  & n13831 ;
  assign n28696 = \wishbone_bd_ram_mem1_reg[73][11]/P0001  & n13456 ;
  assign n28697 = ~n28695 & ~n28696 ;
  assign n28698 = n28694 & n28697 ;
  assign n28699 = \wishbone_bd_ram_mem1_reg[186][11]/P0001  & n13616 ;
  assign n28700 = \wishbone_bd_ram_mem1_reg[25][11]/P0001  & n13742 ;
  assign n28701 = ~n28699 & ~n28700 ;
  assign n28702 = \wishbone_bd_ram_mem1_reg[188][11]/P0001  & n13407 ;
  assign n28703 = \wishbone_bd_ram_mem1_reg[172][11]/P0001  & n13377 ;
  assign n28704 = ~n28702 & ~n28703 ;
  assign n28705 = n28701 & n28704 ;
  assign n28706 = n28698 & n28705 ;
  assign n28707 = n28691 & n28706 ;
  assign n28708 = n28676 & n28707 ;
  assign n28709 = \wishbone_bd_ram_mem1_reg[215][11]/P0001  & n13901 ;
  assign n28710 = \wishbone_bd_ram_mem1_reg[93][11]/P0001  & n13891 ;
  assign n28711 = ~n28709 & ~n28710 ;
  assign n28712 = \wishbone_bd_ram_mem1_reg[120][11]/P0001  & n13550 ;
  assign n28713 = \wishbone_bd_ram_mem1_reg[212][11]/P0001  & n13634 ;
  assign n28714 = ~n28712 & ~n28713 ;
  assign n28715 = n28711 & n28714 ;
  assign n28716 = \wishbone_bd_ram_mem1_reg[227][11]/P0001  & n13388 ;
  assign n28717 = \wishbone_bd_ram_mem1_reg[255][11]/P0001  & n13952 ;
  assign n28718 = ~n28716 & ~n28717 ;
  assign n28719 = \wishbone_bd_ram_mem1_reg[53][11]/P0001  & n13875 ;
  assign n28720 = \wishbone_bd_ram_mem1_reg[169][11]/P0001  & n13541 ;
  assign n28721 = ~n28719 & ~n28720 ;
  assign n28722 = n28718 & n28721 ;
  assign n28723 = n28715 & n28722 ;
  assign n28724 = \wishbone_bd_ram_mem1_reg[72][11]/P0001  & n13582 ;
  assign n28725 = \wishbone_bd_ram_mem1_reg[66][11]/P0001  & n13603 ;
  assign n28726 = ~n28724 & ~n28725 ;
  assign n28727 = \wishbone_bd_ram_mem1_reg[108][11]/P0001  & n13814 ;
  assign n28728 = \wishbone_bd_ram_mem1_reg[243][11]/P0001  & n13575 ;
  assign n28729 = ~n28727 & ~n28728 ;
  assign n28730 = n28726 & n28729 ;
  assign n28731 = \wishbone_bd_ram_mem1_reg[47][11]/P0001  & n13436 ;
  assign n28732 = \wishbone_bd_ram_mem1_reg[117][11]/P0001  & n13557 ;
  assign n28733 = ~n28731 & ~n28732 ;
  assign n28734 = \wishbone_bd_ram_mem1_reg[112][11]/P0001  & n13482 ;
  assign n28735 = \wishbone_bd_ram_mem1_reg[87][11]/P0001  & n13691 ;
  assign n28736 = ~n28734 & ~n28735 ;
  assign n28737 = n28733 & n28736 ;
  assign n28738 = n28730 & n28737 ;
  assign n28739 = n28723 & n28738 ;
  assign n28740 = \wishbone_bd_ram_mem1_reg[223][11]/P0001  & n13335 ;
  assign n28741 = \wishbone_bd_ram_mem1_reg[43][11]/P0001  & n13761 ;
  assign n28742 = ~n28740 & ~n28741 ;
  assign n28743 = \wishbone_bd_ram_mem1_reg[233][11]/P0001  & n13332 ;
  assign n28744 = \wishbone_bd_ram_mem1_reg[152][11]/P0001  & n13912 ;
  assign n28745 = ~n28743 & ~n28744 ;
  assign n28746 = n28742 & n28745 ;
  assign n28747 = \wishbone_bd_ram_mem1_reg[67][11]/P0001  & n13663 ;
  assign n28748 = \wishbone_bd_ram_mem1_reg[9][11]/P0001  & n13580 ;
  assign n28749 = ~n28747 & ~n28748 ;
  assign n28750 = \wishbone_bd_ram_mem1_reg[100][11]/P0001  & n13401 ;
  assign n28751 = \wishbone_bd_ram_mem1_reg[0][11]/P0001  & n13539 ;
  assign n28752 = ~n28750 & ~n28751 ;
  assign n28753 = n28749 & n28752 ;
  assign n28754 = n28746 & n28753 ;
  assign n28755 = \wishbone_bd_ram_mem1_reg[41][11]/P0001  & n14017 ;
  assign n28756 = \wishbone_bd_ram_mem1_reg[89][11]/P0001  & n13910 ;
  assign n28757 = ~n28755 & ~n28756 ;
  assign n28758 = \wishbone_bd_ram_mem1_reg[45][11]/P0001  & n13420 ;
  assign n28759 = \wishbone_bd_ram_mem1_reg[248][11]/P0001  & n13647 ;
  assign n28760 = ~n28758 & ~n28759 ;
  assign n28761 = n28757 & n28760 ;
  assign n28762 = \wishbone_bd_ram_mem1_reg[109][11]/P0001  & n13306 ;
  assign n28763 = \wishbone_bd_ram_mem1_reg[88][11]/P0001  & n13347 ;
  assign n28764 = ~n28762 & ~n28763 ;
  assign n28765 = \wishbone_bd_ram_mem1_reg[3][11]/P0001  & n13354 ;
  assign n28766 = \wishbone_bd_ram_mem1_reg[17][11]/P0001  & n13324 ;
  assign n28767 = ~n28765 & ~n28766 ;
  assign n28768 = n28764 & n28767 ;
  assign n28769 = n28761 & n28768 ;
  assign n28770 = n28754 & n28769 ;
  assign n28771 = n28739 & n28770 ;
  assign n28772 = n28708 & n28771 ;
  assign n28773 = \wishbone_bd_ram_mem1_reg[37][11]/P0001  & n13710 ;
  assign n28774 = \wishbone_bd_ram_mem1_reg[167][11]/P0001  & n13940 ;
  assign n28775 = ~n28773 & ~n28774 ;
  assign n28776 = \wishbone_bd_ram_mem1_reg[254][11]/P0001  & n13283 ;
  assign n28777 = \wishbone_bd_ram_mem1_reg[198][11]/P0001  & n13592 ;
  assign n28778 = ~n28776 & ~n28777 ;
  assign n28779 = n28775 & n28778 ;
  assign n28780 = \wishbone_bd_ram_mem1_reg[50][11]/P0001  & n13686 ;
  assign n28781 = \wishbone_bd_ram_mem1_reg[229][11]/P0001  & n13552 ;
  assign n28782 = ~n28780 & ~n28781 ;
  assign n28783 = \wishbone_bd_ram_mem1_reg[130][11]/P0001  & n13427 ;
  assign n28784 = \wishbone_bd_ram_mem1_reg[187][11]/P0001  & n13756 ;
  assign n28785 = ~n28783 & ~n28784 ;
  assign n28786 = n28782 & n28785 ;
  assign n28787 = n28779 & n28786 ;
  assign n28788 = \wishbone_bd_ram_mem1_reg[22][11]/P0001  & n13744 ;
  assign n28789 = \wishbone_bd_ram_mem1_reg[193][11]/P0001  & n14022 ;
  assign n28790 = ~n28788 & ~n28789 ;
  assign n28791 = \wishbone_bd_ram_mem1_reg[11][11]/P0001  & n13774 ;
  assign n28792 = \wishbone_bd_ram_mem1_reg[145][11]/P0001  & n13715 ;
  assign n28793 = ~n28791 & ~n28792 ;
  assign n28794 = n28790 & n28793 ;
  assign n28795 = \wishbone_bd_ram_mem1_reg[105][11]/P0001  & n13503 ;
  assign n28796 = \wishbone_bd_ram_mem1_reg[52][11]/P0001  & n13988 ;
  assign n28797 = ~n28795 & ~n28796 ;
  assign n28798 = \wishbone_bd_ram_mem1_reg[155][11]/P0001  & n13738 ;
  assign n28799 = \wishbone_bd_ram_mem1_reg[85][11]/P0001  & n13784 ;
  assign n28800 = ~n28798 & ~n28799 ;
  assign n28801 = n28797 & n28800 ;
  assign n28802 = n28794 & n28801 ;
  assign n28803 = n28787 & n28802 ;
  assign n28804 = \wishbone_bd_ram_mem1_reg[24][11]/P0001  & n13970 ;
  assign n28805 = \wishbone_bd_ram_mem1_reg[240][11]/P0001  & n13352 ;
  assign n28806 = ~n28804 & ~n28805 ;
  assign n28807 = \wishbone_bd_ram_mem1_reg[230][11]/P0001  & n13994 ;
  assign n28808 = \wishbone_bd_ram_mem1_reg[126][11]/P0001  & n13786 ;
  assign n28809 = ~n28807 & ~n28808 ;
  assign n28810 = n28806 & n28809 ;
  assign n28811 = \wishbone_bd_ram_mem1_reg[39][11]/P0001  & n13893 ;
  assign n28812 = \wishbone_bd_ram_mem1_reg[133][11]/P0001  & n13492 ;
  assign n28813 = ~n28811 & ~n28812 ;
  assign n28814 = \wishbone_bd_ram_mem1_reg[159][11]/P0001  & n13627 ;
  assign n28815 = \wishbone_bd_ram_mem1_reg[139][11]/P0001  & n13566 ;
  assign n28816 = ~n28814 & ~n28815 ;
  assign n28817 = n28813 & n28816 ;
  assign n28818 = n28810 & n28817 ;
  assign n28819 = \wishbone_bd_ram_mem1_reg[60][11]/P0001  & n13790 ;
  assign n28820 = \wishbone_bd_ram_mem1_reg[228][11]/P0001  & n13497 ;
  assign n28821 = ~n28819 & ~n28820 ;
  assign n28822 = \wishbone_bd_ram_mem1_reg[92][11]/P0001  & n13859 ;
  assign n28823 = \wishbone_bd_ram_mem1_reg[13][11]/P0001  & n13844 ;
  assign n28824 = ~n28822 & ~n28823 ;
  assign n28825 = n28821 & n28824 ;
  assign n28826 = \wishbone_bd_ram_mem1_reg[5][11]/P0001  & n13243 ;
  assign n28827 = \wishbone_bd_ram_mem1_reg[143][11]/P0001  & n13461 ;
  assign n28828 = ~n28826 & ~n28827 ;
  assign n28829 = \wishbone_bd_ram_mem1_reg[226][11]/P0001  & n13668 ;
  assign n28830 = \wishbone_bd_ram_mem1_reg[70][11]/P0001  & n13339 ;
  assign n28831 = ~n28829 & ~n28830 ;
  assign n28832 = n28828 & n28831 ;
  assign n28833 = n28825 & n28832 ;
  assign n28834 = n28818 & n28833 ;
  assign n28835 = n28803 & n28834 ;
  assign n28836 = \wishbone_bd_ram_mem1_reg[235][11]/P0001  & n13518 ;
  assign n28837 = \wishbone_bd_ram_mem1_reg[135][11]/P0001  & n13672 ;
  assign n28838 = ~n28836 & ~n28837 ;
  assign n28839 = \wishbone_bd_ram_mem1_reg[149][11]/P0001  & n13469 ;
  assign n28840 = \wishbone_bd_ram_mem1_reg[63][11]/P0001  & n13327 ;
  assign n28841 = ~n28839 & ~n28840 ;
  assign n28842 = n28838 & n28841 ;
  assign n28843 = \wishbone_bd_ram_mem1_reg[156][11]/P0001  & n13769 ;
  assign n28844 = \wishbone_bd_ram_mem1_reg[225][11]/P0001  & n13719 ;
  assign n28845 = ~n28843 & ~n28844 ;
  assign n28846 = \wishbone_bd_ram_mem1_reg[238][11]/P0001  & n13819 ;
  assign n28847 = \wishbone_bd_ram_mem1_reg[57][11]/P0001  & n13731 ;
  assign n28848 = ~n28846 & ~n28847 ;
  assign n28849 = n28845 & n28848 ;
  assign n28850 = n28842 & n28849 ;
  assign n28851 = \wishbone_bd_ram_mem1_reg[86][11]/P0001  & n13485 ;
  assign n28852 = \wishbone_bd_ram_mem1_reg[19][11]/P0001  & n13886 ;
  assign n28853 = ~n28851 & ~n28852 ;
  assign n28854 = \wishbone_bd_ram_mem1_reg[166][11]/P0001  & n13999 ;
  assign n28855 = \wishbone_bd_ram_mem1_reg[34][11]/P0001  & n13450 ;
  assign n28856 = ~n28854 & ~n28855 ;
  assign n28857 = n28853 & n28856 ;
  assign n28858 = \wishbone_bd_ram_mem1_reg[251][11]/P0001  & n14019 ;
  assign n28859 = \wishbone_bd_ram_mem1_reg[77][11]/P0001  & n13935 ;
  assign n28860 = ~n28858 & ~n28859 ;
  assign n28861 = \wishbone_bd_ram_mem1_reg[165][11]/P0001  & n14028 ;
  assign n28862 = \wishbone_bd_ram_mem1_reg[244][11]/P0001  & n13474 ;
  assign n28863 = ~n28861 & ~n28862 ;
  assign n28864 = n28860 & n28863 ;
  assign n28865 = n28857 & n28864 ;
  assign n28866 = n28850 & n28865 ;
  assign n28867 = \wishbone_bd_ram_mem1_reg[102][11]/P0001  & n13534 ;
  assign n28868 = \wishbone_bd_ram_mem1_reg[158][11]/P0001  & n13294 ;
  assign n28869 = ~n28867 & ~n28868 ;
  assign n28870 = \wishbone_bd_ram_mem1_reg[140][11]/P0001  & n13287 ;
  assign n28871 = \wishbone_bd_ram_mem1_reg[137][11]/P0001  & n13808 ;
  assign n28872 = ~n28870 & ~n28871 ;
  assign n28873 = n28869 & n28872 ;
  assign n28874 = \wishbone_bd_ram_mem1_reg[116][11]/P0001  & n13865 ;
  assign n28875 = \wishbone_bd_ram_mem1_reg[29][11]/P0001  & n13412 ;
  assign n28876 = ~n28874 & ~n28875 ;
  assign n28877 = \wishbone_bd_ram_mem1_reg[59][11]/P0001  & n13613 ;
  assign n28878 = \wishbone_bd_ram_mem1_reg[204][11]/P0001  & n13821 ;
  assign n28879 = ~n28877 & ~n28878 ;
  assign n28880 = n28876 & n28879 ;
  assign n28881 = n28873 & n28880 ;
  assign n28882 = \wishbone_bd_ram_mem1_reg[15][11]/P0001  & n13797 ;
  assign n28883 = \wishbone_bd_ram_mem1_reg[97][11]/P0001  & n13724 ;
  assign n28884 = ~n28882 & ~n28883 ;
  assign n28885 = \wishbone_bd_ram_mem1_reg[94][11]/P0001  & n13833 ;
  assign n28886 = \wishbone_bd_ram_mem1_reg[195][11]/P0001  & n13700 ;
  assign n28887 = ~n28885 & ~n28886 ;
  assign n28888 = n28884 & n28887 ;
  assign n28889 = \wishbone_bd_ram_mem1_reg[23][11]/P0001  & n13857 ;
  assign n28890 = \wishbone_bd_ram_mem1_reg[249][11]/P0001  & n13431 ;
  assign n28891 = ~n28889 & ~n28890 ;
  assign n28892 = \wishbone_bd_ram_mem1_reg[1][11]/P0001  & n13888 ;
  assign n28893 = \wishbone_bd_ram_mem1_reg[209][11]/P0001  & n13689 ;
  assign n28894 = ~n28892 & ~n28893 ;
  assign n28895 = n28891 & n28894 ;
  assign n28896 = n28888 & n28895 ;
  assign n28897 = n28881 & n28896 ;
  assign n28898 = n28866 & n28897 ;
  assign n28899 = n28835 & n28898 ;
  assign n28900 = n28772 & n28899 ;
  assign n28901 = n28645 & n28900 ;
  assign n28902 = ~wb_rst_i_pad & ~n28389 ;
  assign n28903 = ~n28901 & n28902 ;
  assign n28904 = ~n28390 & ~n28903 ;
  assign n28905 = ~\wishbone_TxLength_reg[10]/NET0131  & n14053 ;
  assign n28906 = n14057 & n28905 ;
  assign n28907 = ~n17918 & n28906 ;
  assign n28908 = \wishbone_TxLength_reg[11]/NET0131  & n28907 ;
  assign n28909 = ~\wishbone_TxLength_reg[11]/NET0131  & ~n28907 ;
  assign n28910 = n19277 & ~n28909 ;
  assign n28911 = ~n28908 & n28910 ;
  assign n28912 = ~n21644 & ~n28911 ;
  assign n28913 = \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  & n23737 ;
  assign n28914 = \ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131  & n23743 ;
  assign n28915 = n23747 & n28914 ;
  assign n28916 = \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  & n25084 ;
  assign n28917 = ~n28915 & ~n28916 ;
  assign n28918 = \ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131  & n23743 ;
  assign n28919 = n23741 & n28918 ;
  assign n28920 = \ethreg1_IPGT_0_DataOut_reg[2]/NET0131  & n25090 ;
  assign n28921 = ~n28919 & ~n28920 ;
  assign n28922 = n28917 & n28921 ;
  assign n28923 = \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131  & n25079 ;
  assign n28924 = \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  & n23751 ;
  assign n28925 = n23747 & n28924 ;
  assign n28926 = ~n28923 & ~n28925 ;
  assign n28927 = \ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131  & n23782 ;
  assign n28928 = \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131  & n25088 ;
  assign n28929 = ~n28927 & ~n28928 ;
  assign n28930 = n28926 & n28929 ;
  assign n28931 = n28922 & n28930 ;
  assign n28932 = ~n28913 & n28931 ;
  assign n28933 = \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  & n23751 ;
  assign n28934 = n23741 & n28933 ;
  assign n28935 = \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131  & n23794 ;
  assign n28936 = n23741 & n28935 ;
  assign n28937 = ~n28934 & ~n28936 ;
  assign n28938 = \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131  & n25069 ;
  assign n28939 = n23801 & n25063 ;
  assign n28940 = \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  & n28939 ;
  assign n28941 = ~n28938 & ~n28940 ;
  assign n28942 = n28937 & n28941 ;
  assign n28943 = n23730 & n28942 ;
  assign n28944 = \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131  & n23802 ;
  assign n28945 = n23781 & n23812 ;
  assign n28946 = \miim1_Nvalid_reg/NET0131  & n28945 ;
  assign n28947 = ~n28944 & ~n28946 ;
  assign n28948 = n23781 & n25063 ;
  assign n28949 = \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131  & n28948 ;
  assign n28950 = \ethreg1_irq_rxb_reg/NET0131  & n25064 ;
  assign n28951 = ~n28949 & ~n28950 ;
  assign n28952 = n28947 & n28951 ;
  assign n28953 = \ethreg1_MODER_0_DataOut_reg[2]/NET0131  & n23808 ;
  assign n28954 = \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131  & n23813 ;
  assign n28955 = ~n28953 & ~n28954 ;
  assign n28956 = n23812 & n25078 ;
  assign n28957 = \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  & n28956 ;
  assign n28958 = \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131  & n25082 ;
  assign n28959 = ~n28957 & ~n28958 ;
  assign n28960 = n28955 & n28959 ;
  assign n28961 = n28952 & n28960 ;
  assign n28962 = n28943 & n28961 ;
  assign n28963 = n28932 & n28962 ;
  assign n28964 = n23730 & ~n28963 ;
  assign n28965 = \wishbone_bd_ram_mem0_reg[43][2]/P0001  & n13761 ;
  assign n28966 = \wishbone_bd_ram_mem0_reg[13][2]/P0001  & n13844 ;
  assign n28967 = ~n28965 & ~n28966 ;
  assign n28968 = \wishbone_bd_ram_mem0_reg[50][2]/P0001  & n13686 ;
  assign n28969 = \wishbone_bd_ram_mem0_reg[87][2]/P0001  & n13691 ;
  assign n28970 = ~n28968 & ~n28969 ;
  assign n28971 = n28967 & n28970 ;
  assign n28972 = \wishbone_bd_ram_mem0_reg[91][2]/P0001  & n13954 ;
  assign n28973 = \wishbone_bd_ram_mem0_reg[193][2]/P0001  & n14022 ;
  assign n28974 = ~n28972 & ~n28973 ;
  assign n28975 = \wishbone_bd_ram_mem0_reg[160][2]/P0001  & n13271 ;
  assign n28976 = \wishbone_bd_ram_mem0_reg[236][2]/P0001  & n13480 ;
  assign n28977 = ~n28975 & ~n28976 ;
  assign n28978 = n28974 & n28977 ;
  assign n28979 = n28971 & n28978 ;
  assign n28980 = \wishbone_bd_ram_mem0_reg[240][2]/P0001  & n13352 ;
  assign n28981 = \wishbone_bd_ram_mem0_reg[179][2]/P0001  & n14035 ;
  assign n28982 = ~n28980 & ~n28981 ;
  assign n28983 = \wishbone_bd_ram_mem0_reg[34][2]/P0001  & n13450 ;
  assign n28984 = \wishbone_bd_ram_mem0_reg[186][2]/P0001  & n13616 ;
  assign n28985 = ~n28983 & ~n28984 ;
  assign n28986 = n28982 & n28985 ;
  assign n28987 = \wishbone_bd_ram_mem0_reg[28][2]/P0001  & n13810 ;
  assign n28988 = \wishbone_bd_ram_mem0_reg[248][2]/P0001  & n13647 ;
  assign n28989 = ~n28987 & ~n28988 ;
  assign n28990 = \wishbone_bd_ram_mem0_reg[11][2]/P0001  & n13774 ;
  assign n28991 = \wishbone_bd_ram_mem0_reg[231][2]/P0001  & n13363 ;
  assign n28992 = ~n28990 & ~n28991 ;
  assign n28993 = n28989 & n28992 ;
  assign n28994 = n28986 & n28993 ;
  assign n28995 = n28979 & n28994 ;
  assign n28996 = \wishbone_bd_ram_mem0_reg[104][2]/P0001  & n13684 ;
  assign n28997 = \wishbone_bd_ram_mem0_reg[153][2]/P0001  & n13309 ;
  assign n28998 = ~n28996 & ~n28997 ;
  assign n28999 = \wishbone_bd_ram_mem0_reg[44][2]/P0001  & n13291 ;
  assign n29000 = \wishbone_bd_ram_mem0_reg[59][2]/P0001  & n13613 ;
  assign n29001 = ~n28999 & ~n29000 ;
  assign n29002 = n28998 & n29001 ;
  assign n29003 = \wishbone_bd_ram_mem0_reg[233][2]/P0001  & n13332 ;
  assign n29004 = \wishbone_bd_ram_mem0_reg[183][2]/P0001  & n13645 ;
  assign n29005 = ~n29003 & ~n29004 ;
  assign n29006 = \wishbone_bd_ram_mem0_reg[70][2]/P0001  & n13339 ;
  assign n29007 = \wishbone_bd_ram_mem0_reg[2][2]/P0001  & n13975 ;
  assign n29008 = ~n29006 & ~n29007 ;
  assign n29009 = n29005 & n29008 ;
  assign n29010 = n29002 & n29009 ;
  assign n29011 = \wishbone_bd_ram_mem0_reg[166][2]/P0001  & n13999 ;
  assign n29012 = \wishbone_bd_ram_mem0_reg[207][2]/P0001  & n13826 ;
  assign n29013 = ~n29011 & ~n29012 ;
  assign n29014 = \wishbone_bd_ram_mem0_reg[178][2]/P0001  & n13301 ;
  assign n29015 = \wishbone_bd_ram_mem0_reg[118][2]/P0001  & n13589 ;
  assign n29016 = ~n29014 & ~n29015 ;
  assign n29017 = n29013 & n29016 ;
  assign n29018 = \wishbone_bd_ram_mem0_reg[1][2]/P0001  & n13888 ;
  assign n29019 = \wishbone_bd_ram_mem0_reg[170][2]/P0001  & n14007 ;
  assign n29020 = ~n29018 & ~n29019 ;
  assign n29021 = \wishbone_bd_ram_mem0_reg[103][2]/P0001  & n13320 ;
  assign n29022 = \wishbone_bd_ram_mem0_reg[194][2]/P0001  & n13624 ;
  assign n29023 = ~n29021 & ~n29022 ;
  assign n29024 = n29020 & n29023 ;
  assign n29025 = n29017 & n29024 ;
  assign n29026 = n29010 & n29025 ;
  assign n29027 = n28995 & n29026 ;
  assign n29028 = \wishbone_bd_ram_mem0_reg[88][2]/P0001  & n13347 ;
  assign n29029 = \wishbone_bd_ram_mem0_reg[82][2]/P0001  & n13374 ;
  assign n29030 = ~n29028 & ~n29029 ;
  assign n29031 = \wishbone_bd_ram_mem0_reg[169][2]/P0001  & n13541 ;
  assign n29032 = \wishbone_bd_ram_mem0_reg[84][2]/P0001  & n13385 ;
  assign n29033 = ~n29031 & ~n29032 ;
  assign n29034 = n29030 & n29033 ;
  assign n29035 = \wishbone_bd_ram_mem0_reg[199][2]/P0001  & n13499 ;
  assign n29036 = \wishbone_bd_ram_mem0_reg[164][2]/P0001  & n13236 ;
  assign n29037 = ~n29035 & ~n29036 ;
  assign n29038 = \wishbone_bd_ram_mem0_reg[249][2]/P0001  & n13431 ;
  assign n29039 = \wishbone_bd_ram_mem0_reg[98][2]/P0001  & n13569 ;
  assign n29040 = ~n29038 & ~n29039 ;
  assign n29041 = n29037 & n29040 ;
  assign n29042 = n29034 & n29041 ;
  assign n29043 = \wishbone_bd_ram_mem0_reg[143][2]/P0001  & n13461 ;
  assign n29044 = \wishbone_bd_ram_mem0_reg[7][2]/P0001  & n13546 ;
  assign n29045 = ~n29043 & ~n29044 ;
  assign n29046 = \wishbone_bd_ram_mem0_reg[142][2]/P0001  & n13448 ;
  assign n29047 = \wishbone_bd_ram_mem0_reg[237][2]/P0001  & n13924 ;
  assign n29048 = ~n29046 & ~n29047 ;
  assign n29049 = n29045 & n29048 ;
  assign n29050 = \wishbone_bd_ram_mem0_reg[112][2]/P0001  & n13482 ;
  assign n29051 = \wishbone_bd_ram_mem0_reg[245][2]/P0001  & n13877 ;
  assign n29052 = ~n29050 & ~n29051 ;
  assign n29053 = \wishbone_bd_ram_mem0_reg[57][2]/P0001  & n13731 ;
  assign n29054 = \wishbone_bd_ram_mem0_reg[206][2]/P0001  & n13414 ;
  assign n29055 = ~n29053 & ~n29054 ;
  assign n29056 = n29052 & n29055 ;
  assign n29057 = n29049 & n29056 ;
  assign n29058 = n29042 & n29057 ;
  assign n29059 = \wishbone_bd_ram_mem0_reg[214][2]/P0001  & n13938 ;
  assign n29060 = \wishbone_bd_ram_mem0_reg[174][2]/P0001  & n13899 ;
  assign n29061 = ~n29059 & ~n29060 ;
  assign n29062 = \wishbone_bd_ram_mem0_reg[96][2]/P0001  & n13425 ;
  assign n29063 = \wishbone_bd_ram_mem0_reg[189][2]/P0001  & n14001 ;
  assign n29064 = ~n29062 & ~n29063 ;
  assign n29065 = n29061 & n29064 ;
  assign n29066 = \wishbone_bd_ram_mem0_reg[190][2]/P0001  & n13365 ;
  assign n29067 = \wishbone_bd_ram_mem0_reg[140][2]/P0001  & n13287 ;
  assign n29068 = ~n29066 & ~n29067 ;
  assign n29069 = \wishbone_bd_ram_mem0_reg[149][2]/P0001  & n13469 ;
  assign n29070 = \wishbone_bd_ram_mem0_reg[24][2]/P0001  & n13970 ;
  assign n29071 = ~n29069 & ~n29070 ;
  assign n29072 = n29068 & n29071 ;
  assign n29073 = n29065 & n29072 ;
  assign n29074 = \wishbone_bd_ram_mem0_reg[210][2]/P0001  & n13443 ;
  assign n29075 = \wishbone_bd_ram_mem0_reg[47][2]/P0001  & n13436 ;
  assign n29076 = ~n29074 & ~n29075 ;
  assign n29077 = \wishbone_bd_ram_mem0_reg[195][2]/P0001  & n13700 ;
  assign n29078 = \wishbone_bd_ram_mem0_reg[39][2]/P0001  & n13893 ;
  assign n29079 = ~n29077 & ~n29078 ;
  assign n29080 = n29076 & n29079 ;
  assign n29081 = \wishbone_bd_ram_mem0_reg[163][2]/P0001  & n13255 ;
  assign n29082 = \wishbone_bd_ram_mem0_reg[73][2]/P0001  & n13456 ;
  assign n29083 = ~n29081 & ~n29082 ;
  assign n29084 = \wishbone_bd_ram_mem0_reg[64][2]/P0001  & n13904 ;
  assign n29085 = \wishbone_bd_ram_mem0_reg[145][2]/P0001  & n13715 ;
  assign n29086 = ~n29084 & ~n29085 ;
  assign n29087 = n29083 & n29086 ;
  assign n29088 = n29080 & n29087 ;
  assign n29089 = n29073 & n29088 ;
  assign n29090 = n29058 & n29089 ;
  assign n29091 = n29027 & n29090 ;
  assign n29092 = \wishbone_bd_ram_mem0_reg[157][2]/P0001  & n13445 ;
  assign n29093 = \wishbone_bd_ram_mem0_reg[124][2]/P0001  & n14024 ;
  assign n29094 = ~n29092 & ~n29093 ;
  assign n29095 = \wishbone_bd_ram_mem0_reg[113][2]/P0001  & n13882 ;
  assign n29096 = \wishbone_bd_ram_mem0_reg[146][2]/P0001  & n13958 ;
  assign n29097 = ~n29095 & ~n29096 ;
  assign n29098 = n29094 & n29097 ;
  assign n29099 = \wishbone_bd_ram_mem0_reg[212][2]/P0001  & n13634 ;
  assign n29100 = \wishbone_bd_ram_mem0_reg[25][2]/P0001  & n13742 ;
  assign n29101 = ~n29099 & ~n29100 ;
  assign n29102 = \wishbone_bd_ram_mem0_reg[85][2]/P0001  & n13784 ;
  assign n29103 = \wishbone_bd_ram_mem0_reg[72][2]/P0001  & n13582 ;
  assign n29104 = ~n29102 & ~n29103 ;
  assign n29105 = n29101 & n29104 ;
  assign n29106 = n29098 & n29105 ;
  assign n29107 = \wishbone_bd_ram_mem0_reg[196][2]/P0001  & n13977 ;
  assign n29108 = \wishbone_bd_ram_mem0_reg[100][2]/P0001  & n13401 ;
  assign n29109 = ~n29107 & ~n29108 ;
  assign n29110 = \wishbone_bd_ram_mem0_reg[198][2]/P0001  & n13592 ;
  assign n29111 = \wishbone_bd_ram_mem0_reg[224][2]/P0001  & n13433 ;
  assign n29112 = ~n29110 & ~n29111 ;
  assign n29113 = n29109 & n29112 ;
  assign n29114 = \wishbone_bd_ram_mem0_reg[188][2]/P0001  & n13407 ;
  assign n29115 = \wishbone_bd_ram_mem0_reg[26][2]/P0001  & n13521 ;
  assign n29116 = ~n29114 & ~n29115 ;
  assign n29117 = \wishbone_bd_ram_mem0_reg[108][2]/P0001  & n13814 ;
  assign n29118 = \wishbone_bd_ram_mem0_reg[228][2]/P0001  & n13497 ;
  assign n29119 = ~n29117 & ~n29118 ;
  assign n29120 = n29116 & n29119 ;
  assign n29121 = n29113 & n29120 ;
  assign n29122 = n29106 & n29121 ;
  assign n29123 = \wishbone_bd_ram_mem0_reg[80][2]/P0001  & n13516 ;
  assign n29124 = \wishbone_bd_ram_mem0_reg[235][2]/P0001  & n13518 ;
  assign n29125 = ~n29123 & ~n29124 ;
  assign n29126 = \wishbone_bd_ram_mem0_reg[135][2]/P0001  & n13672 ;
  assign n29127 = \wishbone_bd_ram_mem0_reg[31][2]/P0001  & n13758 ;
  assign n29128 = ~n29126 & ~n29127 ;
  assign n29129 = n29125 & n29128 ;
  assign n29130 = \wishbone_bd_ram_mem0_reg[8][2]/P0001  & n13459 ;
  assign n29131 = \wishbone_bd_ram_mem0_reg[60][2]/P0001  & n13790 ;
  assign n29132 = ~n29130 & ~n29131 ;
  assign n29133 = \wishbone_bd_ram_mem0_reg[42][2]/P0001  & n13341 ;
  assign n29134 = \wishbone_bd_ram_mem0_reg[95][2]/P0001  & n13317 ;
  assign n29135 = ~n29133 & ~n29134 ;
  assign n29136 = n29132 & n29135 ;
  assign n29137 = n29129 & n29136 ;
  assign n29138 = \wishbone_bd_ram_mem0_reg[16][2]/P0001  & n13695 ;
  assign n29139 = \wishbone_bd_ram_mem0_reg[219][2]/P0001  & n13577 ;
  assign n29140 = ~n29138 & ~n29139 ;
  assign n29141 = \wishbone_bd_ram_mem0_reg[38][2]/P0001  & n13828 ;
  assign n29142 = \wishbone_bd_ram_mem0_reg[23][2]/P0001  & n13857 ;
  assign n29143 = ~n29141 & ~n29142 ;
  assign n29144 = n29140 & n29143 ;
  assign n29145 = \wishbone_bd_ram_mem0_reg[121][2]/P0001  & n13983 ;
  assign n29146 = \wishbone_bd_ram_mem0_reg[246][2]/P0001  & n13981 ;
  assign n29147 = ~n29145 & ~n29146 ;
  assign n29148 = \wishbone_bd_ram_mem0_reg[200][2]/P0001  & n13922 ;
  assign n29149 = \wishbone_bd_ram_mem0_reg[136][2]/P0001  & n13963 ;
  assign n29150 = ~n29148 & ~n29149 ;
  assign n29151 = n29147 & n29150 ;
  assign n29152 = n29144 & n29151 ;
  assign n29153 = n29137 & n29152 ;
  assign n29154 = n29122 & n29153 ;
  assign n29155 = \wishbone_bd_ram_mem0_reg[76][2]/P0001  & n13831 ;
  assign n29156 = \wishbone_bd_ram_mem0_reg[132][2]/P0001  & n13927 ;
  assign n29157 = ~n29155 & ~n29156 ;
  assign n29158 = \wishbone_bd_ram_mem0_reg[102][2]/P0001  & n13534 ;
  assign n29159 = \wishbone_bd_ram_mem0_reg[114][2]/P0001  & n13763 ;
  assign n29160 = ~n29158 & ~n29159 ;
  assign n29161 = n29157 & n29160 ;
  assign n29162 = \wishbone_bd_ram_mem0_reg[242][2]/P0001  & n13383 ;
  assign n29163 = \wishbone_bd_ram_mem0_reg[238][2]/P0001  & n13819 ;
  assign n29164 = ~n29162 & ~n29163 ;
  assign n29165 = \wishbone_bd_ram_mem0_reg[223][2]/P0001  & n13335 ;
  assign n29166 = \wishbone_bd_ram_mem0_reg[86][2]/P0001  & n13485 ;
  assign n29167 = ~n29165 & ~n29166 ;
  assign n29168 = n29164 & n29167 ;
  assign n29169 = n29161 & n29168 ;
  assign n29170 = \wishbone_bd_ram_mem0_reg[221][2]/P0001  & n13641 ;
  assign n29171 = \wishbone_bd_ram_mem0_reg[131][2]/P0001  & n13358 ;
  assign n29172 = ~n29170 & ~n29171 ;
  assign n29173 = \wishbone_bd_ram_mem0_reg[222][2]/P0001  & n13721 ;
  assign n29174 = \wishbone_bd_ram_mem0_reg[255][2]/P0001  & n13952 ;
  assign n29175 = ~n29173 & ~n29174 ;
  assign n29176 = n29172 & n29175 ;
  assign n29177 = \wishbone_bd_ram_mem0_reg[192][2]/P0001  & n13390 ;
  assign n29178 = \wishbone_bd_ram_mem0_reg[62][2]/P0001  & n13529 ;
  assign n29179 = ~n29177 & ~n29178 ;
  assign n29180 = \wishbone_bd_ram_mem0_reg[137][2]/P0001  & n13808 ;
  assign n29181 = \wishbone_bd_ram_mem0_reg[93][2]/P0001  & n13891 ;
  assign n29182 = ~n29180 & ~n29181 ;
  assign n29183 = n29179 & n29182 ;
  assign n29184 = n29176 & n29183 ;
  assign n29185 = n29169 & n29184 ;
  assign n29186 = \wishbone_bd_ram_mem0_reg[3][2]/P0001  & n13354 ;
  assign n29187 = \wishbone_bd_ram_mem0_reg[10][2]/P0001  & n13837 ;
  assign n29188 = ~n29186 & ~n29187 ;
  assign n29189 = \wishbone_bd_ram_mem0_reg[12][2]/P0001  & n13733 ;
  assign n29190 = \wishbone_bd_ram_mem0_reg[109][2]/P0001  & n13306 ;
  assign n29191 = ~n29189 & ~n29190 ;
  assign n29192 = n29188 & n29191 ;
  assign n29193 = \wishbone_bd_ram_mem0_reg[150][2]/P0001  & n13666 ;
  assign n29194 = \wishbone_bd_ram_mem0_reg[253][2]/P0001  & n13708 ;
  assign n29195 = ~n29193 & ~n29194 ;
  assign n29196 = \wishbone_bd_ram_mem0_reg[159][2]/P0001  & n13627 ;
  assign n29197 = \wishbone_bd_ram_mem0_reg[138][2]/P0001  & n13398 ;
  assign n29198 = ~n29196 & ~n29197 ;
  assign n29199 = n29195 & n29198 ;
  assign n29200 = n29192 & n29199 ;
  assign n29201 = \wishbone_bd_ram_mem0_reg[175][2]/P0001  & n13674 ;
  assign n29202 = \wishbone_bd_ram_mem0_reg[229][2]/P0001  & n13552 ;
  assign n29203 = ~n29201 & ~n29202 ;
  assign n29204 = \wishbone_bd_ram_mem0_reg[51][2]/P0001  & n13880 ;
  assign n29205 = \wishbone_bd_ram_mem0_reg[250][2]/P0001  & n13677 ;
  assign n29206 = ~n29204 & ~n29205 ;
  assign n29207 = n29203 & n29206 ;
  assign n29208 = \wishbone_bd_ram_mem0_reg[191][2]/P0001  & n14012 ;
  assign n29209 = \wishbone_bd_ram_mem0_reg[202][2]/P0001  & n13268 ;
  assign n29210 = ~n29208 & ~n29209 ;
  assign n29211 = \wishbone_bd_ram_mem0_reg[180][2]/P0001  & n13650 ;
  assign n29212 = \wishbone_bd_ram_mem0_reg[119][2]/P0001  & n14033 ;
  assign n29213 = ~n29211 & ~n29212 ;
  assign n29214 = n29210 & n29213 ;
  assign n29215 = n29207 & n29214 ;
  assign n29216 = n29200 & n29215 ;
  assign n29217 = n29185 & n29216 ;
  assign n29218 = n29154 & n29217 ;
  assign n29219 = n29091 & n29218 ;
  assign n29220 = \wishbone_bd_ram_mem0_reg[9][2]/P0001  & n13580 ;
  assign n29221 = \wishbone_bd_ram_mem0_reg[69][2]/P0001  & n13487 ;
  assign n29222 = ~n29220 & ~n29221 ;
  assign n29223 = \wishbone_bd_ram_mem0_reg[218][2]/P0001  & n13792 ;
  assign n29224 = \wishbone_bd_ram_mem0_reg[225][2]/P0001  & n13719 ;
  assign n29225 = ~n29223 & ~n29224 ;
  assign n29226 = n29222 & n29225 ;
  assign n29227 = \wishbone_bd_ram_mem0_reg[20][2]/P0001  & n13839 ;
  assign n29228 = \wishbone_bd_ram_mem0_reg[67][2]/P0001  & n13663 ;
  assign n29229 = ~n29227 & ~n29228 ;
  assign n29230 = \wishbone_bd_ram_mem0_reg[181][2]/P0001  & n13587 ;
  assign n29231 = \wishbone_bd_ram_mem0_reg[155][2]/P0001  & n13738 ;
  assign n29232 = ~n29230 & ~n29231 ;
  assign n29233 = n29229 & n29232 ;
  assign n29234 = n29226 & n29233 ;
  assign n29235 = \wishbone_bd_ram_mem0_reg[144][2]/P0001  & n13508 ;
  assign n29236 = \wishbone_bd_ram_mem0_reg[33][2]/P0001  & n13933 ;
  assign n29237 = ~n29235 & ~n29236 ;
  assign n29238 = \wishbone_bd_ram_mem0_reg[209][2]/P0001  & n13689 ;
  assign n29239 = \wishbone_bd_ram_mem0_reg[165][2]/P0001  & n14028 ;
  assign n29240 = ~n29238 & ~n29239 ;
  assign n29241 = n29237 & n29240 ;
  assign n29242 = \wishbone_bd_ram_mem0_reg[128][2]/P0001  & n13652 ;
  assign n29243 = \wishbone_bd_ram_mem0_reg[182][2]/P0001  & n13598 ;
  assign n29244 = ~n29242 & ~n29243 ;
  assign n29245 = \wishbone_bd_ram_mem0_reg[158][2]/P0001  & n13294 ;
  assign n29246 = \wishbone_bd_ram_mem0_reg[148][2]/P0001  & n13868 ;
  assign n29247 = ~n29245 & ~n29246 ;
  assign n29248 = n29244 & n29247 ;
  assign n29249 = n29241 & n29248 ;
  assign n29250 = n29234 & n29249 ;
  assign n29251 = \wishbone_bd_ram_mem0_reg[252][2]/P0001  & n13986 ;
  assign n29252 = \wishbone_bd_ram_mem0_reg[152][2]/P0001  & n13912 ;
  assign n29253 = ~n29251 & ~n29252 ;
  assign n29254 = \wishbone_bd_ram_mem0_reg[5][2]/P0001  & n13243 ;
  assign n29255 = \wishbone_bd_ram_mem0_reg[120][2]/P0001  & n13550 ;
  assign n29256 = ~n29254 & ~n29255 ;
  assign n29257 = n29253 & n29256 ;
  assign n29258 = \wishbone_bd_ram_mem0_reg[226][2]/P0001  & n13668 ;
  assign n29259 = \wishbone_bd_ram_mem0_reg[139][2]/P0001  & n13566 ;
  assign n29260 = ~n29258 & ~n29259 ;
  assign n29261 = \wishbone_bd_ram_mem0_reg[105][2]/P0001  & n13503 ;
  assign n29262 = \wishbone_bd_ram_mem0_reg[162][2]/P0001  & n13726 ;
  assign n29263 = ~n29261 & ~n29262 ;
  assign n29264 = n29260 & n29263 ;
  assign n29265 = n29257 & n29264 ;
  assign n29266 = \wishbone_bd_ram_mem0_reg[161][2]/P0001  & n13505 ;
  assign n29267 = \wishbone_bd_ram_mem0_reg[40][2]/P0001  & n13661 ;
  assign n29268 = ~n29266 & ~n29267 ;
  assign n29269 = \wishbone_bd_ram_mem0_reg[14][2]/P0001  & n13972 ;
  assign n29270 = \wishbone_bd_ram_mem0_reg[6][2]/P0001  & n13915 ;
  assign n29271 = ~n29269 & ~n29270 ;
  assign n29272 = n29268 & n29271 ;
  assign n29273 = \wishbone_bd_ram_mem0_reg[66][2]/P0001  & n13603 ;
  assign n29274 = \wishbone_bd_ram_mem0_reg[55][2]/P0001  & n13618 ;
  assign n29275 = ~n29273 & ~n29274 ;
  assign n29276 = \wishbone_bd_ram_mem0_reg[15][2]/P0001  & n13797 ;
  assign n29277 = \wishbone_bd_ram_mem0_reg[116][2]/P0001  & n13865 ;
  assign n29278 = ~n29276 & ~n29277 ;
  assign n29279 = n29275 & n29278 ;
  assign n29280 = n29272 & n29279 ;
  assign n29281 = n29265 & n29280 ;
  assign n29282 = n29250 & n29281 ;
  assign n29283 = \wishbone_bd_ram_mem0_reg[172][2]/P0001  & n13377 ;
  assign n29284 = \wishbone_bd_ram_mem0_reg[83][2]/P0001  & n13454 ;
  assign n29285 = ~n29283 & ~n29284 ;
  assign n29286 = \wishbone_bd_ram_mem0_reg[21][2]/P0001  & n13438 ;
  assign n29287 = \wishbone_bd_ram_mem0_reg[127][2]/P0001  & n13803 ;
  assign n29288 = ~n29286 & ~n29287 ;
  assign n29289 = n29285 & n29288 ;
  assign n29290 = \wishbone_bd_ram_mem0_reg[217][2]/P0001  & n13767 ;
  assign n29291 = \wishbone_bd_ram_mem0_reg[147][2]/P0001  & n13702 ;
  assign n29292 = ~n29290 & ~n29291 ;
  assign n29293 = \wishbone_bd_ram_mem0_reg[208][2]/P0001  & n14010 ;
  assign n29294 = \wishbone_bd_ram_mem0_reg[115][2]/P0001  & n13747 ;
  assign n29295 = ~n29293 & ~n29294 ;
  assign n29296 = n29292 & n29295 ;
  assign n29297 = n29289 & n29296 ;
  assign n29298 = \wishbone_bd_ram_mem0_reg[68][2]/P0001  & n13379 ;
  assign n29299 = \wishbone_bd_ram_mem0_reg[176][2]/P0001  & n13262 ;
  assign n29300 = ~n29298 & ~n29299 ;
  assign n29301 = \wishbone_bd_ram_mem0_reg[78][2]/P0001  & n13277 ;
  assign n29302 = \wishbone_bd_ram_mem0_reg[151][2]/P0001  & n13697 ;
  assign n29303 = ~n29301 & ~n29302 ;
  assign n29304 = n29300 & n29303 ;
  assign n29305 = \wishbone_bd_ram_mem0_reg[141][2]/P0001  & n13852 ;
  assign n29306 = \wishbone_bd_ram_mem0_reg[54][2]/P0001  & n13622 ;
  assign n29307 = ~n29305 & ~n29306 ;
  assign n29308 = \wishbone_bd_ram_mem0_reg[81][2]/P0001  & n13409 ;
  assign n29309 = \wishbone_bd_ram_mem0_reg[22][2]/P0001  & n13744 ;
  assign n29310 = ~n29308 & ~n29309 ;
  assign n29311 = n29307 & n29310 ;
  assign n29312 = n29304 & n29311 ;
  assign n29313 = n29297 & n29312 ;
  assign n29314 = \wishbone_bd_ram_mem0_reg[126][2]/P0001  & n13786 ;
  assign n29315 = \wishbone_bd_ram_mem0_reg[211][2]/P0001  & n13805 ;
  assign n29316 = ~n29314 & ~n29315 ;
  assign n29317 = \wishbone_bd_ram_mem0_reg[63][2]/P0001  & n13327 ;
  assign n29318 = \wishbone_bd_ram_mem0_reg[239][2]/P0001  & n13349 ;
  assign n29319 = ~n29317 & ~n29318 ;
  assign n29320 = n29316 & n29319 ;
  assign n29321 = \wishbone_bd_ram_mem0_reg[17][2]/P0001  & n13324 ;
  assign n29322 = \wishbone_bd_ram_mem0_reg[205][2]/P0001  & n13947 ;
  assign n29323 = ~n29321 & ~n29322 ;
  assign n29324 = \wishbone_bd_ram_mem0_reg[187][2]/P0001  & n13756 ;
  assign n29325 = \wishbone_bd_ram_mem0_reg[204][2]/P0001  & n13821 ;
  assign n29326 = ~n29324 & ~n29325 ;
  assign n29327 = n29323 & n29326 ;
  assign n29328 = n29320 & n29327 ;
  assign n29329 = \wishbone_bd_ram_mem0_reg[201][2]/P0001  & n13600 ;
  assign n29330 = \wishbone_bd_ram_mem0_reg[173][2]/P0001  & n13360 ;
  assign n29331 = ~n29329 & ~n29330 ;
  assign n29332 = \wishbone_bd_ram_mem0_reg[75][2]/P0001  & n13605 ;
  assign n29333 = \wishbone_bd_ram_mem0_reg[94][2]/P0001  & n13833 ;
  assign n29334 = ~n29332 & ~n29333 ;
  assign n29335 = n29331 & n29334 ;
  assign n29336 = \wishbone_bd_ram_mem0_reg[122][2]/P0001  & n13679 ;
  assign n29337 = \wishbone_bd_ram_mem0_reg[29][2]/P0001  & n13412 ;
  assign n29338 = ~n29336 & ~n29337 ;
  assign n29339 = \wishbone_bd_ram_mem0_reg[65][2]/P0001  & n13842 ;
  assign n29340 = \wishbone_bd_ram_mem0_reg[18][2]/P0001  & n13532 ;
  assign n29341 = ~n29339 & ~n29340 ;
  assign n29342 = n29338 & n29341 ;
  assign n29343 = n29335 & n29342 ;
  assign n29344 = n29328 & n29343 ;
  assign n29345 = n29313 & n29344 ;
  assign n29346 = n29282 & n29345 ;
  assign n29347 = \wishbone_bd_ram_mem0_reg[134][2]/P0001  & n13494 ;
  assign n29348 = \wishbone_bd_ram_mem0_reg[111][2]/P0001  & n13471 ;
  assign n29349 = ~n29347 & ~n29348 ;
  assign n29350 = \wishbone_bd_ram_mem0_reg[129][2]/P0001  & n13629 ;
  assign n29351 = \wishbone_bd_ram_mem0_reg[92][2]/P0001  & n13859 ;
  assign n29352 = ~n29350 & ~n29351 ;
  assign n29353 = n29349 & n29352 ;
  assign n29354 = \wishbone_bd_ram_mem0_reg[107][2]/P0001  & n13476 ;
  assign n29355 = \wishbone_bd_ram_mem0_reg[101][2]/P0001  & n13772 ;
  assign n29356 = ~n29354 & ~n29355 ;
  assign n29357 = \wishbone_bd_ram_mem0_reg[184][2]/P0001  & n13960 ;
  assign n29358 = \wishbone_bd_ram_mem0_reg[215][2]/P0001  & n13901 ;
  assign n29359 = ~n29357 & ~n29358 ;
  assign n29360 = n29356 & n29359 ;
  assign n29361 = n29353 & n29360 ;
  assign n29362 = \wishbone_bd_ram_mem0_reg[99][2]/P0001  & n13996 ;
  assign n29363 = \wishbone_bd_ram_mem0_reg[213][2]/P0001  & n13870 ;
  assign n29364 = ~n29362 & ~n29363 ;
  assign n29365 = \wishbone_bd_ram_mem0_reg[41][2]/P0001  & n14017 ;
  assign n29366 = \wishbone_bd_ram_mem0_reg[220][2]/P0001  & n13965 ;
  assign n29367 = ~n29365 & ~n29366 ;
  assign n29368 = n29364 & n29367 ;
  assign n29369 = \wishbone_bd_ram_mem0_reg[46][2]/P0001  & n13298 ;
  assign n29370 = \wishbone_bd_ram_mem0_reg[4][2]/P0001  & n13527 ;
  assign n29371 = ~n29369 & ~n29370 ;
  assign n29372 = \wishbone_bd_ram_mem0_reg[168][2]/P0001  & n13795 ;
  assign n29373 = \wishbone_bd_ram_mem0_reg[56][2]/P0001  & n13611 ;
  assign n29374 = ~n29372 & ~n29373 ;
  assign n29375 = n29371 & n29374 ;
  assign n29376 = n29368 & n29375 ;
  assign n29377 = n29361 & n29376 ;
  assign n29378 = \wishbone_bd_ram_mem0_reg[89][2]/P0001  & n13910 ;
  assign n29379 = \wishbone_bd_ram_mem0_reg[74][2]/P0001  & n13564 ;
  assign n29380 = ~n29378 & ~n29379 ;
  assign n29381 = \wishbone_bd_ram_mem0_reg[203][2]/P0001  & n13816 ;
  assign n29382 = \wishbone_bd_ram_mem0_reg[90][2]/P0001  & n13906 ;
  assign n29383 = ~n29381 & ~n29382 ;
  assign n29384 = n29380 & n29383 ;
  assign n29385 = \wishbone_bd_ram_mem0_reg[171][2]/P0001  & n13422 ;
  assign n29386 = \wishbone_bd_ram_mem0_reg[156][2]/P0001  & n13769 ;
  assign n29387 = ~n29385 & ~n29386 ;
  assign n29388 = \wishbone_bd_ram_mem0_reg[32][2]/P0001  & n13736 ;
  assign n29389 = \wishbone_bd_ram_mem0_reg[35][2]/P0001  & n13523 ;
  assign n29390 = ~n29388 & ~n29389 ;
  assign n29391 = n29387 & n29390 ;
  assign n29392 = n29384 & n29391 ;
  assign n29393 = \wishbone_bd_ram_mem0_reg[185][2]/P0001  & n13372 ;
  assign n29394 = \wishbone_bd_ram_mem0_reg[110][2]/P0001  & n14030 ;
  assign n29395 = ~n29393 & ~n29394 ;
  assign n29396 = \wishbone_bd_ram_mem0_reg[232][2]/P0001  & n13510 ;
  assign n29397 = \wishbone_bd_ram_mem0_reg[61][2]/P0001  & n13544 ;
  assign n29398 = ~n29396 & ~n29397 ;
  assign n29399 = n29395 & n29398 ;
  assign n29400 = \wishbone_bd_ram_mem0_reg[27][2]/P0001  & n13251 ;
  assign n29401 = \wishbone_bd_ram_mem0_reg[77][2]/P0001  & n13935 ;
  assign n29402 = ~n29400 & ~n29401 ;
  assign n29403 = \wishbone_bd_ram_mem0_reg[216][2]/P0001  & n14005 ;
  assign n29404 = \wishbone_bd_ram_mem0_reg[167][2]/P0001  & n13940 ;
  assign n29405 = ~n29403 & ~n29404 ;
  assign n29406 = n29402 & n29405 ;
  assign n29407 = n29399 & n29406 ;
  assign n29408 = n29392 & n29407 ;
  assign n29409 = n29377 & n29408 ;
  assign n29410 = \wishbone_bd_ram_mem0_reg[247][2]/P0001  & n13571 ;
  assign n29411 = \wishbone_bd_ram_mem0_reg[58][2]/P0001  & n13949 ;
  assign n29412 = ~n29410 & ~n29411 ;
  assign n29413 = \wishbone_bd_ram_mem0_reg[197][2]/P0001  & n13594 ;
  assign n29414 = \wishbone_bd_ram_mem0_reg[234][2]/P0001  & n13781 ;
  assign n29415 = ~n29413 & ~n29414 ;
  assign n29416 = n29412 & n29415 ;
  assign n29417 = \wishbone_bd_ram_mem0_reg[19][2]/P0001  & n13886 ;
  assign n29418 = \wishbone_bd_ram_mem0_reg[37][2]/P0001  & n13710 ;
  assign n29419 = ~n29417 & ~n29418 ;
  assign n29420 = \wishbone_bd_ram_mem0_reg[123][2]/P0001  & n13749 ;
  assign n29421 = \wishbone_bd_ram_mem0_reg[244][2]/P0001  & n13474 ;
  assign n29422 = ~n29420 & ~n29421 ;
  assign n29423 = n29419 & n29422 ;
  assign n29424 = n29416 & n29423 ;
  assign n29425 = \wishbone_bd_ram_mem0_reg[79][2]/P0001  & n13779 ;
  assign n29426 = \wishbone_bd_ram_mem0_reg[71][2]/P0001  & n13636 ;
  assign n29427 = ~n29425 & ~n29426 ;
  assign n29428 = \wishbone_bd_ram_mem0_reg[30][2]/P0001  & n13713 ;
  assign n29429 = \wishbone_bd_ram_mem0_reg[133][2]/P0001  & n13492 ;
  assign n29430 = ~n29428 & ~n29429 ;
  assign n29431 = n29427 & n29430 ;
  assign n29432 = \wishbone_bd_ram_mem0_reg[254][2]/P0001  & n13283 ;
  assign n29433 = \wishbone_bd_ram_mem0_reg[230][2]/P0001  & n13994 ;
  assign n29434 = ~n29432 & ~n29433 ;
  assign n29435 = \wishbone_bd_ram_mem0_reg[227][2]/P0001  & n13388 ;
  assign n29436 = \wishbone_bd_ram_mem0_reg[52][2]/P0001  & n13988 ;
  assign n29437 = ~n29435 & ~n29436 ;
  assign n29438 = n29434 & n29437 ;
  assign n29439 = n29431 & n29438 ;
  assign n29440 = n29424 & n29439 ;
  assign n29441 = \wishbone_bd_ram_mem0_reg[125][2]/P0001  & n13396 ;
  assign n29442 = \wishbone_bd_ram_mem0_reg[45][2]/P0001  & n13420 ;
  assign n29443 = ~n29441 & ~n29442 ;
  assign n29444 = \wishbone_bd_ram_mem0_reg[106][2]/P0001  & n13555 ;
  assign n29445 = \wishbone_bd_ram_mem0_reg[130][2]/P0001  & n13427 ;
  assign n29446 = ~n29444 & ~n29445 ;
  assign n29447 = n29443 & n29446 ;
  assign n29448 = \wishbone_bd_ram_mem0_reg[53][2]/P0001  & n13875 ;
  assign n29449 = \wishbone_bd_ram_mem0_reg[49][2]/P0001  & n13929 ;
  assign n29450 = ~n29448 & ~n29449 ;
  assign n29451 = \wishbone_bd_ram_mem0_reg[117][2]/P0001  & n13557 ;
  assign n29452 = \wishbone_bd_ram_mem0_reg[177][2]/P0001  & n13863 ;
  assign n29453 = ~n29451 & ~n29452 ;
  assign n29454 = n29450 & n29453 ;
  assign n29455 = n29447 & n29454 ;
  assign n29456 = \wishbone_bd_ram_mem0_reg[36][2]/P0001  & n13639 ;
  assign n29457 = \wishbone_bd_ram_mem0_reg[251][2]/P0001  & n14019 ;
  assign n29458 = ~n29456 & ~n29457 ;
  assign n29459 = \wishbone_bd_ram_mem0_reg[241][2]/P0001  & n13854 ;
  assign n29460 = \wishbone_bd_ram_mem0_reg[97][2]/P0001  & n13724 ;
  assign n29461 = ~n29459 & ~n29460 ;
  assign n29462 = n29458 & n29461 ;
  assign n29463 = \wishbone_bd_ram_mem0_reg[48][2]/P0001  & n13917 ;
  assign n29464 = \wishbone_bd_ram_mem0_reg[154][2]/P0001  & n13403 ;
  assign n29465 = ~n29463 & ~n29464 ;
  assign n29466 = \wishbone_bd_ram_mem0_reg[0][2]/P0001  & n13539 ;
  assign n29467 = \wishbone_bd_ram_mem0_reg[243][2]/P0001  & n13575 ;
  assign n29468 = ~n29466 & ~n29467 ;
  assign n29469 = n29465 & n29468 ;
  assign n29470 = n29462 & n29469 ;
  assign n29471 = n29455 & n29470 ;
  assign n29472 = n29440 & n29471 ;
  assign n29473 = n29409 & n29472 ;
  assign n29474 = n29346 & n29473 ;
  assign n29475 = n29219 & n29474 ;
  assign n29476 = ~wb_rst_i_pad & ~n28963 ;
  assign n29477 = ~n29475 & n29476 ;
  assign n29478 = ~n28964 & ~n29477 ;
  assign n29479 = \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  & n23737 ;
  assign n29480 = \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  & n28956 ;
  assign n29481 = \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131  & n25088 ;
  assign n29482 = ~n29480 & ~n29481 ;
  assign n29483 = \ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131  & n25084 ;
  assign n29484 = \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131  & n25079 ;
  assign n29485 = ~n29483 & ~n29484 ;
  assign n29486 = n29482 & n29485 ;
  assign n29487 = \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131  & n23802 ;
  assign n29488 = \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  & n23751 ;
  assign n29489 = n23747 & n29488 ;
  assign n29490 = ~n29487 & ~n29489 ;
  assign n29491 = \miim1_shftrg_LinkFail_reg/NET0131  & n28945 ;
  assign n29492 = \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131  & n23813 ;
  assign n29493 = ~n29491 & ~n29492 ;
  assign n29494 = n29490 & n29493 ;
  assign n29495 = n29486 & n29494 ;
  assign n29496 = ~n29479 & n29495 ;
  assign n29497 = \ethreg1_IPGT_0_DataOut_reg[0]/NET0131  & n25090 ;
  assign n29498 = \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  & n23751 ;
  assign n29499 = n23741 & n29498 ;
  assign n29500 = ~n29497 & ~n29499 ;
  assign n29501 = \ethreg1_IPGR1_0_DataOut_reg[0]/NET0131  & n25069 ;
  assign n29502 = \ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131  & n23782 ;
  assign n29503 = ~n29501 & ~n29502 ;
  assign n29504 = n29500 & n29503 ;
  assign n29505 = n23730 & n29504 ;
  assign n29506 = \ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131  & n23743 ;
  assign n29507 = n23747 & n29506 ;
  assign n29508 = \ethreg1_MODER_0_DataOut_reg[0]/NET0131  & n23808 ;
  assign n29509 = ~n29507 & ~n29508 ;
  assign n29510 = \ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131  & n23743 ;
  assign n29511 = n23741 & n29510 ;
  assign n29512 = \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131  & n25082 ;
  assign n29513 = ~n29511 & ~n29512 ;
  assign n29514 = n29509 & n29513 ;
  assign n29515 = \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131  & n23794 ;
  assign n29516 = n23741 & n29515 ;
  assign n29517 = \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  & n28939 ;
  assign n29518 = ~n29516 & ~n29517 ;
  assign n29519 = \ethreg1_irq_txb_reg/NET0131  & n25064 ;
  assign n29520 = \ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131  & n28948 ;
  assign n29521 = ~n29519 & ~n29520 ;
  assign n29522 = n29518 & n29521 ;
  assign n29523 = n29514 & n29522 ;
  assign n29524 = n29505 & n29523 ;
  assign n29525 = n29496 & n29524 ;
  assign n29526 = n23730 & ~n29525 ;
  assign n29527 = ~wb_rst_i_pad & ~n29525 ;
  assign n29528 = ~n24902 & n29527 ;
  assign n29529 = ~n29526 & ~n29528 ;
  assign n29530 = \ethreg1_irq_txe_reg/NET0131  & n25064 ;
  assign n29531 = \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  & n28939 ;
  assign n29532 = ~n29530 & ~n29531 ;
  assign n29533 = ~\miim1_InProgress_reg/NET0131  & ~\miim1_Nvalid_reg/NET0131  ;
  assign n29534 = ~\miim1_RStatStart_reg/NET0131  & ~\miim1_SyncStatMdcEn_reg/NET0131  ;
  assign n29535 = n29533 & n29534 ;
  assign n29536 = ~\miim1_EndBusy_reg/NET0131  & ~\miim1_WCtrlDataStart_reg/NET0131  ;
  assign n29537 = ~\ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131  & ~\miim1_InProgress_q3_reg/NET0131  ;
  assign n29538 = n29536 & n29537 ;
  assign n29539 = n29535 & n29538 ;
  assign n29540 = n28945 & ~n29539 ;
  assign n29541 = \ethreg1_MODER_0_DataOut_reg[1]/NET0131  & n23808 ;
  assign n29542 = ~n29540 & ~n29541 ;
  assign n29543 = n29532 & n29542 ;
  assign n29544 = \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131  & n25069 ;
  assign n29545 = \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131  & n25079 ;
  assign n29546 = ~n29544 & ~n29545 ;
  assign n29547 = \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  & n23737 ;
  assign n29548 = \ethreg1_IPGT_0_DataOut_reg[1]/NET0131  & n25090 ;
  assign n29549 = ~n29547 & ~n29548 ;
  assign n29550 = n29546 & n29549 ;
  assign n29551 = n29543 & n29550 ;
  assign n29552 = \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131  & n25088 ;
  assign n29553 = \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  & n23751 ;
  assign n29554 = n23741 & n29553 ;
  assign n29555 = ~n29552 & ~n29554 ;
  assign n29556 = \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131  & n25082 ;
  assign n29557 = \ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131  & n23743 ;
  assign n29558 = n23741 & n29557 ;
  assign n29559 = ~n29556 & ~n29558 ;
  assign n29560 = n29555 & n29559 ;
  assign n29561 = ~\wb_adr_i[6]_pad  & n23746 ;
  assign n29562 = n23781 & n29561 ;
  assign n29563 = \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131  & n29562 ;
  assign n29564 = n23730 & ~n29563 ;
  assign n29565 = n29560 & n29564 ;
  assign n29566 = \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131  & n23802 ;
  assign n29567 = \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  & n23751 ;
  assign n29568 = n23747 & n29567 ;
  assign n29569 = ~n29566 & ~n29568 ;
  assign n29570 = \ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131  & n23813 ;
  assign n29571 = \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  & n28956 ;
  assign n29572 = ~n29570 & ~n29571 ;
  assign n29573 = n29569 & n29572 ;
  assign n29574 = \ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131  & n23743 ;
  assign n29575 = n23747 & n29574 ;
  assign n29576 = \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131  & n23794 ;
  assign n29577 = n23741 & n29576 ;
  assign n29578 = ~n29575 & ~n29577 ;
  assign n29579 = \ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131  & n23782 ;
  assign n29580 = \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  & n25084 ;
  assign n29581 = ~n29579 & ~n29580 ;
  assign n29582 = n29578 & n29581 ;
  assign n29583 = n29573 & n29582 ;
  assign n29584 = n29565 & n29583 ;
  assign n29585 = n29551 & n29584 ;
  assign n29586 = n23730 & ~n29585 ;
  assign n29587 = ~wb_rst_i_pad & ~n29585 ;
  assign n29588 = ~n16820 & n29587 ;
  assign n29589 = ~n29586 & ~n29588 ;
  assign n29590 = n14057 & ~n17918 ;
  assign n29591 = \wishbone_TxLength_reg[7]/NET0131  & ~n29590 ;
  assign n29592 = ~n15700 & ~n29591 ;
  assign n29593 = n19277 & ~n29592 ;
  assign n29594 = ~n23203 & ~n29593 ;
  assign n29595 = \wishbone_TxLength_reg[5]/NET0131  & ~n14049 ;
  assign n29596 = ~n14046 & n29595 ;
  assign n29597 = \wishbone_TxLength_reg[5]/NET0131  & ~n14055 ;
  assign n29598 = ~n24357 & ~n29597 ;
  assign n29599 = ~\wishbone_TxLength_reg[5]/NET0131  & \wishbone_TxPointerLSB_rst_reg[0]/NET0131  ;
  assign n29600 = n17365 & n29599 ;
  assign n29601 = ~\wishbone_TxPointerLSB_rst_reg[1]/NET0131  & ~n29600 ;
  assign n29602 = ~n29598 & n29601 ;
  assign n29603 = \wishbone_TxLength_reg[5]/NET0131  & n17367 ;
  assign n29604 = n17365 & n29603 ;
  assign n29605 = ~n29602 & ~n29604 ;
  assign n29606 = n17372 & n24357 ;
  assign n29607 = n17371 & n29606 ;
  assign n29608 = \wishbone_TxLength_reg[5]/NET0131  & n17371 ;
  assign n29609 = ~n17375 & n29608 ;
  assign n29610 = ~n29607 & ~n29609 ;
  assign n29611 = \wishbone_TxLength_reg[5]/NET0131  & n17381 ;
  assign n29612 = ~n17383 & n29611 ;
  assign n29613 = ~\wishbone_TxLength_reg[5]/NET0131  & n17381 ;
  assign n29614 = n17383 & n29613 ;
  assign n29615 = ~n29612 & ~n29614 ;
  assign n29616 = n29610 & n29615 ;
  assign n29617 = n29605 & n29616 ;
  assign n29618 = ~n14046 & n17360 ;
  assign n29619 = ~n29617 & n29618 ;
  assign n29620 = ~n29596 & ~n29619 ;
  assign n29621 = ~n22689 & n29620 ;
  assign n29622 = \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131  & n23794 ;
  assign n29623 = n23741 & n29622 ;
  assign n29624 = \ethreg1_MODER_2_DataOut_reg[0]/NET0131  & n23808 ;
  assign n29625 = \ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131  & n23743 ;
  assign n29626 = n23741 & n29625 ;
  assign n29627 = ~n29624 & ~n29626 ;
  assign n29628 = ~n29623 & n29627 ;
  assign n29629 = \ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131  & n23743 ;
  assign n29630 = n23747 & n29629 ;
  assign n29631 = \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  & n23751 ;
  assign n29632 = n23741 & n29631 ;
  assign n29633 = ~n29630 & ~n29632 ;
  assign n29634 = \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131  & n25059 ;
  assign n29635 = \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  & n23737 ;
  assign n29636 = ~n29634 & ~n29635 ;
  assign n29637 = n29633 & n29636 ;
  assign n29638 = n29628 & n29637 ;
  assign n29639 = n23730 & ~n29638 ;
  assign n29640 = ~wb_rst_i_pad & ~n23730 ;
  assign n29641 = ~n19794 & n29640 ;
  assign n29642 = ~n29639 & ~n29641 ;
  assign n29643 = \ethreg1_IPGT_0_DataOut_reg[6]/NET0131  & n25090 ;
  assign n29644 = \ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131  & n23743 ;
  assign n29645 = n23747 & n29644 ;
  assign n29646 = ~n29643 & ~n29645 ;
  assign n29647 = \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131  & n25082 ;
  assign n29648 = \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  & n25084 ;
  assign n29649 = ~n29647 & ~n29648 ;
  assign n29650 = n29646 & n29649 ;
  assign n29651 = n23730 & n29650 ;
  assign n29652 = \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131  & n25069 ;
  assign n29653 = \ethreg1_MODER_0_DataOut_reg[6]/NET0131  & n23808 ;
  assign n29654 = ~n29652 & ~n29653 ;
  assign n29655 = \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131  & n25088 ;
  assign n29656 = \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  & n23751 ;
  assign n29657 = n23747 & n29656 ;
  assign n29658 = ~n29655 & ~n29657 ;
  assign n29659 = n29654 & n29658 ;
  assign n29660 = \ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131  & n23743 ;
  assign n29661 = n23741 & n29660 ;
  assign n29662 = \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131  & n25079 ;
  assign n29663 = ~n29661 & ~n29662 ;
  assign n29664 = \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  & n23751 ;
  assign n29665 = n23741 & n29664 ;
  assign n29666 = \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131  & n23794 ;
  assign n29667 = n23741 & n29666 ;
  assign n29668 = ~n29665 & ~n29667 ;
  assign n29669 = n29663 & n29668 ;
  assign n29670 = n29659 & n29669 ;
  assign n29671 = \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131  & n23813 ;
  assign n29672 = \ethreg1_irq_rxc_reg/NET0131  & n25064 ;
  assign n29673 = ~n29671 & ~n29672 ;
  assign n29674 = \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  & n23737 ;
  assign n29675 = \ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131  & n23782 ;
  assign n29676 = ~n29674 & ~n29675 ;
  assign n29677 = n29673 & n29676 ;
  assign n29678 = n29670 & n29677 ;
  assign n29679 = n29651 & n29678 ;
  assign n29680 = n23730 & ~n29679 ;
  assign n29681 = \wishbone_bd_ram_mem0_reg[80][6]/P0001  & n13516 ;
  assign n29682 = \wishbone_bd_ram_mem0_reg[33][6]/P0001  & n13933 ;
  assign n29683 = ~n29681 & ~n29682 ;
  assign n29684 = \wishbone_bd_ram_mem0_reg[21][6]/P0001  & n13438 ;
  assign n29685 = \wishbone_bd_ram_mem0_reg[73][6]/P0001  & n13456 ;
  assign n29686 = ~n29684 & ~n29685 ;
  assign n29687 = n29683 & n29686 ;
  assign n29688 = \wishbone_bd_ram_mem0_reg[210][6]/P0001  & n13443 ;
  assign n29689 = \wishbone_bd_ram_mem0_reg[121][6]/P0001  & n13983 ;
  assign n29690 = ~n29688 & ~n29689 ;
  assign n29691 = \wishbone_bd_ram_mem0_reg[149][6]/P0001  & n13469 ;
  assign n29692 = \wishbone_bd_ram_mem0_reg[183][6]/P0001  & n13645 ;
  assign n29693 = ~n29691 & ~n29692 ;
  assign n29694 = n29690 & n29693 ;
  assign n29695 = n29687 & n29694 ;
  assign n29696 = \wishbone_bd_ram_mem0_reg[249][6]/P0001  & n13431 ;
  assign n29697 = \wishbone_bd_ram_mem0_reg[255][6]/P0001  & n13952 ;
  assign n29698 = ~n29696 & ~n29697 ;
  assign n29699 = \wishbone_bd_ram_mem0_reg[84][6]/P0001  & n13385 ;
  assign n29700 = \wishbone_bd_ram_mem0_reg[237][6]/P0001  & n13924 ;
  assign n29701 = ~n29699 & ~n29700 ;
  assign n29702 = n29698 & n29701 ;
  assign n29703 = \wishbone_bd_ram_mem0_reg[51][6]/P0001  & n13880 ;
  assign n29704 = \wishbone_bd_ram_mem0_reg[252][6]/P0001  & n13986 ;
  assign n29705 = ~n29703 & ~n29704 ;
  assign n29706 = \wishbone_bd_ram_mem0_reg[32][6]/P0001  & n13736 ;
  assign n29707 = \wishbone_bd_ram_mem0_reg[144][6]/P0001  & n13508 ;
  assign n29708 = ~n29706 & ~n29707 ;
  assign n29709 = n29705 & n29708 ;
  assign n29710 = n29702 & n29709 ;
  assign n29711 = n29695 & n29710 ;
  assign n29712 = \wishbone_bd_ram_mem0_reg[89][6]/P0001  & n13910 ;
  assign n29713 = \wishbone_bd_ram_mem0_reg[104][6]/P0001  & n13684 ;
  assign n29714 = ~n29712 & ~n29713 ;
  assign n29715 = \wishbone_bd_ram_mem0_reg[194][6]/P0001  & n13624 ;
  assign n29716 = \wishbone_bd_ram_mem0_reg[92][6]/P0001  & n13859 ;
  assign n29717 = ~n29715 & ~n29716 ;
  assign n29718 = n29714 & n29717 ;
  assign n29719 = \wishbone_bd_ram_mem0_reg[221][6]/P0001  & n13641 ;
  assign n29720 = \wishbone_bd_ram_mem0_reg[127][6]/P0001  & n13803 ;
  assign n29721 = ~n29719 & ~n29720 ;
  assign n29722 = \wishbone_bd_ram_mem0_reg[74][6]/P0001  & n13564 ;
  assign n29723 = \wishbone_bd_ram_mem0_reg[4][6]/P0001  & n13527 ;
  assign n29724 = ~n29722 & ~n29723 ;
  assign n29725 = n29721 & n29724 ;
  assign n29726 = n29718 & n29725 ;
  assign n29727 = \wishbone_bd_ram_mem0_reg[174][6]/P0001  & n13899 ;
  assign n29728 = \wishbone_bd_ram_mem0_reg[178][6]/P0001  & n13301 ;
  assign n29729 = ~n29727 & ~n29728 ;
  assign n29730 = \wishbone_bd_ram_mem0_reg[217][6]/P0001  & n13767 ;
  assign n29731 = \wishbone_bd_ram_mem0_reg[72][6]/P0001  & n13582 ;
  assign n29732 = ~n29730 & ~n29731 ;
  assign n29733 = n29729 & n29732 ;
  assign n29734 = \wishbone_bd_ram_mem0_reg[79][6]/P0001  & n13779 ;
  assign n29735 = \wishbone_bd_ram_mem0_reg[212][6]/P0001  & n13634 ;
  assign n29736 = ~n29734 & ~n29735 ;
  assign n29737 = \wishbone_bd_ram_mem0_reg[151][6]/P0001  & n13697 ;
  assign n29738 = \wishbone_bd_ram_mem0_reg[225][6]/P0001  & n13719 ;
  assign n29739 = ~n29737 & ~n29738 ;
  assign n29740 = n29736 & n29739 ;
  assign n29741 = n29733 & n29740 ;
  assign n29742 = n29726 & n29741 ;
  assign n29743 = n29711 & n29742 ;
  assign n29744 = \wishbone_bd_ram_mem0_reg[197][6]/P0001  & n13594 ;
  assign n29745 = \wishbone_bd_ram_mem0_reg[208][6]/P0001  & n14010 ;
  assign n29746 = ~n29744 & ~n29745 ;
  assign n29747 = \wishbone_bd_ram_mem0_reg[176][6]/P0001  & n13262 ;
  assign n29748 = \wishbone_bd_ram_mem0_reg[65][6]/P0001  & n13842 ;
  assign n29749 = ~n29747 & ~n29748 ;
  assign n29750 = n29746 & n29749 ;
  assign n29751 = \wishbone_bd_ram_mem0_reg[3][6]/P0001  & n13354 ;
  assign n29752 = \wishbone_bd_ram_mem0_reg[85][6]/P0001  & n13784 ;
  assign n29753 = ~n29751 & ~n29752 ;
  assign n29754 = \wishbone_bd_ram_mem0_reg[9][6]/P0001  & n13580 ;
  assign n29755 = \wishbone_bd_ram_mem0_reg[145][6]/P0001  & n13715 ;
  assign n29756 = ~n29754 & ~n29755 ;
  assign n29757 = n29753 & n29756 ;
  assign n29758 = n29750 & n29757 ;
  assign n29759 = \wishbone_bd_ram_mem0_reg[64][6]/P0001  & n13904 ;
  assign n29760 = \wishbone_bd_ram_mem0_reg[147][6]/P0001  & n13702 ;
  assign n29761 = ~n29759 & ~n29760 ;
  assign n29762 = \wishbone_bd_ram_mem0_reg[218][6]/P0001  & n13792 ;
  assign n29763 = \wishbone_bd_ram_mem0_reg[188][6]/P0001  & n13407 ;
  assign n29764 = ~n29762 & ~n29763 ;
  assign n29765 = n29761 & n29764 ;
  assign n29766 = \wishbone_bd_ram_mem0_reg[139][6]/P0001  & n13566 ;
  assign n29767 = \wishbone_bd_ram_mem0_reg[207][6]/P0001  & n13826 ;
  assign n29768 = ~n29766 & ~n29767 ;
  assign n29769 = \wishbone_bd_ram_mem0_reg[128][6]/P0001  & n13652 ;
  assign n29770 = \wishbone_bd_ram_mem0_reg[216][6]/P0001  & n14005 ;
  assign n29771 = ~n29769 & ~n29770 ;
  assign n29772 = n29768 & n29771 ;
  assign n29773 = n29765 & n29772 ;
  assign n29774 = n29758 & n29773 ;
  assign n29775 = \wishbone_bd_ram_mem0_reg[138][6]/P0001  & n13398 ;
  assign n29776 = \wishbone_bd_ram_mem0_reg[177][6]/P0001  & n13863 ;
  assign n29777 = ~n29775 & ~n29776 ;
  assign n29778 = \wishbone_bd_ram_mem0_reg[171][6]/P0001  & n13422 ;
  assign n29779 = \wishbone_bd_ram_mem0_reg[182][6]/P0001  & n13598 ;
  assign n29780 = ~n29778 & ~n29779 ;
  assign n29781 = n29777 & n29780 ;
  assign n29782 = \wishbone_bd_ram_mem0_reg[181][6]/P0001  & n13587 ;
  assign n29783 = \wishbone_bd_ram_mem0_reg[113][6]/P0001  & n13882 ;
  assign n29784 = ~n29782 & ~n29783 ;
  assign n29785 = \wishbone_bd_ram_mem0_reg[49][6]/P0001  & n13929 ;
  assign n29786 = \wishbone_bd_ram_mem0_reg[13][6]/P0001  & n13844 ;
  assign n29787 = ~n29785 & ~n29786 ;
  assign n29788 = n29784 & n29787 ;
  assign n29789 = n29781 & n29788 ;
  assign n29790 = \wishbone_bd_ram_mem0_reg[154][6]/P0001  & n13403 ;
  assign n29791 = \wishbone_bd_ram_mem0_reg[118][6]/P0001  & n13589 ;
  assign n29792 = ~n29790 & ~n29791 ;
  assign n29793 = \wishbone_bd_ram_mem0_reg[137][6]/P0001  & n13808 ;
  assign n29794 = \wishbone_bd_ram_mem0_reg[20][6]/P0001  & n13839 ;
  assign n29795 = ~n29793 & ~n29794 ;
  assign n29796 = n29792 & n29795 ;
  assign n29797 = \wishbone_bd_ram_mem0_reg[76][6]/P0001  & n13831 ;
  assign n29798 = \wishbone_bd_ram_mem0_reg[109][6]/P0001  & n13306 ;
  assign n29799 = ~n29797 & ~n29798 ;
  assign n29800 = \wishbone_bd_ram_mem0_reg[2][6]/P0001  & n13975 ;
  assign n29801 = \wishbone_bd_ram_mem0_reg[186][6]/P0001  & n13616 ;
  assign n29802 = ~n29800 & ~n29801 ;
  assign n29803 = n29799 & n29802 ;
  assign n29804 = n29796 & n29803 ;
  assign n29805 = n29789 & n29804 ;
  assign n29806 = n29774 & n29805 ;
  assign n29807 = n29743 & n29806 ;
  assign n29808 = \wishbone_bd_ram_mem0_reg[61][6]/P0001  & n13544 ;
  assign n29809 = \wishbone_bd_ram_mem0_reg[162][6]/P0001  & n13726 ;
  assign n29810 = ~n29808 & ~n29809 ;
  assign n29811 = \wishbone_bd_ram_mem0_reg[203][6]/P0001  & n13816 ;
  assign n29812 = \wishbone_bd_ram_mem0_reg[231][6]/P0001  & n13363 ;
  assign n29813 = ~n29811 & ~n29812 ;
  assign n29814 = n29810 & n29813 ;
  assign n29815 = \wishbone_bd_ram_mem0_reg[223][6]/P0001  & n13335 ;
  assign n29816 = \wishbone_bd_ram_mem0_reg[196][6]/P0001  & n13977 ;
  assign n29817 = ~n29815 & ~n29816 ;
  assign n29818 = \wishbone_bd_ram_mem0_reg[62][6]/P0001  & n13529 ;
  assign n29819 = \wishbone_bd_ram_mem0_reg[52][6]/P0001  & n13988 ;
  assign n29820 = ~n29818 & ~n29819 ;
  assign n29821 = n29817 & n29820 ;
  assign n29822 = n29814 & n29821 ;
  assign n29823 = \wishbone_bd_ram_mem0_reg[193][6]/P0001  & n14022 ;
  assign n29824 = \wishbone_bd_ram_mem0_reg[59][6]/P0001  & n13613 ;
  assign n29825 = ~n29823 & ~n29824 ;
  assign n29826 = \wishbone_bd_ram_mem0_reg[71][6]/P0001  & n13636 ;
  assign n29827 = \wishbone_bd_ram_mem0_reg[191][6]/P0001  & n14012 ;
  assign n29828 = ~n29826 & ~n29827 ;
  assign n29829 = n29825 & n29828 ;
  assign n29830 = \wishbone_bd_ram_mem0_reg[198][6]/P0001  & n13592 ;
  assign n29831 = \wishbone_bd_ram_mem0_reg[98][6]/P0001  & n13569 ;
  assign n29832 = ~n29830 & ~n29831 ;
  assign n29833 = \wishbone_bd_ram_mem0_reg[120][6]/P0001  & n13550 ;
  assign n29834 = \wishbone_bd_ram_mem0_reg[63][6]/P0001  & n13327 ;
  assign n29835 = ~n29833 & ~n29834 ;
  assign n29836 = n29832 & n29835 ;
  assign n29837 = n29829 & n29836 ;
  assign n29838 = n29822 & n29837 ;
  assign n29839 = \wishbone_bd_ram_mem0_reg[161][6]/P0001  & n13505 ;
  assign n29840 = \wishbone_bd_ram_mem0_reg[243][6]/P0001  & n13575 ;
  assign n29841 = ~n29839 & ~n29840 ;
  assign n29842 = \wishbone_bd_ram_mem0_reg[38][6]/P0001  & n13828 ;
  assign n29843 = \wishbone_bd_ram_mem0_reg[22][6]/P0001  & n13744 ;
  assign n29844 = ~n29842 & ~n29843 ;
  assign n29845 = n29841 & n29844 ;
  assign n29846 = \wishbone_bd_ram_mem0_reg[58][6]/P0001  & n13949 ;
  assign n29847 = \wishbone_bd_ram_mem0_reg[56][6]/P0001  & n13611 ;
  assign n29848 = ~n29846 & ~n29847 ;
  assign n29849 = \wishbone_bd_ram_mem0_reg[126][6]/P0001  & n13786 ;
  assign n29850 = \wishbone_bd_ram_mem0_reg[125][6]/P0001  & n13396 ;
  assign n29851 = ~n29849 & ~n29850 ;
  assign n29852 = n29848 & n29851 ;
  assign n29853 = n29845 & n29852 ;
  assign n29854 = \wishbone_bd_ram_mem0_reg[44][6]/P0001  & n13291 ;
  assign n29855 = \wishbone_bd_ram_mem0_reg[94][6]/P0001  & n13833 ;
  assign n29856 = ~n29854 & ~n29855 ;
  assign n29857 = \wishbone_bd_ram_mem0_reg[29][6]/P0001  & n13412 ;
  assign n29858 = \wishbone_bd_ram_mem0_reg[66][6]/P0001  & n13603 ;
  assign n29859 = ~n29857 & ~n29858 ;
  assign n29860 = n29856 & n29859 ;
  assign n29861 = \wishbone_bd_ram_mem0_reg[130][6]/P0001  & n13427 ;
  assign n29862 = \wishbone_bd_ram_mem0_reg[18][6]/P0001  & n13532 ;
  assign n29863 = ~n29861 & ~n29862 ;
  assign n29864 = \wishbone_bd_ram_mem0_reg[199][6]/P0001  & n13499 ;
  assign n29865 = \wishbone_bd_ram_mem0_reg[45][6]/P0001  & n13420 ;
  assign n29866 = ~n29864 & ~n29865 ;
  assign n29867 = n29863 & n29866 ;
  assign n29868 = n29860 & n29867 ;
  assign n29869 = n29853 & n29868 ;
  assign n29870 = n29838 & n29869 ;
  assign n29871 = \wishbone_bd_ram_mem0_reg[19][6]/P0001  & n13886 ;
  assign n29872 = \wishbone_bd_ram_mem0_reg[133][6]/P0001  & n13492 ;
  assign n29873 = ~n29871 & ~n29872 ;
  assign n29874 = \wishbone_bd_ram_mem0_reg[96][6]/P0001  & n13425 ;
  assign n29875 = \wishbone_bd_ram_mem0_reg[224][6]/P0001  & n13433 ;
  assign n29876 = ~n29874 & ~n29875 ;
  assign n29877 = n29873 & n29876 ;
  assign n29878 = \wishbone_bd_ram_mem0_reg[114][6]/P0001  & n13763 ;
  assign n29879 = \wishbone_bd_ram_mem0_reg[227][6]/P0001  & n13388 ;
  assign n29880 = ~n29878 & ~n29879 ;
  assign n29881 = \wishbone_bd_ram_mem0_reg[1][6]/P0001  & n13888 ;
  assign n29882 = \wishbone_bd_ram_mem0_reg[60][6]/P0001  & n13790 ;
  assign n29883 = ~n29881 & ~n29882 ;
  assign n29884 = n29880 & n29883 ;
  assign n29885 = n29877 & n29884 ;
  assign n29886 = \wishbone_bd_ram_mem0_reg[219][6]/P0001  & n13577 ;
  assign n29887 = \wishbone_bd_ram_mem0_reg[179][6]/P0001  & n14035 ;
  assign n29888 = ~n29886 & ~n29887 ;
  assign n29889 = \wishbone_bd_ram_mem0_reg[146][6]/P0001  & n13958 ;
  assign n29890 = \wishbone_bd_ram_mem0_reg[204][6]/P0001  & n13821 ;
  assign n29891 = ~n29889 & ~n29890 ;
  assign n29892 = n29888 & n29891 ;
  assign n29893 = \wishbone_bd_ram_mem0_reg[88][6]/P0001  & n13347 ;
  assign n29894 = \wishbone_bd_ram_mem0_reg[254][6]/P0001  & n13283 ;
  assign n29895 = ~n29893 & ~n29894 ;
  assign n29896 = \wishbone_bd_ram_mem0_reg[87][6]/P0001  & n13691 ;
  assign n29897 = \wishbone_bd_ram_mem0_reg[100][6]/P0001  & n13401 ;
  assign n29898 = ~n29896 & ~n29897 ;
  assign n29899 = n29895 & n29898 ;
  assign n29900 = n29892 & n29899 ;
  assign n29901 = n29885 & n29900 ;
  assign n29902 = \wishbone_bd_ram_mem0_reg[26][6]/P0001  & n13521 ;
  assign n29903 = \wishbone_bd_ram_mem0_reg[117][6]/P0001  & n13557 ;
  assign n29904 = ~n29902 & ~n29903 ;
  assign n29905 = \wishbone_bd_ram_mem0_reg[241][6]/P0001  & n13854 ;
  assign n29906 = \wishbone_bd_ram_mem0_reg[248][6]/P0001  & n13647 ;
  assign n29907 = ~n29905 & ~n29906 ;
  assign n29908 = n29904 & n29907 ;
  assign n29909 = \wishbone_bd_ram_mem0_reg[53][6]/P0001  & n13875 ;
  assign n29910 = \wishbone_bd_ram_mem0_reg[187][6]/P0001  & n13756 ;
  assign n29911 = ~n29909 & ~n29910 ;
  assign n29912 = \wishbone_bd_ram_mem0_reg[36][6]/P0001  & n13639 ;
  assign n29913 = \wishbone_bd_ram_mem0_reg[155][6]/P0001  & n13738 ;
  assign n29914 = ~n29912 & ~n29913 ;
  assign n29915 = n29911 & n29914 ;
  assign n29916 = n29908 & n29915 ;
  assign n29917 = \wishbone_bd_ram_mem0_reg[211][6]/P0001  & n13805 ;
  assign n29918 = \wishbone_bd_ram_mem0_reg[81][6]/P0001  & n13409 ;
  assign n29919 = ~n29917 & ~n29918 ;
  assign n29920 = \wishbone_bd_ram_mem0_reg[35][6]/P0001  & n13523 ;
  assign n29921 = \wishbone_bd_ram_mem0_reg[238][6]/P0001  & n13819 ;
  assign n29922 = ~n29920 & ~n29921 ;
  assign n29923 = n29919 & n29922 ;
  assign n29924 = \wishbone_bd_ram_mem0_reg[244][6]/P0001  & n13474 ;
  assign n29925 = \wishbone_bd_ram_mem0_reg[215][6]/P0001  & n13901 ;
  assign n29926 = ~n29924 & ~n29925 ;
  assign n29927 = \wishbone_bd_ram_mem0_reg[153][6]/P0001  & n13309 ;
  assign n29928 = \wishbone_bd_ram_mem0_reg[131][6]/P0001  & n13358 ;
  assign n29929 = ~n29927 & ~n29928 ;
  assign n29930 = n29926 & n29929 ;
  assign n29931 = n29923 & n29930 ;
  assign n29932 = n29916 & n29931 ;
  assign n29933 = n29901 & n29932 ;
  assign n29934 = n29870 & n29933 ;
  assign n29935 = n29807 & n29934 ;
  assign n29936 = \wishbone_bd_ram_mem0_reg[50][6]/P0001  & n13686 ;
  assign n29937 = \wishbone_bd_ram_mem0_reg[12][6]/P0001  & n13733 ;
  assign n29938 = ~n29936 & ~n29937 ;
  assign n29939 = \wishbone_bd_ram_mem0_reg[99][6]/P0001  & n13996 ;
  assign n29940 = \wishbone_bd_ram_mem0_reg[206][6]/P0001  & n13414 ;
  assign n29941 = ~n29939 & ~n29940 ;
  assign n29942 = n29938 & n29941 ;
  assign n29943 = \wishbone_bd_ram_mem0_reg[141][6]/P0001  & n13852 ;
  assign n29944 = \wishbone_bd_ram_mem0_reg[40][6]/P0001  & n13661 ;
  assign n29945 = ~n29943 & ~n29944 ;
  assign n29946 = \wishbone_bd_ram_mem0_reg[229][6]/P0001  & n13552 ;
  assign n29947 = \wishbone_bd_ram_mem0_reg[57][6]/P0001  & n13731 ;
  assign n29948 = ~n29946 & ~n29947 ;
  assign n29949 = n29945 & n29948 ;
  assign n29950 = n29942 & n29949 ;
  assign n29951 = \wishbone_bd_ram_mem0_reg[143][6]/P0001  & n13461 ;
  assign n29952 = \wishbone_bd_ram_mem0_reg[17][6]/P0001  & n13324 ;
  assign n29953 = ~n29951 & ~n29952 ;
  assign n29954 = \wishbone_bd_ram_mem0_reg[236][6]/P0001  & n13480 ;
  assign n29955 = \wishbone_bd_ram_mem0_reg[168][6]/P0001  & n13795 ;
  assign n29956 = ~n29954 & ~n29955 ;
  assign n29957 = n29953 & n29956 ;
  assign n29958 = \wishbone_bd_ram_mem0_reg[148][6]/P0001  & n13868 ;
  assign n29959 = \wishbone_bd_ram_mem0_reg[132][6]/P0001  & n13927 ;
  assign n29960 = ~n29958 & ~n29959 ;
  assign n29961 = \wishbone_bd_ram_mem0_reg[124][6]/P0001  & n14024 ;
  assign n29962 = \wishbone_bd_ram_mem0_reg[163][6]/P0001  & n13255 ;
  assign n29963 = ~n29961 & ~n29962 ;
  assign n29964 = n29960 & n29963 ;
  assign n29965 = n29957 & n29964 ;
  assign n29966 = n29950 & n29965 ;
  assign n29967 = \wishbone_bd_ram_mem0_reg[240][6]/P0001  & n13352 ;
  assign n29968 = \wishbone_bd_ram_mem0_reg[68][6]/P0001  & n13379 ;
  assign n29969 = ~n29967 & ~n29968 ;
  assign n29970 = \wishbone_bd_ram_mem0_reg[28][6]/P0001  & n13810 ;
  assign n29971 = \wishbone_bd_ram_mem0_reg[103][6]/P0001  & n13320 ;
  assign n29972 = ~n29970 & ~n29971 ;
  assign n29973 = n29969 & n29972 ;
  assign n29974 = \wishbone_bd_ram_mem0_reg[246][6]/P0001  & n13981 ;
  assign n29975 = \wishbone_bd_ram_mem0_reg[110][6]/P0001  & n14030 ;
  assign n29976 = ~n29974 & ~n29975 ;
  assign n29977 = \wishbone_bd_ram_mem0_reg[91][6]/P0001  & n13954 ;
  assign n29978 = \wishbone_bd_ram_mem0_reg[234][6]/P0001  & n13781 ;
  assign n29979 = ~n29977 & ~n29978 ;
  assign n29980 = n29976 & n29979 ;
  assign n29981 = n29973 & n29980 ;
  assign n29982 = \wishbone_bd_ram_mem0_reg[95][6]/P0001  & n13317 ;
  assign n29983 = \wishbone_bd_ram_mem0_reg[8][6]/P0001  & n13459 ;
  assign n29984 = ~n29982 & ~n29983 ;
  assign n29985 = \wishbone_bd_ram_mem0_reg[70][6]/P0001  & n13339 ;
  assign n29986 = \wishbone_bd_ram_mem0_reg[83][6]/P0001  & n13454 ;
  assign n29987 = ~n29985 & ~n29986 ;
  assign n29988 = n29984 & n29987 ;
  assign n29989 = \wishbone_bd_ram_mem0_reg[101][6]/P0001  & n13772 ;
  assign n29990 = \wishbone_bd_ram_mem0_reg[7][6]/P0001  & n13546 ;
  assign n29991 = ~n29989 & ~n29990 ;
  assign n29992 = \wishbone_bd_ram_mem0_reg[142][6]/P0001  & n13448 ;
  assign n29993 = \wishbone_bd_ram_mem0_reg[54][6]/P0001  & n13622 ;
  assign n29994 = ~n29992 & ~n29993 ;
  assign n29995 = n29991 & n29994 ;
  assign n29996 = n29988 & n29995 ;
  assign n29997 = n29981 & n29996 ;
  assign n29998 = n29966 & n29997 ;
  assign n29999 = \wishbone_bd_ram_mem0_reg[226][6]/P0001  & n13668 ;
  assign n30000 = \wishbone_bd_ram_mem0_reg[23][6]/P0001  & n13857 ;
  assign n30001 = ~n29999 & ~n30000 ;
  assign n30002 = \wishbone_bd_ram_mem0_reg[30][6]/P0001  & n13713 ;
  assign n30003 = \wishbone_bd_ram_mem0_reg[209][6]/P0001  & n13689 ;
  assign n30004 = ~n30002 & ~n30003 ;
  assign n30005 = n30001 & n30004 ;
  assign n30006 = \wishbone_bd_ram_mem0_reg[245][6]/P0001  & n13877 ;
  assign n30007 = \wishbone_bd_ram_mem0_reg[166][6]/P0001  & n13999 ;
  assign n30008 = ~n30006 & ~n30007 ;
  assign n30009 = \wishbone_bd_ram_mem0_reg[97][6]/P0001  & n13724 ;
  assign n30010 = \wishbone_bd_ram_mem0_reg[31][6]/P0001  & n13758 ;
  assign n30011 = ~n30009 & ~n30010 ;
  assign n30012 = n30008 & n30011 ;
  assign n30013 = n30005 & n30012 ;
  assign n30014 = \wishbone_bd_ram_mem0_reg[69][6]/P0001  & n13487 ;
  assign n30015 = \wishbone_bd_ram_mem0_reg[195][6]/P0001  & n13700 ;
  assign n30016 = ~n30014 & ~n30015 ;
  assign n30017 = \wishbone_bd_ram_mem0_reg[160][6]/P0001  & n13271 ;
  assign n30018 = \wishbone_bd_ram_mem0_reg[175][6]/P0001  & n13674 ;
  assign n30019 = ~n30017 & ~n30018 ;
  assign n30020 = n30016 & n30019 ;
  assign n30021 = \wishbone_bd_ram_mem0_reg[157][6]/P0001  & n13445 ;
  assign n30022 = \wishbone_bd_ram_mem0_reg[122][6]/P0001  & n13679 ;
  assign n30023 = ~n30021 & ~n30022 ;
  assign n30024 = \wishbone_bd_ram_mem0_reg[167][6]/P0001  & n13940 ;
  assign n30025 = \wishbone_bd_ram_mem0_reg[41][6]/P0001  & n14017 ;
  assign n30026 = ~n30024 & ~n30025 ;
  assign n30027 = n30023 & n30026 ;
  assign n30028 = n30020 & n30027 ;
  assign n30029 = n30013 & n30028 ;
  assign n30030 = \wishbone_bd_ram_mem0_reg[242][6]/P0001  & n13383 ;
  assign n30031 = \wishbone_bd_ram_mem0_reg[220][6]/P0001  & n13965 ;
  assign n30032 = ~n30030 & ~n30031 ;
  assign n30033 = \wishbone_bd_ram_mem0_reg[123][6]/P0001  & n13749 ;
  assign n30034 = \wishbone_bd_ram_mem0_reg[6][6]/P0001  & n13915 ;
  assign n30035 = ~n30033 & ~n30034 ;
  assign n30036 = n30032 & n30035 ;
  assign n30037 = \wishbone_bd_ram_mem0_reg[189][6]/P0001  & n14001 ;
  assign n30038 = \wishbone_bd_ram_mem0_reg[55][6]/P0001  & n13618 ;
  assign n30039 = ~n30037 & ~n30038 ;
  assign n30040 = \wishbone_bd_ram_mem0_reg[190][6]/P0001  & n13365 ;
  assign n30041 = \wishbone_bd_ram_mem0_reg[170][6]/P0001  & n14007 ;
  assign n30042 = ~n30040 & ~n30041 ;
  assign n30043 = n30039 & n30042 ;
  assign n30044 = n30036 & n30043 ;
  assign n30045 = \wishbone_bd_ram_mem0_reg[250][6]/P0001  & n13677 ;
  assign n30046 = \wishbone_bd_ram_mem0_reg[119][6]/P0001  & n14033 ;
  assign n30047 = ~n30045 & ~n30046 ;
  assign n30048 = \wishbone_bd_ram_mem0_reg[159][6]/P0001  & n13627 ;
  assign n30049 = \wishbone_bd_ram_mem0_reg[232][6]/P0001  & n13510 ;
  assign n30050 = ~n30048 & ~n30049 ;
  assign n30051 = n30047 & n30050 ;
  assign n30052 = \wishbone_bd_ram_mem0_reg[75][6]/P0001  & n13605 ;
  assign n30053 = \wishbone_bd_ram_mem0_reg[47][6]/P0001  & n13436 ;
  assign n30054 = ~n30052 & ~n30053 ;
  assign n30055 = \wishbone_bd_ram_mem0_reg[42][6]/P0001  & n13341 ;
  assign n30056 = \wishbone_bd_ram_mem0_reg[0][6]/P0001  & n13539 ;
  assign n30057 = ~n30055 & ~n30056 ;
  assign n30058 = n30054 & n30057 ;
  assign n30059 = n30051 & n30058 ;
  assign n30060 = n30044 & n30059 ;
  assign n30061 = n30029 & n30060 ;
  assign n30062 = n29998 & n30061 ;
  assign n30063 = \wishbone_bd_ram_mem0_reg[34][6]/P0001  & n13450 ;
  assign n30064 = \wishbone_bd_ram_mem0_reg[222][6]/P0001  & n13721 ;
  assign n30065 = ~n30063 & ~n30064 ;
  assign n30066 = \wishbone_bd_ram_mem0_reg[152][6]/P0001  & n13912 ;
  assign n30067 = \wishbone_bd_ram_mem0_reg[93][6]/P0001  & n13891 ;
  assign n30068 = ~n30066 & ~n30067 ;
  assign n30069 = n30065 & n30068 ;
  assign n30070 = \wishbone_bd_ram_mem0_reg[102][6]/P0001  & n13534 ;
  assign n30071 = \wishbone_bd_ram_mem0_reg[129][6]/P0001  & n13629 ;
  assign n30072 = ~n30070 & ~n30071 ;
  assign n30073 = \wishbone_bd_ram_mem0_reg[164][6]/P0001  & n13236 ;
  assign n30074 = \wishbone_bd_ram_mem0_reg[233][6]/P0001  & n13332 ;
  assign n30075 = ~n30073 & ~n30074 ;
  assign n30076 = n30072 & n30075 ;
  assign n30077 = n30069 & n30076 ;
  assign n30078 = \wishbone_bd_ram_mem0_reg[136][6]/P0001  & n13963 ;
  assign n30079 = \wishbone_bd_ram_mem0_reg[239][6]/P0001  & n13349 ;
  assign n30080 = ~n30078 & ~n30079 ;
  assign n30081 = \wishbone_bd_ram_mem0_reg[25][6]/P0001  & n13742 ;
  assign n30082 = \wishbone_bd_ram_mem0_reg[106][6]/P0001  & n13555 ;
  assign n30083 = ~n30081 & ~n30082 ;
  assign n30084 = n30080 & n30083 ;
  assign n30085 = \wishbone_bd_ram_mem0_reg[14][6]/P0001  & n13972 ;
  assign n30086 = \wishbone_bd_ram_mem0_reg[5][6]/P0001  & n13243 ;
  assign n30087 = ~n30085 & ~n30086 ;
  assign n30088 = \wishbone_bd_ram_mem0_reg[134][6]/P0001  & n13494 ;
  assign n30089 = \wishbone_bd_ram_mem0_reg[77][6]/P0001  & n13935 ;
  assign n30090 = ~n30088 & ~n30089 ;
  assign n30091 = n30087 & n30090 ;
  assign n30092 = n30084 & n30091 ;
  assign n30093 = n30077 & n30092 ;
  assign n30094 = \wishbone_bd_ram_mem0_reg[180][6]/P0001  & n13650 ;
  assign n30095 = \wishbone_bd_ram_mem0_reg[46][6]/P0001  & n13298 ;
  assign n30096 = ~n30094 & ~n30095 ;
  assign n30097 = \wishbone_bd_ram_mem0_reg[78][6]/P0001  & n13277 ;
  assign n30098 = \wishbone_bd_ram_mem0_reg[230][6]/P0001  & n13994 ;
  assign n30099 = ~n30097 & ~n30098 ;
  assign n30100 = n30096 & n30099 ;
  assign n30101 = \wishbone_bd_ram_mem0_reg[107][6]/P0001  & n13476 ;
  assign n30102 = \wishbone_bd_ram_mem0_reg[165][6]/P0001  & n14028 ;
  assign n30103 = ~n30101 & ~n30102 ;
  assign n30104 = \wishbone_bd_ram_mem0_reg[15][6]/P0001  & n13797 ;
  assign n30105 = \wishbone_bd_ram_mem0_reg[115][6]/P0001  & n13747 ;
  assign n30106 = ~n30104 & ~n30105 ;
  assign n30107 = n30103 & n30106 ;
  assign n30108 = n30100 & n30107 ;
  assign n30109 = \wishbone_bd_ram_mem0_reg[140][6]/P0001  & n13287 ;
  assign n30110 = \wishbone_bd_ram_mem0_reg[202][6]/P0001  & n13268 ;
  assign n30111 = ~n30109 & ~n30110 ;
  assign n30112 = \wishbone_bd_ram_mem0_reg[112][6]/P0001  & n13482 ;
  assign n30113 = \wishbone_bd_ram_mem0_reg[135][6]/P0001  & n13672 ;
  assign n30114 = ~n30112 & ~n30113 ;
  assign n30115 = n30111 & n30114 ;
  assign n30116 = \wishbone_bd_ram_mem0_reg[43][6]/P0001  & n13761 ;
  assign n30117 = \wishbone_bd_ram_mem0_reg[86][6]/P0001  & n13485 ;
  assign n30118 = ~n30116 & ~n30117 ;
  assign n30119 = \wishbone_bd_ram_mem0_reg[213][6]/P0001  & n13870 ;
  assign n30120 = \wishbone_bd_ram_mem0_reg[150][6]/P0001  & n13666 ;
  assign n30121 = ~n30119 & ~n30120 ;
  assign n30122 = n30118 & n30121 ;
  assign n30123 = n30115 & n30122 ;
  assign n30124 = n30108 & n30123 ;
  assign n30125 = n30093 & n30124 ;
  assign n30126 = \wishbone_bd_ram_mem0_reg[173][6]/P0001  & n13360 ;
  assign n30127 = \wishbone_bd_ram_mem0_reg[67][6]/P0001  & n13663 ;
  assign n30128 = ~n30126 & ~n30127 ;
  assign n30129 = \wishbone_bd_ram_mem0_reg[205][6]/P0001  & n13947 ;
  assign n30130 = \wishbone_bd_ram_mem0_reg[158][6]/P0001  & n13294 ;
  assign n30131 = ~n30129 & ~n30130 ;
  assign n30132 = n30128 & n30131 ;
  assign n30133 = \wishbone_bd_ram_mem0_reg[192][6]/P0001  & n13390 ;
  assign n30134 = \wishbone_bd_ram_mem0_reg[169][6]/P0001  & n13541 ;
  assign n30135 = ~n30133 & ~n30134 ;
  assign n30136 = \wishbone_bd_ram_mem0_reg[201][6]/P0001  & n13600 ;
  assign n30137 = \wishbone_bd_ram_mem0_reg[200][6]/P0001  & n13922 ;
  assign n30138 = ~n30136 & ~n30137 ;
  assign n30139 = n30135 & n30138 ;
  assign n30140 = n30132 & n30139 ;
  assign n30141 = \wishbone_bd_ram_mem0_reg[16][6]/P0001  & n13695 ;
  assign n30142 = \wishbone_bd_ram_mem0_reg[11][6]/P0001  & n13774 ;
  assign n30143 = ~n30141 & ~n30142 ;
  assign n30144 = \wishbone_bd_ram_mem0_reg[24][6]/P0001  & n13970 ;
  assign n30145 = \wishbone_bd_ram_mem0_reg[184][6]/P0001  & n13960 ;
  assign n30146 = ~n30144 & ~n30145 ;
  assign n30147 = n30143 & n30146 ;
  assign n30148 = \wishbone_bd_ram_mem0_reg[214][6]/P0001  & n13938 ;
  assign n30149 = \wishbone_bd_ram_mem0_reg[108][6]/P0001  & n13814 ;
  assign n30150 = ~n30148 & ~n30149 ;
  assign n30151 = \wishbone_bd_ram_mem0_reg[10][6]/P0001  & n13837 ;
  assign n30152 = \wishbone_bd_ram_mem0_reg[27][6]/P0001  & n13251 ;
  assign n30153 = ~n30151 & ~n30152 ;
  assign n30154 = n30150 & n30153 ;
  assign n30155 = n30147 & n30154 ;
  assign n30156 = n30140 & n30155 ;
  assign n30157 = \wishbone_bd_ram_mem0_reg[39][6]/P0001  & n13893 ;
  assign n30158 = \wishbone_bd_ram_mem0_reg[116][6]/P0001  & n13865 ;
  assign n30159 = ~n30157 & ~n30158 ;
  assign n30160 = \wishbone_bd_ram_mem0_reg[90][6]/P0001  & n13906 ;
  assign n30161 = \wishbone_bd_ram_mem0_reg[156][6]/P0001  & n13769 ;
  assign n30162 = ~n30160 & ~n30161 ;
  assign n30163 = n30159 & n30162 ;
  assign n30164 = \wishbone_bd_ram_mem0_reg[251][6]/P0001  & n14019 ;
  assign n30165 = \wishbone_bd_ram_mem0_reg[235][6]/P0001  & n13518 ;
  assign n30166 = ~n30164 & ~n30165 ;
  assign n30167 = \wishbone_bd_ram_mem0_reg[111][6]/P0001  & n13471 ;
  assign n30168 = \wishbone_bd_ram_mem0_reg[247][6]/P0001  & n13571 ;
  assign n30169 = ~n30167 & ~n30168 ;
  assign n30170 = n30166 & n30169 ;
  assign n30171 = n30163 & n30170 ;
  assign n30172 = \wishbone_bd_ram_mem0_reg[48][6]/P0001  & n13917 ;
  assign n30173 = \wishbone_bd_ram_mem0_reg[253][6]/P0001  & n13708 ;
  assign n30174 = ~n30172 & ~n30173 ;
  assign n30175 = \wishbone_bd_ram_mem0_reg[172][6]/P0001  & n13377 ;
  assign n30176 = \wishbone_bd_ram_mem0_reg[228][6]/P0001  & n13497 ;
  assign n30177 = ~n30175 & ~n30176 ;
  assign n30178 = n30174 & n30177 ;
  assign n30179 = \wishbone_bd_ram_mem0_reg[82][6]/P0001  & n13374 ;
  assign n30180 = \wishbone_bd_ram_mem0_reg[105][6]/P0001  & n13503 ;
  assign n30181 = ~n30179 & ~n30180 ;
  assign n30182 = \wishbone_bd_ram_mem0_reg[37][6]/P0001  & n13710 ;
  assign n30183 = \wishbone_bd_ram_mem0_reg[185][6]/P0001  & n13372 ;
  assign n30184 = ~n30182 & ~n30183 ;
  assign n30185 = n30181 & n30184 ;
  assign n30186 = n30178 & n30185 ;
  assign n30187 = n30171 & n30186 ;
  assign n30188 = n30156 & n30187 ;
  assign n30189 = n30125 & n30188 ;
  assign n30190 = n30062 & n30189 ;
  assign n30191 = n29935 & n30190 ;
  assign n30192 = ~wb_rst_i_pad & ~n29679 ;
  assign n30193 = ~n30191 & n30192 ;
  assign n30194 = ~n29680 & ~n30193 ;
  assign n30195 = \ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131  & n23743 ;
  assign n30196 = n23747 & n30195 ;
  assign n30197 = \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  & n23751 ;
  assign n30198 = n23741 & n30197 ;
  assign n30199 = ~n30196 & ~n30198 ;
  assign n30200 = \ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131  & n23743 ;
  assign n30201 = n23741 & n30200 ;
  assign n30202 = n23730 & ~n30201 ;
  assign n30203 = n30199 & n30202 ;
  assign n30204 = \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131  & n25059 ;
  assign n30205 = \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  & n23737 ;
  assign n30206 = ~n30204 & ~n30205 ;
  assign n30207 = n30203 & n30206 ;
  assign n30208 = n23730 & ~n30207 ;
  assign n30209 = ~wb_rst_i_pad & ~n30207 ;
  assign n30210 = ~n20833 & n30209 ;
  assign n30211 = ~n30208 & ~n30210 ;
  assign n30212 = \ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131  & n23743 ;
  assign n30213 = n23747 & n30212 ;
  assign n30214 = \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  & n23751 ;
  assign n30215 = n23741 & n30214 ;
  assign n30216 = ~n30213 & ~n30215 ;
  assign n30217 = \ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131  & n23743 ;
  assign n30218 = n23741 & n30217 ;
  assign n30219 = n23730 & ~n30218 ;
  assign n30220 = n30216 & n30219 ;
  assign n30221 = \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131  & n25059 ;
  assign n30222 = \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  & n23737 ;
  assign n30223 = ~n30221 & ~n30222 ;
  assign n30224 = n30220 & n30223 ;
  assign n30225 = n23730 & ~n30224 ;
  assign n30226 = ~wb_rst_i_pad & ~n30224 ;
  assign n30227 = ~n19273 & n30226 ;
  assign n30228 = ~n30225 & ~n30227 ;
  assign n30229 = \ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131  & n23743 ;
  assign n30230 = n23747 & n30229 ;
  assign n30231 = \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  & n23751 ;
  assign n30232 = n23741 & n30231 ;
  assign n30233 = ~n30230 & ~n30232 ;
  assign n30234 = \ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131  & n23743 ;
  assign n30235 = n23741 & n30234 ;
  assign n30236 = n23730 & ~n30235 ;
  assign n30237 = n30233 & n30236 ;
  assign n30238 = \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131  & n25059 ;
  assign n30239 = \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  & n23737 ;
  assign n30240 = ~n30238 & ~n30239 ;
  assign n30241 = n30237 & n30240 ;
  assign n30242 = n23730 & ~n30241 ;
  assign n30243 = ~wb_rst_i_pad & ~n30241 ;
  assign n30244 = ~n22172 & n30243 ;
  assign n30245 = ~n30242 & ~n30244 ;
  assign n30246 = n18507 & ~n22172 ;
  assign n30247 = \wishbone_RxPointerMSB_reg[15]/NET0131  & \wishbone_RxPointerMSB_reg[17]/NET0131  ;
  assign n30248 = \wishbone_RxPointerMSB_reg[16]/NET0131  & n30247 ;
  assign n30249 = n18521 & n30248 ;
  assign n30250 = \wishbone_RxPointerMSB_reg[18]/NET0131  & n30249 ;
  assign n30251 = ~\wishbone_RxPointerMSB_reg[19]/NET0131  & ~n30250 ;
  assign n30252 = \wishbone_RxPointerMSB_reg[15]/NET0131  & n18524 ;
  assign n30253 = n18521 & n30252 ;
  assign n30254 = ~n16305 & ~n30253 ;
  assign n30255 = ~n30251 & n30254 ;
  assign n30256 = ~n30246 & ~n30255 ;
  assign n30257 = ~\wishbone_RxPointerMSB_reg[20]/NET0131  & ~n30253 ;
  assign n30258 = ~n16305 & ~n18527 ;
  assign n30259 = ~n30257 & n30258 ;
  assign n30260 = ~n17358 & n18507 ;
  assign n30261 = ~n30259 & ~n30260 ;
  assign n30262 = \wishbone_RxPointerMSB_reg[21]/NET0131  & ~n16305 ;
  assign n30263 = ~n18527 & n30262 ;
  assign n30264 = ~\wishbone_RxPointerMSB_reg[21]/NET0131  & ~n16305 ;
  assign n30265 = n18527 & n30264 ;
  assign n30266 = ~n30263 & ~n30265 ;
  assign n30267 = n18507 & ~n22688 ;
  assign n30268 = n30266 & ~n30267 ;
  assign n30269 = n18507 & ~n23718 ;
  assign n30270 = \wishbone_RxPointerMSB_reg[21]/NET0131  & n18527 ;
  assign n30271 = ~\wishbone_RxPointerMSB_reg[22]/NET0131  & ~n30270 ;
  assign n30272 = n18527 & n18528 ;
  assign n30273 = ~n16305 & ~n30272 ;
  assign n30274 = ~n30271 & n30273 ;
  assign n30275 = ~n30269 & ~n30274 ;
  assign n30276 = ~\wishbone_RxPointerMSB_reg[23]/NET0131  & ~n30272 ;
  assign n30277 = \wishbone_RxPointerMSB_reg[23]/NET0131  & n18528 ;
  assign n30278 = n18527 & n30277 ;
  assign n30279 = ~n16305 & ~n30278 ;
  assign n30280 = ~n30276 & n30279 ;
  assign n30281 = n18507 & ~n23202 ;
  assign n30282 = ~n30280 & ~n30281 ;
  assign n30283 = ~\wishbone_RxPointerMSB_reg[24]/NET0131  & ~n30278 ;
  assign n30284 = ~n16305 & ~n18531 ;
  assign n30285 = ~n30283 & n30284 ;
  assign n30286 = ~n15695 & n18507 ;
  assign n30287 = ~n30285 & ~n30286 ;
  assign n30288 = \wishbone_RxPointerMSB_reg[25]/NET0131  & ~n16305 ;
  assign n30289 = ~n18531 & n30288 ;
  assign n30290 = ~\wishbone_RxPointerMSB_reg[25]/NET0131  & ~n16305 ;
  assign n30291 = n18531 & n30290 ;
  assign n30292 = ~n30289 & ~n30291 ;
  assign n30293 = ~n18434 & n18507 ;
  assign n30294 = n30292 & ~n30293 ;
  assign n30295 = \wishbone_RxPointerMSB_reg[25]/NET0131  & \wishbone_RxPointerMSB_reg[26]/NET0131  ;
  assign n30296 = n18531 & n30295 ;
  assign n30297 = n18531 & n30288 ;
  assign n30298 = \wishbone_RxPointerMSB_reg[26]/NET0131  & ~n16305 ;
  assign n30299 = ~n30297 & ~n30298 ;
  assign n30300 = ~n30296 & ~n30299 ;
  assign n30301 = ~n17905 & n18507 ;
  assign n30302 = ~n30300 & ~n30301 ;
  assign n30303 = ~\wishbone_RxPointerMSB_reg[27]/NET0131  & ~n30296 ;
  assign n30304 = \wishbone_RxPointerMSB_reg[25]/NET0131  & \wishbone_RxPointerMSB_reg[27]/NET0131  ;
  assign n30305 = \wishbone_RxPointerMSB_reg[26]/NET0131  & n30304 ;
  assign n30306 = n18531 & n30305 ;
  assign n30307 = ~n16305 & ~n30306 ;
  assign n30308 = ~n30303 & n30307 ;
  assign n30309 = n18507 & ~n21643 ;
  assign n30310 = ~n30308 & ~n30309 ;
  assign n30311 = ~n14044 & n18507 ;
  assign n30312 = ~\wishbone_RxPointerMSB_reg[28]/NET0131  & ~n30306 ;
  assign n30313 = \wishbone_RxPointerMSB_reg[25]/NET0131  & n18533 ;
  assign n30314 = n18531 & n30313 ;
  assign n30315 = ~n16305 & ~n30314 ;
  assign n30316 = ~n30312 & n30315 ;
  assign n30317 = ~n30311 & ~n30316 ;
  assign n30318 = ~\wishbone_RxPointerMSB_reg[29]/NET0131  & ~n30314 ;
  assign n30319 = ~n16305 & ~n18536 ;
  assign n30320 = ~n30318 & n30319 ;
  assign n30321 = ~n14593 & n18507 ;
  assign n30322 = ~n30320 & ~n30321 ;
  assign n30323 = ~\wishbone_RxPointerMSB_reg[31]/NET0131  & ~n16305 ;
  assign n30324 = ~n18541 & n30323 ;
  assign n30325 = \wishbone_RxPointerMSB_reg[31]/NET0131  & ~n16305 ;
  assign n30326 = n18541 & n30325 ;
  assign n30327 = ~n30324 & ~n30326 ;
  assign n30328 = ~n16305 & n30327 ;
  assign n30329 = ~wb_rst_i_pad & n30327 ;
  assign n30330 = ~n20314 & n30329 ;
  assign n30331 = ~n30328 & ~n30330 ;
  assign n30332 = n18507 & ~n28346 ;
  assign n30333 = \wishbone_RxPointerMSB_reg[7]/NET0131  & \wishbone_RxPointerMSB_reg[8]/NET0131  ;
  assign n30334 = n18513 & n30333 ;
  assign n30335 = ~\wishbone_RxPointerMSB_reg[9]/NET0131  & ~n30334 ;
  assign n30336 = \wishbone_RxPointerMSB_reg[7]/NET0131  & n18514 ;
  assign n30337 = n18513 & n30336 ;
  assign n30338 = ~n16305 & ~n30337 ;
  assign n30339 = ~n30335 & n30338 ;
  assign n30340 = ~n30332 & ~n30339 ;
  assign n30341 = \wishbone_TxPointerMSB_reg[18]/NET0131  & \wishbone_TxPointerMSB_reg[19]/NET0131  ;
  assign n30342 = n18562 & n30341 ;
  assign n30343 = \wishbone_TxPointerMSB_reg[19]/NET0131  & ~n18545 ;
  assign n30344 = \wishbone_TxPointerMSB_reg[18]/NET0131  & ~n18545 ;
  assign n30345 = n18562 & n30344 ;
  assign n30346 = ~n30343 & ~n30345 ;
  assign n30347 = ~n30342 & ~n30346 ;
  assign n30348 = ~n22172 & n24387 ;
  assign n30349 = ~n30347 & ~n30348 ;
  assign n30350 = ~n17358 & n24387 ;
  assign n30351 = ~\wishbone_TxPointerMSB_reg[20]/NET0131  & ~n30342 ;
  assign n30352 = n18562 & n18564 ;
  assign n30353 = ~n18545 & ~n30352 ;
  assign n30354 = ~n30351 & n30353 ;
  assign n30355 = ~n30350 & ~n30354 ;
  assign n30356 = ~\wishbone_TxPointerMSB_reg[21]/NET0131  & ~n30352 ;
  assign n30357 = \wishbone_TxPointerMSB_reg[18]/NET0131  & \wishbone_TxPointerMSB_reg[21]/NET0131  ;
  assign n30358 = n18563 & n30357 ;
  assign n30359 = n18562 & n30358 ;
  assign n30360 = ~n18545 & ~n30359 ;
  assign n30361 = ~n30356 & n30360 ;
  assign n30362 = ~n22688 & n24387 ;
  assign n30363 = ~n30361 & ~n30362 ;
  assign n30364 = ~n23718 & n24387 ;
  assign n30365 = ~\wishbone_TxPointerMSB_reg[22]/NET0131  & ~n30359 ;
  assign n30366 = ~n18545 & ~n18567 ;
  assign n30367 = ~n30365 & n30366 ;
  assign n30368 = ~n30364 & ~n30367 ;
  assign n30369 = \wishbone_TxPointerMSB_reg[23]/NET0131  & ~n18545 ;
  assign n30370 = ~n18567 & n30369 ;
  assign n30371 = ~\wishbone_TxPointerMSB_reg[23]/NET0131  & ~n18545 ;
  assign n30372 = n18567 & n30371 ;
  assign n30373 = ~n30370 & ~n30372 ;
  assign n30374 = ~n23202 & n24387 ;
  assign n30375 = n30373 & ~n30374 ;
  assign n30376 = ~n15695 & n24387 ;
  assign n30377 = \wishbone_TxPointerMSB_reg[23]/NET0131  & n18567 ;
  assign n30378 = ~\wishbone_TxPointerMSB_reg[24]/NET0131  & ~n30377 ;
  assign n30379 = n18567 & n18570 ;
  assign n30380 = ~n18545 & ~n30379 ;
  assign n30381 = ~n30378 & n30380 ;
  assign n30382 = ~n30376 & ~n30381 ;
  assign n30383 = \wishbone_TxPointerMSB_reg[25]/NET0131  & n18570 ;
  assign n30384 = n18567 & n30383 ;
  assign n30385 = \wishbone_TxPointerMSB_reg[25]/NET0131  & ~n18545 ;
  assign n30386 = ~n18545 & n18570 ;
  assign n30387 = n18567 & n30386 ;
  assign n30388 = ~n30385 & ~n30387 ;
  assign n30389 = ~n30384 & ~n30388 ;
  assign n30390 = ~n18434 & n24387 ;
  assign n30391 = ~n30389 & ~n30390 ;
  assign n30392 = ~n17905 & n24387 ;
  assign n30393 = ~\wishbone_TxPointerMSB_reg[26]/NET0131  & ~n30384 ;
  assign n30394 = n18568 & n18570 ;
  assign n30395 = n18567 & n30394 ;
  assign n30396 = ~n18545 & ~n30395 ;
  assign n30397 = ~n30393 & n30396 ;
  assign n30398 = ~n30392 & ~n30397 ;
  assign n30399 = ~\wishbone_TxPointerMSB_reg[27]/NET0131  & ~n30395 ;
  assign n30400 = \wishbone_TxPointerMSB_reg[27]/NET0131  & n18570 ;
  assign n30401 = n18568 & n30400 ;
  assign n30402 = n18567 & n30401 ;
  assign n30403 = ~n18545 & ~n30402 ;
  assign n30404 = ~n30399 & n30403 ;
  assign n30405 = ~n21643 & n24387 ;
  assign n30406 = ~n30404 & ~n30405 ;
  assign n30407 = \wishbone_TxPointerMSB_reg[29]/NET0131  & ~n18545 ;
  assign n30408 = ~n18573 & n30407 ;
  assign n30409 = ~\wishbone_TxPointerMSB_reg[29]/NET0131  & ~n18545 ;
  assign n30410 = n18573 & n30409 ;
  assign n30411 = ~n30408 & ~n30410 ;
  assign n30412 = ~n14593 & n24387 ;
  assign n30413 = n30411 & ~n30412 ;
  assign n30414 = ~n14044 & n24387 ;
  assign n30415 = ~\wishbone_TxPointerMSB_reg[28]/NET0131  & ~n30402 ;
  assign n30416 = ~n18545 & ~n18573 ;
  assign n30417 = ~n30415 & n30416 ;
  assign n30418 = ~n30414 & ~n30417 ;
  assign n30419 = n18569 & n18574 ;
  assign n30420 = n30394 & n30419 ;
  assign n30421 = n18567 & n30420 ;
  assign n30422 = \wishbone_TxPointerMSB_reg[31]/NET0131  & ~n18545 ;
  assign n30423 = ~n30421 & n30422 ;
  assign n30424 = ~\wishbone_TxPointerMSB_reg[31]/NET0131  & ~n18545 ;
  assign n30425 = n30421 & n30424 ;
  assign n30426 = ~n30423 & ~n30425 ;
  assign n30427 = ~n20314 & n24387 ;
  assign n30428 = n30426 & ~n30427 ;
  assign n30429 = \wishbone_TxPointerMSB_reg[7]/NET0131  & \wishbone_TxPointerMSB_reg[8]/NET0131  ;
  assign n30430 = n18551 & n30429 ;
  assign n30431 = ~\wishbone_TxPointerMSB_reg[9]/NET0131  & ~n30430 ;
  assign n30432 = ~n18545 & ~n18554 ;
  assign n30433 = ~n30431 & n30432 ;
  assign n30434 = n24387 & ~n28346 ;
  assign n30435 = ~n30433 & ~n30434 ;
  assign n30436 = \ethreg1_MODER_1_DataOut_reg[5]/NET0131  & n23808 ;
  assign n30437 = \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131  & n23794 ;
  assign n30438 = n23741 & n30437 ;
  assign n30439 = ~n30436 & ~n30438 ;
  assign n30440 = \ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131  & n23743 ;
  assign n30441 = n23741 & n30440 ;
  assign n30442 = \ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131  & n23743 ;
  assign n30443 = n23747 & n30442 ;
  assign n30444 = ~n30441 & ~n30443 ;
  assign n30445 = n30439 & n30444 ;
  assign n30446 = n23730 & n30445 ;
  assign n30447 = \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  & n23737 ;
  assign n30448 = \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131  & n23813 ;
  assign n30449 = \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  & n23751 ;
  assign n30450 = n23741 & n30449 ;
  assign n30451 = ~n30448 & ~n30450 ;
  assign n30452 = \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  & n23751 ;
  assign n30453 = n23747 & n30452 ;
  assign n30454 = \ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131  & n23782 ;
  assign n30455 = ~n30453 & ~n30454 ;
  assign n30456 = n30451 & n30455 ;
  assign n30457 = ~n30447 & n30456 ;
  assign n30458 = n30446 & n30457 ;
  assign n30459 = n23730 & ~n30458 ;
  assign n30460 = \wishbone_bd_ram_mem1_reg[65][13]/P0001  & n13842 ;
  assign n30461 = \wishbone_bd_ram_mem1_reg[126][13]/P0001  & n13786 ;
  assign n30462 = ~n30460 & ~n30461 ;
  assign n30463 = \wishbone_bd_ram_mem1_reg[57][13]/P0001  & n13731 ;
  assign n30464 = \wishbone_bd_ram_mem1_reg[82][13]/P0001  & n13374 ;
  assign n30465 = ~n30463 & ~n30464 ;
  assign n30466 = n30462 & n30465 ;
  assign n30467 = \wishbone_bd_ram_mem1_reg[188][13]/P0001  & n13407 ;
  assign n30468 = \wishbone_bd_ram_mem1_reg[134][13]/P0001  & n13494 ;
  assign n30469 = ~n30467 & ~n30468 ;
  assign n30470 = \wishbone_bd_ram_mem1_reg[37][13]/P0001  & n13710 ;
  assign n30471 = \wishbone_bd_ram_mem1_reg[203][13]/P0001  & n13816 ;
  assign n30472 = ~n30470 & ~n30471 ;
  assign n30473 = n30469 & n30472 ;
  assign n30474 = n30466 & n30473 ;
  assign n30475 = \wishbone_bd_ram_mem1_reg[201][13]/P0001  & n13600 ;
  assign n30476 = \wishbone_bd_ram_mem1_reg[209][13]/P0001  & n13689 ;
  assign n30477 = ~n30475 & ~n30476 ;
  assign n30478 = \wishbone_bd_ram_mem1_reg[29][13]/P0001  & n13412 ;
  assign n30479 = \wishbone_bd_ram_mem1_reg[36][13]/P0001  & n13639 ;
  assign n30480 = ~n30478 & ~n30479 ;
  assign n30481 = n30477 & n30480 ;
  assign n30482 = \wishbone_bd_ram_mem1_reg[154][13]/P0001  & n13403 ;
  assign n30483 = \wishbone_bd_ram_mem1_reg[233][13]/P0001  & n13332 ;
  assign n30484 = ~n30482 & ~n30483 ;
  assign n30485 = \wishbone_bd_ram_mem1_reg[87][13]/P0001  & n13691 ;
  assign n30486 = \wishbone_bd_ram_mem1_reg[179][13]/P0001  & n14035 ;
  assign n30487 = ~n30485 & ~n30486 ;
  assign n30488 = n30484 & n30487 ;
  assign n30489 = n30481 & n30488 ;
  assign n30490 = n30474 & n30489 ;
  assign n30491 = \wishbone_bd_ram_mem1_reg[90][13]/P0001  & n13906 ;
  assign n30492 = \wishbone_bd_ram_mem1_reg[255][13]/P0001  & n13952 ;
  assign n30493 = ~n30491 & ~n30492 ;
  assign n30494 = \wishbone_bd_ram_mem1_reg[177][13]/P0001  & n13863 ;
  assign n30495 = \wishbone_bd_ram_mem1_reg[213][13]/P0001  & n13870 ;
  assign n30496 = ~n30494 & ~n30495 ;
  assign n30497 = n30493 & n30496 ;
  assign n30498 = \wishbone_bd_ram_mem1_reg[184][13]/P0001  & n13960 ;
  assign n30499 = \wishbone_bd_ram_mem1_reg[47][13]/P0001  & n13436 ;
  assign n30500 = ~n30498 & ~n30499 ;
  assign n30501 = \wishbone_bd_ram_mem1_reg[74][13]/P0001  & n13564 ;
  assign n30502 = \wishbone_bd_ram_mem1_reg[84][13]/P0001  & n13385 ;
  assign n30503 = ~n30501 & ~n30502 ;
  assign n30504 = n30500 & n30503 ;
  assign n30505 = n30497 & n30504 ;
  assign n30506 = \wishbone_bd_ram_mem1_reg[30][13]/P0001  & n13713 ;
  assign n30507 = \wishbone_bd_ram_mem1_reg[54][13]/P0001  & n13622 ;
  assign n30508 = ~n30506 & ~n30507 ;
  assign n30509 = \wishbone_bd_ram_mem1_reg[176][13]/P0001  & n13262 ;
  assign n30510 = \wishbone_bd_ram_mem1_reg[175][13]/P0001  & n13674 ;
  assign n30511 = ~n30509 & ~n30510 ;
  assign n30512 = n30508 & n30511 ;
  assign n30513 = \wishbone_bd_ram_mem1_reg[13][13]/P0001  & n13844 ;
  assign n30514 = \wishbone_bd_ram_mem1_reg[143][13]/P0001  & n13461 ;
  assign n30515 = ~n30513 & ~n30514 ;
  assign n30516 = \wishbone_bd_ram_mem1_reg[5][13]/P0001  & n13243 ;
  assign n30517 = \wishbone_bd_ram_mem1_reg[217][13]/P0001  & n13767 ;
  assign n30518 = ~n30516 & ~n30517 ;
  assign n30519 = n30515 & n30518 ;
  assign n30520 = n30512 & n30519 ;
  assign n30521 = n30505 & n30520 ;
  assign n30522 = n30490 & n30521 ;
  assign n30523 = \wishbone_bd_ram_mem1_reg[78][13]/P0001  & n13277 ;
  assign n30524 = \wishbone_bd_ram_mem1_reg[137][13]/P0001  & n13808 ;
  assign n30525 = ~n30523 & ~n30524 ;
  assign n30526 = \wishbone_bd_ram_mem1_reg[115][13]/P0001  & n13747 ;
  assign n30527 = \wishbone_bd_ram_mem1_reg[80][13]/P0001  & n13516 ;
  assign n30528 = ~n30526 & ~n30527 ;
  assign n30529 = n30525 & n30528 ;
  assign n30530 = \wishbone_bd_ram_mem1_reg[182][13]/P0001  & n13598 ;
  assign n30531 = \wishbone_bd_ram_mem1_reg[199][13]/P0001  & n13499 ;
  assign n30532 = ~n30530 & ~n30531 ;
  assign n30533 = \wishbone_bd_ram_mem1_reg[216][13]/P0001  & n14005 ;
  assign n30534 = \wishbone_bd_ram_mem1_reg[146][13]/P0001  & n13958 ;
  assign n30535 = ~n30533 & ~n30534 ;
  assign n30536 = n30532 & n30535 ;
  assign n30537 = n30529 & n30536 ;
  assign n30538 = \wishbone_bd_ram_mem1_reg[44][13]/P0001  & n13291 ;
  assign n30539 = \wishbone_bd_ram_mem1_reg[219][13]/P0001  & n13577 ;
  assign n30540 = ~n30538 & ~n30539 ;
  assign n30541 = \wishbone_bd_ram_mem1_reg[150][13]/P0001  & n13666 ;
  assign n30542 = \wishbone_bd_ram_mem1_reg[194][13]/P0001  & n13624 ;
  assign n30543 = ~n30541 & ~n30542 ;
  assign n30544 = n30540 & n30543 ;
  assign n30545 = \wishbone_bd_ram_mem1_reg[100][13]/P0001  & n13401 ;
  assign n30546 = \wishbone_bd_ram_mem1_reg[229][13]/P0001  & n13552 ;
  assign n30547 = ~n30545 & ~n30546 ;
  assign n30548 = \wishbone_bd_ram_mem1_reg[96][13]/P0001  & n13425 ;
  assign n30549 = \wishbone_bd_ram_mem1_reg[252][13]/P0001  & n13986 ;
  assign n30550 = ~n30548 & ~n30549 ;
  assign n30551 = n30547 & n30550 ;
  assign n30552 = n30544 & n30551 ;
  assign n30553 = n30537 & n30552 ;
  assign n30554 = \wishbone_bd_ram_mem1_reg[232][13]/P0001  & n13510 ;
  assign n30555 = \wishbone_bd_ram_mem1_reg[56][13]/P0001  & n13611 ;
  assign n30556 = ~n30554 & ~n30555 ;
  assign n30557 = \wishbone_bd_ram_mem1_reg[171][13]/P0001  & n13422 ;
  assign n30558 = \wishbone_bd_ram_mem1_reg[38][13]/P0001  & n13828 ;
  assign n30559 = ~n30557 & ~n30558 ;
  assign n30560 = n30556 & n30559 ;
  assign n30561 = \wishbone_bd_ram_mem1_reg[97][13]/P0001  & n13724 ;
  assign n30562 = \wishbone_bd_ram_mem1_reg[95][13]/P0001  & n13317 ;
  assign n30563 = ~n30561 & ~n30562 ;
  assign n30564 = \wishbone_bd_ram_mem1_reg[130][13]/P0001  & n13427 ;
  assign n30565 = \wishbone_bd_ram_mem1_reg[107][13]/P0001  & n13476 ;
  assign n30566 = ~n30564 & ~n30565 ;
  assign n30567 = n30563 & n30566 ;
  assign n30568 = n30560 & n30567 ;
  assign n30569 = \wishbone_bd_ram_mem1_reg[152][13]/P0001  & n13912 ;
  assign n30570 = \wishbone_bd_ram_mem1_reg[145][13]/P0001  & n13715 ;
  assign n30571 = ~n30569 & ~n30570 ;
  assign n30572 = \wishbone_bd_ram_mem1_reg[218][13]/P0001  & n13792 ;
  assign n30573 = \wishbone_bd_ram_mem1_reg[141][13]/P0001  & n13852 ;
  assign n30574 = ~n30572 & ~n30573 ;
  assign n30575 = n30571 & n30574 ;
  assign n30576 = \wishbone_bd_ram_mem1_reg[136][13]/P0001  & n13963 ;
  assign n30577 = \wishbone_bd_ram_mem1_reg[6][13]/P0001  & n13915 ;
  assign n30578 = ~n30576 & ~n30577 ;
  assign n30579 = \wishbone_bd_ram_mem1_reg[180][13]/P0001  & n13650 ;
  assign n30580 = \wishbone_bd_ram_mem1_reg[166][13]/P0001  & n13999 ;
  assign n30581 = ~n30579 & ~n30580 ;
  assign n30582 = n30578 & n30581 ;
  assign n30583 = n30575 & n30582 ;
  assign n30584 = n30568 & n30583 ;
  assign n30585 = n30553 & n30584 ;
  assign n30586 = n30522 & n30585 ;
  assign n30587 = \wishbone_bd_ram_mem1_reg[18][13]/P0001  & n13532 ;
  assign n30588 = \wishbone_bd_ram_mem1_reg[76][13]/P0001  & n13831 ;
  assign n30589 = ~n30587 & ~n30588 ;
  assign n30590 = \wishbone_bd_ram_mem1_reg[224][13]/P0001  & n13433 ;
  assign n30591 = \wishbone_bd_ram_mem1_reg[27][13]/P0001  & n13251 ;
  assign n30592 = ~n30590 & ~n30591 ;
  assign n30593 = n30589 & n30592 ;
  assign n30594 = \wishbone_bd_ram_mem1_reg[102][13]/P0001  & n13534 ;
  assign n30595 = \wishbone_bd_ram_mem1_reg[75][13]/P0001  & n13605 ;
  assign n30596 = ~n30594 & ~n30595 ;
  assign n30597 = \wishbone_bd_ram_mem1_reg[8][13]/P0001  & n13459 ;
  assign n30598 = \wishbone_bd_ram_mem1_reg[21][13]/P0001  & n13438 ;
  assign n30599 = ~n30597 & ~n30598 ;
  assign n30600 = n30596 & n30599 ;
  assign n30601 = n30593 & n30600 ;
  assign n30602 = \wishbone_bd_ram_mem1_reg[45][13]/P0001  & n13420 ;
  assign n30603 = \wishbone_bd_ram_mem1_reg[110][13]/P0001  & n14030 ;
  assign n30604 = ~n30602 & ~n30603 ;
  assign n30605 = \wishbone_bd_ram_mem1_reg[66][13]/P0001  & n13603 ;
  assign n30606 = \wishbone_bd_ram_mem1_reg[170][13]/P0001  & n14007 ;
  assign n30607 = ~n30605 & ~n30606 ;
  assign n30608 = n30604 & n30607 ;
  assign n30609 = \wishbone_bd_ram_mem1_reg[208][13]/P0001  & n14010 ;
  assign n30610 = \wishbone_bd_ram_mem1_reg[79][13]/P0001  & n13779 ;
  assign n30611 = ~n30609 & ~n30610 ;
  assign n30612 = \wishbone_bd_ram_mem1_reg[60][13]/P0001  & n13790 ;
  assign n30613 = \wishbone_bd_ram_mem1_reg[214][13]/P0001  & n13938 ;
  assign n30614 = ~n30612 & ~n30613 ;
  assign n30615 = n30611 & n30614 ;
  assign n30616 = n30608 & n30615 ;
  assign n30617 = n30601 & n30616 ;
  assign n30618 = \wishbone_bd_ram_mem1_reg[34][13]/P0001  & n13450 ;
  assign n30619 = \wishbone_bd_ram_mem1_reg[247][13]/P0001  & n13571 ;
  assign n30620 = ~n30618 & ~n30619 ;
  assign n30621 = \wishbone_bd_ram_mem1_reg[131][13]/P0001  & n13358 ;
  assign n30622 = \wishbone_bd_ram_mem1_reg[158][13]/P0001  & n13294 ;
  assign n30623 = ~n30621 & ~n30622 ;
  assign n30624 = n30620 & n30623 ;
  assign n30625 = \wishbone_bd_ram_mem1_reg[85][13]/P0001  & n13784 ;
  assign n30626 = \wishbone_bd_ram_mem1_reg[103][13]/P0001  & n13320 ;
  assign n30627 = ~n30625 & ~n30626 ;
  assign n30628 = \wishbone_bd_ram_mem1_reg[114][13]/P0001  & n13763 ;
  assign n30629 = \wishbone_bd_ram_mem1_reg[52][13]/P0001  & n13988 ;
  assign n30630 = ~n30628 & ~n30629 ;
  assign n30631 = n30627 & n30630 ;
  assign n30632 = n30624 & n30631 ;
  assign n30633 = \wishbone_bd_ram_mem1_reg[24][13]/P0001  & n13970 ;
  assign n30634 = \wishbone_bd_ram_mem1_reg[138][13]/P0001  & n13398 ;
  assign n30635 = ~n30633 & ~n30634 ;
  assign n30636 = \wishbone_bd_ram_mem1_reg[40][13]/P0001  & n13661 ;
  assign n30637 = \wishbone_bd_ram_mem1_reg[31][13]/P0001  & n13758 ;
  assign n30638 = ~n30636 & ~n30637 ;
  assign n30639 = n30635 & n30638 ;
  assign n30640 = \wishbone_bd_ram_mem1_reg[77][13]/P0001  & n13935 ;
  assign n30641 = \wishbone_bd_ram_mem1_reg[239][13]/P0001  & n13349 ;
  assign n30642 = ~n30640 & ~n30641 ;
  assign n30643 = \wishbone_bd_ram_mem1_reg[42][13]/P0001  & n13341 ;
  assign n30644 = \wishbone_bd_ram_mem1_reg[155][13]/P0001  & n13738 ;
  assign n30645 = ~n30643 & ~n30644 ;
  assign n30646 = n30642 & n30645 ;
  assign n30647 = n30639 & n30646 ;
  assign n30648 = n30632 & n30647 ;
  assign n30649 = n30617 & n30648 ;
  assign n30650 = \wishbone_bd_ram_mem1_reg[178][13]/P0001  & n13301 ;
  assign n30651 = \wishbone_bd_ram_mem1_reg[92][13]/P0001  & n13859 ;
  assign n30652 = ~n30650 & ~n30651 ;
  assign n30653 = \wishbone_bd_ram_mem1_reg[69][13]/P0001  & n13487 ;
  assign n30654 = \wishbone_bd_ram_mem1_reg[191][13]/P0001  & n14012 ;
  assign n30655 = ~n30653 & ~n30654 ;
  assign n30656 = n30652 & n30655 ;
  assign n30657 = \wishbone_bd_ram_mem1_reg[88][13]/P0001  & n13347 ;
  assign n30658 = \wishbone_bd_ram_mem1_reg[109][13]/P0001  & n13306 ;
  assign n30659 = ~n30657 & ~n30658 ;
  assign n30660 = \wishbone_bd_ram_mem1_reg[50][13]/P0001  & n13686 ;
  assign n30661 = \wishbone_bd_ram_mem1_reg[118][13]/P0001  & n13589 ;
  assign n30662 = ~n30660 & ~n30661 ;
  assign n30663 = n30659 & n30662 ;
  assign n30664 = n30656 & n30663 ;
  assign n30665 = \wishbone_bd_ram_mem1_reg[7][13]/P0001  & n13546 ;
  assign n30666 = \wishbone_bd_ram_mem1_reg[12][13]/P0001  & n13733 ;
  assign n30667 = ~n30665 & ~n30666 ;
  assign n30668 = \wishbone_bd_ram_mem1_reg[169][13]/P0001  & n13541 ;
  assign n30669 = \wishbone_bd_ram_mem1_reg[49][13]/P0001  & n13929 ;
  assign n30670 = ~n30668 & ~n30669 ;
  assign n30671 = n30667 & n30670 ;
  assign n30672 = \wishbone_bd_ram_mem1_reg[120][13]/P0001  & n13550 ;
  assign n30673 = \wishbone_bd_ram_mem1_reg[237][13]/P0001  & n13924 ;
  assign n30674 = ~n30672 & ~n30673 ;
  assign n30675 = \wishbone_bd_ram_mem1_reg[116][13]/P0001  & n13865 ;
  assign n30676 = \wishbone_bd_ram_mem1_reg[122][13]/P0001  & n13679 ;
  assign n30677 = ~n30675 & ~n30676 ;
  assign n30678 = n30674 & n30677 ;
  assign n30679 = n30671 & n30678 ;
  assign n30680 = n30664 & n30679 ;
  assign n30681 = \wishbone_bd_ram_mem1_reg[160][13]/P0001  & n13271 ;
  assign n30682 = \wishbone_bd_ram_mem1_reg[167][13]/P0001  & n13940 ;
  assign n30683 = ~n30681 & ~n30682 ;
  assign n30684 = \wishbone_bd_ram_mem1_reg[250][13]/P0001  & n13677 ;
  assign n30685 = \wishbone_bd_ram_mem1_reg[240][13]/P0001  & n13352 ;
  assign n30686 = ~n30684 & ~n30685 ;
  assign n30687 = n30683 & n30686 ;
  assign n30688 = \wishbone_bd_ram_mem1_reg[133][13]/P0001  & n13492 ;
  assign n30689 = \wishbone_bd_ram_mem1_reg[111][13]/P0001  & n13471 ;
  assign n30690 = ~n30688 & ~n30689 ;
  assign n30691 = \wishbone_bd_ram_mem1_reg[206][13]/P0001  & n13414 ;
  assign n30692 = \wishbone_bd_ram_mem1_reg[112][13]/P0001  & n13482 ;
  assign n30693 = ~n30691 & ~n30692 ;
  assign n30694 = n30690 & n30693 ;
  assign n30695 = n30687 & n30694 ;
  assign n30696 = \wishbone_bd_ram_mem1_reg[200][13]/P0001  & n13922 ;
  assign n30697 = \wishbone_bd_ram_mem1_reg[91][13]/P0001  & n13954 ;
  assign n30698 = ~n30696 & ~n30697 ;
  assign n30699 = \wishbone_bd_ram_mem1_reg[101][13]/P0001  & n13772 ;
  assign n30700 = \wishbone_bd_ram_mem1_reg[132][13]/P0001  & n13927 ;
  assign n30701 = ~n30699 & ~n30700 ;
  assign n30702 = n30698 & n30701 ;
  assign n30703 = \wishbone_bd_ram_mem1_reg[220][13]/P0001  & n13965 ;
  assign n30704 = \wishbone_bd_ram_mem1_reg[251][13]/P0001  & n14019 ;
  assign n30705 = ~n30703 & ~n30704 ;
  assign n30706 = \wishbone_bd_ram_mem1_reg[148][13]/P0001  & n13868 ;
  assign n30707 = \wishbone_bd_ram_mem1_reg[108][13]/P0001  & n13814 ;
  assign n30708 = ~n30706 & ~n30707 ;
  assign n30709 = n30705 & n30708 ;
  assign n30710 = n30702 & n30709 ;
  assign n30711 = n30695 & n30710 ;
  assign n30712 = n30680 & n30711 ;
  assign n30713 = n30649 & n30712 ;
  assign n30714 = n30586 & n30713 ;
  assign n30715 = \wishbone_bd_ram_mem1_reg[153][13]/P0001  & n13309 ;
  assign n30716 = \wishbone_bd_ram_mem1_reg[127][13]/P0001  & n13803 ;
  assign n30717 = ~n30715 & ~n30716 ;
  assign n30718 = \wishbone_bd_ram_mem1_reg[55][13]/P0001  & n13618 ;
  assign n30719 = \wishbone_bd_ram_mem1_reg[53][13]/P0001  & n13875 ;
  assign n30720 = ~n30718 & ~n30719 ;
  assign n30721 = n30717 & n30720 ;
  assign n30722 = \wishbone_bd_ram_mem1_reg[68][13]/P0001  & n13379 ;
  assign n30723 = \wishbone_bd_ram_mem1_reg[17][13]/P0001  & n13324 ;
  assign n30724 = ~n30722 & ~n30723 ;
  assign n30725 = \wishbone_bd_ram_mem1_reg[249][13]/P0001  & n13431 ;
  assign n30726 = \wishbone_bd_ram_mem1_reg[19][13]/P0001  & n13886 ;
  assign n30727 = ~n30725 & ~n30726 ;
  assign n30728 = n30724 & n30727 ;
  assign n30729 = n30721 & n30728 ;
  assign n30730 = \wishbone_bd_ram_mem1_reg[161][13]/P0001  & n13505 ;
  assign n30731 = \wishbone_bd_ram_mem1_reg[20][13]/P0001  & n13839 ;
  assign n30732 = ~n30730 & ~n30731 ;
  assign n30733 = \wishbone_bd_ram_mem1_reg[86][13]/P0001  & n13485 ;
  assign n30734 = \wishbone_bd_ram_mem1_reg[227][13]/P0001  & n13388 ;
  assign n30735 = ~n30733 & ~n30734 ;
  assign n30736 = n30732 & n30735 ;
  assign n30737 = \wishbone_bd_ram_mem1_reg[104][13]/P0001  & n13684 ;
  assign n30738 = \wishbone_bd_ram_mem1_reg[62][13]/P0001  & n13529 ;
  assign n30739 = ~n30737 & ~n30738 ;
  assign n30740 = \wishbone_bd_ram_mem1_reg[41][13]/P0001  & n14017 ;
  assign n30741 = \wishbone_bd_ram_mem1_reg[117][13]/P0001  & n13557 ;
  assign n30742 = ~n30740 & ~n30741 ;
  assign n30743 = n30739 & n30742 ;
  assign n30744 = n30736 & n30743 ;
  assign n30745 = n30729 & n30744 ;
  assign n30746 = \wishbone_bd_ram_mem1_reg[172][13]/P0001  & n13377 ;
  assign n30747 = \wishbone_bd_ram_mem1_reg[26][13]/P0001  & n13521 ;
  assign n30748 = ~n30746 & ~n30747 ;
  assign n30749 = \wishbone_bd_ram_mem1_reg[164][13]/P0001  & n13236 ;
  assign n30750 = \wishbone_bd_ram_mem1_reg[3][13]/P0001  & n13354 ;
  assign n30751 = ~n30749 & ~n30750 ;
  assign n30752 = n30748 & n30751 ;
  assign n30753 = \wishbone_bd_ram_mem1_reg[187][13]/P0001  & n13756 ;
  assign n30754 = \wishbone_bd_ram_mem1_reg[10][13]/P0001  & n13837 ;
  assign n30755 = ~n30753 & ~n30754 ;
  assign n30756 = \wishbone_bd_ram_mem1_reg[94][13]/P0001  & n13833 ;
  assign n30757 = \wishbone_bd_ram_mem1_reg[234][13]/P0001  & n13781 ;
  assign n30758 = ~n30756 & ~n30757 ;
  assign n30759 = n30755 & n30758 ;
  assign n30760 = n30752 & n30759 ;
  assign n30761 = \wishbone_bd_ram_mem1_reg[39][13]/P0001  & n13893 ;
  assign n30762 = \wishbone_bd_ram_mem1_reg[113][13]/P0001  & n13882 ;
  assign n30763 = ~n30761 & ~n30762 ;
  assign n30764 = \wishbone_bd_ram_mem1_reg[168][13]/P0001  & n13795 ;
  assign n30765 = \wishbone_bd_ram_mem1_reg[22][13]/P0001  & n13744 ;
  assign n30766 = ~n30764 & ~n30765 ;
  assign n30767 = n30763 & n30766 ;
  assign n30768 = \wishbone_bd_ram_mem1_reg[195][13]/P0001  & n13700 ;
  assign n30769 = \wishbone_bd_ram_mem1_reg[70][13]/P0001  & n13339 ;
  assign n30770 = ~n30768 & ~n30769 ;
  assign n30771 = \wishbone_bd_ram_mem1_reg[165][13]/P0001  & n14028 ;
  assign n30772 = \wishbone_bd_ram_mem1_reg[71][13]/P0001  & n13636 ;
  assign n30773 = ~n30771 & ~n30772 ;
  assign n30774 = n30770 & n30773 ;
  assign n30775 = n30767 & n30774 ;
  assign n30776 = n30760 & n30775 ;
  assign n30777 = n30745 & n30776 ;
  assign n30778 = \wishbone_bd_ram_mem1_reg[81][13]/P0001  & n13409 ;
  assign n30779 = \wishbone_bd_ram_mem1_reg[253][13]/P0001  & n13708 ;
  assign n30780 = ~n30778 & ~n30779 ;
  assign n30781 = \wishbone_bd_ram_mem1_reg[197][13]/P0001  & n13594 ;
  assign n30782 = \wishbone_bd_ram_mem1_reg[174][13]/P0001  & n13899 ;
  assign n30783 = ~n30781 & ~n30782 ;
  assign n30784 = n30780 & n30783 ;
  assign n30785 = \wishbone_bd_ram_mem1_reg[93][13]/P0001  & n13891 ;
  assign n30786 = \wishbone_bd_ram_mem1_reg[125][13]/P0001  & n13396 ;
  assign n30787 = ~n30785 & ~n30786 ;
  assign n30788 = \wishbone_bd_ram_mem1_reg[63][13]/P0001  & n13327 ;
  assign n30789 = \wishbone_bd_ram_mem1_reg[246][13]/P0001  & n13981 ;
  assign n30790 = ~n30788 & ~n30789 ;
  assign n30791 = n30787 & n30790 ;
  assign n30792 = n30784 & n30791 ;
  assign n30793 = \wishbone_bd_ram_mem1_reg[135][13]/P0001  & n13672 ;
  assign n30794 = \wishbone_bd_ram_mem1_reg[59][13]/P0001  & n13613 ;
  assign n30795 = ~n30793 & ~n30794 ;
  assign n30796 = \wishbone_bd_ram_mem1_reg[61][13]/P0001  & n13544 ;
  assign n30797 = \wishbone_bd_ram_mem1_reg[235][13]/P0001  & n13518 ;
  assign n30798 = ~n30796 & ~n30797 ;
  assign n30799 = n30795 & n30798 ;
  assign n30800 = \wishbone_bd_ram_mem1_reg[149][13]/P0001  & n13469 ;
  assign n30801 = \wishbone_bd_ram_mem1_reg[222][13]/P0001  & n13721 ;
  assign n30802 = ~n30800 & ~n30801 ;
  assign n30803 = \wishbone_bd_ram_mem1_reg[99][13]/P0001  & n13996 ;
  assign n30804 = \wishbone_bd_ram_mem1_reg[248][13]/P0001  & n13647 ;
  assign n30805 = ~n30803 & ~n30804 ;
  assign n30806 = n30802 & n30805 ;
  assign n30807 = n30799 & n30806 ;
  assign n30808 = n30792 & n30807 ;
  assign n30809 = \wishbone_bd_ram_mem1_reg[211][13]/P0001  & n13805 ;
  assign n30810 = \wishbone_bd_ram_mem1_reg[156][13]/P0001  & n13769 ;
  assign n30811 = ~n30809 & ~n30810 ;
  assign n30812 = \wishbone_bd_ram_mem1_reg[142][13]/P0001  & n13448 ;
  assign n30813 = \wishbone_bd_ram_mem1_reg[51][13]/P0001  & n13880 ;
  assign n30814 = ~n30812 & ~n30813 ;
  assign n30815 = n30811 & n30814 ;
  assign n30816 = \wishbone_bd_ram_mem1_reg[72][13]/P0001  & n13582 ;
  assign n30817 = \wishbone_bd_ram_mem1_reg[223][13]/P0001  & n13335 ;
  assign n30818 = ~n30816 & ~n30817 ;
  assign n30819 = \wishbone_bd_ram_mem1_reg[207][13]/P0001  & n13826 ;
  assign n30820 = \wishbone_bd_ram_mem1_reg[242][13]/P0001  & n13383 ;
  assign n30821 = ~n30819 & ~n30820 ;
  assign n30822 = n30818 & n30821 ;
  assign n30823 = n30815 & n30822 ;
  assign n30824 = \wishbone_bd_ram_mem1_reg[221][13]/P0001  & n13641 ;
  assign n30825 = \wishbone_bd_ram_mem1_reg[230][13]/P0001  & n13994 ;
  assign n30826 = ~n30824 & ~n30825 ;
  assign n30827 = \wishbone_bd_ram_mem1_reg[35][13]/P0001  & n13523 ;
  assign n30828 = \wishbone_bd_ram_mem1_reg[241][13]/P0001  & n13854 ;
  assign n30829 = ~n30827 & ~n30828 ;
  assign n30830 = n30826 & n30829 ;
  assign n30831 = \wishbone_bd_ram_mem1_reg[215][13]/P0001  & n13901 ;
  assign n30832 = \wishbone_bd_ram_mem1_reg[64][13]/P0001  & n13904 ;
  assign n30833 = ~n30831 & ~n30832 ;
  assign n30834 = \wishbone_bd_ram_mem1_reg[1][13]/P0001  & n13888 ;
  assign n30835 = \wishbone_bd_ram_mem1_reg[58][13]/P0001  & n13949 ;
  assign n30836 = ~n30834 & ~n30835 ;
  assign n30837 = n30833 & n30836 ;
  assign n30838 = n30830 & n30837 ;
  assign n30839 = n30823 & n30838 ;
  assign n30840 = n30808 & n30839 ;
  assign n30841 = n30777 & n30840 ;
  assign n30842 = \wishbone_bd_ram_mem1_reg[157][13]/P0001  & n13445 ;
  assign n30843 = \wishbone_bd_ram_mem1_reg[186][13]/P0001  & n13616 ;
  assign n30844 = ~n30842 & ~n30843 ;
  assign n30845 = \wishbone_bd_ram_mem1_reg[105][13]/P0001  & n13503 ;
  assign n30846 = \wishbone_bd_ram_mem1_reg[245][13]/P0001  & n13877 ;
  assign n30847 = ~n30845 & ~n30846 ;
  assign n30848 = n30844 & n30847 ;
  assign n30849 = \wishbone_bd_ram_mem1_reg[33][13]/P0001  & n13933 ;
  assign n30850 = \wishbone_bd_ram_mem1_reg[162][13]/P0001  & n13726 ;
  assign n30851 = ~n30849 & ~n30850 ;
  assign n30852 = \wishbone_bd_ram_mem1_reg[2][13]/P0001  & n13975 ;
  assign n30853 = \wishbone_bd_ram_mem1_reg[238][13]/P0001  & n13819 ;
  assign n30854 = ~n30852 & ~n30853 ;
  assign n30855 = n30851 & n30854 ;
  assign n30856 = n30848 & n30855 ;
  assign n30857 = \wishbone_bd_ram_mem1_reg[23][13]/P0001  & n13857 ;
  assign n30858 = \wishbone_bd_ram_mem1_reg[124][13]/P0001  & n14024 ;
  assign n30859 = ~n30857 & ~n30858 ;
  assign n30860 = \wishbone_bd_ram_mem1_reg[123][13]/P0001  & n13749 ;
  assign n30861 = \wishbone_bd_ram_mem1_reg[0][13]/P0001  & n13539 ;
  assign n30862 = ~n30860 & ~n30861 ;
  assign n30863 = n30859 & n30862 ;
  assign n30864 = \wishbone_bd_ram_mem1_reg[181][13]/P0001  & n13587 ;
  assign n30865 = \wishbone_bd_ram_mem1_reg[9][13]/P0001  & n13580 ;
  assign n30866 = ~n30864 & ~n30865 ;
  assign n30867 = \wishbone_bd_ram_mem1_reg[14][13]/P0001  & n13972 ;
  assign n30868 = \wishbone_bd_ram_mem1_reg[212][13]/P0001  & n13634 ;
  assign n30869 = ~n30867 & ~n30868 ;
  assign n30870 = n30866 & n30869 ;
  assign n30871 = n30863 & n30870 ;
  assign n30872 = n30856 & n30871 ;
  assign n30873 = \wishbone_bd_ram_mem1_reg[144][13]/P0001  & n13508 ;
  assign n30874 = \wishbone_bd_ram_mem1_reg[25][13]/P0001  & n13742 ;
  assign n30875 = ~n30873 & ~n30874 ;
  assign n30876 = \wishbone_bd_ram_mem1_reg[89][13]/P0001  & n13910 ;
  assign n30877 = \wishbone_bd_ram_mem1_reg[192][13]/P0001  & n13390 ;
  assign n30878 = ~n30876 & ~n30877 ;
  assign n30879 = n30875 & n30878 ;
  assign n30880 = \wishbone_bd_ram_mem1_reg[151][13]/P0001  & n13697 ;
  assign n30881 = \wishbone_bd_ram_mem1_reg[11][13]/P0001  & n13774 ;
  assign n30882 = ~n30880 & ~n30881 ;
  assign n30883 = \wishbone_bd_ram_mem1_reg[28][13]/P0001  & n13810 ;
  assign n30884 = \wishbone_bd_ram_mem1_reg[226][13]/P0001  & n13668 ;
  assign n30885 = ~n30883 & ~n30884 ;
  assign n30886 = n30882 & n30885 ;
  assign n30887 = n30879 & n30886 ;
  assign n30888 = \wishbone_bd_ram_mem1_reg[183][13]/P0001  & n13645 ;
  assign n30889 = \wishbone_bd_ram_mem1_reg[15][13]/P0001  & n13797 ;
  assign n30890 = ~n30888 & ~n30889 ;
  assign n30891 = \wishbone_bd_ram_mem1_reg[32][13]/P0001  & n13736 ;
  assign n30892 = \wishbone_bd_ram_mem1_reg[16][13]/P0001  & n13695 ;
  assign n30893 = ~n30891 & ~n30892 ;
  assign n30894 = n30890 & n30893 ;
  assign n30895 = \wishbone_bd_ram_mem1_reg[128][13]/P0001  & n13652 ;
  assign n30896 = \wishbone_bd_ram_mem1_reg[236][13]/P0001  & n13480 ;
  assign n30897 = ~n30895 & ~n30896 ;
  assign n30898 = \wishbone_bd_ram_mem1_reg[198][13]/P0001  & n13592 ;
  assign n30899 = \wishbone_bd_ram_mem1_reg[147][13]/P0001  & n13702 ;
  assign n30900 = ~n30898 & ~n30899 ;
  assign n30901 = n30897 & n30900 ;
  assign n30902 = n30894 & n30901 ;
  assign n30903 = n30887 & n30902 ;
  assign n30904 = n30872 & n30903 ;
  assign n30905 = \wishbone_bd_ram_mem1_reg[140][13]/P0001  & n13287 ;
  assign n30906 = \wishbone_bd_ram_mem1_reg[67][13]/P0001  & n13663 ;
  assign n30907 = ~n30905 & ~n30906 ;
  assign n30908 = \wishbone_bd_ram_mem1_reg[185][13]/P0001  & n13372 ;
  assign n30909 = \wishbone_bd_ram_mem1_reg[202][13]/P0001  & n13268 ;
  assign n30910 = ~n30908 & ~n30909 ;
  assign n30911 = n30907 & n30910 ;
  assign n30912 = \wishbone_bd_ram_mem1_reg[244][13]/P0001  & n13474 ;
  assign n30913 = \wishbone_bd_ram_mem1_reg[228][13]/P0001  & n13497 ;
  assign n30914 = ~n30912 & ~n30913 ;
  assign n30915 = \wishbone_bd_ram_mem1_reg[163][13]/P0001  & n13255 ;
  assign n30916 = \wishbone_bd_ram_mem1_reg[121][13]/P0001  & n13983 ;
  assign n30917 = ~n30915 & ~n30916 ;
  assign n30918 = n30914 & n30917 ;
  assign n30919 = n30911 & n30918 ;
  assign n30920 = \wishbone_bd_ram_mem1_reg[243][13]/P0001  & n13575 ;
  assign n30921 = \wishbone_bd_ram_mem1_reg[210][13]/P0001  & n13443 ;
  assign n30922 = ~n30920 & ~n30921 ;
  assign n30923 = \wishbone_bd_ram_mem1_reg[205][13]/P0001  & n13947 ;
  assign n30924 = \wishbone_bd_ram_mem1_reg[48][13]/P0001  & n13917 ;
  assign n30925 = ~n30923 & ~n30924 ;
  assign n30926 = n30922 & n30925 ;
  assign n30927 = \wishbone_bd_ram_mem1_reg[190][13]/P0001  & n13365 ;
  assign n30928 = \wishbone_bd_ram_mem1_reg[4][13]/P0001  & n13527 ;
  assign n30929 = ~n30927 & ~n30928 ;
  assign n30930 = \wishbone_bd_ram_mem1_reg[193][13]/P0001  & n14022 ;
  assign n30931 = \wishbone_bd_ram_mem1_reg[204][13]/P0001  & n13821 ;
  assign n30932 = ~n30930 & ~n30931 ;
  assign n30933 = n30929 & n30932 ;
  assign n30934 = n30926 & n30933 ;
  assign n30935 = n30919 & n30934 ;
  assign n30936 = \wishbone_bd_ram_mem1_reg[173][13]/P0001  & n13360 ;
  assign n30937 = \wishbone_bd_ram_mem1_reg[46][13]/P0001  & n13298 ;
  assign n30938 = ~n30936 & ~n30937 ;
  assign n30939 = \wishbone_bd_ram_mem1_reg[119][13]/P0001  & n14033 ;
  assign n30940 = \wishbone_bd_ram_mem1_reg[43][13]/P0001  & n13761 ;
  assign n30941 = ~n30939 & ~n30940 ;
  assign n30942 = n30938 & n30941 ;
  assign n30943 = \wishbone_bd_ram_mem1_reg[196][13]/P0001  & n13977 ;
  assign n30944 = \wishbone_bd_ram_mem1_reg[189][13]/P0001  & n14001 ;
  assign n30945 = ~n30943 & ~n30944 ;
  assign n30946 = \wishbone_bd_ram_mem1_reg[83][13]/P0001  & n13454 ;
  assign n30947 = \wishbone_bd_ram_mem1_reg[231][13]/P0001  & n13363 ;
  assign n30948 = ~n30946 & ~n30947 ;
  assign n30949 = n30945 & n30948 ;
  assign n30950 = n30942 & n30949 ;
  assign n30951 = \wishbone_bd_ram_mem1_reg[129][13]/P0001  & n13629 ;
  assign n30952 = \wishbone_bd_ram_mem1_reg[254][13]/P0001  & n13283 ;
  assign n30953 = ~n30951 & ~n30952 ;
  assign n30954 = \wishbone_bd_ram_mem1_reg[139][13]/P0001  & n13566 ;
  assign n30955 = \wishbone_bd_ram_mem1_reg[159][13]/P0001  & n13627 ;
  assign n30956 = ~n30954 & ~n30955 ;
  assign n30957 = n30953 & n30956 ;
  assign n30958 = \wishbone_bd_ram_mem1_reg[73][13]/P0001  & n13456 ;
  assign n30959 = \wishbone_bd_ram_mem1_reg[225][13]/P0001  & n13719 ;
  assign n30960 = ~n30958 & ~n30959 ;
  assign n30961 = \wishbone_bd_ram_mem1_reg[106][13]/P0001  & n13555 ;
  assign n30962 = \wishbone_bd_ram_mem1_reg[98][13]/P0001  & n13569 ;
  assign n30963 = ~n30961 & ~n30962 ;
  assign n30964 = n30960 & n30963 ;
  assign n30965 = n30957 & n30964 ;
  assign n30966 = n30950 & n30965 ;
  assign n30967 = n30935 & n30966 ;
  assign n30968 = n30904 & n30967 ;
  assign n30969 = n30841 & n30968 ;
  assign n30970 = n30714 & n30969 ;
  assign n30971 = ~wb_rst_i_pad & ~n30458 ;
  assign n30972 = ~n30970 & n30971 ;
  assign n30973 = ~n30459 & ~n30972 ;
  assign n30974 = \ethreg1_MODER_1_DataOut_reg[6]/NET0131  & n23808 ;
  assign n30975 = \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131  & n23794 ;
  assign n30976 = n23741 & n30975 ;
  assign n30977 = ~n30974 & ~n30976 ;
  assign n30978 = \ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131  & n23743 ;
  assign n30979 = n23741 & n30978 ;
  assign n30980 = \ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131  & n23743 ;
  assign n30981 = n23747 & n30980 ;
  assign n30982 = ~n30979 & ~n30981 ;
  assign n30983 = n30977 & n30982 ;
  assign n30984 = n23730 & n30983 ;
  assign n30985 = \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  & n23737 ;
  assign n30986 = \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131  & n23813 ;
  assign n30987 = \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  & n23751 ;
  assign n30988 = n23741 & n30987 ;
  assign n30989 = ~n30986 & ~n30988 ;
  assign n30990 = \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  & n23751 ;
  assign n30991 = n23747 & n30990 ;
  assign n30992 = \ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131  & n23782 ;
  assign n30993 = ~n30991 & ~n30992 ;
  assign n30994 = n30989 & n30993 ;
  assign n30995 = ~n30985 & n30994 ;
  assign n30996 = n30984 & n30995 ;
  assign n30997 = n23730 & ~n30996 ;
  assign n30998 = \wishbone_bd_ram_mem1_reg[107][14]/P0001  & n13476 ;
  assign n30999 = \wishbone_bd_ram_mem1_reg[95][14]/P0001  & n13317 ;
  assign n31000 = ~n30998 & ~n30999 ;
  assign n31001 = \wishbone_bd_ram_mem1_reg[164][14]/P0001  & n13236 ;
  assign n31002 = \wishbone_bd_ram_mem1_reg[207][14]/P0001  & n13826 ;
  assign n31003 = ~n31001 & ~n31002 ;
  assign n31004 = n31000 & n31003 ;
  assign n31005 = \wishbone_bd_ram_mem1_reg[198][14]/P0001  & n13592 ;
  assign n31006 = \wishbone_bd_ram_mem1_reg[137][14]/P0001  & n13808 ;
  assign n31007 = ~n31005 & ~n31006 ;
  assign n31008 = \wishbone_bd_ram_mem1_reg[4][14]/P0001  & n13527 ;
  assign n31009 = \wishbone_bd_ram_mem1_reg[220][14]/P0001  & n13965 ;
  assign n31010 = ~n31008 & ~n31009 ;
  assign n31011 = n31007 & n31010 ;
  assign n31012 = n31004 & n31011 ;
  assign n31013 = \wishbone_bd_ram_mem1_reg[206][14]/P0001  & n13414 ;
  assign n31014 = \wishbone_bd_ram_mem1_reg[140][14]/P0001  & n13287 ;
  assign n31015 = ~n31013 & ~n31014 ;
  assign n31016 = \wishbone_bd_ram_mem1_reg[2][14]/P0001  & n13975 ;
  assign n31017 = \wishbone_bd_ram_mem1_reg[112][14]/P0001  & n13482 ;
  assign n31018 = ~n31016 & ~n31017 ;
  assign n31019 = n31015 & n31018 ;
  assign n31020 = \wishbone_bd_ram_mem1_reg[45][14]/P0001  & n13420 ;
  assign n31021 = \wishbone_bd_ram_mem1_reg[202][14]/P0001  & n13268 ;
  assign n31022 = ~n31020 & ~n31021 ;
  assign n31023 = \wishbone_bd_ram_mem1_reg[76][14]/P0001  & n13831 ;
  assign n31024 = \wishbone_bd_ram_mem1_reg[170][14]/P0001  & n14007 ;
  assign n31025 = ~n31023 & ~n31024 ;
  assign n31026 = n31022 & n31025 ;
  assign n31027 = n31019 & n31026 ;
  assign n31028 = n31012 & n31027 ;
  assign n31029 = \wishbone_bd_ram_mem1_reg[0][14]/P0001  & n13539 ;
  assign n31030 = \wishbone_bd_ram_mem1_reg[56][14]/P0001  & n13611 ;
  assign n31031 = ~n31029 & ~n31030 ;
  assign n31032 = \wishbone_bd_ram_mem1_reg[247][14]/P0001  & n13571 ;
  assign n31033 = \wishbone_bd_ram_mem1_reg[101][14]/P0001  & n13772 ;
  assign n31034 = ~n31032 & ~n31033 ;
  assign n31035 = n31031 & n31034 ;
  assign n31036 = \wishbone_bd_ram_mem1_reg[114][14]/P0001  & n13763 ;
  assign n31037 = \wishbone_bd_ram_mem1_reg[209][14]/P0001  & n13689 ;
  assign n31038 = ~n31036 & ~n31037 ;
  assign n31039 = \wishbone_bd_ram_mem1_reg[28][14]/P0001  & n13810 ;
  assign n31040 = \wishbone_bd_ram_mem1_reg[69][14]/P0001  & n13487 ;
  assign n31041 = ~n31039 & ~n31040 ;
  assign n31042 = n31038 & n31041 ;
  assign n31043 = n31035 & n31042 ;
  assign n31044 = \wishbone_bd_ram_mem1_reg[177][14]/P0001  & n13863 ;
  assign n31045 = \wishbone_bd_ram_mem1_reg[217][14]/P0001  & n13767 ;
  assign n31046 = ~n31044 & ~n31045 ;
  assign n31047 = \wishbone_bd_ram_mem1_reg[194][14]/P0001  & n13624 ;
  assign n31048 = \wishbone_bd_ram_mem1_reg[255][14]/P0001  & n13952 ;
  assign n31049 = ~n31047 & ~n31048 ;
  assign n31050 = n31046 & n31049 ;
  assign n31051 = \wishbone_bd_ram_mem1_reg[242][14]/P0001  & n13383 ;
  assign n31052 = \wishbone_bd_ram_mem1_reg[223][14]/P0001  & n13335 ;
  assign n31053 = ~n31051 & ~n31052 ;
  assign n31054 = \wishbone_bd_ram_mem1_reg[214][14]/P0001  & n13938 ;
  assign n31055 = \wishbone_bd_ram_mem1_reg[190][14]/P0001  & n13365 ;
  assign n31056 = ~n31054 & ~n31055 ;
  assign n31057 = n31053 & n31056 ;
  assign n31058 = n31050 & n31057 ;
  assign n31059 = n31043 & n31058 ;
  assign n31060 = n31028 & n31059 ;
  assign n31061 = \wishbone_bd_ram_mem1_reg[224][14]/P0001  & n13433 ;
  assign n31062 = \wishbone_bd_ram_mem1_reg[41][14]/P0001  & n14017 ;
  assign n31063 = ~n31061 & ~n31062 ;
  assign n31064 = \wishbone_bd_ram_mem1_reg[195][14]/P0001  & n13700 ;
  assign n31065 = \wishbone_bd_ram_mem1_reg[183][14]/P0001  & n13645 ;
  assign n31066 = ~n31064 & ~n31065 ;
  assign n31067 = n31063 & n31066 ;
  assign n31068 = \wishbone_bd_ram_mem1_reg[205][14]/P0001  & n13947 ;
  assign n31069 = \wishbone_bd_ram_mem1_reg[12][14]/P0001  & n13733 ;
  assign n31070 = ~n31068 & ~n31069 ;
  assign n31071 = \wishbone_bd_ram_mem1_reg[253][14]/P0001  & n13708 ;
  assign n31072 = \wishbone_bd_ram_mem1_reg[156][14]/P0001  & n13769 ;
  assign n31073 = ~n31071 & ~n31072 ;
  assign n31074 = n31070 & n31073 ;
  assign n31075 = n31067 & n31074 ;
  assign n31076 = \wishbone_bd_ram_mem1_reg[131][14]/P0001  & n13358 ;
  assign n31077 = \wishbone_bd_ram_mem1_reg[73][14]/P0001  & n13456 ;
  assign n31078 = ~n31076 & ~n31077 ;
  assign n31079 = \wishbone_bd_ram_mem1_reg[31][14]/P0001  & n13758 ;
  assign n31080 = \wishbone_bd_ram_mem1_reg[216][14]/P0001  & n14005 ;
  assign n31081 = ~n31079 & ~n31080 ;
  assign n31082 = n31078 & n31081 ;
  assign n31083 = \wishbone_bd_ram_mem1_reg[231][14]/P0001  & n13363 ;
  assign n31084 = \wishbone_bd_ram_mem1_reg[221][14]/P0001  & n13641 ;
  assign n31085 = ~n31083 & ~n31084 ;
  assign n31086 = \wishbone_bd_ram_mem1_reg[13][14]/P0001  & n13844 ;
  assign n31087 = \wishbone_bd_ram_mem1_reg[238][14]/P0001  & n13819 ;
  assign n31088 = ~n31086 & ~n31087 ;
  assign n31089 = n31085 & n31088 ;
  assign n31090 = n31082 & n31089 ;
  assign n31091 = n31075 & n31090 ;
  assign n31092 = \wishbone_bd_ram_mem1_reg[123][14]/P0001  & n13749 ;
  assign n31093 = \wishbone_bd_ram_mem1_reg[189][14]/P0001  & n14001 ;
  assign n31094 = ~n31092 & ~n31093 ;
  assign n31095 = \wishbone_bd_ram_mem1_reg[146][14]/P0001  & n13958 ;
  assign n31096 = \wishbone_bd_ram_mem1_reg[72][14]/P0001  & n13582 ;
  assign n31097 = ~n31095 & ~n31096 ;
  assign n31098 = n31094 & n31097 ;
  assign n31099 = \wishbone_bd_ram_mem1_reg[248][14]/P0001  & n13647 ;
  assign n31100 = \wishbone_bd_ram_mem1_reg[126][14]/P0001  & n13786 ;
  assign n31101 = ~n31099 & ~n31100 ;
  assign n31102 = \wishbone_bd_ram_mem1_reg[8][14]/P0001  & n13459 ;
  assign n31103 = \wishbone_bd_ram_mem1_reg[218][14]/P0001  & n13792 ;
  assign n31104 = ~n31102 & ~n31103 ;
  assign n31105 = n31101 & n31104 ;
  assign n31106 = n31098 & n31105 ;
  assign n31107 = \wishbone_bd_ram_mem1_reg[98][14]/P0001  & n13569 ;
  assign n31108 = \wishbone_bd_ram_mem1_reg[172][14]/P0001  & n13377 ;
  assign n31109 = ~n31107 & ~n31108 ;
  assign n31110 = \wishbone_bd_ram_mem1_reg[53][14]/P0001  & n13875 ;
  assign n31111 = \wishbone_bd_ram_mem1_reg[148][14]/P0001  & n13868 ;
  assign n31112 = ~n31110 & ~n31111 ;
  assign n31113 = n31109 & n31112 ;
  assign n31114 = \wishbone_bd_ram_mem1_reg[134][14]/P0001  & n13494 ;
  assign n31115 = \wishbone_bd_ram_mem1_reg[54][14]/P0001  & n13622 ;
  assign n31116 = ~n31114 & ~n31115 ;
  assign n31117 = \wishbone_bd_ram_mem1_reg[203][14]/P0001  & n13816 ;
  assign n31118 = \wishbone_bd_ram_mem1_reg[230][14]/P0001  & n13994 ;
  assign n31119 = ~n31117 & ~n31118 ;
  assign n31120 = n31116 & n31119 ;
  assign n31121 = n31113 & n31120 ;
  assign n31122 = n31106 & n31121 ;
  assign n31123 = n31091 & n31122 ;
  assign n31124 = n31060 & n31123 ;
  assign n31125 = \wishbone_bd_ram_mem1_reg[68][14]/P0001  & n13379 ;
  assign n31126 = \wishbone_bd_ram_mem1_reg[132][14]/P0001  & n13927 ;
  assign n31127 = ~n31125 & ~n31126 ;
  assign n31128 = \wishbone_bd_ram_mem1_reg[87][14]/P0001  & n13691 ;
  assign n31129 = \wishbone_bd_ram_mem1_reg[108][14]/P0001  & n13814 ;
  assign n31130 = ~n31128 & ~n31129 ;
  assign n31131 = n31127 & n31130 ;
  assign n31132 = \wishbone_bd_ram_mem1_reg[197][14]/P0001  & n13594 ;
  assign n31133 = \wishbone_bd_ram_mem1_reg[222][14]/P0001  & n13721 ;
  assign n31134 = ~n31132 & ~n31133 ;
  assign n31135 = \wishbone_bd_ram_mem1_reg[16][14]/P0001  & n13695 ;
  assign n31136 = \wishbone_bd_ram_mem1_reg[135][14]/P0001  & n13672 ;
  assign n31137 = ~n31135 & ~n31136 ;
  assign n31138 = n31134 & n31137 ;
  assign n31139 = n31131 & n31138 ;
  assign n31140 = \wishbone_bd_ram_mem1_reg[75][14]/P0001  & n13605 ;
  assign n31141 = \wishbone_bd_ram_mem1_reg[70][14]/P0001  & n13339 ;
  assign n31142 = ~n31140 & ~n31141 ;
  assign n31143 = \wishbone_bd_ram_mem1_reg[155][14]/P0001  & n13738 ;
  assign n31144 = \wishbone_bd_ram_mem1_reg[243][14]/P0001  & n13575 ;
  assign n31145 = ~n31143 & ~n31144 ;
  assign n31146 = n31142 & n31145 ;
  assign n31147 = \wishbone_bd_ram_mem1_reg[210][14]/P0001  & n13443 ;
  assign n31148 = \wishbone_bd_ram_mem1_reg[85][14]/P0001  & n13784 ;
  assign n31149 = ~n31147 & ~n31148 ;
  assign n31150 = \wishbone_bd_ram_mem1_reg[50][14]/P0001  & n13686 ;
  assign n31151 = \wishbone_bd_ram_mem1_reg[176][14]/P0001  & n13262 ;
  assign n31152 = ~n31150 & ~n31151 ;
  assign n31153 = n31149 & n31152 ;
  assign n31154 = n31146 & n31153 ;
  assign n31155 = n31139 & n31154 ;
  assign n31156 = \wishbone_bd_ram_mem1_reg[33][14]/P0001  & n13933 ;
  assign n31157 = \wishbone_bd_ram_mem1_reg[113][14]/P0001  & n13882 ;
  assign n31158 = ~n31156 & ~n31157 ;
  assign n31159 = \wishbone_bd_ram_mem1_reg[44][14]/P0001  & n13291 ;
  assign n31160 = \wishbone_bd_ram_mem1_reg[237][14]/P0001  & n13924 ;
  assign n31161 = ~n31159 & ~n31160 ;
  assign n31162 = n31158 & n31161 ;
  assign n31163 = \wishbone_bd_ram_mem1_reg[18][14]/P0001  & n13532 ;
  assign n31164 = \wishbone_bd_ram_mem1_reg[58][14]/P0001  & n13949 ;
  assign n31165 = ~n31163 & ~n31164 ;
  assign n31166 = \wishbone_bd_ram_mem1_reg[171][14]/P0001  & n13422 ;
  assign n31167 = \wishbone_bd_ram_mem1_reg[118][14]/P0001  & n13589 ;
  assign n31168 = ~n31166 & ~n31167 ;
  assign n31169 = n31165 & n31168 ;
  assign n31170 = n31162 & n31169 ;
  assign n31171 = \wishbone_bd_ram_mem1_reg[78][14]/P0001  & n13277 ;
  assign n31172 = \wishbone_bd_ram_mem1_reg[46][14]/P0001  & n13298 ;
  assign n31173 = ~n31171 & ~n31172 ;
  assign n31174 = \wishbone_bd_ram_mem1_reg[157][14]/P0001  & n13445 ;
  assign n31175 = \wishbone_bd_ram_mem1_reg[81][14]/P0001  & n13409 ;
  assign n31176 = ~n31174 & ~n31175 ;
  assign n31177 = n31173 & n31176 ;
  assign n31178 = \wishbone_bd_ram_mem1_reg[29][14]/P0001  & n13412 ;
  assign n31179 = \wishbone_bd_ram_mem1_reg[241][14]/P0001  & n13854 ;
  assign n31180 = ~n31178 & ~n31179 ;
  assign n31181 = \wishbone_bd_ram_mem1_reg[211][14]/P0001  & n13805 ;
  assign n31182 = \wishbone_bd_ram_mem1_reg[66][14]/P0001  & n13603 ;
  assign n31183 = ~n31181 & ~n31182 ;
  assign n31184 = n31180 & n31183 ;
  assign n31185 = n31177 & n31184 ;
  assign n31186 = n31170 & n31185 ;
  assign n31187 = n31155 & n31186 ;
  assign n31188 = \wishbone_bd_ram_mem1_reg[138][14]/P0001  & n13398 ;
  assign n31189 = \wishbone_bd_ram_mem1_reg[116][14]/P0001  & n13865 ;
  assign n31190 = ~n31188 & ~n31189 ;
  assign n31191 = \wishbone_bd_ram_mem1_reg[121][14]/P0001  & n13983 ;
  assign n31192 = \wishbone_bd_ram_mem1_reg[204][14]/P0001  & n13821 ;
  assign n31193 = ~n31191 & ~n31192 ;
  assign n31194 = n31190 & n31193 ;
  assign n31195 = \wishbone_bd_ram_mem1_reg[212][14]/P0001  & n13634 ;
  assign n31196 = \wishbone_bd_ram_mem1_reg[233][14]/P0001  & n13332 ;
  assign n31197 = ~n31195 & ~n31196 ;
  assign n31198 = \wishbone_bd_ram_mem1_reg[43][14]/P0001  & n13761 ;
  assign n31199 = \wishbone_bd_ram_mem1_reg[27][14]/P0001  & n13251 ;
  assign n31200 = ~n31198 & ~n31199 ;
  assign n31201 = n31197 & n31200 ;
  assign n31202 = n31194 & n31201 ;
  assign n31203 = \wishbone_bd_ram_mem1_reg[178][14]/P0001  & n13301 ;
  assign n31204 = \wishbone_bd_ram_mem1_reg[1][14]/P0001  & n13888 ;
  assign n31205 = ~n31203 & ~n31204 ;
  assign n31206 = \wishbone_bd_ram_mem1_reg[232][14]/P0001  & n13510 ;
  assign n31207 = \wishbone_bd_ram_mem1_reg[235][14]/P0001  & n13518 ;
  assign n31208 = ~n31206 & ~n31207 ;
  assign n31209 = n31205 & n31208 ;
  assign n31210 = \wishbone_bd_ram_mem1_reg[125][14]/P0001  & n13396 ;
  assign n31211 = \wishbone_bd_ram_mem1_reg[219][14]/P0001  & n13577 ;
  assign n31212 = ~n31210 & ~n31211 ;
  assign n31213 = \wishbone_bd_ram_mem1_reg[11][14]/P0001  & n13774 ;
  assign n31214 = \wishbone_bd_ram_mem1_reg[36][14]/P0001  & n13639 ;
  assign n31215 = ~n31213 & ~n31214 ;
  assign n31216 = n31212 & n31215 ;
  assign n31217 = n31209 & n31216 ;
  assign n31218 = n31202 & n31217 ;
  assign n31219 = \wishbone_bd_ram_mem1_reg[17][14]/P0001  & n13324 ;
  assign n31220 = \wishbone_bd_ram_mem1_reg[25][14]/P0001  & n13742 ;
  assign n31221 = ~n31219 & ~n31220 ;
  assign n31222 = \wishbone_bd_ram_mem1_reg[105][14]/P0001  & n13503 ;
  assign n31223 = \wishbone_bd_ram_mem1_reg[234][14]/P0001  & n13781 ;
  assign n31224 = ~n31222 & ~n31223 ;
  assign n31225 = n31221 & n31224 ;
  assign n31226 = \wishbone_bd_ram_mem1_reg[14][14]/P0001  & n13972 ;
  assign n31227 = \wishbone_bd_ram_mem1_reg[93][14]/P0001  & n13891 ;
  assign n31228 = ~n31226 & ~n31227 ;
  assign n31229 = \wishbone_bd_ram_mem1_reg[32][14]/P0001  & n13736 ;
  assign n31230 = \wishbone_bd_ram_mem1_reg[215][14]/P0001  & n13901 ;
  assign n31231 = ~n31229 & ~n31230 ;
  assign n31232 = n31228 & n31231 ;
  assign n31233 = n31225 & n31232 ;
  assign n31234 = \wishbone_bd_ram_mem1_reg[199][14]/P0001  & n13499 ;
  assign n31235 = \wishbone_bd_ram_mem1_reg[133][14]/P0001  & n13492 ;
  assign n31236 = ~n31234 & ~n31235 ;
  assign n31237 = \wishbone_bd_ram_mem1_reg[165][14]/P0001  & n14028 ;
  assign n31238 = \wishbone_bd_ram_mem1_reg[169][14]/P0001  & n13541 ;
  assign n31239 = ~n31237 & ~n31238 ;
  assign n31240 = n31236 & n31239 ;
  assign n31241 = \wishbone_bd_ram_mem1_reg[185][14]/P0001  & n13372 ;
  assign n31242 = \wishbone_bd_ram_mem1_reg[129][14]/P0001  & n13629 ;
  assign n31243 = ~n31241 & ~n31242 ;
  assign n31244 = \wishbone_bd_ram_mem1_reg[240][14]/P0001  & n13352 ;
  assign n31245 = \wishbone_bd_ram_mem1_reg[175][14]/P0001  & n13674 ;
  assign n31246 = ~n31244 & ~n31245 ;
  assign n31247 = n31243 & n31246 ;
  assign n31248 = n31240 & n31247 ;
  assign n31249 = n31233 & n31248 ;
  assign n31250 = n31218 & n31249 ;
  assign n31251 = n31187 & n31250 ;
  assign n31252 = n31124 & n31251 ;
  assign n31253 = \wishbone_bd_ram_mem1_reg[38][14]/P0001  & n13828 ;
  assign n31254 = \wishbone_bd_ram_mem1_reg[119][14]/P0001  & n14033 ;
  assign n31255 = ~n31253 & ~n31254 ;
  assign n31256 = \wishbone_bd_ram_mem1_reg[163][14]/P0001  & n13255 ;
  assign n31257 = \wishbone_bd_ram_mem1_reg[251][14]/P0001  & n14019 ;
  assign n31258 = ~n31256 & ~n31257 ;
  assign n31259 = n31255 & n31258 ;
  assign n31260 = \wishbone_bd_ram_mem1_reg[161][14]/P0001  & n13505 ;
  assign n31261 = \wishbone_bd_ram_mem1_reg[153][14]/P0001  & n13309 ;
  assign n31262 = ~n31260 & ~n31261 ;
  assign n31263 = \wishbone_bd_ram_mem1_reg[84][14]/P0001  & n13385 ;
  assign n31264 = \wishbone_bd_ram_mem1_reg[6][14]/P0001  & n13915 ;
  assign n31265 = ~n31263 & ~n31264 ;
  assign n31266 = n31262 & n31265 ;
  assign n31267 = n31259 & n31266 ;
  assign n31268 = \wishbone_bd_ram_mem1_reg[180][14]/P0001  & n13650 ;
  assign n31269 = \wishbone_bd_ram_mem1_reg[173][14]/P0001  & n13360 ;
  assign n31270 = ~n31268 & ~n31269 ;
  assign n31271 = \wishbone_bd_ram_mem1_reg[191][14]/P0001  & n14012 ;
  assign n31272 = \wishbone_bd_ram_mem1_reg[19][14]/P0001  & n13886 ;
  assign n31273 = ~n31271 & ~n31272 ;
  assign n31274 = n31270 & n31273 ;
  assign n31275 = \wishbone_bd_ram_mem1_reg[80][14]/P0001  & n13516 ;
  assign n31276 = \wishbone_bd_ram_mem1_reg[34][14]/P0001  & n13450 ;
  assign n31277 = ~n31275 & ~n31276 ;
  assign n31278 = \wishbone_bd_ram_mem1_reg[92][14]/P0001  & n13859 ;
  assign n31279 = \wishbone_bd_ram_mem1_reg[188][14]/P0001  & n13407 ;
  assign n31280 = ~n31278 & ~n31279 ;
  assign n31281 = n31277 & n31280 ;
  assign n31282 = n31274 & n31281 ;
  assign n31283 = n31267 & n31282 ;
  assign n31284 = \wishbone_bd_ram_mem1_reg[213][14]/P0001  & n13870 ;
  assign n31285 = \wishbone_bd_ram_mem1_reg[144][14]/P0001  & n13508 ;
  assign n31286 = ~n31284 & ~n31285 ;
  assign n31287 = \wishbone_bd_ram_mem1_reg[42][14]/P0001  & n13341 ;
  assign n31288 = \wishbone_bd_ram_mem1_reg[64][14]/P0001  & n13904 ;
  assign n31289 = ~n31287 & ~n31288 ;
  assign n31290 = n31286 & n31289 ;
  assign n31291 = \wishbone_bd_ram_mem1_reg[91][14]/P0001  & n13954 ;
  assign n31292 = \wishbone_bd_ram_mem1_reg[71][14]/P0001  & n13636 ;
  assign n31293 = ~n31291 & ~n31292 ;
  assign n31294 = \wishbone_bd_ram_mem1_reg[7][14]/P0001  & n13546 ;
  assign n31295 = \wishbone_bd_ram_mem1_reg[186][14]/P0001  & n13616 ;
  assign n31296 = ~n31294 & ~n31295 ;
  assign n31297 = n31293 & n31296 ;
  assign n31298 = n31290 & n31297 ;
  assign n31299 = \wishbone_bd_ram_mem1_reg[236][14]/P0001  & n13480 ;
  assign n31300 = \wishbone_bd_ram_mem1_reg[96][14]/P0001  & n13425 ;
  assign n31301 = ~n31299 & ~n31300 ;
  assign n31302 = \wishbone_bd_ram_mem1_reg[55][14]/P0001  & n13618 ;
  assign n31303 = \wishbone_bd_ram_mem1_reg[252][14]/P0001  & n13986 ;
  assign n31304 = ~n31302 & ~n31303 ;
  assign n31305 = n31301 & n31304 ;
  assign n31306 = \wishbone_bd_ram_mem1_reg[254][14]/P0001  & n13283 ;
  assign n31307 = \wishbone_bd_ram_mem1_reg[139][14]/P0001  & n13566 ;
  assign n31308 = ~n31306 & ~n31307 ;
  assign n31309 = \wishbone_bd_ram_mem1_reg[109][14]/P0001  & n13306 ;
  assign n31310 = \wishbone_bd_ram_mem1_reg[10][14]/P0001  & n13837 ;
  assign n31311 = ~n31309 & ~n31310 ;
  assign n31312 = n31308 & n31311 ;
  assign n31313 = n31305 & n31312 ;
  assign n31314 = n31298 & n31313 ;
  assign n31315 = n31283 & n31314 ;
  assign n31316 = \wishbone_bd_ram_mem1_reg[249][14]/P0001  & n13431 ;
  assign n31317 = \wishbone_bd_ram_mem1_reg[15][14]/P0001  & n13797 ;
  assign n31318 = ~n31316 & ~n31317 ;
  assign n31319 = \wishbone_bd_ram_mem1_reg[52][14]/P0001  & n13988 ;
  assign n31320 = \wishbone_bd_ram_mem1_reg[179][14]/P0001  & n14035 ;
  assign n31321 = ~n31319 & ~n31320 ;
  assign n31322 = n31318 & n31321 ;
  assign n31323 = \wishbone_bd_ram_mem1_reg[201][14]/P0001  & n13600 ;
  assign n31324 = \wishbone_bd_ram_mem1_reg[61][14]/P0001  & n13544 ;
  assign n31325 = ~n31323 & ~n31324 ;
  assign n31326 = \wishbone_bd_ram_mem1_reg[245][14]/P0001  & n13877 ;
  assign n31327 = \wishbone_bd_ram_mem1_reg[193][14]/P0001  & n14022 ;
  assign n31328 = ~n31326 & ~n31327 ;
  assign n31329 = n31325 & n31328 ;
  assign n31330 = n31322 & n31329 ;
  assign n31331 = \wishbone_bd_ram_mem1_reg[62][14]/P0001  & n13529 ;
  assign n31332 = \wishbone_bd_ram_mem1_reg[196][14]/P0001  & n13977 ;
  assign n31333 = ~n31331 & ~n31332 ;
  assign n31334 = \wishbone_bd_ram_mem1_reg[30][14]/P0001  & n13713 ;
  assign n31335 = \wishbone_bd_ram_mem1_reg[128][14]/P0001  & n13652 ;
  assign n31336 = ~n31334 & ~n31335 ;
  assign n31337 = n31333 & n31336 ;
  assign n31338 = \wishbone_bd_ram_mem1_reg[24][14]/P0001  & n13970 ;
  assign n31339 = \wishbone_bd_ram_mem1_reg[88][14]/P0001  & n13347 ;
  assign n31340 = ~n31338 & ~n31339 ;
  assign n31341 = \wishbone_bd_ram_mem1_reg[115][14]/P0001  & n13747 ;
  assign n31342 = \wishbone_bd_ram_mem1_reg[97][14]/P0001  & n13724 ;
  assign n31343 = ~n31341 & ~n31342 ;
  assign n31344 = n31340 & n31343 ;
  assign n31345 = n31337 & n31344 ;
  assign n31346 = n31330 & n31345 ;
  assign n31347 = \wishbone_bd_ram_mem1_reg[151][14]/P0001  & n13697 ;
  assign n31348 = \wishbone_bd_ram_mem1_reg[39][14]/P0001  & n13893 ;
  assign n31349 = ~n31347 & ~n31348 ;
  assign n31350 = \wishbone_bd_ram_mem1_reg[152][14]/P0001  & n13912 ;
  assign n31351 = \wishbone_bd_ram_mem1_reg[48][14]/P0001  & n13917 ;
  assign n31352 = ~n31350 & ~n31351 ;
  assign n31353 = n31349 & n31352 ;
  assign n31354 = \wishbone_bd_ram_mem1_reg[145][14]/P0001  & n13715 ;
  assign n31355 = \wishbone_bd_ram_mem1_reg[192][14]/P0001  & n13390 ;
  assign n31356 = ~n31354 & ~n31355 ;
  assign n31357 = \wishbone_bd_ram_mem1_reg[51][14]/P0001  & n13880 ;
  assign n31358 = \wishbone_bd_ram_mem1_reg[200][14]/P0001  & n13922 ;
  assign n31359 = ~n31357 & ~n31358 ;
  assign n31360 = n31356 & n31359 ;
  assign n31361 = n31353 & n31360 ;
  assign n31362 = \wishbone_bd_ram_mem1_reg[187][14]/P0001  & n13756 ;
  assign n31363 = \wishbone_bd_ram_mem1_reg[20][14]/P0001  & n13839 ;
  assign n31364 = ~n31362 & ~n31363 ;
  assign n31365 = \wishbone_bd_ram_mem1_reg[136][14]/P0001  & n13963 ;
  assign n31366 = \wishbone_bd_ram_mem1_reg[110][14]/P0001  & n14030 ;
  assign n31367 = ~n31365 & ~n31366 ;
  assign n31368 = n31364 & n31367 ;
  assign n31369 = \wishbone_bd_ram_mem1_reg[225][14]/P0001  & n13719 ;
  assign n31370 = \wishbone_bd_ram_mem1_reg[3][14]/P0001  & n13354 ;
  assign n31371 = ~n31369 & ~n31370 ;
  assign n31372 = \wishbone_bd_ram_mem1_reg[47][14]/P0001  & n13436 ;
  assign n31373 = \wishbone_bd_ram_mem1_reg[120][14]/P0001  & n13550 ;
  assign n31374 = ~n31372 & ~n31373 ;
  assign n31375 = n31371 & n31374 ;
  assign n31376 = n31368 & n31375 ;
  assign n31377 = n31361 & n31376 ;
  assign n31378 = n31346 & n31377 ;
  assign n31379 = n31315 & n31378 ;
  assign n31380 = \wishbone_bd_ram_mem1_reg[49][14]/P0001  & n13929 ;
  assign n31381 = \wishbone_bd_ram_mem1_reg[184][14]/P0001  & n13960 ;
  assign n31382 = ~n31380 & ~n31381 ;
  assign n31383 = \wishbone_bd_ram_mem1_reg[82][14]/P0001  & n13374 ;
  assign n31384 = \wishbone_bd_ram_mem1_reg[142][14]/P0001  & n13448 ;
  assign n31385 = ~n31383 & ~n31384 ;
  assign n31386 = n31382 & n31385 ;
  assign n31387 = \wishbone_bd_ram_mem1_reg[77][14]/P0001  & n13935 ;
  assign n31388 = \wishbone_bd_ram_mem1_reg[22][14]/P0001  & n13744 ;
  assign n31389 = ~n31387 & ~n31388 ;
  assign n31390 = \wishbone_bd_ram_mem1_reg[21][14]/P0001  & n13438 ;
  assign n31391 = \wishbone_bd_ram_mem1_reg[227][14]/P0001  & n13388 ;
  assign n31392 = ~n31390 & ~n31391 ;
  assign n31393 = n31389 & n31392 ;
  assign n31394 = n31386 & n31393 ;
  assign n31395 = \wishbone_bd_ram_mem1_reg[167][14]/P0001  & n13940 ;
  assign n31396 = \wishbone_bd_ram_mem1_reg[226][14]/P0001  & n13668 ;
  assign n31397 = ~n31395 & ~n31396 ;
  assign n31398 = \wishbone_bd_ram_mem1_reg[83][14]/P0001  & n13454 ;
  assign n31399 = \wishbone_bd_ram_mem1_reg[127][14]/P0001  & n13803 ;
  assign n31400 = ~n31398 & ~n31399 ;
  assign n31401 = n31397 & n31400 ;
  assign n31402 = \wishbone_bd_ram_mem1_reg[162][14]/P0001  & n13726 ;
  assign n31403 = \wishbone_bd_ram_mem1_reg[37][14]/P0001  & n13710 ;
  assign n31404 = ~n31402 & ~n31403 ;
  assign n31405 = \wishbone_bd_ram_mem1_reg[23][14]/P0001  & n13857 ;
  assign n31406 = \wishbone_bd_ram_mem1_reg[57][14]/P0001  & n13731 ;
  assign n31407 = ~n31405 & ~n31406 ;
  assign n31408 = n31404 & n31407 ;
  assign n31409 = n31401 & n31408 ;
  assign n31410 = n31394 & n31409 ;
  assign n31411 = \wishbone_bd_ram_mem1_reg[143][14]/P0001  & n13461 ;
  assign n31412 = \wishbone_bd_ram_mem1_reg[154][14]/P0001  & n13403 ;
  assign n31413 = ~n31411 & ~n31412 ;
  assign n31414 = \wishbone_bd_ram_mem1_reg[130][14]/P0001  & n13427 ;
  assign n31415 = \wishbone_bd_ram_mem1_reg[103][14]/P0001  & n13320 ;
  assign n31416 = ~n31414 & ~n31415 ;
  assign n31417 = n31413 & n31416 ;
  assign n31418 = \wishbone_bd_ram_mem1_reg[149][14]/P0001  & n13469 ;
  assign n31419 = \wishbone_bd_ram_mem1_reg[35][14]/P0001  & n13523 ;
  assign n31420 = ~n31418 & ~n31419 ;
  assign n31421 = \wishbone_bd_ram_mem1_reg[147][14]/P0001  & n13702 ;
  assign n31422 = \wishbone_bd_ram_mem1_reg[159][14]/P0001  & n13627 ;
  assign n31423 = ~n31421 & ~n31422 ;
  assign n31424 = n31420 & n31423 ;
  assign n31425 = n31417 & n31424 ;
  assign n31426 = \wishbone_bd_ram_mem1_reg[250][14]/P0001  & n13677 ;
  assign n31427 = \wishbone_bd_ram_mem1_reg[79][14]/P0001  & n13779 ;
  assign n31428 = ~n31426 & ~n31427 ;
  assign n31429 = \wishbone_bd_ram_mem1_reg[74][14]/P0001  & n13564 ;
  assign n31430 = \wishbone_bd_ram_mem1_reg[160][14]/P0001  & n13271 ;
  assign n31431 = ~n31429 & ~n31430 ;
  assign n31432 = n31428 & n31431 ;
  assign n31433 = \wishbone_bd_ram_mem1_reg[102][14]/P0001  & n13534 ;
  assign n31434 = \wishbone_bd_ram_mem1_reg[141][14]/P0001  & n13852 ;
  assign n31435 = ~n31433 & ~n31434 ;
  assign n31436 = \wishbone_bd_ram_mem1_reg[239][14]/P0001  & n13349 ;
  assign n31437 = \wishbone_bd_ram_mem1_reg[63][14]/P0001  & n13327 ;
  assign n31438 = ~n31436 & ~n31437 ;
  assign n31439 = n31435 & n31438 ;
  assign n31440 = n31432 & n31439 ;
  assign n31441 = n31425 & n31440 ;
  assign n31442 = n31410 & n31441 ;
  assign n31443 = \wishbone_bd_ram_mem1_reg[26][14]/P0001  & n13521 ;
  assign n31444 = \wishbone_bd_ram_mem1_reg[9][14]/P0001  & n13580 ;
  assign n31445 = ~n31443 & ~n31444 ;
  assign n31446 = \wishbone_bd_ram_mem1_reg[89][14]/P0001  & n13910 ;
  assign n31447 = \wishbone_bd_ram_mem1_reg[150][14]/P0001  & n13666 ;
  assign n31448 = ~n31446 & ~n31447 ;
  assign n31449 = n31445 & n31448 ;
  assign n31450 = \wishbone_bd_ram_mem1_reg[104][14]/P0001  & n13684 ;
  assign n31451 = \wishbone_bd_ram_mem1_reg[99][14]/P0001  & n13996 ;
  assign n31452 = ~n31450 & ~n31451 ;
  assign n31453 = \wishbone_bd_ram_mem1_reg[208][14]/P0001  & n14010 ;
  assign n31454 = \wishbone_bd_ram_mem1_reg[166][14]/P0001  & n13999 ;
  assign n31455 = ~n31453 & ~n31454 ;
  assign n31456 = n31452 & n31455 ;
  assign n31457 = n31449 & n31456 ;
  assign n31458 = \wishbone_bd_ram_mem1_reg[5][14]/P0001  & n13243 ;
  assign n31459 = \wishbone_bd_ram_mem1_reg[229][14]/P0001  & n13552 ;
  assign n31460 = ~n31458 & ~n31459 ;
  assign n31461 = \wishbone_bd_ram_mem1_reg[182][14]/P0001  & n13598 ;
  assign n31462 = \wishbone_bd_ram_mem1_reg[94][14]/P0001  & n13833 ;
  assign n31463 = ~n31461 & ~n31462 ;
  assign n31464 = n31460 & n31463 ;
  assign n31465 = \wishbone_bd_ram_mem1_reg[117][14]/P0001  & n13557 ;
  assign n31466 = \wishbone_bd_ram_mem1_reg[67][14]/P0001  & n13663 ;
  assign n31467 = ~n31465 & ~n31466 ;
  assign n31468 = \wishbone_bd_ram_mem1_reg[246][14]/P0001  & n13981 ;
  assign n31469 = \wishbone_bd_ram_mem1_reg[111][14]/P0001  & n13471 ;
  assign n31470 = ~n31468 & ~n31469 ;
  assign n31471 = n31467 & n31470 ;
  assign n31472 = n31464 & n31471 ;
  assign n31473 = n31457 & n31472 ;
  assign n31474 = \wishbone_bd_ram_mem1_reg[174][14]/P0001  & n13899 ;
  assign n31475 = \wishbone_bd_ram_mem1_reg[244][14]/P0001  & n13474 ;
  assign n31476 = ~n31474 & ~n31475 ;
  assign n31477 = \wishbone_bd_ram_mem1_reg[40][14]/P0001  & n13661 ;
  assign n31478 = \wishbone_bd_ram_mem1_reg[90][14]/P0001  & n13906 ;
  assign n31479 = ~n31477 & ~n31478 ;
  assign n31480 = n31476 & n31479 ;
  assign n31481 = \wishbone_bd_ram_mem1_reg[100][14]/P0001  & n13401 ;
  assign n31482 = \wishbone_bd_ram_mem1_reg[60][14]/P0001  & n13790 ;
  assign n31483 = ~n31481 & ~n31482 ;
  assign n31484 = \wishbone_bd_ram_mem1_reg[168][14]/P0001  & n13795 ;
  assign n31485 = \wishbone_bd_ram_mem1_reg[106][14]/P0001  & n13555 ;
  assign n31486 = ~n31484 & ~n31485 ;
  assign n31487 = n31483 & n31486 ;
  assign n31488 = n31480 & n31487 ;
  assign n31489 = \wishbone_bd_ram_mem1_reg[124][14]/P0001  & n14024 ;
  assign n31490 = \wishbone_bd_ram_mem1_reg[181][14]/P0001  & n13587 ;
  assign n31491 = ~n31489 & ~n31490 ;
  assign n31492 = \wishbone_bd_ram_mem1_reg[228][14]/P0001  & n13497 ;
  assign n31493 = \wishbone_bd_ram_mem1_reg[122][14]/P0001  & n13679 ;
  assign n31494 = ~n31492 & ~n31493 ;
  assign n31495 = n31491 & n31494 ;
  assign n31496 = \wishbone_bd_ram_mem1_reg[158][14]/P0001  & n13294 ;
  assign n31497 = \wishbone_bd_ram_mem1_reg[59][14]/P0001  & n13613 ;
  assign n31498 = ~n31496 & ~n31497 ;
  assign n31499 = \wishbone_bd_ram_mem1_reg[65][14]/P0001  & n13842 ;
  assign n31500 = \wishbone_bd_ram_mem1_reg[86][14]/P0001  & n13485 ;
  assign n31501 = ~n31499 & ~n31500 ;
  assign n31502 = n31498 & n31501 ;
  assign n31503 = n31495 & n31502 ;
  assign n31504 = n31488 & n31503 ;
  assign n31505 = n31473 & n31504 ;
  assign n31506 = n31442 & n31505 ;
  assign n31507 = n31379 & n31506 ;
  assign n31508 = n31252 & n31507 ;
  assign n31509 = ~wb_rst_i_pad & ~n30996 ;
  assign n31510 = ~n31508 & n31509 ;
  assign n31511 = ~n30997 & ~n31510 ;
  assign n31512 = \ethreg1_MODER_1_DataOut_reg[7]/NET0131  & n23808 ;
  assign n31513 = \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131  & n23794 ;
  assign n31514 = n23741 & n31513 ;
  assign n31515 = ~n31512 & ~n31514 ;
  assign n31516 = \ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131  & n23743 ;
  assign n31517 = n23741 & n31516 ;
  assign n31518 = \ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131  & n23743 ;
  assign n31519 = n23747 & n31518 ;
  assign n31520 = ~n31517 & ~n31519 ;
  assign n31521 = n31515 & n31520 ;
  assign n31522 = n23730 & n31521 ;
  assign n31523 = \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  & n23737 ;
  assign n31524 = \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131  & n23813 ;
  assign n31525 = \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  & n23751 ;
  assign n31526 = n23741 & n31525 ;
  assign n31527 = ~n31524 & ~n31526 ;
  assign n31528 = \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  & n23751 ;
  assign n31529 = n23747 & n31528 ;
  assign n31530 = \ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131  & n23782 ;
  assign n31531 = ~n31529 & ~n31530 ;
  assign n31532 = n31527 & n31531 ;
  assign n31533 = ~n31523 & n31532 ;
  assign n31534 = n31522 & n31533 ;
  assign n31535 = n23730 & ~n31534 ;
  assign n31536 = ~wb_rst_i_pad & ~n31534 ;
  assign n31537 = ~n16296 & n31536 ;
  assign n31538 = ~n31535 & ~n31537 ;
  assign n31539 = \wishbone_RxPointerMSB_reg[11]/NET0131  & n18517 ;
  assign n31540 = ~\wishbone_RxPointerMSB_reg[12]/NET0131  & ~n31539 ;
  assign n31541 = \wishbone_RxPointerMSB_reg[11]/NET0131  & \wishbone_RxPointerMSB_reg[12]/NET0131  ;
  assign n31542 = n18517 & n31541 ;
  assign n31543 = ~n16305 & ~n31542 ;
  assign n31544 = ~n31540 & n31543 ;
  assign n31545 = n18507 & ~n24329 ;
  assign n31546 = ~n31544 & ~n31545 ;
  assign n31547 = \wishbone_RxPointerMSB_reg[11]/NET0131  & n18518 ;
  assign n31548 = n18517 & n31547 ;
  assign n31549 = ~\wishbone_RxPointerMSB_reg[14]/NET0131  & ~n31548 ;
  assign n31550 = ~n16305 & ~n18521 ;
  assign n31551 = ~n31549 & n31550 ;
  assign n31552 = n18507 & ~n31508 ;
  assign n31553 = ~n31551 & ~n31552 ;
  assign n31554 = ~\wishbone_RxPointerMSB_reg[4]/NET0131  & ~n18510 ;
  assign n31555 = \wishbone_RxPointerMSB_reg[4]/NET0131  & n18510 ;
  assign n31556 = ~n16305 & ~n31555 ;
  assign n31557 = ~n31554 & n31556 ;
  assign n31558 = n18507 & ~n26168 ;
  assign n31559 = ~n31557 & ~n31558 ;
  assign n31560 = ~\wishbone_RxPointerMSB_reg[5]/NET0131  & ~n31555 ;
  assign n31561 = \wishbone_RxPointerMSB_reg[4]/NET0131  & \wishbone_RxPointerMSB_reg[5]/NET0131  ;
  assign n31562 = n18510 & n31561 ;
  assign n31563 = ~n16305 & ~n31562 ;
  assign n31564 = ~n31560 & n31563 ;
  assign n31565 = n18507 & ~n26722 ;
  assign n31566 = ~n31564 & ~n31565 ;
  assign n31567 = \wishbone_RxPointerMSB_reg[7]/NET0131  & ~n16305 ;
  assign n31568 = ~n18513 & n31567 ;
  assign n31569 = ~\wishbone_RxPointerMSB_reg[7]/NET0131  & ~n16305 ;
  assign n31570 = n18513 & n31569 ;
  assign n31571 = ~n31568 & ~n31570 ;
  assign n31572 = n18507 & ~n27264 ;
  assign n31573 = n31571 & ~n31572 ;
  assign n31574 = ~\wishbone_RxPointerMSB_reg[6]/NET0131  & ~n31562 ;
  assign n31575 = ~n16305 & ~n18513 ;
  assign n31576 = ~n31574 & n31575 ;
  assign n31577 = n18507 & ~n30191 ;
  assign n31578 = ~n31576 & ~n31577 ;
  assign n31579 = \wishbone_TxPointerMSB_reg[10]/NET0131  & \wishbone_TxPointerMSB_reg[11]/NET0131  ;
  assign n31580 = n18554 & n31579 ;
  assign n31581 = ~\wishbone_TxPointerMSB_reg[12]/NET0131  & ~n31580 ;
  assign n31582 = ~n18545 & ~n18557 ;
  assign n31583 = ~n31581 & n31582 ;
  assign n31584 = ~n24329 & n24387 ;
  assign n31585 = ~n31583 & ~n31584 ;
  assign n31586 = n24387 & ~n31508 ;
  assign n31587 = \wishbone_TxPointerMSB_reg[13]/NET0131  & n18557 ;
  assign n31588 = ~\wishbone_TxPointerMSB_reg[14]/NET0131  & ~n31587 ;
  assign n31589 = n18557 & n18559 ;
  assign n31590 = ~n18545 & ~n31589 ;
  assign n31591 = ~n31588 & n31590 ;
  assign n31592 = ~n31586 & ~n31591 ;
  assign n31593 = ~\wishbone_TxPointerMSB_reg[4]/NET0131  & ~n18548 ;
  assign n31594 = \wishbone_TxPointerMSB_reg[4]/NET0131  & n18548 ;
  assign n31595 = ~n18545 & ~n31594 ;
  assign n31596 = ~n31593 & n31595 ;
  assign n31597 = n24387 & ~n26168 ;
  assign n31598 = ~n31596 & ~n31597 ;
  assign n31599 = ~\wishbone_TxPointerMSB_reg[5]/NET0131  & ~n31594 ;
  assign n31600 = \wishbone_TxPointerMSB_reg[4]/NET0131  & \wishbone_TxPointerMSB_reg[5]/NET0131  ;
  assign n31601 = n18548 & n31600 ;
  assign n31602 = ~n18545 & ~n31601 ;
  assign n31603 = ~n31599 & n31602 ;
  assign n31604 = n24387 & ~n26722 ;
  assign n31605 = ~n31603 & ~n31604 ;
  assign n31606 = ~\wishbone_TxPointerMSB_reg[6]/NET0131  & ~n31601 ;
  assign n31607 = ~n18545 & ~n18551 ;
  assign n31608 = ~n31606 & n31607 ;
  assign n31609 = n24387 & ~n30191 ;
  assign n31610 = ~n31608 & ~n31609 ;
  assign n31611 = \wishbone_TxPointerMSB_reg[7]/NET0131  & ~n18545 ;
  assign n31612 = ~n18551 & n31611 ;
  assign n31613 = ~\wishbone_TxPointerMSB_reg[7]/NET0131  & ~n18545 ;
  assign n31614 = n18551 & n31613 ;
  assign n31615 = ~n31612 & ~n31614 ;
  assign n31616 = n24387 & ~n27264 ;
  assign n31617 = n31615 & ~n31616 ;
  assign n31618 = \wishbone_RxPointerMSB_reg[11]/NET0131  & ~n16305 ;
  assign n31619 = ~n18517 & n31618 ;
  assign n31620 = ~\wishbone_RxPointerMSB_reg[11]/NET0131  & ~n16305 ;
  assign n31621 = n18517 & n31620 ;
  assign n31622 = ~n31619 & ~n31621 ;
  assign n31623 = n18507 & ~n28901 ;
  assign n31624 = n31622 & ~n31623 ;
  assign n31625 = n18507 & ~n30970 ;
  assign n31626 = ~\wishbone_RxPointerMSB_reg[13]/NET0131  & ~n31542 ;
  assign n31627 = ~n16305 & ~n31548 ;
  assign n31628 = ~n31626 & n31627 ;
  assign n31629 = ~n31625 & ~n31628 ;
  assign n31630 = \wishbone_RxPointerMSB_reg[15]/NET0131  & ~n16305 ;
  assign n31631 = ~n18521 & n31630 ;
  assign n31632 = ~\wishbone_RxPointerMSB_reg[15]/NET0131  & ~n16305 ;
  assign n31633 = n18521 & n31632 ;
  assign n31634 = ~n31631 & ~n31633 ;
  assign n31635 = ~n16296 & n18507 ;
  assign n31636 = n31634 & ~n31635 ;
  assign n31637 = \wishbone_RxPointerMSB_reg[15]/NET0131  & n18521 ;
  assign n31638 = ~\wishbone_RxPointerMSB_reg[16]/NET0131  & ~n31637 ;
  assign n31639 = \wishbone_RxPointerMSB_reg[15]/NET0131  & \wishbone_RxPointerMSB_reg[16]/NET0131  ;
  assign n31640 = n18521 & n31639 ;
  assign n31641 = ~n16305 & ~n31640 ;
  assign n31642 = ~n31638 & n31641 ;
  assign n31643 = n18507 & ~n19794 ;
  assign n31644 = ~n31642 & ~n31643 ;
  assign n31645 = ~\wishbone_RxPointerMSB_reg[17]/NET0131  & ~n31640 ;
  assign n31646 = ~n16305 & ~n30249 ;
  assign n31647 = ~n31645 & n31646 ;
  assign n31648 = n18507 & ~n20833 ;
  assign n31649 = ~n31647 & ~n31648 ;
  assign n31650 = \wishbone_RxPointerMSB_reg[18]/NET0131  & ~n16305 ;
  assign n31651 = ~n30249 & n31650 ;
  assign n31652 = ~\wishbone_RxPointerMSB_reg[18]/NET0131  & ~n16305 ;
  assign n31653 = n30249 & n31652 ;
  assign n31654 = ~n31651 & ~n31653 ;
  assign n31655 = n18507 & ~n19273 ;
  assign n31656 = n31654 & ~n31655 ;
  assign n31657 = ~\wishbone_RxPointerMSB_reg[2]/NET0131  & ~n16307 ;
  assign n31658 = \wishbone_RxPointerMSB_reg[2]/NET0131  & n16307 ;
  assign n31659 = ~n16305 & ~n31658 ;
  assign n31660 = ~n31657 & n31659 ;
  assign n31661 = n18507 & ~n29475 ;
  assign n31662 = ~n31660 & ~n31661 ;
  assign n31663 = ~\wishbone_RxPointerMSB_reg[3]/NET0131  & ~n31658 ;
  assign n31664 = ~n16305 & ~n18510 ;
  assign n31665 = ~n31663 & n31664 ;
  assign n31666 = n18507 & ~n25612 ;
  assign n31667 = ~n31665 & ~n31666 ;
  assign n31668 = \wishbone_RxPointerMSB_reg[7]/NET0131  & n18513 ;
  assign n31669 = ~\wishbone_RxPointerMSB_reg[8]/NET0131  & ~n31668 ;
  assign n31670 = ~n16305 & ~n30334 ;
  assign n31671 = ~n31669 & n31670 ;
  assign n31672 = n18507 & ~n27806 ;
  assign n31673 = ~n31671 & ~n31672 ;
  assign n31674 = \wishbone_TxPointerMSB_reg[10]/NET0131  & ~n18545 ;
  assign n31675 = ~n18554 & n31674 ;
  assign n31676 = ~\wishbone_TxPointerMSB_reg[10]/NET0131  & ~n18545 ;
  assign n31677 = n18554 & n31676 ;
  assign n31678 = ~n31675 & ~n31677 ;
  assign n31679 = \wishbone_bd_ram_mem1_reg[20][10]/P0001  & n13839 ;
  assign n31680 = \wishbone_bd_ram_mem1_reg[88][10]/P0001  & n13347 ;
  assign n31681 = ~n31679 & ~n31680 ;
  assign n31682 = \wishbone_bd_ram_mem1_reg[33][10]/P0001  & n13933 ;
  assign n31683 = \wishbone_bd_ram_mem1_reg[222][10]/P0001  & n13721 ;
  assign n31684 = ~n31682 & ~n31683 ;
  assign n31685 = n31681 & n31684 ;
  assign n31686 = \wishbone_bd_ram_mem1_reg[134][10]/P0001  & n13494 ;
  assign n31687 = \wishbone_bd_ram_mem1_reg[199][10]/P0001  & n13499 ;
  assign n31688 = ~n31686 & ~n31687 ;
  assign n31689 = \wishbone_bd_ram_mem1_reg[112][10]/P0001  & n13482 ;
  assign n31690 = \wishbone_bd_ram_mem1_reg[78][10]/P0001  & n13277 ;
  assign n31691 = ~n31689 & ~n31690 ;
  assign n31692 = n31688 & n31691 ;
  assign n31693 = n31685 & n31692 ;
  assign n31694 = \wishbone_bd_ram_mem1_reg[208][10]/P0001  & n14010 ;
  assign n31695 = \wishbone_bd_ram_mem1_reg[107][10]/P0001  & n13476 ;
  assign n31696 = ~n31694 & ~n31695 ;
  assign n31697 = \wishbone_bd_ram_mem1_reg[118][10]/P0001  & n13589 ;
  assign n31698 = \wishbone_bd_ram_mem1_reg[155][10]/P0001  & n13738 ;
  assign n31699 = ~n31697 & ~n31698 ;
  assign n31700 = n31696 & n31699 ;
  assign n31701 = \wishbone_bd_ram_mem1_reg[193][10]/P0001  & n14022 ;
  assign n31702 = \wishbone_bd_ram_mem1_reg[116][10]/P0001  & n13865 ;
  assign n31703 = ~n31701 & ~n31702 ;
  assign n31704 = \wishbone_bd_ram_mem1_reg[251][10]/P0001  & n14019 ;
  assign n31705 = \wishbone_bd_ram_mem1_reg[113][10]/P0001  & n13882 ;
  assign n31706 = ~n31704 & ~n31705 ;
  assign n31707 = n31703 & n31706 ;
  assign n31708 = n31700 & n31707 ;
  assign n31709 = n31693 & n31708 ;
  assign n31710 = \wishbone_bd_ram_mem1_reg[200][10]/P0001  & n13922 ;
  assign n31711 = \wishbone_bd_ram_mem1_reg[148][10]/P0001  & n13868 ;
  assign n31712 = ~n31710 & ~n31711 ;
  assign n31713 = \wishbone_bd_ram_mem1_reg[230][10]/P0001  & n13994 ;
  assign n31714 = \wishbone_bd_ram_mem1_reg[14][10]/P0001  & n13972 ;
  assign n31715 = ~n31713 & ~n31714 ;
  assign n31716 = n31712 & n31715 ;
  assign n31717 = \wishbone_bd_ram_mem1_reg[38][10]/P0001  & n13828 ;
  assign n31718 = \wishbone_bd_ram_mem1_reg[64][10]/P0001  & n13904 ;
  assign n31719 = ~n31717 & ~n31718 ;
  assign n31720 = \wishbone_bd_ram_mem1_reg[132][10]/P0001  & n13927 ;
  assign n31721 = \wishbone_bd_ram_mem1_reg[235][10]/P0001  & n13518 ;
  assign n31722 = ~n31720 & ~n31721 ;
  assign n31723 = n31719 & n31722 ;
  assign n31724 = n31716 & n31723 ;
  assign n31725 = \wishbone_bd_ram_mem1_reg[255][10]/P0001  & n13952 ;
  assign n31726 = \wishbone_bd_ram_mem1_reg[71][10]/P0001  & n13636 ;
  assign n31727 = ~n31725 & ~n31726 ;
  assign n31728 = \wishbone_bd_ram_mem1_reg[127][10]/P0001  & n13803 ;
  assign n31729 = \wishbone_bd_ram_mem1_reg[21][10]/P0001  & n13438 ;
  assign n31730 = ~n31728 & ~n31729 ;
  assign n31731 = n31727 & n31730 ;
  assign n31732 = \wishbone_bd_ram_mem1_reg[17][10]/P0001  & n13324 ;
  assign n31733 = \wishbone_bd_ram_mem1_reg[0][10]/P0001  & n13539 ;
  assign n31734 = ~n31732 & ~n31733 ;
  assign n31735 = \wishbone_bd_ram_mem1_reg[27][10]/P0001  & n13251 ;
  assign n31736 = \wishbone_bd_ram_mem1_reg[158][10]/P0001  & n13294 ;
  assign n31737 = ~n31735 & ~n31736 ;
  assign n31738 = n31734 & n31737 ;
  assign n31739 = n31731 & n31738 ;
  assign n31740 = n31724 & n31739 ;
  assign n31741 = n31709 & n31740 ;
  assign n31742 = \wishbone_bd_ram_mem1_reg[247][10]/P0001  & n13571 ;
  assign n31743 = \wishbone_bd_ram_mem1_reg[180][10]/P0001  & n13650 ;
  assign n31744 = ~n31742 & ~n31743 ;
  assign n31745 = \wishbone_bd_ram_mem1_reg[225][10]/P0001  & n13719 ;
  assign n31746 = \wishbone_bd_ram_mem1_reg[145][10]/P0001  & n13715 ;
  assign n31747 = ~n31745 & ~n31746 ;
  assign n31748 = n31744 & n31747 ;
  assign n31749 = \wishbone_bd_ram_mem1_reg[49][10]/P0001  & n13929 ;
  assign n31750 = \wishbone_bd_ram_mem1_reg[128][10]/P0001  & n13652 ;
  assign n31751 = ~n31749 & ~n31750 ;
  assign n31752 = \wishbone_bd_ram_mem1_reg[245][10]/P0001  & n13877 ;
  assign n31753 = \wishbone_bd_ram_mem1_reg[120][10]/P0001  & n13550 ;
  assign n31754 = ~n31752 & ~n31753 ;
  assign n31755 = n31751 & n31754 ;
  assign n31756 = n31748 & n31755 ;
  assign n31757 = \wishbone_bd_ram_mem1_reg[106][10]/P0001  & n13555 ;
  assign n31758 = \wishbone_bd_ram_mem1_reg[212][10]/P0001  & n13634 ;
  assign n31759 = ~n31757 & ~n31758 ;
  assign n31760 = \wishbone_bd_ram_mem1_reg[246][10]/P0001  & n13981 ;
  assign n31761 = \wishbone_bd_ram_mem1_reg[181][10]/P0001  & n13587 ;
  assign n31762 = ~n31760 & ~n31761 ;
  assign n31763 = n31759 & n31762 ;
  assign n31764 = \wishbone_bd_ram_mem1_reg[196][10]/P0001  & n13977 ;
  assign n31765 = \wishbone_bd_ram_mem1_reg[81][10]/P0001  & n13409 ;
  assign n31766 = ~n31764 & ~n31765 ;
  assign n31767 = \wishbone_bd_ram_mem1_reg[183][10]/P0001  & n13645 ;
  assign n31768 = \wishbone_bd_ram_mem1_reg[250][10]/P0001  & n13677 ;
  assign n31769 = ~n31767 & ~n31768 ;
  assign n31770 = n31766 & n31769 ;
  assign n31771 = n31763 & n31770 ;
  assign n31772 = n31756 & n31771 ;
  assign n31773 = \wishbone_bd_ram_mem1_reg[241][10]/P0001  & n13854 ;
  assign n31774 = \wishbone_bd_ram_mem1_reg[146][10]/P0001  & n13958 ;
  assign n31775 = ~n31773 & ~n31774 ;
  assign n31776 = \wishbone_bd_ram_mem1_reg[18][10]/P0001  & n13532 ;
  assign n31777 = \wishbone_bd_ram_mem1_reg[58][10]/P0001  & n13949 ;
  assign n31778 = ~n31776 & ~n31777 ;
  assign n31779 = n31775 & n31778 ;
  assign n31780 = \wishbone_bd_ram_mem1_reg[83][10]/P0001  & n13454 ;
  assign n31781 = \wishbone_bd_ram_mem1_reg[79][10]/P0001  & n13779 ;
  assign n31782 = ~n31780 & ~n31781 ;
  assign n31783 = \wishbone_bd_ram_mem1_reg[204][10]/P0001  & n13821 ;
  assign n31784 = \wishbone_bd_ram_mem1_reg[243][10]/P0001  & n13575 ;
  assign n31785 = ~n31783 & ~n31784 ;
  assign n31786 = n31782 & n31785 ;
  assign n31787 = n31779 & n31786 ;
  assign n31788 = \wishbone_bd_ram_mem1_reg[24][10]/P0001  & n13970 ;
  assign n31789 = \wishbone_bd_ram_mem1_reg[149][10]/P0001  & n13469 ;
  assign n31790 = ~n31788 & ~n31789 ;
  assign n31791 = \wishbone_bd_ram_mem1_reg[32][10]/P0001  & n13736 ;
  assign n31792 = \wishbone_bd_ram_mem1_reg[42][10]/P0001  & n13341 ;
  assign n31793 = ~n31791 & ~n31792 ;
  assign n31794 = n31790 & n31793 ;
  assign n31795 = \wishbone_bd_ram_mem1_reg[133][10]/P0001  & n13492 ;
  assign n31796 = \wishbone_bd_ram_mem1_reg[52][10]/P0001  & n13988 ;
  assign n31797 = ~n31795 & ~n31796 ;
  assign n31798 = \wishbone_bd_ram_mem1_reg[136][10]/P0001  & n13963 ;
  assign n31799 = \wishbone_bd_ram_mem1_reg[86][10]/P0001  & n13485 ;
  assign n31800 = ~n31798 & ~n31799 ;
  assign n31801 = n31797 & n31800 ;
  assign n31802 = n31794 & n31801 ;
  assign n31803 = n31787 & n31802 ;
  assign n31804 = n31772 & n31803 ;
  assign n31805 = n31741 & n31804 ;
  assign n31806 = \wishbone_bd_ram_mem1_reg[103][10]/P0001  & n13320 ;
  assign n31807 = \wishbone_bd_ram_mem1_reg[56][10]/P0001  & n13611 ;
  assign n31808 = ~n31806 & ~n31807 ;
  assign n31809 = \wishbone_bd_ram_mem1_reg[220][10]/P0001  & n13965 ;
  assign n31810 = \wishbone_bd_ram_mem1_reg[131][10]/P0001  & n13358 ;
  assign n31811 = ~n31809 & ~n31810 ;
  assign n31812 = n31808 & n31811 ;
  assign n31813 = \wishbone_bd_ram_mem1_reg[141][10]/P0001  & n13852 ;
  assign n31814 = \wishbone_bd_ram_mem1_reg[137][10]/P0001  & n13808 ;
  assign n31815 = ~n31813 & ~n31814 ;
  assign n31816 = \wishbone_bd_ram_mem1_reg[191][10]/P0001  & n14012 ;
  assign n31817 = \wishbone_bd_ram_mem1_reg[177][10]/P0001  & n13863 ;
  assign n31818 = ~n31816 & ~n31817 ;
  assign n31819 = n31815 & n31818 ;
  assign n31820 = n31812 & n31819 ;
  assign n31821 = \wishbone_bd_ram_mem1_reg[70][10]/P0001  & n13339 ;
  assign n31822 = \wishbone_bd_ram_mem1_reg[10][10]/P0001  & n13837 ;
  assign n31823 = ~n31821 & ~n31822 ;
  assign n31824 = \wishbone_bd_ram_mem1_reg[219][10]/P0001  & n13577 ;
  assign n31825 = \wishbone_bd_ram_mem1_reg[236][10]/P0001  & n13480 ;
  assign n31826 = ~n31824 & ~n31825 ;
  assign n31827 = n31823 & n31826 ;
  assign n31828 = \wishbone_bd_ram_mem1_reg[228][10]/P0001  & n13497 ;
  assign n31829 = \wishbone_bd_ram_mem1_reg[65][10]/P0001  & n13842 ;
  assign n31830 = ~n31828 & ~n31829 ;
  assign n31831 = \wishbone_bd_ram_mem1_reg[189][10]/P0001  & n14001 ;
  assign n31832 = \wishbone_bd_ram_mem1_reg[82][10]/P0001  & n13374 ;
  assign n31833 = ~n31831 & ~n31832 ;
  assign n31834 = n31830 & n31833 ;
  assign n31835 = n31827 & n31834 ;
  assign n31836 = n31820 & n31835 ;
  assign n31837 = \wishbone_bd_ram_mem1_reg[210][10]/P0001  & n13443 ;
  assign n31838 = \wishbone_bd_ram_mem1_reg[159][10]/P0001  & n13627 ;
  assign n31839 = ~n31837 & ~n31838 ;
  assign n31840 = \wishbone_bd_ram_mem1_reg[43][10]/P0001  & n13761 ;
  assign n31841 = \wishbone_bd_ram_mem1_reg[253][10]/P0001  & n13708 ;
  assign n31842 = ~n31840 & ~n31841 ;
  assign n31843 = n31839 & n31842 ;
  assign n31844 = \wishbone_bd_ram_mem1_reg[124][10]/P0001  & n14024 ;
  assign n31845 = \wishbone_bd_ram_mem1_reg[3][10]/P0001  & n13354 ;
  assign n31846 = ~n31844 & ~n31845 ;
  assign n31847 = \wishbone_bd_ram_mem1_reg[164][10]/P0001  & n13236 ;
  assign n31848 = \wishbone_bd_ram_mem1_reg[29][10]/P0001  & n13412 ;
  assign n31849 = ~n31847 & ~n31848 ;
  assign n31850 = n31846 & n31849 ;
  assign n31851 = n31843 & n31850 ;
  assign n31852 = \wishbone_bd_ram_mem1_reg[77][10]/P0001  & n13935 ;
  assign n31853 = \wishbone_bd_ram_mem1_reg[249][10]/P0001  & n13431 ;
  assign n31854 = ~n31852 & ~n31853 ;
  assign n31855 = \wishbone_bd_ram_mem1_reg[119][10]/P0001  & n14033 ;
  assign n31856 = \wishbone_bd_ram_mem1_reg[92][10]/P0001  & n13859 ;
  assign n31857 = ~n31855 & ~n31856 ;
  assign n31858 = n31854 & n31857 ;
  assign n31859 = \wishbone_bd_ram_mem1_reg[60][10]/P0001  & n13790 ;
  assign n31860 = \wishbone_bd_ram_mem1_reg[30][10]/P0001  & n13713 ;
  assign n31861 = ~n31859 & ~n31860 ;
  assign n31862 = \wishbone_bd_ram_mem1_reg[242][10]/P0001  & n13383 ;
  assign n31863 = \wishbone_bd_ram_mem1_reg[48][10]/P0001  & n13917 ;
  assign n31864 = ~n31862 & ~n31863 ;
  assign n31865 = n31861 & n31864 ;
  assign n31866 = n31858 & n31865 ;
  assign n31867 = n31851 & n31866 ;
  assign n31868 = n31836 & n31867 ;
  assign n31869 = \wishbone_bd_ram_mem1_reg[28][10]/P0001  & n13810 ;
  assign n31870 = \wishbone_bd_ram_mem1_reg[100][10]/P0001  & n13401 ;
  assign n31871 = ~n31869 & ~n31870 ;
  assign n31872 = \wishbone_bd_ram_mem1_reg[102][10]/P0001  & n13534 ;
  assign n31873 = \wishbone_bd_ram_mem1_reg[161][10]/P0001  & n13505 ;
  assign n31874 = ~n31872 & ~n31873 ;
  assign n31875 = n31871 & n31874 ;
  assign n31876 = \wishbone_bd_ram_mem1_reg[90][10]/P0001  & n13906 ;
  assign n31877 = \wishbone_bd_ram_mem1_reg[252][10]/P0001  & n13986 ;
  assign n31878 = ~n31876 & ~n31877 ;
  assign n31879 = \wishbone_bd_ram_mem1_reg[39][10]/P0001  & n13893 ;
  assign n31880 = \wishbone_bd_ram_mem1_reg[175][10]/P0001  & n13674 ;
  assign n31881 = ~n31879 & ~n31880 ;
  assign n31882 = n31878 & n31881 ;
  assign n31883 = n31875 & n31882 ;
  assign n31884 = \wishbone_bd_ram_mem1_reg[184][10]/P0001  & n13960 ;
  assign n31885 = \wishbone_bd_ram_mem1_reg[139][10]/P0001  & n13566 ;
  assign n31886 = ~n31884 & ~n31885 ;
  assign n31887 = \wishbone_bd_ram_mem1_reg[93][10]/P0001  & n13891 ;
  assign n31888 = \wishbone_bd_ram_mem1_reg[76][10]/P0001  & n13831 ;
  assign n31889 = ~n31887 & ~n31888 ;
  assign n31890 = n31886 & n31889 ;
  assign n31891 = \wishbone_bd_ram_mem1_reg[151][10]/P0001  & n13697 ;
  assign n31892 = \wishbone_bd_ram_mem1_reg[240][10]/P0001  & n13352 ;
  assign n31893 = ~n31891 & ~n31892 ;
  assign n31894 = \wishbone_bd_ram_mem1_reg[122][10]/P0001  & n13679 ;
  assign n31895 = \wishbone_bd_ram_mem1_reg[215][10]/P0001  & n13901 ;
  assign n31896 = ~n31894 & ~n31895 ;
  assign n31897 = n31893 & n31896 ;
  assign n31898 = n31890 & n31897 ;
  assign n31899 = n31883 & n31898 ;
  assign n31900 = \wishbone_bd_ram_mem1_reg[22][10]/P0001  & n13744 ;
  assign n31901 = \wishbone_bd_ram_mem1_reg[140][10]/P0001  & n13287 ;
  assign n31902 = ~n31900 & ~n31901 ;
  assign n31903 = \wishbone_bd_ram_mem1_reg[111][10]/P0001  & n13471 ;
  assign n31904 = \wishbone_bd_ram_mem1_reg[165][10]/P0001  & n14028 ;
  assign n31905 = ~n31903 & ~n31904 ;
  assign n31906 = n31902 & n31905 ;
  assign n31907 = \wishbone_bd_ram_mem1_reg[206][10]/P0001  & n13414 ;
  assign n31908 = \wishbone_bd_ram_mem1_reg[163][10]/P0001  & n13255 ;
  assign n31909 = ~n31907 & ~n31908 ;
  assign n31910 = \wishbone_bd_ram_mem1_reg[187][10]/P0001  & n13756 ;
  assign n31911 = \wishbone_bd_ram_mem1_reg[162][10]/P0001  & n13726 ;
  assign n31912 = ~n31910 & ~n31911 ;
  assign n31913 = n31909 & n31912 ;
  assign n31914 = n31906 & n31913 ;
  assign n31915 = \wishbone_bd_ram_mem1_reg[12][10]/P0001  & n13733 ;
  assign n31916 = \wishbone_bd_ram_mem1_reg[99][10]/P0001  & n13996 ;
  assign n31917 = ~n31915 & ~n31916 ;
  assign n31918 = \wishbone_bd_ram_mem1_reg[41][10]/P0001  & n14017 ;
  assign n31919 = \wishbone_bd_ram_mem1_reg[54][10]/P0001  & n13622 ;
  assign n31920 = ~n31918 & ~n31919 ;
  assign n31921 = n31917 & n31920 ;
  assign n31922 = \wishbone_bd_ram_mem1_reg[44][10]/P0001  & n13291 ;
  assign n31923 = \wishbone_bd_ram_mem1_reg[188][10]/P0001  & n13407 ;
  assign n31924 = ~n31922 & ~n31923 ;
  assign n31925 = \wishbone_bd_ram_mem1_reg[31][10]/P0001  & n13758 ;
  assign n31926 = \wishbone_bd_ram_mem1_reg[96][10]/P0001  & n13425 ;
  assign n31927 = ~n31925 & ~n31926 ;
  assign n31928 = n31924 & n31927 ;
  assign n31929 = n31921 & n31928 ;
  assign n31930 = n31914 & n31929 ;
  assign n31931 = n31899 & n31930 ;
  assign n31932 = n31868 & n31931 ;
  assign n31933 = n31805 & n31932 ;
  assign n31934 = \wishbone_bd_ram_mem1_reg[182][10]/P0001  & n13598 ;
  assign n31935 = \wishbone_bd_ram_mem1_reg[9][10]/P0001  & n13580 ;
  assign n31936 = ~n31934 & ~n31935 ;
  assign n31937 = \wishbone_bd_ram_mem1_reg[110][10]/P0001  & n14030 ;
  assign n31938 = \wishbone_bd_ram_mem1_reg[85][10]/P0001  & n13784 ;
  assign n31939 = ~n31937 & ~n31938 ;
  assign n31940 = n31936 & n31939 ;
  assign n31941 = \wishbone_bd_ram_mem1_reg[171][10]/P0001  & n13422 ;
  assign n31942 = \wishbone_bd_ram_mem1_reg[72][10]/P0001  & n13582 ;
  assign n31943 = ~n31941 & ~n31942 ;
  assign n31944 = \wishbone_bd_ram_mem1_reg[221][10]/P0001  & n13641 ;
  assign n31945 = \wishbone_bd_ram_mem1_reg[227][10]/P0001  & n13388 ;
  assign n31946 = ~n31944 & ~n31945 ;
  assign n31947 = n31943 & n31946 ;
  assign n31948 = n31940 & n31947 ;
  assign n31949 = \wishbone_bd_ram_mem1_reg[125][10]/P0001  & n13396 ;
  assign n31950 = \wishbone_bd_ram_mem1_reg[153][10]/P0001  & n13309 ;
  assign n31951 = ~n31949 & ~n31950 ;
  assign n31952 = \wishbone_bd_ram_mem1_reg[179][10]/P0001  & n14035 ;
  assign n31953 = \wishbone_bd_ram_mem1_reg[129][10]/P0001  & n13629 ;
  assign n31954 = ~n31952 & ~n31953 ;
  assign n31955 = n31951 & n31954 ;
  assign n31956 = \wishbone_bd_ram_mem1_reg[168][10]/P0001  & n13795 ;
  assign n31957 = \wishbone_bd_ram_mem1_reg[143][10]/P0001  & n13461 ;
  assign n31958 = ~n31956 & ~n31957 ;
  assign n31959 = \wishbone_bd_ram_mem1_reg[248][10]/P0001  & n13647 ;
  assign n31960 = \wishbone_bd_ram_mem1_reg[51][10]/P0001  & n13880 ;
  assign n31961 = ~n31959 & ~n31960 ;
  assign n31962 = n31958 & n31961 ;
  assign n31963 = n31955 & n31962 ;
  assign n31964 = n31948 & n31963 ;
  assign n31965 = \wishbone_bd_ram_mem1_reg[94][10]/P0001  & n13833 ;
  assign n31966 = \wishbone_bd_ram_mem1_reg[50][10]/P0001  & n13686 ;
  assign n31967 = ~n31965 & ~n31966 ;
  assign n31968 = \wishbone_bd_ram_mem1_reg[67][10]/P0001  & n13663 ;
  assign n31969 = \wishbone_bd_ram_mem1_reg[84][10]/P0001  & n13385 ;
  assign n31970 = ~n31968 & ~n31969 ;
  assign n31971 = n31967 & n31970 ;
  assign n31972 = \wishbone_bd_ram_mem1_reg[217][10]/P0001  & n13767 ;
  assign n31973 = \wishbone_bd_ram_mem1_reg[87][10]/P0001  & n13691 ;
  assign n31974 = ~n31972 & ~n31973 ;
  assign n31975 = \wishbone_bd_ram_mem1_reg[238][10]/P0001  & n13819 ;
  assign n31976 = \wishbone_bd_ram_mem1_reg[55][10]/P0001  & n13618 ;
  assign n31977 = ~n31975 & ~n31976 ;
  assign n31978 = n31974 & n31977 ;
  assign n31979 = n31971 & n31978 ;
  assign n31980 = \wishbone_bd_ram_mem1_reg[166][10]/P0001  & n13999 ;
  assign n31981 = \wishbone_bd_ram_mem1_reg[95][10]/P0001  & n13317 ;
  assign n31982 = ~n31980 & ~n31981 ;
  assign n31983 = \wishbone_bd_ram_mem1_reg[178][10]/P0001  & n13301 ;
  assign n31984 = \wishbone_bd_ram_mem1_reg[25][10]/P0001  & n13742 ;
  assign n31985 = ~n31983 & ~n31984 ;
  assign n31986 = n31982 & n31985 ;
  assign n31987 = \wishbone_bd_ram_mem1_reg[232][10]/P0001  & n13510 ;
  assign n31988 = \wishbone_bd_ram_mem1_reg[46][10]/P0001  & n13298 ;
  assign n31989 = ~n31987 & ~n31988 ;
  assign n31990 = \wishbone_bd_ram_mem1_reg[74][10]/P0001  & n13564 ;
  assign n31991 = \wishbone_bd_ram_mem1_reg[214][10]/P0001  & n13938 ;
  assign n31992 = ~n31990 & ~n31991 ;
  assign n31993 = n31989 & n31992 ;
  assign n31994 = n31986 & n31993 ;
  assign n31995 = n31979 & n31994 ;
  assign n31996 = n31964 & n31995 ;
  assign n31997 = \wishbone_bd_ram_mem1_reg[254][10]/P0001  & n13283 ;
  assign n31998 = \wishbone_bd_ram_mem1_reg[6][10]/P0001  & n13915 ;
  assign n31999 = ~n31997 & ~n31998 ;
  assign n32000 = \wishbone_bd_ram_mem1_reg[2][10]/P0001  & n13975 ;
  assign n32001 = \wishbone_bd_ram_mem1_reg[8][10]/P0001  & n13459 ;
  assign n32002 = ~n32000 & ~n32001 ;
  assign n32003 = n31999 & n32002 ;
  assign n32004 = \wishbone_bd_ram_mem1_reg[194][10]/P0001  & n13624 ;
  assign n32005 = \wishbone_bd_ram_mem1_reg[231][10]/P0001  & n13363 ;
  assign n32006 = ~n32004 & ~n32005 ;
  assign n32007 = \wishbone_bd_ram_mem1_reg[169][10]/P0001  & n13541 ;
  assign n32008 = \wishbone_bd_ram_mem1_reg[105][10]/P0001  & n13503 ;
  assign n32009 = ~n32007 & ~n32008 ;
  assign n32010 = n32006 & n32009 ;
  assign n32011 = n32003 & n32010 ;
  assign n32012 = \wishbone_bd_ram_mem1_reg[130][10]/P0001  & n13427 ;
  assign n32013 = \wishbone_bd_ram_mem1_reg[186][10]/P0001  & n13616 ;
  assign n32014 = ~n32012 & ~n32013 ;
  assign n32015 = \wishbone_bd_ram_mem1_reg[223][10]/P0001  & n13335 ;
  assign n32016 = \wishbone_bd_ram_mem1_reg[144][10]/P0001  & n13508 ;
  assign n32017 = ~n32015 & ~n32016 ;
  assign n32018 = n32014 & n32017 ;
  assign n32019 = \wishbone_bd_ram_mem1_reg[205][10]/P0001  & n13947 ;
  assign n32020 = \wishbone_bd_ram_mem1_reg[150][10]/P0001  & n13666 ;
  assign n32021 = ~n32019 & ~n32020 ;
  assign n32022 = \wishbone_bd_ram_mem1_reg[239][10]/P0001  & n13349 ;
  assign n32023 = \wishbone_bd_ram_mem1_reg[172][10]/P0001  & n13377 ;
  assign n32024 = ~n32022 & ~n32023 ;
  assign n32025 = n32021 & n32024 ;
  assign n32026 = n32018 & n32025 ;
  assign n32027 = n32011 & n32026 ;
  assign n32028 = \wishbone_bd_ram_mem1_reg[13][10]/P0001  & n13844 ;
  assign n32029 = \wishbone_bd_ram_mem1_reg[45][10]/P0001  & n13420 ;
  assign n32030 = ~n32028 & ~n32029 ;
  assign n32031 = \wishbone_bd_ram_mem1_reg[109][10]/P0001  & n13306 ;
  assign n32032 = \wishbone_bd_ram_mem1_reg[63][10]/P0001  & n13327 ;
  assign n32033 = ~n32031 & ~n32032 ;
  assign n32034 = n32030 & n32033 ;
  assign n32035 = \wishbone_bd_ram_mem1_reg[34][10]/P0001  & n13450 ;
  assign n32036 = \wishbone_bd_ram_mem1_reg[198][10]/P0001  & n13592 ;
  assign n32037 = ~n32035 & ~n32036 ;
  assign n32038 = \wishbone_bd_ram_mem1_reg[226][10]/P0001  & n13668 ;
  assign n32039 = \wishbone_bd_ram_mem1_reg[244][10]/P0001  & n13474 ;
  assign n32040 = ~n32038 & ~n32039 ;
  assign n32041 = n32037 & n32040 ;
  assign n32042 = n32034 & n32041 ;
  assign n32043 = \wishbone_bd_ram_mem1_reg[66][10]/P0001  & n13603 ;
  assign n32044 = \wishbone_bd_ram_mem1_reg[192][10]/P0001  & n13390 ;
  assign n32045 = ~n32043 & ~n32044 ;
  assign n32046 = \wishbone_bd_ram_mem1_reg[195][10]/P0001  & n13700 ;
  assign n32047 = \wishbone_bd_ram_mem1_reg[160][10]/P0001  & n13271 ;
  assign n32048 = ~n32046 & ~n32047 ;
  assign n32049 = n32045 & n32048 ;
  assign n32050 = \wishbone_bd_ram_mem1_reg[35][10]/P0001  & n13523 ;
  assign n32051 = \wishbone_bd_ram_mem1_reg[173][10]/P0001  & n13360 ;
  assign n32052 = ~n32050 & ~n32051 ;
  assign n32053 = \wishbone_bd_ram_mem1_reg[233][10]/P0001  & n13332 ;
  assign n32054 = \wishbone_bd_ram_mem1_reg[40][10]/P0001  & n13661 ;
  assign n32055 = ~n32053 & ~n32054 ;
  assign n32056 = n32052 & n32055 ;
  assign n32057 = n32049 & n32056 ;
  assign n32058 = n32042 & n32057 ;
  assign n32059 = n32027 & n32058 ;
  assign n32060 = n31996 & n32059 ;
  assign n32061 = \wishbone_bd_ram_mem1_reg[4][10]/P0001  & n13527 ;
  assign n32062 = \wishbone_bd_ram_mem1_reg[190][10]/P0001  & n13365 ;
  assign n32063 = ~n32061 & ~n32062 ;
  assign n32064 = \wishbone_bd_ram_mem1_reg[213][10]/P0001  & n13870 ;
  assign n32065 = \wishbone_bd_ram_mem1_reg[101][10]/P0001  & n13772 ;
  assign n32066 = ~n32064 & ~n32065 ;
  assign n32067 = n32063 & n32066 ;
  assign n32068 = \wishbone_bd_ram_mem1_reg[126][10]/P0001  & n13786 ;
  assign n32069 = \wishbone_bd_ram_mem1_reg[207][10]/P0001  & n13826 ;
  assign n32070 = ~n32068 & ~n32069 ;
  assign n32071 = \wishbone_bd_ram_mem1_reg[157][10]/P0001  & n13445 ;
  assign n32072 = \wishbone_bd_ram_mem1_reg[19][10]/P0001  & n13886 ;
  assign n32073 = ~n32071 & ~n32072 ;
  assign n32074 = n32070 & n32073 ;
  assign n32075 = n32067 & n32074 ;
  assign n32076 = \wishbone_bd_ram_mem1_reg[117][10]/P0001  & n13557 ;
  assign n32077 = \wishbone_bd_ram_mem1_reg[142][10]/P0001  & n13448 ;
  assign n32078 = ~n32076 & ~n32077 ;
  assign n32079 = \wishbone_bd_ram_mem1_reg[154][10]/P0001  & n13403 ;
  assign n32080 = \wishbone_bd_ram_mem1_reg[156][10]/P0001  & n13769 ;
  assign n32081 = ~n32079 & ~n32080 ;
  assign n32082 = n32078 & n32081 ;
  assign n32083 = \wishbone_bd_ram_mem1_reg[97][10]/P0001  & n13724 ;
  assign n32084 = \wishbone_bd_ram_mem1_reg[16][10]/P0001  & n13695 ;
  assign n32085 = ~n32083 & ~n32084 ;
  assign n32086 = \wishbone_bd_ram_mem1_reg[201][10]/P0001  & n13600 ;
  assign n32087 = \wishbone_bd_ram_mem1_reg[59][10]/P0001  & n13613 ;
  assign n32088 = ~n32086 & ~n32087 ;
  assign n32089 = n32085 & n32088 ;
  assign n32090 = n32082 & n32089 ;
  assign n32091 = n32075 & n32090 ;
  assign n32092 = \wishbone_bd_ram_mem1_reg[62][10]/P0001  & n13529 ;
  assign n32093 = \wishbone_bd_ram_mem1_reg[75][10]/P0001  & n13605 ;
  assign n32094 = ~n32092 & ~n32093 ;
  assign n32095 = \wishbone_bd_ram_mem1_reg[61][10]/P0001  & n13544 ;
  assign n32096 = \wishbone_bd_ram_mem1_reg[211][10]/P0001  & n13805 ;
  assign n32097 = ~n32095 & ~n32096 ;
  assign n32098 = n32094 & n32097 ;
  assign n32099 = \wishbone_bd_ram_mem1_reg[89][10]/P0001  & n13910 ;
  assign n32100 = \wishbone_bd_ram_mem1_reg[218][10]/P0001  & n13792 ;
  assign n32101 = ~n32099 & ~n32100 ;
  assign n32102 = \wishbone_bd_ram_mem1_reg[23][10]/P0001  & n13857 ;
  assign n32103 = \wishbone_bd_ram_mem1_reg[11][10]/P0001  & n13774 ;
  assign n32104 = ~n32102 & ~n32103 ;
  assign n32105 = n32101 & n32104 ;
  assign n32106 = n32098 & n32105 ;
  assign n32107 = \wishbone_bd_ram_mem1_reg[197][10]/P0001  & n13594 ;
  assign n32108 = \wishbone_bd_ram_mem1_reg[36][10]/P0001  & n13639 ;
  assign n32109 = ~n32107 & ~n32108 ;
  assign n32110 = \wishbone_bd_ram_mem1_reg[216][10]/P0001  & n14005 ;
  assign n32111 = \wishbone_bd_ram_mem1_reg[26][10]/P0001  & n13521 ;
  assign n32112 = ~n32110 & ~n32111 ;
  assign n32113 = n32109 & n32112 ;
  assign n32114 = \wishbone_bd_ram_mem1_reg[37][10]/P0001  & n13710 ;
  assign n32115 = \wishbone_bd_ram_mem1_reg[57][10]/P0001  & n13731 ;
  assign n32116 = ~n32114 & ~n32115 ;
  assign n32117 = \wishbone_bd_ram_mem1_reg[7][10]/P0001  & n13546 ;
  assign n32118 = \wishbone_bd_ram_mem1_reg[108][10]/P0001  & n13814 ;
  assign n32119 = ~n32117 & ~n32118 ;
  assign n32120 = n32116 & n32119 ;
  assign n32121 = n32113 & n32120 ;
  assign n32122 = n32106 & n32121 ;
  assign n32123 = n32091 & n32122 ;
  assign n32124 = \wishbone_bd_ram_mem1_reg[203][10]/P0001  & n13816 ;
  assign n32125 = \wishbone_bd_ram_mem1_reg[121][10]/P0001  & n13983 ;
  assign n32126 = ~n32124 & ~n32125 ;
  assign n32127 = \wishbone_bd_ram_mem1_reg[209][10]/P0001  & n13689 ;
  assign n32128 = \wishbone_bd_ram_mem1_reg[91][10]/P0001  & n13954 ;
  assign n32129 = ~n32127 & ~n32128 ;
  assign n32130 = n32126 & n32129 ;
  assign n32131 = \wishbone_bd_ram_mem1_reg[98][10]/P0001  & n13569 ;
  assign n32132 = \wishbone_bd_ram_mem1_reg[237][10]/P0001  & n13924 ;
  assign n32133 = ~n32131 & ~n32132 ;
  assign n32134 = \wishbone_bd_ram_mem1_reg[234][10]/P0001  & n13781 ;
  assign n32135 = \wishbone_bd_ram_mem1_reg[47][10]/P0001  & n13436 ;
  assign n32136 = ~n32134 & ~n32135 ;
  assign n32137 = n32133 & n32136 ;
  assign n32138 = n32130 & n32137 ;
  assign n32139 = \wishbone_bd_ram_mem1_reg[1][10]/P0001  & n13888 ;
  assign n32140 = \wishbone_bd_ram_mem1_reg[135][10]/P0001  & n13672 ;
  assign n32141 = ~n32139 & ~n32140 ;
  assign n32142 = \wishbone_bd_ram_mem1_reg[104][10]/P0001  & n13684 ;
  assign n32143 = \wishbone_bd_ram_mem1_reg[176][10]/P0001  & n13262 ;
  assign n32144 = ~n32142 & ~n32143 ;
  assign n32145 = n32141 & n32144 ;
  assign n32146 = \wishbone_bd_ram_mem1_reg[229][10]/P0001  & n13552 ;
  assign n32147 = \wishbone_bd_ram_mem1_reg[170][10]/P0001  & n14007 ;
  assign n32148 = ~n32146 & ~n32147 ;
  assign n32149 = \wishbone_bd_ram_mem1_reg[53][10]/P0001  & n13875 ;
  assign n32150 = \wishbone_bd_ram_mem1_reg[185][10]/P0001  & n13372 ;
  assign n32151 = ~n32149 & ~n32150 ;
  assign n32152 = n32148 & n32151 ;
  assign n32153 = n32145 & n32152 ;
  assign n32154 = n32138 & n32153 ;
  assign n32155 = \wishbone_bd_ram_mem1_reg[80][10]/P0001  & n13516 ;
  assign n32156 = \wishbone_bd_ram_mem1_reg[138][10]/P0001  & n13398 ;
  assign n32157 = ~n32155 & ~n32156 ;
  assign n32158 = \wishbone_bd_ram_mem1_reg[224][10]/P0001  & n13433 ;
  assign n32159 = \wishbone_bd_ram_mem1_reg[174][10]/P0001  & n13899 ;
  assign n32160 = ~n32158 & ~n32159 ;
  assign n32161 = n32157 & n32160 ;
  assign n32162 = \wishbone_bd_ram_mem1_reg[15][10]/P0001  & n13797 ;
  assign n32163 = \wishbone_bd_ram_mem1_reg[5][10]/P0001  & n13243 ;
  assign n32164 = ~n32162 & ~n32163 ;
  assign n32165 = \wishbone_bd_ram_mem1_reg[73][10]/P0001  & n13456 ;
  assign n32166 = \wishbone_bd_ram_mem1_reg[114][10]/P0001  & n13763 ;
  assign n32167 = ~n32165 & ~n32166 ;
  assign n32168 = n32164 & n32167 ;
  assign n32169 = n32161 & n32168 ;
  assign n32170 = \wishbone_bd_ram_mem1_reg[147][10]/P0001  & n13702 ;
  assign n32171 = \wishbone_bd_ram_mem1_reg[167][10]/P0001  & n13940 ;
  assign n32172 = ~n32170 & ~n32171 ;
  assign n32173 = \wishbone_bd_ram_mem1_reg[202][10]/P0001  & n13268 ;
  assign n32174 = \wishbone_bd_ram_mem1_reg[115][10]/P0001  & n13747 ;
  assign n32175 = ~n32173 & ~n32174 ;
  assign n32176 = n32172 & n32175 ;
  assign n32177 = \wishbone_bd_ram_mem1_reg[123][10]/P0001  & n13749 ;
  assign n32178 = \wishbone_bd_ram_mem1_reg[152][10]/P0001  & n13912 ;
  assign n32179 = ~n32177 & ~n32178 ;
  assign n32180 = \wishbone_bd_ram_mem1_reg[69][10]/P0001  & n13487 ;
  assign n32181 = \wishbone_bd_ram_mem1_reg[68][10]/P0001  & n13379 ;
  assign n32182 = ~n32180 & ~n32181 ;
  assign n32183 = n32179 & n32182 ;
  assign n32184 = n32176 & n32183 ;
  assign n32185 = n32169 & n32184 ;
  assign n32186 = n32154 & n32185 ;
  assign n32187 = n32123 & n32186 ;
  assign n32188 = n32060 & n32187 ;
  assign n32189 = n31933 & n32188 ;
  assign n32190 = n24387 & ~n32189 ;
  assign n32191 = n31678 & ~n32190 ;
  assign n32192 = \wishbone_TxPointerMSB_reg[10]/NET0131  & n18554 ;
  assign n32193 = ~\wishbone_TxPointerMSB_reg[11]/NET0131  & ~n32192 ;
  assign n32194 = ~n18545 & ~n31580 ;
  assign n32195 = ~n32193 & n32194 ;
  assign n32196 = n24387 & ~n28901 ;
  assign n32197 = ~n32195 & ~n32196 ;
  assign n32198 = \wishbone_TxPointerMSB_reg[13]/NET0131  & ~n18545 ;
  assign n32199 = ~n18557 & n32198 ;
  assign n32200 = ~\wishbone_TxPointerMSB_reg[13]/NET0131  & ~n18545 ;
  assign n32201 = n18557 & n32200 ;
  assign n32202 = ~n32199 & ~n32201 ;
  assign n32203 = n24387 & ~n30970 ;
  assign n32204 = n32202 & ~n32203 ;
  assign n32205 = ~\wishbone_TxPointerMSB_reg[15]/NET0131  & ~n31589 ;
  assign n32206 = \wishbone_TxPointerMSB_reg[15]/NET0131  & n18559 ;
  assign n32207 = n18557 & n32206 ;
  assign n32208 = ~n18545 & ~n32207 ;
  assign n32209 = ~n32205 & n32208 ;
  assign n32210 = ~n16296 & n24387 ;
  assign n32211 = ~n32209 & ~n32210 ;
  assign n32212 = ~n19794 & n24387 ;
  assign n32213 = ~\wishbone_TxPointerMSB_reg[16]/NET0131  & ~n32207 ;
  assign n32214 = n18558 & n18559 ;
  assign n32215 = n18557 & n32214 ;
  assign n32216 = ~n18545 & ~n32215 ;
  assign n32217 = ~n32213 & n32216 ;
  assign n32218 = ~n32212 & ~n32217 ;
  assign n32219 = ~\wishbone_TxPointerMSB_reg[17]/NET0131  & ~n32215 ;
  assign n32220 = ~n18545 & ~n18562 ;
  assign n32221 = ~n32219 & n32220 ;
  assign n32222 = ~n20833 & n24387 ;
  assign n32223 = ~n32221 & ~n32222 ;
  assign n32224 = ~n18562 & n30344 ;
  assign n32225 = ~\wishbone_TxPointerMSB_reg[18]/NET0131  & ~n18545 ;
  assign n32226 = n18562 & n32225 ;
  assign n32227 = ~n32224 & ~n32226 ;
  assign n32228 = ~n19273 & n24387 ;
  assign n32229 = n32227 & ~n32228 ;
  assign n32230 = ~\wishbone_TxPointerMSB_reg[2]/NET0131  & ~n18546 ;
  assign n32231 = \wishbone_TxPointerMSB_reg[2]/NET0131  & n18546 ;
  assign n32232 = ~n18545 & ~n32231 ;
  assign n32233 = ~n32230 & n32232 ;
  assign n32234 = n24387 & ~n29475 ;
  assign n32235 = ~n32233 & ~n32234 ;
  assign n32236 = ~\wishbone_TxPointerMSB_reg[3]/NET0131  & ~n32231 ;
  assign n32237 = ~n18545 & ~n18548 ;
  assign n32238 = ~n32236 & n32237 ;
  assign n32239 = n24387 & ~n25612 ;
  assign n32240 = ~n32238 & ~n32239 ;
  assign n32241 = \wishbone_TxPointerMSB_reg[7]/NET0131  & n18551 ;
  assign n32242 = ~\wishbone_TxPointerMSB_reg[8]/NET0131  & ~n32241 ;
  assign n32243 = ~n18545 & ~n30430 ;
  assign n32244 = ~n32242 & n32243 ;
  assign n32245 = n24387 & ~n27806 ;
  assign n32246 = ~n32244 & ~n32245 ;
  assign n32247 = ~\miim1_clkgen_Counter_reg[0]/NET0131  & ~\miim1_clkgen_Counter_reg[1]/NET0131  ;
  assign n32248 = ~\miim1_clkgen_Counter_reg[2]/NET0131  & ~\miim1_clkgen_Counter_reg[3]/NET0131  ;
  assign n32249 = n32247 & n32248 ;
  assign n32250 = ~\miim1_clkgen_Counter_reg[4]/NET0131  & n32249 ;
  assign n32251 = \miim1_clkgen_Counter_reg[4]/NET0131  & ~n32249 ;
  assign n32252 = ~n32250 & ~n32251 ;
  assign n32253 = ~\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  & ~\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  ;
  assign n32254 = ~\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  & ~\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  ;
  assign n32255 = n32253 & n32254 ;
  assign n32256 = ~\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  & ~\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  ;
  assign n32257 = ~\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  & n32256 ;
  assign n32258 = ~n32255 & n32257 ;
  assign n32259 = ~\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  & n32258 ;
  assign n32260 = \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  & ~n32259 ;
  assign n32261 = n32253 & n32258 ;
  assign n32262 = ~\miim1_clkgen_Counter_reg[4]/NET0131  & ~\miim1_clkgen_Counter_reg[6]/NET0131  ;
  assign n32263 = ~\miim1_clkgen_Counter_reg[5]/NET0131  & n32262 ;
  assign n32264 = n32249 & n32263 ;
  assign n32265 = ~n32261 & n32264 ;
  assign n32266 = ~n32260 & n32265 ;
  assign n32267 = ~n32252 & ~n32266 ;
  assign n32268 = \wishbone_RxReady_reg/NET0131  & n15726 ;
  assign n32269 = \wishbone_LastByteIn_reg/NET0131  & \wishbone_RxByteCnt_reg[0]/NET0131  ;
  assign n32270 = \rxethmac1_RxValid_reg/NET0131  & \wishbone_RxReady_reg/NET0131  ;
  assign n32271 = \wishbone_RxByteCnt_reg[0]/NET0131  & \wishbone_RxEnableWindow_reg/NET0131  ;
  assign n32272 = n32270 & n32271 ;
  assign n32273 = ~n32269 & ~n32272 ;
  assign n32274 = \wishbone_RxEnableWindow_reg/NET0131  & n32270 ;
  assign n32275 = ~\wishbone_LastByteIn_reg/NET0131  & ~\wishbone_RxByteCnt_reg[0]/NET0131  ;
  assign n32276 = ~n32274 & n32275 ;
  assign n32277 = n32273 & ~n32276 ;
  assign n32278 = ~n32268 & ~n32277 ;
  assign n32279 = ~\RxAbort_wb_reg/NET0131  & ~\wishbone_ShiftEnded_rck_reg/NET0131  ;
  assign n32280 = ~n15728 & n32279 ;
  assign n32281 = ~n32278 & n32280 ;
  assign n32282 = ~\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  & ~n15151 ;
  assign n32283 = \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  & n15151 ;
  assign n32284 = n15162 & ~n32283 ;
  assign n32285 = ~n32282 & n32284 ;
  assign n32286 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & ~\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131  ;
  assign n32287 = n12266 & ~n32286 ;
  assign n32288 = \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  ;
  assign n32289 = n32287 & n32288 ;
  assign n32290 = \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  & \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n32291 = n32289 & n32290 ;
  assign n32292 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  & ~n32291 ;
  assign n32293 = \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  & \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  ;
  assign n32294 = \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  & n32293 ;
  assign n32295 = n32289 & n32294 ;
  assign n32296 = ~\rxethmac1_RxEndFrm_reg/NET0131  & ~n32295 ;
  assign n32297 = ~n32292 & n32296 ;
  assign n32298 = ~\wishbone_RxByteCnt_reg[1]/NET0131  & ~n32268 ;
  assign n32299 = n32273 & n32298 ;
  assign n32300 = \wishbone_RxByteCnt_reg[1]/NET0131  & ~n32268 ;
  assign n32301 = ~n32273 & n32300 ;
  assign n32302 = ~n32299 & ~n32301 ;
  assign n32303 = \wishbone_RxPointerLSB_rst_reg[0]/NET0131  & ~\wishbone_RxPointerLSB_rst_reg[1]/NET0131  ;
  assign n32304 = ~\wishbone_RxPointerLSB_rst_reg[0]/NET0131  & \wishbone_RxPointerLSB_rst_reg[1]/NET0131  ;
  assign n32305 = ~n32303 & ~n32304 ;
  assign n32306 = n32268 & n32305 ;
  assign n32307 = n32279 & ~n32306 ;
  assign n32308 = n32302 & n32307 ;
  assign n32309 = \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  & n12265 ;
  assign n32310 = n12266 & n13225 ;
  assign n32311 = n32309 & n32310 ;
  assign n32312 = n32287 & ~n32311 ;
  assign n32313 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & ~n32312 ;
  assign n32314 = \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  & n32287 ;
  assign n32315 = ~\rxethmac1_RxEndFrm_reg/NET0131  & ~n32314 ;
  assign n32316 = ~n32313 & n32315 ;
  assign n32317 = \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  & ~\rxethmac1_RxEndFrm_reg/NET0131  ;
  assign n32318 = ~n32289 & n32317 ;
  assign n32319 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  & ~\rxethmac1_RxEndFrm_reg/NET0131  ;
  assign n32320 = n32289 & n32319 ;
  assign n32321 = ~n32318 & ~n32320 ;
  assign n32322 = \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  & n32289 ;
  assign n32323 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  & ~n32322 ;
  assign n32324 = ~\rxethmac1_RxEndFrm_reg/NET0131  & ~n32291 ;
  assign n32325 = ~n32323 & n32324 ;
  assign n32326 = \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  & n15162 ;
  assign n32327 = ~n15157 & n32326 ;
  assign n32328 = ~\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  & n15162 ;
  assign n32329 = n15157 & n32328 ;
  assign n32330 = ~n32327 & ~n32329 ;
  assign n32331 = ~\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  & ~n20854 ;
  assign n32332 = \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  ;
  assign n32333 = \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  & n32332 ;
  assign n32334 = n15157 & n32333 ;
  assign n32335 = n15162 & ~n32334 ;
  assign n32336 = ~n32331 & n32335 ;
  assign n32337 = \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  & n15145 ;
  assign n32338 = n15151 & n32337 ;
  assign n32339 = ~\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  & ~n32338 ;
  assign n32340 = \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  & n32337 ;
  assign n32341 = n15151 & n32340 ;
  assign n32342 = n15162 & ~n32341 ;
  assign n32343 = ~n32339 & n32342 ;
  assign n32344 = ~\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  & ~n32341 ;
  assign n32345 = \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  ;
  assign n32346 = n32337 & n32345 ;
  assign n32347 = n15151 & n32346 ;
  assign n32348 = n15162 & ~n32347 ;
  assign n32349 = ~n32344 & n32348 ;
  assign n32350 = ~\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  & ~n32283 ;
  assign n32351 = n15139 & n15151 ;
  assign n32352 = n15162 & ~n32351 ;
  assign n32353 = ~n32350 & n32352 ;
  assign n32354 = ~\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  & ~n32351 ;
  assign n32355 = ~n15154 & n15162 ;
  assign n32356 = ~n32354 & n32355 ;
  assign n32357 = \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  & n15161 ;
  assign n32358 = ~n11392 & n32357 ;
  assign n32359 = ~n15154 & n32358 ;
  assign n32360 = ~\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  & n15161 ;
  assign n32361 = ~n11392 & n32360 ;
  assign n32362 = n15154 & n32361 ;
  assign n32363 = ~n32359 & ~n32362 ;
  assign n32364 = \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  & n15154 ;
  assign n32365 = ~\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  & ~n32364 ;
  assign n32366 = \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n32367 = n15154 & n32366 ;
  assign n32368 = n15162 & ~n32367 ;
  assign n32369 = ~n32365 & n32368 ;
  assign n32370 = ~\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  & ~n32367 ;
  assign n32371 = \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n32372 = \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  & n32371 ;
  assign n32373 = n15154 & n32372 ;
  assign n32374 = n15162 & ~n32373 ;
  assign n32375 = ~n32370 & n32374 ;
  assign n32376 = \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  & n15162 ;
  assign n32377 = ~n32373 & n32376 ;
  assign n32378 = ~\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  & n15162 ;
  assign n32379 = n32373 & n32378 ;
  assign n32380 = ~n32377 & ~n32379 ;
  assign n32381 = \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  & n32373 ;
  assign n32382 = ~\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  & ~n32381 ;
  assign n32383 = n15135 & n32373 ;
  assign n32384 = n15162 & ~n32383 ;
  assign n32385 = ~n32382 & n32384 ;
  assign n32386 = ~\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  & ~n32383 ;
  assign n32387 = \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  & n15138 ;
  assign n32388 = n15154 & n32387 ;
  assign n32389 = n15162 & ~n32388 ;
  assign n32390 = ~n32386 & n32389 ;
  assign n32391 = n15138 & n15141 ;
  assign n32392 = n15151 & n32391 ;
  assign n32393 = ~\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  & ~n32392 ;
  assign n32394 = \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  & n15141 ;
  assign n32395 = n15138 & n32394 ;
  assign n32396 = n15151 & n32395 ;
  assign n32397 = n15162 & ~n32396 ;
  assign n32398 = ~n32393 & n32397 ;
  assign n32399 = ~\txethmac1_txcrc_Crc_reg[3]/NET0131  & n12974 ;
  assign n32400 = n12961 & n32399 ;
  assign n32401 = ~\txethmac1_txcrc_Crc_reg[3]/NET0131  & n11464 ;
  assign n32402 = ~n12979 & ~n32401 ;
  assign n32403 = ~n32400 & ~n32402 ;
  assign n32404 = ~\txethmac1_txcrc_Crc_reg[2]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n32405 = n11626 & n32404 ;
  assign n32406 = ~\txethmac1_txcrc_Crc_reg[2]/NET0131  & n11464 ;
  assign n32407 = ~\txethmac1_txstatem1_StateFCS_reg/NET0131  & n11464 ;
  assign n32408 = n11626 & n32407 ;
  assign n32409 = ~n32406 & ~n32408 ;
  assign n32410 = ~n32405 & ~n32409 ;
  assign n32411 = ~\wishbone_cyc_cleared_reg/NET0131  & ~n13131 ;
  assign n32412 = ~n13182 & ~n32411 ;
  assign n32413 = n13128 & ~n13147 ;
  assign n32414 = n13127 & n32413 ;
  assign n32415 = ~n32412 & n32414 ;
  assign n32416 = ~n13177 & ~n13184 ;
  assign n32417 = ~n32415 & n32416 ;
  assign n32418 = n13178 & n32414 ;
  assign n32419 = ~n13176 & n32412 ;
  assign n32420 = ~n32418 & ~n32419 ;
  assign n32421 = ~n32417 & n32420 ;
  assign n32422 = \wishbone_MasterWbRX_reg/NET0131  & \wishbone_rx_burst_en_reg/NET0131  ;
  assign n32423 = ~n13129 & n32422 ;
  assign n32424 = ~\wishbone_MasterWbRX_reg/NET0131  & \wishbone_tx_burst_en_reg/NET0131  ;
  assign n32425 = n13147 & n32424 ;
  assign n32426 = n13184 & n32411 ;
  assign n32427 = ~n32425 & n32426 ;
  assign n32428 = ~n32414 & n32427 ;
  assign n32429 = ~n32423 & n32428 ;
  assign n32430 = ~n32415 & ~n32429 ;
  assign n32431 = n32421 & n32430 ;
  assign n32432 = \m_wb_sel_o[0]_pad  & ~n32431 ;
  assign n32433 = n13197 & ~n32432 ;
  assign n32434 = \macstatus1_InvalidSymbol_reg/NET0131  & ~\macstatus1_LoadRxStatus_reg/NET0131  ;
  assign n32435 = \ethreg1_MODER_0_DataOut_reg[7]/NET0131  & mtxerr_pad_o_pad ;
  assign n32436 = \RxEnSync_reg/NET0131  & ~\ethreg1_MODER_0_DataOut_reg[7]/NET0131  ;
  assign n32437 = mrxerr_pad_i_pad & n32436 ;
  assign n32438 = ~n32435 & ~n32437 ;
  assign n32439 = ~n10653 & ~n32438 ;
  assign n32440 = ~n10671 & ~n11356 ;
  assign n32441 = n12207 & n32440 ;
  assign n32442 = n32439 & n32441 ;
  assign n32443 = ~n32434 & ~n32442 ;
  assign n32444 = \wishbone_ShiftEndedSync_c1_reg/NET0131  & \wishbone_ShiftEndedSync_c2_reg/NET0131  ;
  assign n32445 = \wishbone_ShiftEnded_rck_reg/NET0131  & ~n32444 ;
  assign n32446 = \rxethmac1_RxEndFrm_reg/NET0131  & \rxethmac1_RxValid_reg/NET0131  ;
  assign n32447 = \wishbone_RxByteCnt_reg[1]/NET0131  & \wishbone_RxEnableWindow_reg/NET0131  ;
  assign n32448 = \wishbone_RxByteCnt_reg[0]/NET0131  & n32447 ;
  assign n32449 = n32446 & n32448 ;
  assign n32450 = ~\wishbone_LastByteIn_reg/NET0131  & ~n32449 ;
  assign n32451 = ~n32445 & n32450 ;
  assign n32452 = ~n15737 & ~n32445 ;
  assign n32453 = n15735 & n32452 ;
  assign n32454 = ~n32451 & ~n32453 ;
  assign n32455 = ~\RxAbort_wb_reg/NET0131  & n32454 ;
  assign n32456 = ~\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  & ~n32314 ;
  assign n32457 = ~\rxethmac1_RxEndFrm_reg/NET0131  & ~n32289 ;
  assign n32458 = ~n32456 & n32457 ;
  assign n32459 = m_wb_stb_o_pad & ~n32421 ;
  assign n32460 = n13197 & ~n32459 ;
  assign n32461 = \wishbone_tx_burst_cnt_reg[0]/NET0131  & \wishbone_tx_burst_cnt_reg[1]/NET0131  ;
  assign n32462 = ~\wishbone_tx_burst_cnt_reg[2]/NET0131  & n32461 ;
  assign n32463 = ~n13166 & ~n32462 ;
  assign n32464 = ~n13164 & n32463 ;
  assign n32465 = \wishbone_tx_burst_en_reg/NET0131  & n32464 ;
  assign n32466 = ~n32418 & ~n32429 ;
  assign n32467 = \wishbone_tx_burst_en_reg/NET0131  & ~n13174 ;
  assign n32468 = n32466 & n32467 ;
  assign n32469 = ~n32465 & ~n32468 ;
  assign n32470 = \wishbone_TxLength_reg[3]/NET0131  & \wishbone_TxLength_reg[4]/NET0131  ;
  assign n32471 = \wishbone_TxLength_reg[2]/NET0131  & \wishbone_TxLength_reg[4]/NET0131  ;
  assign n32472 = ~n17372 & n32471 ;
  assign n32473 = ~n32470 & ~n32472 ;
  assign n32474 = n14053 & n14056 ;
  assign n32475 = n14063 & n32474 ;
  assign n32476 = n32473 & n32475 ;
  assign n32477 = \wishbone_tx_fifo_cnt_reg[2]/NET0131  & \wishbone_tx_fifo_cnt_reg[3]/NET0131  ;
  assign n32478 = ~\wishbone_tx_fifo_cnt_reg[4]/NET0131  & ~n32477 ;
  assign n32479 = ~n32476 & n32478 ;
  assign n32480 = ~n32466 & n32479 ;
  assign n32481 = n32469 & ~n32480 ;
  assign n32482 = \wishbone_IncrTxPointer_reg/NET0131  & ~n32421 ;
  assign n32483 = n13189 & ~n32482 ;
  assign n32484 = n13175 & n13185 ;
  assign n32485 = ~n13181 & n32484 ;
  assign n32486 = ~n13191 & ~n32485 ;
  assign n32487 = n13192 & n13193 ;
  assign n32488 = \wishbone_cyc_cleared_reg/NET0131  & ~n32415 ;
  assign n32489 = ~n32487 & n32488 ;
  assign n32490 = ~n13174 & n32489 ;
  assign n32491 = n32486 & n32490 ;
  assign n32492 = ~n32429 & ~n32491 ;
  assign n32493 = n11182 & n11402 ;
  assign n32494 = ~\txethmac1_StatusLatch_reg/NET0131  & ~\txethmac1_txstatem1_StateIdle_reg/NET0131  ;
  assign n32495 = ~n32493 & n32494 ;
  assign n32496 = ~n11186 & ~n32495 ;
  assign n32497 = ~\rxethmac1_rxstatem1_StatePreamble_reg/NET0131  & ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n32498 = n10649 & n32497 ;
  assign n32499 = ~n12540 & n32498 ;
  assign n32500 = n32439 & ~n32499 ;
  assign n32501 = ~\wishbone_WriteRxDataToFifoSync2_reg/NET0131  & \wishbone_WriteRxDataToFifo_reg/NET0131  ;
  assign n32502 = ~n15737 & ~n32501 ;
  assign n32503 = n15735 & n32502 ;
  assign n32504 = ~\RxAbort_wb_reg/NET0131  & ~n32503 ;
  assign n32505 = \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  & ~n32258 ;
  assign n32506 = ~n32259 & n32264 ;
  assign n32507 = ~n32505 & n32506 ;
  assign n32508 = ~\miim1_clkgen_Counter_reg[2]/NET0131  & n32247 ;
  assign n32509 = \miim1_clkgen_Counter_reg[3]/NET0131  & ~n32508 ;
  assign n32510 = ~n32249 & ~n32509 ;
  assign n32511 = ~n32264 & n32510 ;
  assign n32512 = ~n32507 & ~n32511 ;
  assign n32513 = mdc_pad_o_pad & n32264 ;
  assign n32514 = \miim1_shftrg_ShiftReg_reg[1]/NET0131  & ~n32513 ;
  assign n32515 = ~n32513 & ~n32514 ;
  assign n32516 = \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131  & ~\miim1_BitCounter_reg[2]/NET0131  ;
  assign n32517 = ~\miim1_BitCounter_reg[3]/NET0131  & ~\miim1_BitCounter_reg[4]/NET0131  ;
  assign n32518 = n32516 & n32517 ;
  assign n32519 = ~\miim1_BitCounter_reg[0]/NET0131  & ~\miim1_BitCounter_reg[1]/NET0131  ;
  assign n32520 = ~\miim1_BitCounter_reg[5]/NET0131  & ~\miim1_BitCounter_reg[6]/NET0131  ;
  assign n32521 = n32519 & n32520 ;
  assign n32522 = n32518 & n32521 ;
  assign n32523 = \miim1_InProgress_reg/NET0131  & n32522 ;
  assign n32524 = ~\miim1_BitCounter_reg[2]/NET0131  & \miim1_BitCounter_reg[5]/NET0131  ;
  assign n32525 = n32519 & n32524 ;
  assign n32526 = ~\miim1_BitCounter_reg[6]/NET0131  & \miim1_InProgress_reg/NET0131  ;
  assign n32527 = ~\miim1_BitCounter_reg[4]/NET0131  & n32526 ;
  assign n32528 = ~\ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n32529 = n32527 & n32528 ;
  assign n32530 = n32525 & n32529 ;
  assign n32531 = ~n32523 & ~n32530 ;
  assign n32532 = \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131  & ~n32531 ;
  assign n32533 = \miim1_BitCounter_reg[3]/NET0131  & ~\miim1_BitCounter_reg[4]/NET0131  ;
  assign n32534 = n32526 & n32533 ;
  assign n32535 = n32525 & n32534 ;
  assign n32536 = \miim1_BitCounter_reg[4]/NET0131  & \miim1_WriteOp_reg/NET0131  ;
  assign n32537 = n32526 & n32536 ;
  assign n32538 = n32525 & n32537 ;
  assign n32539 = ~\ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n32540 = ~\ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n32541 = ~n32539 & ~n32540 ;
  assign n32542 = n32538 & n32541 ;
  assign n32543 = ~n32535 & ~n32542 ;
  assign n32544 = ~n32532 & n32543 ;
  assign n32545 = ~n32535 & ~n32538 ;
  assign n32546 = \miim1_shftrg_ShiftReg_reg[0]/NET0131  & n32545 ;
  assign n32547 = n32531 & n32546 ;
  assign n32548 = ~n32514 & ~n32547 ;
  assign n32549 = n32544 & n32548 ;
  assign n32550 = ~n32515 & ~n32549 ;
  assign n32551 = \miim1_shftrg_ShiftReg_reg[2]/NET0131  & ~n32513 ;
  assign n32552 = ~n32513 & ~n32551 ;
  assign n32553 = \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131  & ~n32531 ;
  assign n32554 = \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n32555 = n32538 & n32554 ;
  assign n32556 = \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n32557 = n32538 & n32556 ;
  assign n32558 = \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131  & n32535 ;
  assign n32559 = ~n32557 & ~n32558 ;
  assign n32560 = ~n32555 & n32559 ;
  assign n32561 = ~n32553 & n32560 ;
  assign n32562 = \miim1_shftrg_ShiftReg_reg[1]/NET0131  & n32545 ;
  assign n32563 = n32531 & n32562 ;
  assign n32564 = ~n32551 & ~n32563 ;
  assign n32565 = n32561 & n32564 ;
  assign n32566 = ~n32552 & ~n32565 ;
  assign n32567 = \miim1_shftrg_ShiftReg_reg[3]/NET0131  & ~n32513 ;
  assign n32568 = ~n32513 & ~n32567 ;
  assign n32569 = \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131  & ~n32531 ;
  assign n32570 = \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n32571 = n32538 & n32570 ;
  assign n32572 = \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n32573 = n32538 & n32572 ;
  assign n32574 = \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131  & n32535 ;
  assign n32575 = ~n32573 & ~n32574 ;
  assign n32576 = ~n32571 & n32575 ;
  assign n32577 = ~n32569 & n32576 ;
  assign n32578 = \miim1_shftrg_ShiftReg_reg[2]/NET0131  & n32545 ;
  assign n32579 = n32531 & n32578 ;
  assign n32580 = ~n32567 & ~n32579 ;
  assign n32581 = n32577 & n32580 ;
  assign n32582 = ~n32568 & ~n32581 ;
  assign n32583 = \miim1_shftrg_ShiftReg_reg[4]/NET0131  & ~n32513 ;
  assign n32584 = ~n32513 & ~n32583 ;
  assign n32585 = \miim1_WriteOp_reg/NET0131  & ~n32531 ;
  assign n32586 = \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n32587 = n32538 & n32586 ;
  assign n32588 = \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n32589 = n32538 & n32588 ;
  assign n32590 = \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131  & n32535 ;
  assign n32591 = ~n32589 & ~n32590 ;
  assign n32592 = ~n32587 & n32591 ;
  assign n32593 = ~n32585 & n32592 ;
  assign n32594 = \miim1_shftrg_ShiftReg_reg[3]/NET0131  & n32545 ;
  assign n32595 = n32531 & n32594 ;
  assign n32596 = ~n32583 & ~n32595 ;
  assign n32597 = n32593 & n32596 ;
  assign n32598 = ~n32584 & ~n32597 ;
  assign n32599 = \miim1_shftrg_ShiftReg_reg[5]/NET0131  & ~n32513 ;
  assign n32600 = ~n32513 & ~n32599 ;
  assign n32601 = ~\miim1_WriteOp_reg/NET0131  & ~n32531 ;
  assign n32602 = \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n32603 = n32538 & n32602 ;
  assign n32604 = \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n32605 = n32538 & n32604 ;
  assign n32606 = \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131  & n32535 ;
  assign n32607 = ~n32605 & ~n32606 ;
  assign n32608 = ~n32603 & n32607 ;
  assign n32609 = ~n32601 & n32608 ;
  assign n32610 = \miim1_shftrg_ShiftReg_reg[4]/NET0131  & n32545 ;
  assign n32611 = n32531 & n32610 ;
  assign n32612 = ~n32599 & ~n32611 ;
  assign n32613 = n32609 & n32612 ;
  assign n32614 = ~n32600 & ~n32613 ;
  assign n32615 = \miim1_shftrg_ShiftReg_reg[6]/NET0131  & ~n32513 ;
  assign n32616 = \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131  & n32535 ;
  assign n32617 = \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n32618 = n32538 & n32617 ;
  assign n32619 = ~n32616 & ~n32618 ;
  assign n32620 = n32531 & n32619 ;
  assign n32621 = \miim1_shftrg_ShiftReg_reg[5]/NET0131  & n32545 ;
  assign n32622 = \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n32623 = n32538 & n32622 ;
  assign n32624 = ~n32621 & ~n32623 ;
  assign n32625 = n32620 & n32624 ;
  assign n32626 = n32513 & ~n32625 ;
  assign n32627 = ~n32615 & ~n32626 ;
  assign n32628 = ~\txethmac1_TxAbort_reg/NET0131  & n11558 ;
  assign n32629 = n11551 & n32628 ;
  assign n32630 = ~n11567 & ~n32493 ;
  assign n32631 = ~n32629 & ~n32630 ;
  assign n32632 = ~\ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32633 = \rxethmac1_CrcHash_reg[3]/P0001  & ~\rxethmac1_CrcHash_reg[4]/P0001  ;
  assign n32634 = ~\ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32635 = n32633 & ~n32634 ;
  assign n32636 = ~n32632 & n32635 ;
  assign n32637 = ~\rxethmac1_CrcHash_reg[0]/P0001  & ~n32636 ;
  assign n32638 = ~\ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32639 = ~\rxethmac1_CrcHash_reg[3]/P0001  & ~\rxethmac1_CrcHash_reg[4]/P0001  ;
  assign n32640 = ~\ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32641 = n32639 & ~n32640 ;
  assign n32642 = ~n32638 & n32641 ;
  assign n32643 = ~\ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32644 = \rxethmac1_CrcHash_reg[3]/P0001  & \rxethmac1_CrcHash_reg[4]/P0001  ;
  assign n32645 = ~\ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32646 = n32644 & ~n32645 ;
  assign n32647 = ~n32643 & n32646 ;
  assign n32648 = ~\ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32649 = ~\rxethmac1_CrcHash_reg[3]/P0001  & \rxethmac1_CrcHash_reg[4]/P0001  ;
  assign n32650 = ~\ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32651 = n32649 & ~n32650 ;
  assign n32652 = ~n32648 & n32651 ;
  assign n32653 = ~n32647 & ~n32652 ;
  assign n32654 = ~n32642 & n32653 ;
  assign n32655 = n32637 & n32654 ;
  assign n32656 = ~\ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32657 = ~\ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32658 = n32633 & ~n32657 ;
  assign n32659 = ~n32656 & n32658 ;
  assign n32660 = \rxethmac1_CrcHash_reg[0]/P0001  & ~n32659 ;
  assign n32661 = ~\ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32662 = ~\ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32663 = n32639 & ~n32662 ;
  assign n32664 = ~n32661 & n32663 ;
  assign n32665 = ~\ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32666 = ~\ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32667 = n32649 & ~n32666 ;
  assign n32668 = ~n32665 & n32667 ;
  assign n32669 = ~\ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32670 = ~\ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32671 = n32644 & ~n32670 ;
  assign n32672 = ~n32669 & n32671 ;
  assign n32673 = ~n32668 & ~n32672 ;
  assign n32674 = ~n32664 & n32673 ;
  assign n32675 = n32660 & n32674 ;
  assign n32676 = ~n32655 & ~n32675 ;
  assign n32677 = \rxethmac1_CrcHash_reg[1]/P0001  & ~\rxethmac1_CrcHash_reg[2]/P0001  ;
  assign n32678 = n32676 & n32677 ;
  assign n32679 = ~\ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32680 = ~\ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32681 = n32639 & ~n32680 ;
  assign n32682 = ~n32679 & n32681 ;
  assign n32683 = \rxethmac1_CrcHash_reg[0]/P0001  & ~n32682 ;
  assign n32684 = ~\ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32685 = ~\ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32686 = n32649 & ~n32685 ;
  assign n32687 = ~n32684 & n32686 ;
  assign n32688 = ~\ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32689 = ~\ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32690 = n32633 & ~n32689 ;
  assign n32691 = ~n32688 & n32690 ;
  assign n32692 = ~\ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32693 = ~\ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32694 = n32644 & ~n32693 ;
  assign n32695 = ~n32692 & n32694 ;
  assign n32696 = ~n32691 & ~n32695 ;
  assign n32697 = ~n32687 & n32696 ;
  assign n32698 = n32683 & n32697 ;
  assign n32699 = ~\ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32700 = ~\ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32701 = n32644 & ~n32700 ;
  assign n32702 = ~n32699 & n32701 ;
  assign n32703 = ~\rxethmac1_CrcHash_reg[0]/P0001  & ~n32702 ;
  assign n32704 = ~\ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32705 = ~\ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32706 = n32639 & ~n32705 ;
  assign n32707 = ~n32704 & n32706 ;
  assign n32708 = ~\ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32709 = ~\ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32710 = n32649 & ~n32709 ;
  assign n32711 = ~n32708 & n32710 ;
  assign n32712 = ~\ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32713 = ~\ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32714 = n32633 & ~n32713 ;
  assign n32715 = ~n32712 & n32714 ;
  assign n32716 = ~n32711 & ~n32715 ;
  assign n32717 = ~n32707 & n32716 ;
  assign n32718 = n32703 & n32717 ;
  assign n32719 = ~n32698 & ~n32718 ;
  assign n32720 = ~\rxethmac1_CrcHash_reg[1]/P0001  & ~\rxethmac1_CrcHash_reg[2]/P0001  ;
  assign n32721 = n32719 & n32720 ;
  assign n32722 = ~n32678 & ~n32721 ;
  assign n32723 = \rxethmac1_CrcHashGood_reg/P0001  & \rxethmac1_Multicast_reg/NET0131  ;
  assign n32724 = ~\ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32725 = ~\ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32726 = n32639 & ~n32725 ;
  assign n32727 = ~n32724 & n32726 ;
  assign n32728 = ~\rxethmac1_CrcHash_reg[0]/P0001  & ~n32727 ;
  assign n32729 = ~\ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32730 = ~\ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32731 = n32644 & ~n32730 ;
  assign n32732 = ~n32729 & n32731 ;
  assign n32733 = ~\ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32734 = ~\ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32735 = n32633 & ~n32734 ;
  assign n32736 = ~n32733 & n32735 ;
  assign n32737 = ~\ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32738 = ~\ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32739 = n32649 & ~n32738 ;
  assign n32740 = ~n32737 & n32739 ;
  assign n32741 = ~n32736 & ~n32740 ;
  assign n32742 = ~n32732 & n32741 ;
  assign n32743 = n32728 & n32742 ;
  assign n32744 = ~\ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32745 = ~\ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32746 = n32639 & ~n32745 ;
  assign n32747 = ~n32744 & n32746 ;
  assign n32748 = \rxethmac1_CrcHash_reg[0]/P0001  & ~n32747 ;
  assign n32749 = ~\ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32750 = ~\ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32751 = n32633 & ~n32750 ;
  assign n32752 = ~n32749 & n32751 ;
  assign n32753 = ~\ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32754 = ~\ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32755 = n32649 & ~n32754 ;
  assign n32756 = ~n32753 & n32755 ;
  assign n32757 = ~\ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32758 = ~\ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32759 = n32644 & ~n32758 ;
  assign n32760 = ~n32757 & n32759 ;
  assign n32761 = ~n32756 & ~n32760 ;
  assign n32762 = ~n32752 & n32761 ;
  assign n32763 = n32748 & n32762 ;
  assign n32764 = ~n32743 & ~n32763 ;
  assign n32765 = \rxethmac1_CrcHash_reg[1]/P0001  & \rxethmac1_CrcHash_reg[2]/P0001  ;
  assign n32766 = n32764 & n32765 ;
  assign n32767 = ~\ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32768 = ~\ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32769 = n32644 & ~n32768 ;
  assign n32770 = ~n32767 & n32769 ;
  assign n32771 = \rxethmac1_CrcHash_reg[0]/P0001  & ~n32770 ;
  assign n32772 = ~\ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32773 = ~\ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32774 = n32633 & ~n32773 ;
  assign n32775 = ~n32772 & n32774 ;
  assign n32776 = ~\ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32777 = ~\ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32778 = n32649 & ~n32777 ;
  assign n32779 = ~n32776 & n32778 ;
  assign n32780 = ~\ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32781 = ~\ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32782 = n32639 & ~n32781 ;
  assign n32783 = ~n32780 & n32782 ;
  assign n32784 = ~n32779 & ~n32783 ;
  assign n32785 = ~n32775 & n32784 ;
  assign n32786 = n32771 & n32785 ;
  assign n32787 = ~\ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32788 = ~\ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32789 = n32639 & ~n32788 ;
  assign n32790 = ~n32787 & n32789 ;
  assign n32791 = ~\rxethmac1_CrcHash_reg[0]/P0001  & ~n32790 ;
  assign n32792 = ~\ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32793 = ~\ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32794 = n32644 & ~n32793 ;
  assign n32795 = ~n32792 & n32794 ;
  assign n32796 = ~\ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32797 = ~\ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32798 = n32633 & ~n32797 ;
  assign n32799 = ~n32796 & n32798 ;
  assign n32800 = ~\ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131  & \rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32801 = ~\ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131  & ~\rxethmac1_CrcHash_reg[5]/P0001  ;
  assign n32802 = n32649 & ~n32801 ;
  assign n32803 = ~n32800 & n32802 ;
  assign n32804 = ~n32799 & ~n32803 ;
  assign n32805 = ~n32795 & n32804 ;
  assign n32806 = n32791 & n32805 ;
  assign n32807 = ~n32786 & ~n32806 ;
  assign n32808 = ~\rxethmac1_CrcHash_reg[1]/P0001  & \rxethmac1_CrcHash_reg[2]/P0001  ;
  assign n32809 = n32807 & n32808 ;
  assign n32810 = ~n32766 & ~n32809 ;
  assign n32811 = n32723 & n32810 ;
  assign n32812 = n32722 & n32811 ;
  assign n32813 = ~\rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131  & ~n32723 ;
  assign n32814 = n13019 & ~n32813 ;
  assign n32815 = ~n32812 & n32814 ;
  assign n32816 = ~\wb_adr_i[11]_pad  & \wb_sel_i[0]_pad  ;
  assign n32817 = n23726 & n32816 ;
  assign n32818 = ~n23725 & n32817 ;
  assign n32819 = ~\wb_adr_i[10]_pad  & wb_we_i_pad ;
  assign n32820 = n32818 & n32819 ;
  assign n32821 = ~\wb_adr_i[4]_pad  & \wb_adr_i[5]_pad  ;
  assign n32822 = ~\wb_adr_i[2]_pad  & ~\wb_adr_i[3]_pad  ;
  assign n32823 = ~\wb_adr_i[6]_pad  & ~\wb_dat_i[10]_pad  ;
  assign n32824 = n32822 & n32823 ;
  assign n32825 = n32821 & n32824 ;
  assign n32826 = ~\wb_dat_i[15]_pad  & ~\wb_dat_i[16]_pad  ;
  assign n32827 = ~\wb_dat_i[17]_pad  & ~\wb_dat_i[18]_pad  ;
  assign n32828 = n32826 & n32827 ;
  assign n32829 = ~\wb_dat_i[11]_pad  & ~\wb_dat_i[12]_pad  ;
  assign n32830 = ~\wb_dat_i[13]_pad  & ~\wb_dat_i[14]_pad  ;
  assign n32831 = n32829 & n32830 ;
  assign n32832 = n32828 & n32831 ;
  assign n32833 = ~\wb_dat_i[23]_pad  & ~\wb_dat_i[24]_pad  ;
  assign n32834 = ~\wb_dat_i[25]_pad  & ~\wb_dat_i[26]_pad  ;
  assign n32835 = n32833 & n32834 ;
  assign n32836 = ~\wb_dat_i[19]_pad  & ~\wb_dat_i[20]_pad  ;
  assign n32837 = ~\wb_dat_i[21]_pad  & ~\wb_dat_i[22]_pad  ;
  assign n32838 = n32836 & n32837 ;
  assign n32839 = n32835 & n32838 ;
  assign n32840 = n32832 & n32839 ;
  assign n32841 = n32825 & n32840 ;
  assign n32842 = ~\wb_dat_i[4]_pad  & ~\wb_dat_i[5]_pad  ;
  assign n32843 = ~\wb_dat_i[6]_pad  & n32842 ;
  assign n32844 = ~\wb_dat_i[0]_pad  & ~\wb_dat_i[1]_pad  ;
  assign n32845 = ~\wb_dat_i[2]_pad  & ~\wb_dat_i[3]_pad  ;
  assign n32846 = n32844 & n32845 ;
  assign n32847 = n32843 & n32846 ;
  assign n32848 = \wb_dat_i[7]_pad  & ~n32847 ;
  assign n32849 = ~\wb_adr_i[8]_pad  & n23731 ;
  assign n32850 = ~\wb_dat_i[31]_pad  & ~\wb_dat_i[8]_pad  ;
  assign n32851 = ~\wb_dat_i[9]_pad  & n32850 ;
  assign n32852 = ~\wb_dat_i[27]_pad  & ~\wb_dat_i[28]_pad  ;
  assign n32853 = ~\wb_dat_i[29]_pad  & ~\wb_dat_i[30]_pad  ;
  assign n32854 = n32852 & n32853 ;
  assign n32855 = n32851 & n32854 ;
  assign n32856 = n32849 & n32855 ;
  assign n32857 = ~n32848 & n32856 ;
  assign n32858 = n32841 & n32857 ;
  assign n32859 = n32820 & n32858 ;
  assign n32860 = ~\rxethmac1_crcrx_Crc_reg[17]/NET0131  & ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n32861 = ~n10582 & n32860 ;
  assign n32862 = ~\rxethmac1_crcrx_Crc_reg[2]/NET0131  & ~n11372 ;
  assign n32863 = n11353 & n32862 ;
  assign n32864 = ~\rxethmac1_crcrx_Crc_reg[2]/NET0131  & n10663 ;
  assign n32865 = n11353 & n11376 ;
  assign n32866 = ~n32864 & ~n32865 ;
  assign n32867 = ~n32863 & ~n32866 ;
  assign n32868 = \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n32869 = \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131  & \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131  ;
  assign n32870 = n12269 & n32869 ;
  assign n32871 = n13217 & n32870 ;
  assign n32872 = \maccontrol1_receivecontrol1_AddressOK_reg/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n32873 = n32871 & n32872 ;
  assign n32874 = ~n32868 & ~n32873 ;
  assign n32875 = ~\txethmac1_txcrc_Crc_reg[0]/NET0131  & n12974 ;
  assign n32876 = n12961 & n32875 ;
  assign n32877 = ~\txethmac1_txcrc_Crc_reg[0]/NET0131  & n11464 ;
  assign n32878 = ~n12979 & ~n32877 ;
  assign n32879 = ~n32876 & ~n32878 ;
  assign n32880 = n12266 & n12347 ;
  assign n32881 = n32309 & n32880 ;
  assign n32882 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32883 = ~n32881 & n32882 ;
  assign n32884 = \rxethmac1_RxData_reg[0]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32885 = n32881 & n32884 ;
  assign n32886 = ~n32883 & ~n32885 ;
  assign n32887 = n12266 & n12269 ;
  assign n32888 = n32309 & n32887 ;
  assign n32889 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32890 = ~n32888 & n32889 ;
  assign n32891 = \rxethmac1_RxData_reg[2]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32892 = n32888 & n32891 ;
  assign n32893 = ~n32890 & ~n32892 ;
  assign n32894 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32895 = ~n32888 & n32894 ;
  assign n32896 = \rxethmac1_RxData_reg[3]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32897 = n32888 & n32896 ;
  assign n32898 = ~n32895 & ~n32897 ;
  assign n32899 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32900 = ~n32888 & n32899 ;
  assign n32901 = \rxethmac1_RxData_reg[4]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32902 = n32888 & n32901 ;
  assign n32903 = ~n32900 & ~n32902 ;
  assign n32904 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32905 = ~n32888 & n32904 ;
  assign n32906 = \rxethmac1_RxData_reg[5]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32907 = n32888 & n32906 ;
  assign n32908 = ~n32905 & ~n32907 ;
  assign n32909 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32910 = ~n32888 & n32909 ;
  assign n32911 = \rxethmac1_RxData_reg[6]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32912 = n32888 & n32911 ;
  assign n32913 = ~n32910 & ~n32912 ;
  assign n32914 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32915 = ~n32888 & n32914 ;
  assign n32916 = \rxethmac1_RxData_reg[7]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32917 = n32888 & n32916 ;
  assign n32918 = ~n32915 & ~n32917 ;
  assign n32919 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32920 = ~n32881 & n32919 ;
  assign n32921 = \rxethmac1_RxData_reg[1]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32922 = n32881 & n32921 ;
  assign n32923 = ~n32920 & ~n32922 ;
  assign n32924 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32925 = ~n32881 & n32924 ;
  assign n32926 = n32881 & n32891 ;
  assign n32927 = ~n32925 & ~n32926 ;
  assign n32928 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32929 = ~n32881 & n32928 ;
  assign n32930 = n32881 & n32896 ;
  assign n32931 = ~n32929 & ~n32930 ;
  assign n32932 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32933 = ~n32881 & n32932 ;
  assign n32934 = n32881 & n32901 ;
  assign n32935 = ~n32933 & ~n32934 ;
  assign n32936 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32937 = ~n32881 & n32936 ;
  assign n32938 = n32881 & n32906 ;
  assign n32939 = ~n32937 & ~n32938 ;
  assign n32940 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32941 = ~n32881 & n32940 ;
  assign n32942 = n32881 & n32911 ;
  assign n32943 = ~n32941 & ~n32942 ;
  assign n32944 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32945 = ~n32881 & n32944 ;
  assign n32946 = n32881 & n32916 ;
  assign n32947 = ~n32945 & ~n32946 ;
  assign n32948 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32949 = ~n32888 & n32948 ;
  assign n32950 = n32884 & n32888 ;
  assign n32951 = ~n32949 & ~n32950 ;
  assign n32952 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131  & ~\rxethmac1_RxStartFrm_reg/NET0131  ;
  assign n32953 = ~n32888 & n32952 ;
  assign n32954 = n32888 & n32921 ;
  assign n32955 = ~n32953 & ~n32954 ;
  assign n32956 = \m_wb_sel_o[1]_pad  & ~n32431 ;
  assign n32957 = n13189 & n13196 ;
  assign n32958 = \wishbone_RxPointerLSB_rst_reg[0]/NET0131  & \wishbone_RxPointerLSB_rst_reg[1]/NET0131  ;
  assign n32959 = n13189 & n32958 ;
  assign n32960 = ~n32957 & ~n32959 ;
  assign n32961 = ~n32956 & ~n32960 ;
  assign n32962 = ~\wishbone_RxPointerLSB_rst_reg[1]/NET0131  & ~n13196 ;
  assign n32963 = n13189 & ~n32962 ;
  assign n32964 = \m_wb_sel_o[2]_pad  & ~n32431 ;
  assign n32965 = n32963 & ~n32964 ;
  assign n32966 = \m_wb_sel_o[3]_pad  & ~n32431 ;
  assign n32967 = ~\wishbone_RxPointerLSB_rst_reg[0]/NET0131  & ~\wishbone_RxPointerLSB_rst_reg[1]/NET0131  ;
  assign n32968 = ~n13196 & n32967 ;
  assign n32969 = n13189 & ~n32968 ;
  assign n32970 = ~n32966 & n32969 ;
  assign n32971 = ~n32417 & ~n32419 ;
  assign n32972 = ~n32429 & n32971 ;
  assign n32973 = \wishbone_MasterWbRX_reg/NET0131  & ~n32972 ;
  assign n32974 = n13196 & ~n32973 ;
  assign n32975 = \wishbone_MasterWbTX_reg/NET0131  & ~n32972 ;
  assign n32976 = n13189 & ~n32975 ;
  assign n32977 = ~\macstatus1_RxColWindow_reg/NET0131  & ~\rxethmac1_rxstatem1_StateIdle_reg/NET0131  ;
  assign n32978 = ~\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  & ~n11760 ;
  assign n32979 = \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  & n11760 ;
  assign n32980 = ~n32978 & ~n32979 ;
  assign n32981 = ~\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  & ~n11754 ;
  assign n32982 = \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  & n11754 ;
  assign n32983 = ~n32981 & ~n32982 ;
  assign n32984 = ~\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n32985 = \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n32986 = ~n32984 & ~n32985 ;
  assign n32987 = ~\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n32988 = \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n32989 = ~mcoll_pad_i_pad & \rxethmac1_rxstatem1_StateData1_reg/NET0131  ;
  assign n32990 = ~n32988 & n32989 ;
  assign n32991 = ~n32987 & n32990 ;
  assign n32992 = ~n32986 & n32991 ;
  assign n32993 = ~n32983 & n32992 ;
  assign n32994 = ~n32980 & n32993 ;
  assign n32995 = ~\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n32996 = ~n11665 & n32995 ;
  assign n32997 = ~\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n32998 = n11665 & n32997 ;
  assign n32999 = ~n32996 & ~n32998 ;
  assign n33000 = \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n33001 = ~n11665 & n33000 ;
  assign n33002 = \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n33003 = n11665 & n33002 ;
  assign n33004 = ~n33001 & ~n33003 ;
  assign n33005 = n32999 & n33004 ;
  assign n33006 = \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n33007 = ~n11758 & n33006 ;
  assign n33008 = \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n33009 = n11758 & n33008 ;
  assign n33010 = ~n33007 & ~n33009 ;
  assign n33011 = ~\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  & ~n11665 ;
  assign n33012 = ~n11766 & n33011 ;
  assign n33013 = n33010 & ~n33012 ;
  assign n33014 = ~n33005 & n33013 ;
  assign n33015 = n32994 & n33014 ;
  assign n33016 = ~n32977 & ~n33015 ;
  assign n33017 = \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  & \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  ;
  assign n33018 = n10579 & ~n33017 ;
  assign n33019 = n10512 & n33018 ;
  assign n33020 = n10525 & n33019 ;
  assign n33021 = \rxethmac1_rxstatem1_StateData0_reg/NET0131  & ~n33020 ;
  assign n33022 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[0]/NET0131  ;
  assign n33023 = ~n33021 & n33022 ;
  assign n33024 = \rxethmac1_LatchedByte_reg[0]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n33025 = ~n33020 & n33024 ;
  assign n33026 = ~n33023 & ~n33025 ;
  assign n33027 = \txethmac1_StopExcessiveDeferOccured_reg/NET0131  & ~n11186 ;
  assign n33028 = n11182 & n11199 ;
  assign n33029 = ~n33027 & ~n33028 ;
  assign n33030 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33031 = n32311 & n33030 ;
  assign n33032 = \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  & n32311 ;
  assign n33033 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33034 = ~n33032 & n33033 ;
  assign n33035 = ~n33031 & ~n33034 ;
  assign n33036 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33037 = n32311 & n33036 ;
  assign n33038 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33039 = ~n33032 & n33038 ;
  assign n33040 = ~n33037 & ~n33039 ;
  assign n33041 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33042 = n32311 & n33041 ;
  assign n33043 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33044 = ~n33032 & n33043 ;
  assign n33045 = ~n33042 & ~n33044 ;
  assign n33046 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33047 = n32311 & n33046 ;
  assign n33048 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33049 = ~n33032 & n33048 ;
  assign n33050 = ~n33047 & ~n33049 ;
  assign n33051 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33052 = n32311 & n33051 ;
  assign n33053 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33054 = ~n33032 & n33053 ;
  assign n33055 = ~n33052 & ~n33054 ;
  assign n33056 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33057 = n32311 & n33056 ;
  assign n33058 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33059 = ~n33032 & n33058 ;
  assign n33060 = ~n33057 & ~n33059 ;
  assign n33061 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33062 = n32311 & n33061 ;
  assign n33063 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33064 = ~n33032 & n33063 ;
  assign n33065 = ~n33062 & ~n33064 ;
  assign n33066 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33067 = n32311 & n33066 ;
  assign n33068 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33069 = ~n33032 & n33068 ;
  assign n33070 = ~n33067 & ~n33069 ;
  assign n33071 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33072 = n32311 & n33071 ;
  assign n33073 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33074 = ~n33032 & n33073 ;
  assign n33075 = ~n33072 & ~n33074 ;
  assign n33076 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33077 = n32311 & n33076 ;
  assign n33078 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33079 = ~n33032 & n33078 ;
  assign n33080 = ~n33077 & ~n33079 ;
  assign n33081 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33082 = n32311 & n33081 ;
  assign n33083 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33084 = ~n33032 & n33083 ;
  assign n33085 = ~n33082 & ~n33084 ;
  assign n33086 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33087 = n32311 & n33086 ;
  assign n33088 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33089 = ~n33032 & n33088 ;
  assign n33090 = ~n33087 & ~n33089 ;
  assign n33091 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33092 = n32311 & n33091 ;
  assign n33093 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33094 = ~n33032 & n33093 ;
  assign n33095 = ~n33092 & ~n33094 ;
  assign n33096 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33097 = n32311 & n33096 ;
  assign n33098 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33099 = ~n33032 & n33098 ;
  assign n33100 = ~n33097 & ~n33099 ;
  assign n33101 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33102 = n32311 & n33101 ;
  assign n33103 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33104 = ~n33032 & n33103 ;
  assign n33105 = ~n33102 & ~n33104 ;
  assign n33106 = \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131  & \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
  assign n33107 = n32311 & n33106 ;
  assign n33108 = \maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n33109 = ~n33032 & n33108 ;
  assign n33110 = ~n33107 & ~n33109 ;
  assign n33111 = ~\wishbone_LastByteIn_reg/NET0131  & \wishbone_RxEnableWindow_reg/NET0131  ;
  assign n33112 = n15730 & n33111 ;
  assign n33113 = ~\wishbone_RxValidBytes_reg[0]/NET0131  & ~n15726 ;
  assign n33114 = ~n33112 & n33113 ;
  assign n33115 = \wishbone_RxValidBytes_reg[0]/NET0131  & ~n15726 ;
  assign n33116 = n33112 & n33115 ;
  assign n33117 = ~n33114 & ~n33116 ;
  assign n33118 = \wishbone_RxPointerLSB_rst_reg[0]/NET0131  & n15726 ;
  assign n33119 = n33117 & ~n33118 ;
  assign n33120 = \wishbone_RxValidBytes_reg[1]/NET0131  & ~n33112 ;
  assign n33121 = n15743 & n33112 ;
  assign n33122 = ~n33120 & ~n33121 ;
  assign n33123 = ~n15726 & ~n33122 ;
  assign n33124 = n15726 & ~n32305 ;
  assign n33125 = ~n33123 & ~n33124 ;
  assign n33126 = \miim1_shftrg_ShiftReg_reg[0]/NET0131  & ~n32513 ;
  assign n33127 = ~n32513 & ~n33126 ;
  assign n33128 = \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131  & ~n32531 ;
  assign n33129 = \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n33130 = n32538 & n33129 ;
  assign n33131 = \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n33132 = n32538 & n33131 ;
  assign n33133 = ~n33130 & ~n33132 ;
  assign n33134 = ~n33128 & n33133 ;
  assign n33135 = md_pad_i_pad & n32545 ;
  assign n33136 = n32531 & n33135 ;
  assign n33137 = ~n33126 & ~n33136 ;
  assign n33138 = n33134 & n33137 ;
  assign n33139 = ~n33127 & ~n33138 ;
  assign n33140 = \miim1_shftrg_ShiftReg_reg[6]/NET0131  & n32545 ;
  assign n33141 = n32531 & n33140 ;
  assign n33142 = \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n33143 = n32538 & n33142 ;
  assign n33144 = \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n33145 = n32538 & n33144 ;
  assign n33146 = \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131  & n32535 ;
  assign n33147 = ~n33145 & ~n33146 ;
  assign n33148 = ~n33143 & n33147 ;
  assign n33149 = ~n33141 & n33148 ;
  assign n33150 = n32513 & ~n33149 ;
  assign n33151 = \miim1_shftrg_ShiftReg_reg[7]/NET0131  & ~n32513 ;
  assign n33152 = ~n33150 & ~n33151 ;
  assign n33153 = ~\wishbone_tx_burst_cnt_reg[0]/NET0131  & n13174 ;
  assign n33154 = \wishbone_tx_burst_cnt_reg[0]/NET0131  & ~n13174 ;
  assign n33155 = n32466 & n33154 ;
  assign n33156 = ~n33153 & ~n33155 ;
  assign n33157 = \wishbone_tx_burst_cnt_reg[2]/NET0131  & ~n32461 ;
  assign n33158 = ~n32462 & ~n33157 ;
  assign n33159 = ~n13166 & ~n33158 ;
  assign n33160 = ~n13164 & n33159 ;
  assign n33161 = \wishbone_tx_burst_cnt_reg[2]/NET0131  & ~n13174 ;
  assign n33162 = n32466 & n33161 ;
  assign n33163 = ~n33160 & ~n33162 ;
  assign n33164 = ~\wishbone_SyncRxStartFrm_q2_reg/NET0131  & \wishbone_SyncRxStartFrm_q_reg/NET0131  ;
  assign n33165 = ~\wishbone_rx_fifo_read_pointer_reg[0]/NET0131  & ~\wishbone_rx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n33166 = ~\wishbone_rx_fifo_read_pointer_reg[2]/NET0131  & ~\wishbone_rx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n33167 = n33165 & n33166 ;
  assign n33168 = ~n33164 & ~n33167 ;
  assign n33169 = \wishbone_rx_fifo_fifo_reg[0][0]/P0001  & ~n33168 ;
  assign n33170 = \wishbone_rx_fifo_read_pointer_reg[0]/NET0131  & \wishbone_rx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n33171 = \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  & \wishbone_rx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n33172 = n33170 & n33171 ;
  assign n33173 = \wishbone_rx_fifo_fifo_reg[15][0]/P0001  & n33172 ;
  assign n33174 = ~\wishbone_rx_fifo_read_pointer_reg[2]/NET0131  & \wishbone_rx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n33175 = \wishbone_rx_fifo_read_pointer_reg[0]/NET0131  & ~\wishbone_rx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n33176 = n33174 & n33175 ;
  assign n33177 = \wishbone_rx_fifo_fifo_reg[9][0]/P0001  & n33176 ;
  assign n33178 = ~n33173 & ~n33177 ;
  assign n33179 = n33165 & n33174 ;
  assign n33180 = \wishbone_rx_fifo_fifo_reg[8][0]/P0001  & n33179 ;
  assign n33181 = n33166 & n33175 ;
  assign n33182 = \wishbone_rx_fifo_fifo_reg[1][0]/P0001  & n33181 ;
  assign n33183 = ~n33180 & ~n33182 ;
  assign n33184 = n33178 & n33183 ;
  assign n33185 = ~\wishbone_rx_fifo_read_pointer_reg[0]/NET0131  & \wishbone_rx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n33186 = \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  & ~\wishbone_rx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n33187 = n33185 & n33186 ;
  assign n33188 = \wishbone_rx_fifo_fifo_reg[6][0]/P0001  & n33187 ;
  assign n33189 = n33174 & n33185 ;
  assign n33190 = \wishbone_rx_fifo_fifo_reg[10][0]/P0001  & n33189 ;
  assign n33191 = ~n33188 & ~n33190 ;
  assign n33192 = n33170 & n33186 ;
  assign n33193 = \wishbone_rx_fifo_fifo_reg[7][0]/P0001  & n33192 ;
  assign n33194 = n33165 & n33186 ;
  assign n33195 = \wishbone_rx_fifo_fifo_reg[4][0]/P0001  & n33194 ;
  assign n33196 = ~n33193 & ~n33195 ;
  assign n33197 = n33191 & n33196 ;
  assign n33198 = n33184 & n33197 ;
  assign n33199 = n33166 & n33170 ;
  assign n33200 = \wishbone_rx_fifo_fifo_reg[3][0]/P0001  & n33199 ;
  assign n33201 = n33171 & n33175 ;
  assign n33202 = \wishbone_rx_fifo_fifo_reg[13][0]/P0001  & n33201 ;
  assign n33203 = n33170 & n33174 ;
  assign n33204 = \wishbone_rx_fifo_fifo_reg[11][0]/P0001  & n33203 ;
  assign n33205 = ~n33202 & ~n33204 ;
  assign n33206 = ~n33200 & n33205 ;
  assign n33207 = n33166 & n33185 ;
  assign n33208 = \wishbone_rx_fifo_fifo_reg[2][0]/P0001  & n33207 ;
  assign n33209 = n33175 & n33186 ;
  assign n33210 = \wishbone_rx_fifo_fifo_reg[5][0]/P0001  & n33209 ;
  assign n33211 = ~n33208 & ~n33210 ;
  assign n33212 = n33171 & n33185 ;
  assign n33213 = \wishbone_rx_fifo_fifo_reg[14][0]/P0001  & n33212 ;
  assign n33214 = n33165 & n33171 ;
  assign n33215 = \wishbone_rx_fifo_fifo_reg[12][0]/P0001  & n33214 ;
  assign n33216 = ~n33213 & ~n33215 ;
  assign n33217 = n33211 & n33216 ;
  assign n33218 = n33206 & n33217 ;
  assign n33219 = n33198 & n33218 ;
  assign n33220 = ~n33164 & ~n33219 ;
  assign n33221 = ~n33169 & ~n33220 ;
  assign n33222 = \wishbone_rx_fifo_fifo_reg[11][10]/P0001  & n33203 ;
  assign n33223 = \wishbone_rx_fifo_fifo_reg[3][10]/P0001  & n33199 ;
  assign n33224 = ~n33222 & ~n33223 ;
  assign n33225 = \wishbone_rx_fifo_fifo_reg[6][10]/P0001  & n33187 ;
  assign n33226 = \wishbone_rx_fifo_fifo_reg[15][10]/P0001  & n33172 ;
  assign n33227 = ~n33225 & ~n33226 ;
  assign n33228 = n33224 & n33227 ;
  assign n33229 = \wishbone_rx_fifo_fifo_reg[5][10]/P0001  & n33209 ;
  assign n33230 = ~n33164 & ~n33229 ;
  assign n33231 = \wishbone_rx_fifo_fifo_reg[7][10]/P0001  & n33192 ;
  assign n33232 = \wishbone_rx_fifo_fifo_reg[1][10]/P0001  & n33181 ;
  assign n33233 = ~n33231 & ~n33232 ;
  assign n33234 = n33230 & n33233 ;
  assign n33235 = n33228 & n33234 ;
  assign n33236 = \wishbone_rx_fifo_fifo_reg[12][10]/P0001  & n33214 ;
  assign n33237 = \wishbone_rx_fifo_fifo_reg[10][10]/P0001  & n33189 ;
  assign n33238 = ~n33236 & ~n33237 ;
  assign n33239 = \wishbone_rx_fifo_fifo_reg[9][10]/P0001  & n33176 ;
  assign n33240 = \wishbone_rx_fifo_fifo_reg[13][10]/P0001  & n33201 ;
  assign n33241 = ~n33239 & ~n33240 ;
  assign n33242 = n33238 & n33241 ;
  assign n33243 = \wishbone_rx_fifo_fifo_reg[14][10]/P0001  & n33212 ;
  assign n33244 = \wishbone_rx_fifo_fifo_reg[2][10]/P0001  & n33207 ;
  assign n33245 = ~n33243 & ~n33244 ;
  assign n33246 = \wishbone_rx_fifo_fifo_reg[8][10]/P0001  & n33179 ;
  assign n33247 = \wishbone_rx_fifo_fifo_reg[4][10]/P0001  & n33194 ;
  assign n33248 = ~n33246 & ~n33247 ;
  assign n33249 = n33245 & n33248 ;
  assign n33250 = n33242 & n33249 ;
  assign n33251 = n33235 & n33250 ;
  assign n33252 = ~\wishbone_rx_fifo_fifo_reg[0][10]/P0001  & n33164 ;
  assign n33253 = ~n33251 & ~n33252 ;
  assign n33254 = \wishbone_rx_fifo_fifo_reg[0][10]/P0001  & n33167 ;
  assign n33255 = ~n33253 & ~n33254 ;
  assign n33256 = \wishbone_rx_fifo_fifo_reg[0][11]/P0001  & ~n33168 ;
  assign n33257 = \wishbone_rx_fifo_fifo_reg[5][11]/P0001  & n33209 ;
  assign n33258 = \wishbone_rx_fifo_fifo_reg[9][11]/P0001  & n33176 ;
  assign n33259 = ~n33257 & ~n33258 ;
  assign n33260 = \wishbone_rx_fifo_fifo_reg[10][11]/P0001  & n33189 ;
  assign n33261 = \wishbone_rx_fifo_fifo_reg[13][11]/P0001  & n33201 ;
  assign n33262 = ~n33260 & ~n33261 ;
  assign n33263 = n33259 & n33262 ;
  assign n33264 = \wishbone_rx_fifo_fifo_reg[6][11]/P0001  & n33187 ;
  assign n33265 = \wishbone_rx_fifo_fifo_reg[12][11]/P0001  & n33214 ;
  assign n33266 = ~n33264 & ~n33265 ;
  assign n33267 = \wishbone_rx_fifo_fifo_reg[8][11]/P0001  & n33179 ;
  assign n33268 = \wishbone_rx_fifo_fifo_reg[11][11]/P0001  & n33203 ;
  assign n33269 = ~n33267 & ~n33268 ;
  assign n33270 = n33266 & n33269 ;
  assign n33271 = n33263 & n33270 ;
  assign n33272 = \wishbone_rx_fifo_fifo_reg[2][11]/P0001  & n33207 ;
  assign n33273 = \wishbone_rx_fifo_fifo_reg[7][11]/P0001  & n33192 ;
  assign n33274 = \wishbone_rx_fifo_fifo_reg[14][11]/P0001  & n33212 ;
  assign n33275 = ~n33273 & ~n33274 ;
  assign n33276 = ~n33272 & n33275 ;
  assign n33277 = \wishbone_rx_fifo_fifo_reg[1][11]/P0001  & n33181 ;
  assign n33278 = \wishbone_rx_fifo_fifo_reg[15][11]/P0001  & n33172 ;
  assign n33279 = ~n33277 & ~n33278 ;
  assign n33280 = \wishbone_rx_fifo_fifo_reg[4][11]/P0001  & n33194 ;
  assign n33281 = \wishbone_rx_fifo_fifo_reg[3][11]/P0001  & n33199 ;
  assign n33282 = ~n33280 & ~n33281 ;
  assign n33283 = n33279 & n33282 ;
  assign n33284 = n33276 & n33283 ;
  assign n33285 = n33271 & n33284 ;
  assign n33286 = ~n33164 & ~n33285 ;
  assign n33287 = ~n33256 & ~n33286 ;
  assign n33288 = \wishbone_rx_fifo_fifo_reg[5][12]/P0001  & n33209 ;
  assign n33289 = \wishbone_rx_fifo_fifo_reg[11][12]/P0001  & n33203 ;
  assign n33290 = ~n33288 & ~n33289 ;
  assign n33291 = \wishbone_rx_fifo_fifo_reg[10][12]/P0001  & n33189 ;
  assign n33292 = \wishbone_rx_fifo_fifo_reg[1][12]/P0001  & n33181 ;
  assign n33293 = ~n33291 & ~n33292 ;
  assign n33294 = n33290 & n33293 ;
  assign n33295 = \wishbone_rx_fifo_fifo_reg[3][12]/P0001  & n33199 ;
  assign n33296 = ~n33164 & ~n33295 ;
  assign n33297 = \wishbone_rx_fifo_fifo_reg[14][12]/P0001  & n33212 ;
  assign n33298 = \wishbone_rx_fifo_fifo_reg[2][12]/P0001  & n33207 ;
  assign n33299 = ~n33297 & ~n33298 ;
  assign n33300 = n33296 & n33299 ;
  assign n33301 = n33294 & n33300 ;
  assign n33302 = \wishbone_rx_fifo_fifo_reg[9][12]/P0001  & n33176 ;
  assign n33303 = \wishbone_rx_fifo_fifo_reg[12][12]/P0001  & n33214 ;
  assign n33304 = ~n33302 & ~n33303 ;
  assign n33305 = \wishbone_rx_fifo_fifo_reg[6][12]/P0001  & n33187 ;
  assign n33306 = \wishbone_rx_fifo_fifo_reg[13][12]/P0001  & n33201 ;
  assign n33307 = ~n33305 & ~n33306 ;
  assign n33308 = n33304 & n33307 ;
  assign n33309 = \wishbone_rx_fifo_fifo_reg[4][12]/P0001  & n33194 ;
  assign n33310 = \wishbone_rx_fifo_fifo_reg[8][12]/P0001  & n33179 ;
  assign n33311 = ~n33309 & ~n33310 ;
  assign n33312 = \wishbone_rx_fifo_fifo_reg[15][12]/P0001  & n33172 ;
  assign n33313 = \wishbone_rx_fifo_fifo_reg[7][12]/P0001  & n33192 ;
  assign n33314 = ~n33312 & ~n33313 ;
  assign n33315 = n33311 & n33314 ;
  assign n33316 = n33308 & n33315 ;
  assign n33317 = n33301 & n33316 ;
  assign n33318 = ~\wishbone_rx_fifo_fifo_reg[0][12]/P0001  & n33164 ;
  assign n33319 = ~n33317 & ~n33318 ;
  assign n33320 = \wishbone_rx_fifo_fifo_reg[0][12]/P0001  & n33167 ;
  assign n33321 = ~n33319 & ~n33320 ;
  assign n33322 = \wishbone_rx_fifo_fifo_reg[0][13]/P0001  & ~n33168 ;
  assign n33323 = \wishbone_rx_fifo_fifo_reg[10][13]/P0001  & n33189 ;
  assign n33324 = \wishbone_rx_fifo_fifo_reg[5][13]/P0001  & n33209 ;
  assign n33325 = ~n33323 & ~n33324 ;
  assign n33326 = \wishbone_rx_fifo_fifo_reg[14][13]/P0001  & n33212 ;
  assign n33327 = \wishbone_rx_fifo_fifo_reg[4][13]/P0001  & n33194 ;
  assign n33328 = ~n33326 & ~n33327 ;
  assign n33329 = n33325 & n33328 ;
  assign n33330 = \wishbone_rx_fifo_fifo_reg[3][13]/P0001  & n33199 ;
  assign n33331 = \wishbone_rx_fifo_fifo_reg[9][13]/P0001  & n33176 ;
  assign n33332 = ~n33330 & ~n33331 ;
  assign n33333 = \wishbone_rx_fifo_fifo_reg[8][13]/P0001  & n33179 ;
  assign n33334 = \wishbone_rx_fifo_fifo_reg[7][13]/P0001  & n33192 ;
  assign n33335 = ~n33333 & ~n33334 ;
  assign n33336 = n33332 & n33335 ;
  assign n33337 = n33329 & n33336 ;
  assign n33338 = \wishbone_rx_fifo_fifo_reg[6][13]/P0001  & n33187 ;
  assign n33339 = \wishbone_rx_fifo_fifo_reg[15][13]/P0001  & n33172 ;
  assign n33340 = \wishbone_rx_fifo_fifo_reg[11][13]/P0001  & n33203 ;
  assign n33341 = ~n33339 & ~n33340 ;
  assign n33342 = ~n33338 & n33341 ;
  assign n33343 = \wishbone_rx_fifo_fifo_reg[1][13]/P0001  & n33181 ;
  assign n33344 = \wishbone_rx_fifo_fifo_reg[13][13]/P0001  & n33201 ;
  assign n33345 = ~n33343 & ~n33344 ;
  assign n33346 = \wishbone_rx_fifo_fifo_reg[2][13]/P0001  & n33207 ;
  assign n33347 = \wishbone_rx_fifo_fifo_reg[12][13]/P0001  & n33214 ;
  assign n33348 = ~n33346 & ~n33347 ;
  assign n33349 = n33345 & n33348 ;
  assign n33350 = n33342 & n33349 ;
  assign n33351 = n33337 & n33350 ;
  assign n33352 = ~n33164 & ~n33351 ;
  assign n33353 = ~n33322 & ~n33352 ;
  assign n33354 = \wishbone_rx_fifo_fifo_reg[11][14]/P0001  & n33203 ;
  assign n33355 = \wishbone_rx_fifo_fifo_reg[3][14]/P0001  & n33199 ;
  assign n33356 = ~n33354 & ~n33355 ;
  assign n33357 = \wishbone_rx_fifo_fifo_reg[6][14]/P0001  & n33187 ;
  assign n33358 = \wishbone_rx_fifo_fifo_reg[8][14]/P0001  & n33179 ;
  assign n33359 = ~n33357 & ~n33358 ;
  assign n33360 = n33356 & n33359 ;
  assign n33361 = \wishbone_rx_fifo_fifo_reg[12][14]/P0001  & n33214 ;
  assign n33362 = ~n33164 & ~n33361 ;
  assign n33363 = \wishbone_rx_fifo_fifo_reg[5][14]/P0001  & n33209 ;
  assign n33364 = \wishbone_rx_fifo_fifo_reg[2][14]/P0001  & n33207 ;
  assign n33365 = ~n33363 & ~n33364 ;
  assign n33366 = n33362 & n33365 ;
  assign n33367 = n33360 & n33366 ;
  assign n33368 = \wishbone_rx_fifo_fifo_reg[1][14]/P0001  & n33181 ;
  assign n33369 = \wishbone_rx_fifo_fifo_reg[10][14]/P0001  & n33189 ;
  assign n33370 = ~n33368 & ~n33369 ;
  assign n33371 = \wishbone_rx_fifo_fifo_reg[9][14]/P0001  & n33176 ;
  assign n33372 = \wishbone_rx_fifo_fifo_reg[4][14]/P0001  & n33194 ;
  assign n33373 = ~n33371 & ~n33372 ;
  assign n33374 = n33370 & n33373 ;
  assign n33375 = \wishbone_rx_fifo_fifo_reg[15][14]/P0001  & n33172 ;
  assign n33376 = \wishbone_rx_fifo_fifo_reg[13][14]/P0001  & n33201 ;
  assign n33377 = ~n33375 & ~n33376 ;
  assign n33378 = \wishbone_rx_fifo_fifo_reg[7][14]/P0001  & n33192 ;
  assign n33379 = \wishbone_rx_fifo_fifo_reg[14][14]/P0001  & n33212 ;
  assign n33380 = ~n33378 & ~n33379 ;
  assign n33381 = n33377 & n33380 ;
  assign n33382 = n33374 & n33381 ;
  assign n33383 = n33367 & n33382 ;
  assign n33384 = ~\wishbone_rx_fifo_fifo_reg[0][14]/P0001  & n33164 ;
  assign n33385 = ~n33383 & ~n33384 ;
  assign n33386 = \wishbone_rx_fifo_fifo_reg[0][14]/P0001  & n33167 ;
  assign n33387 = ~n33385 & ~n33386 ;
  assign n33388 = \wishbone_rx_fifo_fifo_reg[0][15]/P0001  & ~n33168 ;
  assign n33389 = \wishbone_rx_fifo_fifo_reg[14][15]/P0001  & n33212 ;
  assign n33390 = \wishbone_rx_fifo_fifo_reg[6][15]/P0001  & n33187 ;
  assign n33391 = ~n33389 & ~n33390 ;
  assign n33392 = \wishbone_rx_fifo_fifo_reg[1][15]/P0001  & n33181 ;
  assign n33393 = \wishbone_rx_fifo_fifo_reg[10][15]/P0001  & n33189 ;
  assign n33394 = ~n33392 & ~n33393 ;
  assign n33395 = n33391 & n33394 ;
  assign n33396 = \wishbone_rx_fifo_fifo_reg[12][15]/P0001  & n33214 ;
  assign n33397 = \wishbone_rx_fifo_fifo_reg[5][15]/P0001  & n33209 ;
  assign n33398 = ~n33396 & ~n33397 ;
  assign n33399 = \wishbone_rx_fifo_fifo_reg[4][15]/P0001  & n33194 ;
  assign n33400 = \wishbone_rx_fifo_fifo_reg[8][15]/P0001  & n33179 ;
  assign n33401 = ~n33399 & ~n33400 ;
  assign n33402 = n33398 & n33401 ;
  assign n33403 = n33395 & n33402 ;
  assign n33404 = \wishbone_rx_fifo_fifo_reg[11][15]/P0001  & n33203 ;
  assign n33405 = \wishbone_rx_fifo_fifo_reg[15][15]/P0001  & n33172 ;
  assign n33406 = \wishbone_rx_fifo_fifo_reg[3][15]/P0001  & n33199 ;
  assign n33407 = ~n33405 & ~n33406 ;
  assign n33408 = ~n33404 & n33407 ;
  assign n33409 = \wishbone_rx_fifo_fifo_reg[7][15]/P0001  & n33192 ;
  assign n33410 = \wishbone_rx_fifo_fifo_reg[2][15]/P0001  & n33207 ;
  assign n33411 = ~n33409 & ~n33410 ;
  assign n33412 = \wishbone_rx_fifo_fifo_reg[13][15]/P0001  & n33201 ;
  assign n33413 = \wishbone_rx_fifo_fifo_reg[9][15]/P0001  & n33176 ;
  assign n33414 = ~n33412 & ~n33413 ;
  assign n33415 = n33411 & n33414 ;
  assign n33416 = n33408 & n33415 ;
  assign n33417 = n33403 & n33416 ;
  assign n33418 = ~n33164 & ~n33417 ;
  assign n33419 = ~n33388 & ~n33418 ;
  assign n33420 = \wishbone_rx_fifo_fifo_reg[11][16]/P0001  & n33203 ;
  assign n33421 = \wishbone_rx_fifo_fifo_reg[9][16]/P0001  & n33176 ;
  assign n33422 = ~n33420 & ~n33421 ;
  assign n33423 = \wishbone_rx_fifo_fifo_reg[6][16]/P0001  & n33187 ;
  assign n33424 = \wishbone_rx_fifo_fifo_reg[15][16]/P0001  & n33172 ;
  assign n33425 = ~n33423 & ~n33424 ;
  assign n33426 = n33422 & n33425 ;
  assign n33427 = \wishbone_rx_fifo_fifo_reg[12][16]/P0001  & n33214 ;
  assign n33428 = ~n33164 & ~n33427 ;
  assign n33429 = \wishbone_rx_fifo_fifo_reg[3][16]/P0001  & n33199 ;
  assign n33430 = \wishbone_rx_fifo_fifo_reg[1][16]/P0001  & n33181 ;
  assign n33431 = ~n33429 & ~n33430 ;
  assign n33432 = n33428 & n33431 ;
  assign n33433 = n33426 & n33432 ;
  assign n33434 = \wishbone_rx_fifo_fifo_reg[5][16]/P0001  & n33209 ;
  assign n33435 = \wishbone_rx_fifo_fifo_reg[10][16]/P0001  & n33189 ;
  assign n33436 = ~n33434 & ~n33435 ;
  assign n33437 = \wishbone_rx_fifo_fifo_reg[2][16]/P0001  & n33207 ;
  assign n33438 = \wishbone_rx_fifo_fifo_reg[4][16]/P0001  & n33194 ;
  assign n33439 = ~n33437 & ~n33438 ;
  assign n33440 = n33436 & n33439 ;
  assign n33441 = \wishbone_rx_fifo_fifo_reg[7][16]/P0001  & n33192 ;
  assign n33442 = \wishbone_rx_fifo_fifo_reg[8][16]/P0001  & n33179 ;
  assign n33443 = ~n33441 & ~n33442 ;
  assign n33444 = \wishbone_rx_fifo_fifo_reg[13][16]/P0001  & n33201 ;
  assign n33445 = \wishbone_rx_fifo_fifo_reg[14][16]/P0001  & n33212 ;
  assign n33446 = ~n33444 & ~n33445 ;
  assign n33447 = n33443 & n33446 ;
  assign n33448 = n33440 & n33447 ;
  assign n33449 = n33433 & n33448 ;
  assign n33450 = ~\wishbone_rx_fifo_fifo_reg[0][16]/P0001  & n33164 ;
  assign n33451 = ~n33449 & ~n33450 ;
  assign n33452 = \wishbone_rx_fifo_fifo_reg[0][16]/P0001  & n33167 ;
  assign n33453 = ~n33451 & ~n33452 ;
  assign n33454 = \wishbone_rx_fifo_fifo_reg[0][17]/P0001  & ~n33168 ;
  assign n33455 = \wishbone_rx_fifo_fifo_reg[14][17]/P0001  & n33212 ;
  assign n33456 = \wishbone_rx_fifo_fifo_reg[9][17]/P0001  & n33176 ;
  assign n33457 = ~n33455 & ~n33456 ;
  assign n33458 = \wishbone_rx_fifo_fifo_reg[1][17]/P0001  & n33181 ;
  assign n33459 = \wishbone_rx_fifo_fifo_reg[10][17]/P0001  & n33189 ;
  assign n33460 = ~n33458 & ~n33459 ;
  assign n33461 = n33457 & n33460 ;
  assign n33462 = \wishbone_rx_fifo_fifo_reg[12][17]/P0001  & n33214 ;
  assign n33463 = \wishbone_rx_fifo_fifo_reg[5][17]/P0001  & n33209 ;
  assign n33464 = ~n33462 & ~n33463 ;
  assign n33465 = \wishbone_rx_fifo_fifo_reg[4][17]/P0001  & n33194 ;
  assign n33466 = \wishbone_rx_fifo_fifo_reg[8][17]/P0001  & n33179 ;
  assign n33467 = ~n33465 & ~n33466 ;
  assign n33468 = n33464 & n33467 ;
  assign n33469 = n33461 & n33468 ;
  assign n33470 = \wishbone_rx_fifo_fifo_reg[11][17]/P0001  & n33203 ;
  assign n33471 = \wishbone_rx_fifo_fifo_reg[15][17]/P0001  & n33172 ;
  assign n33472 = \wishbone_rx_fifo_fifo_reg[3][17]/P0001  & n33199 ;
  assign n33473 = ~n33471 & ~n33472 ;
  assign n33474 = ~n33470 & n33473 ;
  assign n33475 = \wishbone_rx_fifo_fifo_reg[7][17]/P0001  & n33192 ;
  assign n33476 = \wishbone_rx_fifo_fifo_reg[2][17]/P0001  & n33207 ;
  assign n33477 = ~n33475 & ~n33476 ;
  assign n33478 = \wishbone_rx_fifo_fifo_reg[13][17]/P0001  & n33201 ;
  assign n33479 = \wishbone_rx_fifo_fifo_reg[6][17]/P0001  & n33187 ;
  assign n33480 = ~n33478 & ~n33479 ;
  assign n33481 = n33477 & n33480 ;
  assign n33482 = n33474 & n33481 ;
  assign n33483 = n33469 & n33482 ;
  assign n33484 = ~n33164 & ~n33483 ;
  assign n33485 = ~n33454 & ~n33484 ;
  assign n33486 = \wishbone_rx_fifo_fifo_reg[0][18]/P0001  & ~n33168 ;
  assign n33487 = \wishbone_rx_fifo_fifo_reg[10][18]/P0001  & n33189 ;
  assign n33488 = \wishbone_rx_fifo_fifo_reg[6][18]/P0001  & n33187 ;
  assign n33489 = ~n33487 & ~n33488 ;
  assign n33490 = \wishbone_rx_fifo_fifo_reg[12][18]/P0001  & n33214 ;
  assign n33491 = \wishbone_rx_fifo_fifo_reg[4][18]/P0001  & n33194 ;
  assign n33492 = ~n33490 & ~n33491 ;
  assign n33493 = n33489 & n33492 ;
  assign n33494 = \wishbone_rx_fifo_fifo_reg[3][18]/P0001  & n33199 ;
  assign n33495 = \wishbone_rx_fifo_fifo_reg[9][18]/P0001  & n33176 ;
  assign n33496 = ~n33494 & ~n33495 ;
  assign n33497 = \wishbone_rx_fifo_fifo_reg[5][18]/P0001  & n33209 ;
  assign n33498 = \wishbone_rx_fifo_fifo_reg[7][18]/P0001  & n33192 ;
  assign n33499 = ~n33497 & ~n33498 ;
  assign n33500 = n33496 & n33499 ;
  assign n33501 = n33493 & n33500 ;
  assign n33502 = \wishbone_rx_fifo_fifo_reg[15][18]/P0001  & n33172 ;
  assign n33503 = \wishbone_rx_fifo_fifo_reg[8][18]/P0001  & n33179 ;
  assign n33504 = \wishbone_rx_fifo_fifo_reg[11][18]/P0001  & n33203 ;
  assign n33505 = ~n33503 & ~n33504 ;
  assign n33506 = ~n33502 & n33505 ;
  assign n33507 = \wishbone_rx_fifo_fifo_reg[1][18]/P0001  & n33181 ;
  assign n33508 = \wishbone_rx_fifo_fifo_reg[13][18]/P0001  & n33201 ;
  assign n33509 = ~n33507 & ~n33508 ;
  assign n33510 = \wishbone_rx_fifo_fifo_reg[2][18]/P0001  & n33207 ;
  assign n33511 = \wishbone_rx_fifo_fifo_reg[14][18]/P0001  & n33212 ;
  assign n33512 = ~n33510 & ~n33511 ;
  assign n33513 = n33509 & n33512 ;
  assign n33514 = n33506 & n33513 ;
  assign n33515 = n33501 & n33514 ;
  assign n33516 = ~n33164 & ~n33515 ;
  assign n33517 = ~n33486 & ~n33516 ;
  assign n33518 = \wishbone_rx_fifo_fifo_reg[0][19]/P0001  & ~n33168 ;
  assign n33519 = \wishbone_rx_fifo_fifo_reg[2][19]/P0001  & n33207 ;
  assign n33520 = \wishbone_rx_fifo_fifo_reg[3][19]/P0001  & n33199 ;
  assign n33521 = ~n33519 & ~n33520 ;
  assign n33522 = \wishbone_rx_fifo_fifo_reg[4][19]/P0001  & n33194 ;
  assign n33523 = \wishbone_rx_fifo_fifo_reg[5][19]/P0001  & n33209 ;
  assign n33524 = ~n33522 & ~n33523 ;
  assign n33525 = n33521 & n33524 ;
  assign n33526 = \wishbone_rx_fifo_fifo_reg[9][19]/P0001  & n33176 ;
  assign n33527 = \wishbone_rx_fifo_fifo_reg[8][19]/P0001  & n33179 ;
  assign n33528 = ~n33526 & ~n33527 ;
  assign n33529 = \wishbone_rx_fifo_fifo_reg[12][19]/P0001  & n33214 ;
  assign n33530 = \wishbone_rx_fifo_fifo_reg[13][19]/P0001  & n33201 ;
  assign n33531 = ~n33529 & ~n33530 ;
  assign n33532 = n33528 & n33531 ;
  assign n33533 = n33525 & n33532 ;
  assign n33534 = \wishbone_rx_fifo_fifo_reg[14][19]/P0001  & n33212 ;
  assign n33535 = \wishbone_rx_fifo_fifo_reg[6][19]/P0001  & n33187 ;
  assign n33536 = \wishbone_rx_fifo_fifo_reg[15][19]/P0001  & n33172 ;
  assign n33537 = ~n33535 & ~n33536 ;
  assign n33538 = ~n33534 & n33537 ;
  assign n33539 = \wishbone_rx_fifo_fifo_reg[10][19]/P0001  & n33189 ;
  assign n33540 = \wishbone_rx_fifo_fifo_reg[7][19]/P0001  & n33192 ;
  assign n33541 = ~n33539 & ~n33540 ;
  assign n33542 = \wishbone_rx_fifo_fifo_reg[1][19]/P0001  & n33181 ;
  assign n33543 = \wishbone_rx_fifo_fifo_reg[11][19]/P0001  & n33203 ;
  assign n33544 = ~n33542 & ~n33543 ;
  assign n33545 = n33541 & n33544 ;
  assign n33546 = n33538 & n33545 ;
  assign n33547 = n33533 & n33546 ;
  assign n33548 = ~n33164 & ~n33547 ;
  assign n33549 = ~n33518 & ~n33548 ;
  assign n33550 = \wishbone_rx_fifo_fifo_reg[11][1]/P0001  & n33203 ;
  assign n33551 = \wishbone_rx_fifo_fifo_reg[9][1]/P0001  & n33176 ;
  assign n33552 = ~n33550 & ~n33551 ;
  assign n33553 = \wishbone_rx_fifo_fifo_reg[6][1]/P0001  & n33187 ;
  assign n33554 = \wishbone_rx_fifo_fifo_reg[15][1]/P0001  & n33172 ;
  assign n33555 = ~n33553 & ~n33554 ;
  assign n33556 = n33552 & n33555 ;
  assign n33557 = \wishbone_rx_fifo_fifo_reg[5][1]/P0001  & n33209 ;
  assign n33558 = ~n33164 & ~n33557 ;
  assign n33559 = \wishbone_rx_fifo_fifo_reg[3][1]/P0001  & n33199 ;
  assign n33560 = \wishbone_rx_fifo_fifo_reg[1][1]/P0001  & n33181 ;
  assign n33561 = ~n33559 & ~n33560 ;
  assign n33562 = n33558 & n33561 ;
  assign n33563 = n33556 & n33562 ;
  assign n33564 = \wishbone_rx_fifo_fifo_reg[14][1]/P0001  & n33212 ;
  assign n33565 = \wishbone_rx_fifo_fifo_reg[10][1]/P0001  & n33189 ;
  assign n33566 = ~n33564 & ~n33565 ;
  assign n33567 = \wishbone_rx_fifo_fifo_reg[2][1]/P0001  & n33207 ;
  assign n33568 = \wishbone_rx_fifo_fifo_reg[4][1]/P0001  & n33194 ;
  assign n33569 = ~n33567 & ~n33568 ;
  assign n33570 = n33566 & n33569 ;
  assign n33571 = \wishbone_rx_fifo_fifo_reg[7][1]/P0001  & n33192 ;
  assign n33572 = \wishbone_rx_fifo_fifo_reg[8][1]/P0001  & n33179 ;
  assign n33573 = ~n33571 & ~n33572 ;
  assign n33574 = \wishbone_rx_fifo_fifo_reg[13][1]/P0001  & n33201 ;
  assign n33575 = \wishbone_rx_fifo_fifo_reg[12][1]/P0001  & n33214 ;
  assign n33576 = ~n33574 & ~n33575 ;
  assign n33577 = n33573 & n33576 ;
  assign n33578 = n33570 & n33577 ;
  assign n33579 = n33563 & n33578 ;
  assign n33580 = ~\wishbone_rx_fifo_fifo_reg[0][1]/P0001  & n33164 ;
  assign n33581 = ~n33579 & ~n33580 ;
  assign n33582 = \wishbone_rx_fifo_fifo_reg[0][1]/P0001  & n33167 ;
  assign n33583 = ~n33581 & ~n33582 ;
  assign n33584 = \wishbone_rx_fifo_fifo_reg[14][20]/P0001  & n33212 ;
  assign n33585 = \wishbone_rx_fifo_fifo_reg[1][20]/P0001  & n33181 ;
  assign n33586 = ~n33584 & ~n33585 ;
  assign n33587 = \wishbone_rx_fifo_fifo_reg[2][20]/P0001  & n33207 ;
  assign n33588 = \wishbone_rx_fifo_fifo_reg[6][20]/P0001  & n33187 ;
  assign n33589 = ~n33587 & ~n33588 ;
  assign n33590 = n33586 & n33589 ;
  assign n33591 = \wishbone_rx_fifo_fifo_reg[10][20]/P0001  & n33189 ;
  assign n33592 = ~n33164 & ~n33591 ;
  assign n33593 = \wishbone_rx_fifo_fifo_reg[13][20]/P0001  & n33201 ;
  assign n33594 = \wishbone_rx_fifo_fifo_reg[11][20]/P0001  & n33203 ;
  assign n33595 = ~n33593 & ~n33594 ;
  assign n33596 = n33592 & n33595 ;
  assign n33597 = n33590 & n33596 ;
  assign n33598 = \wishbone_rx_fifo_fifo_reg[5][20]/P0001  & n33209 ;
  assign n33599 = \wishbone_rx_fifo_fifo_reg[15][20]/P0001  & n33172 ;
  assign n33600 = ~n33598 & ~n33599 ;
  assign n33601 = \wishbone_rx_fifo_fifo_reg[12][20]/P0001  & n33214 ;
  assign n33602 = \wishbone_rx_fifo_fifo_reg[8][20]/P0001  & n33179 ;
  assign n33603 = ~n33601 & ~n33602 ;
  assign n33604 = n33600 & n33603 ;
  assign n33605 = \wishbone_rx_fifo_fifo_reg[9][20]/P0001  & n33176 ;
  assign n33606 = \wishbone_rx_fifo_fifo_reg[7][20]/P0001  & n33192 ;
  assign n33607 = ~n33605 & ~n33606 ;
  assign n33608 = \wishbone_rx_fifo_fifo_reg[3][20]/P0001  & n33199 ;
  assign n33609 = \wishbone_rx_fifo_fifo_reg[4][20]/P0001  & n33194 ;
  assign n33610 = ~n33608 & ~n33609 ;
  assign n33611 = n33607 & n33610 ;
  assign n33612 = n33604 & n33611 ;
  assign n33613 = n33597 & n33612 ;
  assign n33614 = ~\wishbone_rx_fifo_fifo_reg[0][20]/P0001  & n33164 ;
  assign n33615 = ~n33613 & ~n33614 ;
  assign n33616 = \wishbone_rx_fifo_fifo_reg[0][20]/P0001  & n33167 ;
  assign n33617 = ~n33615 & ~n33616 ;
  assign n33618 = \wishbone_rx_fifo_fifo_reg[0][21]/P0001  & ~n33168 ;
  assign n33619 = \wishbone_rx_fifo_fifo_reg[7][21]/P0001  & n33192 ;
  assign n33620 = \wishbone_rx_fifo_fifo_reg[5][21]/P0001  & n33209 ;
  assign n33621 = ~n33619 & ~n33620 ;
  assign n33622 = \wishbone_rx_fifo_fifo_reg[2][21]/P0001  & n33207 ;
  assign n33623 = \wishbone_rx_fifo_fifo_reg[13][21]/P0001  & n33201 ;
  assign n33624 = ~n33622 & ~n33623 ;
  assign n33625 = n33621 & n33624 ;
  assign n33626 = \wishbone_rx_fifo_fifo_reg[6][21]/P0001  & n33187 ;
  assign n33627 = \wishbone_rx_fifo_fifo_reg[12][21]/P0001  & n33214 ;
  assign n33628 = ~n33626 & ~n33627 ;
  assign n33629 = \wishbone_rx_fifo_fifo_reg[9][21]/P0001  & n33176 ;
  assign n33630 = \wishbone_rx_fifo_fifo_reg[11][21]/P0001  & n33203 ;
  assign n33631 = ~n33629 & ~n33630 ;
  assign n33632 = n33628 & n33631 ;
  assign n33633 = n33625 & n33632 ;
  assign n33634 = \wishbone_rx_fifo_fifo_reg[3][21]/P0001  & n33199 ;
  assign n33635 = \wishbone_rx_fifo_fifo_reg[10][21]/P0001  & n33189 ;
  assign n33636 = \wishbone_rx_fifo_fifo_reg[1][21]/P0001  & n33181 ;
  assign n33637 = ~n33635 & ~n33636 ;
  assign n33638 = ~n33634 & n33637 ;
  assign n33639 = \wishbone_rx_fifo_fifo_reg[4][21]/P0001  & n33194 ;
  assign n33640 = \wishbone_rx_fifo_fifo_reg[15][21]/P0001  & n33172 ;
  assign n33641 = ~n33639 & ~n33640 ;
  assign n33642 = \wishbone_rx_fifo_fifo_reg[8][21]/P0001  & n33179 ;
  assign n33643 = \wishbone_rx_fifo_fifo_reg[14][21]/P0001  & n33212 ;
  assign n33644 = ~n33642 & ~n33643 ;
  assign n33645 = n33641 & n33644 ;
  assign n33646 = n33638 & n33645 ;
  assign n33647 = n33633 & n33646 ;
  assign n33648 = ~n33164 & ~n33647 ;
  assign n33649 = ~n33618 & ~n33648 ;
  assign n33650 = \wishbone_rx_fifo_fifo_reg[0][22]/P0001  & ~n33168 ;
  assign n33651 = \wishbone_rx_fifo_fifo_reg[7][22]/P0001  & n33192 ;
  assign n33652 = \wishbone_rx_fifo_fifo_reg[5][22]/P0001  & n33209 ;
  assign n33653 = ~n33651 & ~n33652 ;
  assign n33654 = \wishbone_rx_fifo_fifo_reg[2][22]/P0001  & n33207 ;
  assign n33655 = \wishbone_rx_fifo_fifo_reg[13][22]/P0001  & n33201 ;
  assign n33656 = ~n33654 & ~n33655 ;
  assign n33657 = n33653 & n33656 ;
  assign n33658 = \wishbone_rx_fifo_fifo_reg[6][22]/P0001  & n33187 ;
  assign n33659 = \wishbone_rx_fifo_fifo_reg[12][22]/P0001  & n33214 ;
  assign n33660 = ~n33658 & ~n33659 ;
  assign n33661 = \wishbone_rx_fifo_fifo_reg[9][22]/P0001  & n33176 ;
  assign n33662 = \wishbone_rx_fifo_fifo_reg[11][22]/P0001  & n33203 ;
  assign n33663 = ~n33661 & ~n33662 ;
  assign n33664 = n33660 & n33663 ;
  assign n33665 = n33657 & n33664 ;
  assign n33666 = \wishbone_rx_fifo_fifo_reg[3][22]/P0001  & n33199 ;
  assign n33667 = \wishbone_rx_fifo_fifo_reg[10][22]/P0001  & n33189 ;
  assign n33668 = \wishbone_rx_fifo_fifo_reg[1][22]/P0001  & n33181 ;
  assign n33669 = ~n33667 & ~n33668 ;
  assign n33670 = ~n33666 & n33669 ;
  assign n33671 = \wishbone_rx_fifo_fifo_reg[4][22]/P0001  & n33194 ;
  assign n33672 = \wishbone_rx_fifo_fifo_reg[15][22]/P0001  & n33172 ;
  assign n33673 = ~n33671 & ~n33672 ;
  assign n33674 = \wishbone_rx_fifo_fifo_reg[8][22]/P0001  & n33179 ;
  assign n33675 = \wishbone_rx_fifo_fifo_reg[14][22]/P0001  & n33212 ;
  assign n33676 = ~n33674 & ~n33675 ;
  assign n33677 = n33673 & n33676 ;
  assign n33678 = n33670 & n33677 ;
  assign n33679 = n33665 & n33678 ;
  assign n33680 = ~n33164 & ~n33679 ;
  assign n33681 = ~n33650 & ~n33680 ;
  assign n33682 = \wishbone_rx_fifo_fifo_reg[0][23]/P0001  & ~n33168 ;
  assign n33683 = \wishbone_rx_fifo_fifo_reg[7][23]/P0001  & n33192 ;
  assign n33684 = \wishbone_rx_fifo_fifo_reg[5][23]/P0001  & n33209 ;
  assign n33685 = ~n33683 & ~n33684 ;
  assign n33686 = \wishbone_rx_fifo_fifo_reg[2][23]/P0001  & n33207 ;
  assign n33687 = \wishbone_rx_fifo_fifo_reg[13][23]/P0001  & n33201 ;
  assign n33688 = ~n33686 & ~n33687 ;
  assign n33689 = n33685 & n33688 ;
  assign n33690 = \wishbone_rx_fifo_fifo_reg[6][23]/P0001  & n33187 ;
  assign n33691 = \wishbone_rx_fifo_fifo_reg[12][23]/P0001  & n33214 ;
  assign n33692 = ~n33690 & ~n33691 ;
  assign n33693 = \wishbone_rx_fifo_fifo_reg[9][23]/P0001  & n33176 ;
  assign n33694 = \wishbone_rx_fifo_fifo_reg[11][23]/P0001  & n33203 ;
  assign n33695 = ~n33693 & ~n33694 ;
  assign n33696 = n33692 & n33695 ;
  assign n33697 = n33689 & n33696 ;
  assign n33698 = \wishbone_rx_fifo_fifo_reg[3][23]/P0001  & n33199 ;
  assign n33699 = \wishbone_rx_fifo_fifo_reg[10][23]/P0001  & n33189 ;
  assign n33700 = \wishbone_rx_fifo_fifo_reg[1][23]/P0001  & n33181 ;
  assign n33701 = ~n33699 & ~n33700 ;
  assign n33702 = ~n33698 & n33701 ;
  assign n33703 = \wishbone_rx_fifo_fifo_reg[4][23]/P0001  & n33194 ;
  assign n33704 = \wishbone_rx_fifo_fifo_reg[15][23]/P0001  & n33172 ;
  assign n33705 = ~n33703 & ~n33704 ;
  assign n33706 = \wishbone_rx_fifo_fifo_reg[8][23]/P0001  & n33179 ;
  assign n33707 = \wishbone_rx_fifo_fifo_reg[14][23]/P0001  & n33212 ;
  assign n33708 = ~n33706 & ~n33707 ;
  assign n33709 = n33705 & n33708 ;
  assign n33710 = n33702 & n33709 ;
  assign n33711 = n33697 & n33710 ;
  assign n33712 = ~n33164 & ~n33711 ;
  assign n33713 = ~n33682 & ~n33712 ;
  assign n33714 = \wishbone_rx_fifo_fifo_reg[0][24]/P0001  & ~n33168 ;
  assign n33715 = \wishbone_rx_fifo_fifo_reg[2][24]/P0001  & n33207 ;
  assign n33716 = \wishbone_rx_fifo_fifo_reg[3][24]/P0001  & n33199 ;
  assign n33717 = ~n33715 & ~n33716 ;
  assign n33718 = \wishbone_rx_fifo_fifo_reg[4][24]/P0001  & n33194 ;
  assign n33719 = \wishbone_rx_fifo_fifo_reg[5][24]/P0001  & n33209 ;
  assign n33720 = ~n33718 & ~n33719 ;
  assign n33721 = n33717 & n33720 ;
  assign n33722 = \wishbone_rx_fifo_fifo_reg[9][24]/P0001  & n33176 ;
  assign n33723 = \wishbone_rx_fifo_fifo_reg[8][24]/P0001  & n33179 ;
  assign n33724 = ~n33722 & ~n33723 ;
  assign n33725 = \wishbone_rx_fifo_fifo_reg[12][24]/P0001  & n33214 ;
  assign n33726 = \wishbone_rx_fifo_fifo_reg[13][24]/P0001  & n33201 ;
  assign n33727 = ~n33725 & ~n33726 ;
  assign n33728 = n33724 & n33727 ;
  assign n33729 = n33721 & n33728 ;
  assign n33730 = \wishbone_rx_fifo_fifo_reg[14][24]/P0001  & n33212 ;
  assign n33731 = \wishbone_rx_fifo_fifo_reg[6][24]/P0001  & n33187 ;
  assign n33732 = \wishbone_rx_fifo_fifo_reg[15][24]/P0001  & n33172 ;
  assign n33733 = ~n33731 & ~n33732 ;
  assign n33734 = ~n33730 & n33733 ;
  assign n33735 = \wishbone_rx_fifo_fifo_reg[10][24]/P0001  & n33189 ;
  assign n33736 = \wishbone_rx_fifo_fifo_reg[7][24]/P0001  & n33192 ;
  assign n33737 = ~n33735 & ~n33736 ;
  assign n33738 = \wishbone_rx_fifo_fifo_reg[1][24]/P0001  & n33181 ;
  assign n33739 = \wishbone_rx_fifo_fifo_reg[11][24]/P0001  & n33203 ;
  assign n33740 = ~n33738 & ~n33739 ;
  assign n33741 = n33737 & n33740 ;
  assign n33742 = n33734 & n33741 ;
  assign n33743 = n33729 & n33742 ;
  assign n33744 = ~n33164 & ~n33743 ;
  assign n33745 = ~n33714 & ~n33744 ;
  assign n33746 = \wishbone_rx_fifo_fifo_reg[0][25]/P0001  & ~n33168 ;
  assign n33747 = \wishbone_rx_fifo_fifo_reg[15][25]/P0001  & n33172 ;
  assign n33748 = \wishbone_rx_fifo_fifo_reg[9][25]/P0001  & n33176 ;
  assign n33749 = ~n33747 & ~n33748 ;
  assign n33750 = \wishbone_rx_fifo_fifo_reg[8][25]/P0001  & n33179 ;
  assign n33751 = \wishbone_rx_fifo_fifo_reg[3][25]/P0001  & n33199 ;
  assign n33752 = ~n33750 & ~n33751 ;
  assign n33753 = n33749 & n33752 ;
  assign n33754 = \wishbone_rx_fifo_fifo_reg[6][25]/P0001  & n33187 ;
  assign n33755 = \wishbone_rx_fifo_fifo_reg[10][25]/P0001  & n33189 ;
  assign n33756 = ~n33754 & ~n33755 ;
  assign n33757 = \wishbone_rx_fifo_fifo_reg[7][25]/P0001  & n33192 ;
  assign n33758 = \wishbone_rx_fifo_fifo_reg[4][25]/P0001  & n33194 ;
  assign n33759 = ~n33757 & ~n33758 ;
  assign n33760 = n33756 & n33759 ;
  assign n33761 = n33753 & n33760 ;
  assign n33762 = \wishbone_rx_fifo_fifo_reg[1][25]/P0001  & n33181 ;
  assign n33763 = \wishbone_rx_fifo_fifo_reg[13][25]/P0001  & n33201 ;
  assign n33764 = \wishbone_rx_fifo_fifo_reg[2][25]/P0001  & n33207 ;
  assign n33765 = ~n33763 & ~n33764 ;
  assign n33766 = ~n33762 & n33765 ;
  assign n33767 = \wishbone_rx_fifo_fifo_reg[11][25]/P0001  & n33203 ;
  assign n33768 = \wishbone_rx_fifo_fifo_reg[5][25]/P0001  & n33209 ;
  assign n33769 = ~n33767 & ~n33768 ;
  assign n33770 = \wishbone_rx_fifo_fifo_reg[14][25]/P0001  & n33212 ;
  assign n33771 = \wishbone_rx_fifo_fifo_reg[12][25]/P0001  & n33214 ;
  assign n33772 = ~n33770 & ~n33771 ;
  assign n33773 = n33769 & n33772 ;
  assign n33774 = n33766 & n33773 ;
  assign n33775 = n33761 & n33774 ;
  assign n33776 = ~n33164 & ~n33775 ;
  assign n33777 = ~n33746 & ~n33776 ;
  assign n33778 = \wishbone_rx_fifo_fifo_reg[0][26]/P0001  & ~n33168 ;
  assign n33779 = \wishbone_rx_fifo_fifo_reg[8][26]/P0001  & n33179 ;
  assign n33780 = \wishbone_rx_fifo_fifo_reg[5][26]/P0001  & n33209 ;
  assign n33781 = ~n33779 & ~n33780 ;
  assign n33782 = \wishbone_rx_fifo_fifo_reg[13][26]/P0001  & n33201 ;
  assign n33783 = \wishbone_rx_fifo_fifo_reg[4][26]/P0001  & n33194 ;
  assign n33784 = ~n33782 & ~n33783 ;
  assign n33785 = n33781 & n33784 ;
  assign n33786 = \wishbone_rx_fifo_fifo_reg[9][26]/P0001  & n33176 ;
  assign n33787 = \wishbone_rx_fifo_fifo_reg[3][26]/P0001  & n33199 ;
  assign n33788 = ~n33786 & ~n33787 ;
  assign n33789 = \wishbone_rx_fifo_fifo_reg[6][26]/P0001  & n33187 ;
  assign n33790 = \wishbone_rx_fifo_fifo_reg[15][26]/P0001  & n33172 ;
  assign n33791 = ~n33789 & ~n33790 ;
  assign n33792 = n33788 & n33791 ;
  assign n33793 = n33785 & n33792 ;
  assign n33794 = \wishbone_rx_fifo_fifo_reg[11][26]/P0001  & n33203 ;
  assign n33795 = \wishbone_rx_fifo_fifo_reg[1][26]/P0001  & n33181 ;
  assign n33796 = \wishbone_rx_fifo_fifo_reg[10][26]/P0001  & n33189 ;
  assign n33797 = ~n33795 & ~n33796 ;
  assign n33798 = ~n33794 & n33797 ;
  assign n33799 = \wishbone_rx_fifo_fifo_reg[14][26]/P0001  & n33212 ;
  assign n33800 = \wishbone_rx_fifo_fifo_reg[12][26]/P0001  & n33214 ;
  assign n33801 = ~n33799 & ~n33800 ;
  assign n33802 = \wishbone_rx_fifo_fifo_reg[7][26]/P0001  & n33192 ;
  assign n33803 = \wishbone_rx_fifo_fifo_reg[2][26]/P0001  & n33207 ;
  assign n33804 = ~n33802 & ~n33803 ;
  assign n33805 = n33801 & n33804 ;
  assign n33806 = n33798 & n33805 ;
  assign n33807 = n33793 & n33806 ;
  assign n33808 = ~n33164 & ~n33807 ;
  assign n33809 = ~n33778 & ~n33808 ;
  assign n33810 = \wishbone_rx_fifo_fifo_reg[11][27]/P0001  & n33203 ;
  assign n33811 = \wishbone_rx_fifo_fifo_reg[9][27]/P0001  & n33176 ;
  assign n33812 = ~n33810 & ~n33811 ;
  assign n33813 = \wishbone_rx_fifo_fifo_reg[6][27]/P0001  & n33187 ;
  assign n33814 = \wishbone_rx_fifo_fifo_reg[15][27]/P0001  & n33172 ;
  assign n33815 = ~n33813 & ~n33814 ;
  assign n33816 = n33812 & n33815 ;
  assign n33817 = \wishbone_rx_fifo_fifo_reg[12][27]/P0001  & n33214 ;
  assign n33818 = ~n33164 & ~n33817 ;
  assign n33819 = \wishbone_rx_fifo_fifo_reg[3][27]/P0001  & n33199 ;
  assign n33820 = \wishbone_rx_fifo_fifo_reg[1][27]/P0001  & n33181 ;
  assign n33821 = ~n33819 & ~n33820 ;
  assign n33822 = n33818 & n33821 ;
  assign n33823 = n33816 & n33822 ;
  assign n33824 = \wishbone_rx_fifo_fifo_reg[5][27]/P0001  & n33209 ;
  assign n33825 = \wishbone_rx_fifo_fifo_reg[10][27]/P0001  & n33189 ;
  assign n33826 = ~n33824 & ~n33825 ;
  assign n33827 = \wishbone_rx_fifo_fifo_reg[2][27]/P0001  & n33207 ;
  assign n33828 = \wishbone_rx_fifo_fifo_reg[4][27]/P0001  & n33194 ;
  assign n33829 = ~n33827 & ~n33828 ;
  assign n33830 = n33826 & n33829 ;
  assign n33831 = \wishbone_rx_fifo_fifo_reg[7][27]/P0001  & n33192 ;
  assign n33832 = \wishbone_rx_fifo_fifo_reg[8][27]/P0001  & n33179 ;
  assign n33833 = ~n33831 & ~n33832 ;
  assign n33834 = \wishbone_rx_fifo_fifo_reg[13][27]/P0001  & n33201 ;
  assign n33835 = \wishbone_rx_fifo_fifo_reg[14][27]/P0001  & n33212 ;
  assign n33836 = ~n33834 & ~n33835 ;
  assign n33837 = n33833 & n33836 ;
  assign n33838 = n33830 & n33837 ;
  assign n33839 = n33823 & n33838 ;
  assign n33840 = ~\wishbone_rx_fifo_fifo_reg[0][27]/P0001  & n33164 ;
  assign n33841 = ~n33839 & ~n33840 ;
  assign n33842 = \wishbone_rx_fifo_fifo_reg[0][27]/P0001  & n33167 ;
  assign n33843 = ~n33841 & ~n33842 ;
  assign n33844 = \wishbone_rx_fifo_fifo_reg[13][28]/P0001  & n33201 ;
  assign n33845 = \wishbone_rx_fifo_fifo_reg[5][28]/P0001  & n33209 ;
  assign n33846 = ~n33844 & ~n33845 ;
  assign n33847 = \wishbone_rx_fifo_fifo_reg[6][28]/P0001  & n33187 ;
  assign n33848 = \wishbone_rx_fifo_fifo_reg[8][28]/P0001  & n33179 ;
  assign n33849 = ~n33847 & ~n33848 ;
  assign n33850 = n33846 & n33849 ;
  assign n33851 = \wishbone_rx_fifo_fifo_reg[12][28]/P0001  & n33214 ;
  assign n33852 = ~n33164 & ~n33851 ;
  assign n33853 = \wishbone_rx_fifo_fifo_reg[15][28]/P0001  & n33172 ;
  assign n33854 = \wishbone_rx_fifo_fifo_reg[2][28]/P0001  & n33207 ;
  assign n33855 = ~n33853 & ~n33854 ;
  assign n33856 = n33852 & n33855 ;
  assign n33857 = n33850 & n33856 ;
  assign n33858 = \wishbone_rx_fifo_fifo_reg[14][28]/P0001  & n33212 ;
  assign n33859 = \wishbone_rx_fifo_fifo_reg[10][28]/P0001  & n33189 ;
  assign n33860 = ~n33858 & ~n33859 ;
  assign n33861 = \wishbone_rx_fifo_fifo_reg[3][28]/P0001  & n33199 ;
  assign n33862 = \wishbone_rx_fifo_fifo_reg[7][28]/P0001  & n33192 ;
  assign n33863 = ~n33861 & ~n33862 ;
  assign n33864 = n33860 & n33863 ;
  assign n33865 = \wishbone_rx_fifo_fifo_reg[11][28]/P0001  & n33203 ;
  assign n33866 = \wishbone_rx_fifo_fifo_reg[9][28]/P0001  & n33176 ;
  assign n33867 = ~n33865 & ~n33866 ;
  assign n33868 = \wishbone_rx_fifo_fifo_reg[1][28]/P0001  & n33181 ;
  assign n33869 = \wishbone_rx_fifo_fifo_reg[4][28]/P0001  & n33194 ;
  assign n33870 = ~n33868 & ~n33869 ;
  assign n33871 = n33867 & n33870 ;
  assign n33872 = n33864 & n33871 ;
  assign n33873 = n33857 & n33872 ;
  assign n33874 = ~\wishbone_rx_fifo_fifo_reg[0][28]/P0001  & n33164 ;
  assign n33875 = ~n33873 & ~n33874 ;
  assign n33876 = \wishbone_rx_fifo_fifo_reg[0][28]/P0001  & n33167 ;
  assign n33877 = ~n33875 & ~n33876 ;
  assign n33878 = \wishbone_rx_fifo_fifo_reg[1][29]/P0001  & n33181 ;
  assign n33879 = \wishbone_rx_fifo_fifo_reg[5][29]/P0001  & n33209 ;
  assign n33880 = ~n33878 & ~n33879 ;
  assign n33881 = \wishbone_rx_fifo_fifo_reg[8][29]/P0001  & n33179 ;
  assign n33882 = \wishbone_rx_fifo_fifo_reg[6][29]/P0001  & n33187 ;
  assign n33883 = ~n33881 & ~n33882 ;
  assign n33884 = n33880 & n33883 ;
  assign n33885 = \wishbone_rx_fifo_fifo_reg[10][29]/P0001  & n33189 ;
  assign n33886 = ~n33164 & ~n33885 ;
  assign n33887 = \wishbone_rx_fifo_fifo_reg[13][29]/P0001  & n33201 ;
  assign n33888 = \wishbone_rx_fifo_fifo_reg[14][29]/P0001  & n33212 ;
  assign n33889 = ~n33887 & ~n33888 ;
  assign n33890 = n33886 & n33889 ;
  assign n33891 = n33884 & n33890 ;
  assign n33892 = \wishbone_rx_fifo_fifo_reg[3][29]/P0001  & n33199 ;
  assign n33893 = \wishbone_rx_fifo_fifo_reg[15][29]/P0001  & n33172 ;
  assign n33894 = ~n33892 & ~n33893 ;
  assign n33895 = \wishbone_rx_fifo_fifo_reg[11][29]/P0001  & n33203 ;
  assign n33896 = \wishbone_rx_fifo_fifo_reg[2][29]/P0001  & n33207 ;
  assign n33897 = ~n33895 & ~n33896 ;
  assign n33898 = n33894 & n33897 ;
  assign n33899 = \wishbone_rx_fifo_fifo_reg[9][29]/P0001  & n33176 ;
  assign n33900 = \wishbone_rx_fifo_fifo_reg[7][29]/P0001  & n33192 ;
  assign n33901 = ~n33899 & ~n33900 ;
  assign n33902 = \wishbone_rx_fifo_fifo_reg[12][29]/P0001  & n33214 ;
  assign n33903 = \wishbone_rx_fifo_fifo_reg[4][29]/P0001  & n33194 ;
  assign n33904 = ~n33902 & ~n33903 ;
  assign n33905 = n33901 & n33904 ;
  assign n33906 = n33898 & n33905 ;
  assign n33907 = n33891 & n33906 ;
  assign n33908 = ~\wishbone_rx_fifo_fifo_reg[0][29]/P0001  & n33164 ;
  assign n33909 = ~n33907 & ~n33908 ;
  assign n33910 = \wishbone_rx_fifo_fifo_reg[0][29]/P0001  & n33167 ;
  assign n33911 = ~n33909 & ~n33910 ;
  assign n33912 = \wishbone_rx_fifo_fifo_reg[0][2]/P0001  & ~n33168 ;
  assign n33913 = \wishbone_rx_fifo_fifo_reg[10][2]/P0001  & n33189 ;
  assign n33914 = \wishbone_rx_fifo_fifo_reg[6][2]/P0001  & n33187 ;
  assign n33915 = ~n33913 & ~n33914 ;
  assign n33916 = \wishbone_rx_fifo_fifo_reg[12][2]/P0001  & n33214 ;
  assign n33917 = \wishbone_rx_fifo_fifo_reg[4][2]/P0001  & n33194 ;
  assign n33918 = ~n33916 & ~n33917 ;
  assign n33919 = n33915 & n33918 ;
  assign n33920 = \wishbone_rx_fifo_fifo_reg[3][2]/P0001  & n33199 ;
  assign n33921 = \wishbone_rx_fifo_fifo_reg[9][2]/P0001  & n33176 ;
  assign n33922 = ~n33920 & ~n33921 ;
  assign n33923 = \wishbone_rx_fifo_fifo_reg[5][2]/P0001  & n33209 ;
  assign n33924 = \wishbone_rx_fifo_fifo_reg[7][2]/P0001  & n33192 ;
  assign n33925 = ~n33923 & ~n33924 ;
  assign n33926 = n33922 & n33925 ;
  assign n33927 = n33919 & n33926 ;
  assign n33928 = \wishbone_rx_fifo_fifo_reg[15][2]/P0001  & n33172 ;
  assign n33929 = \wishbone_rx_fifo_fifo_reg[8][2]/P0001  & n33179 ;
  assign n33930 = \wishbone_rx_fifo_fifo_reg[11][2]/P0001  & n33203 ;
  assign n33931 = ~n33929 & ~n33930 ;
  assign n33932 = ~n33928 & n33931 ;
  assign n33933 = \wishbone_rx_fifo_fifo_reg[1][2]/P0001  & n33181 ;
  assign n33934 = \wishbone_rx_fifo_fifo_reg[13][2]/P0001  & n33201 ;
  assign n33935 = ~n33933 & ~n33934 ;
  assign n33936 = \wishbone_rx_fifo_fifo_reg[2][2]/P0001  & n33207 ;
  assign n33937 = \wishbone_rx_fifo_fifo_reg[14][2]/P0001  & n33212 ;
  assign n33938 = ~n33936 & ~n33937 ;
  assign n33939 = n33935 & n33938 ;
  assign n33940 = n33932 & n33939 ;
  assign n33941 = n33927 & n33940 ;
  assign n33942 = ~n33164 & ~n33941 ;
  assign n33943 = ~n33912 & ~n33942 ;
  assign n33944 = \wishbone_rx_fifo_fifo_reg[0][30]/P0001  & ~n33168 ;
  assign n33945 = \wishbone_rx_fifo_fifo_reg[13][30]/P0001  & n33201 ;
  assign n33946 = \wishbone_rx_fifo_fifo_reg[9][30]/P0001  & n33176 ;
  assign n33947 = ~n33945 & ~n33946 ;
  assign n33948 = \wishbone_rx_fifo_fifo_reg[8][30]/P0001  & n33179 ;
  assign n33949 = \wishbone_rx_fifo_fifo_reg[14][30]/P0001  & n33212 ;
  assign n33950 = ~n33948 & ~n33949 ;
  assign n33951 = n33947 & n33950 ;
  assign n33952 = \wishbone_rx_fifo_fifo_reg[3][30]/P0001  & n33199 ;
  assign n33953 = \wishbone_rx_fifo_fifo_reg[5][30]/P0001  & n33209 ;
  assign n33954 = ~n33952 & ~n33953 ;
  assign n33955 = \wishbone_rx_fifo_fifo_reg[15][30]/P0001  & n33172 ;
  assign n33956 = \wishbone_rx_fifo_fifo_reg[2][30]/P0001  & n33207 ;
  assign n33957 = ~n33955 & ~n33956 ;
  assign n33958 = n33954 & n33957 ;
  assign n33959 = n33951 & n33958 ;
  assign n33960 = \wishbone_rx_fifo_fifo_reg[1][30]/P0001  & n33181 ;
  assign n33961 = \wishbone_rx_fifo_fifo_reg[4][30]/P0001  & n33194 ;
  assign n33962 = \wishbone_rx_fifo_fifo_reg[6][30]/P0001  & n33187 ;
  assign n33963 = ~n33961 & ~n33962 ;
  assign n33964 = ~n33960 & n33963 ;
  assign n33965 = \wishbone_rx_fifo_fifo_reg[7][30]/P0001  & n33192 ;
  assign n33966 = \wishbone_rx_fifo_fifo_reg[10][30]/P0001  & n33189 ;
  assign n33967 = ~n33965 & ~n33966 ;
  assign n33968 = \wishbone_rx_fifo_fifo_reg[11][30]/P0001  & n33203 ;
  assign n33969 = \wishbone_rx_fifo_fifo_reg[12][30]/P0001  & n33214 ;
  assign n33970 = ~n33968 & ~n33969 ;
  assign n33971 = n33967 & n33970 ;
  assign n33972 = n33964 & n33971 ;
  assign n33973 = n33959 & n33972 ;
  assign n33974 = ~n33164 & ~n33973 ;
  assign n33975 = ~n33944 & ~n33974 ;
  assign n33976 = \wishbone_rx_fifo_fifo_reg[11][31]/P0001  & n33203 ;
  assign n33977 = \wishbone_rx_fifo_fifo_reg[3][31]/P0001  & n33199 ;
  assign n33978 = ~n33976 & ~n33977 ;
  assign n33979 = \wishbone_rx_fifo_fifo_reg[6][31]/P0001  & n33187 ;
  assign n33980 = \wishbone_rx_fifo_fifo_reg[8][31]/P0001  & n33179 ;
  assign n33981 = ~n33979 & ~n33980 ;
  assign n33982 = n33978 & n33981 ;
  assign n33983 = \wishbone_rx_fifo_fifo_reg[12][31]/P0001  & n33214 ;
  assign n33984 = ~n33164 & ~n33983 ;
  assign n33985 = \wishbone_rx_fifo_fifo_reg[5][31]/P0001  & n33209 ;
  assign n33986 = \wishbone_rx_fifo_fifo_reg[2][31]/P0001  & n33207 ;
  assign n33987 = ~n33985 & ~n33986 ;
  assign n33988 = n33984 & n33987 ;
  assign n33989 = n33982 & n33988 ;
  assign n33990 = \wishbone_rx_fifo_fifo_reg[1][31]/P0001  & n33181 ;
  assign n33991 = \wishbone_rx_fifo_fifo_reg[10][31]/P0001  & n33189 ;
  assign n33992 = ~n33990 & ~n33991 ;
  assign n33993 = \wishbone_rx_fifo_fifo_reg[9][31]/P0001  & n33176 ;
  assign n33994 = \wishbone_rx_fifo_fifo_reg[4][31]/P0001  & n33194 ;
  assign n33995 = ~n33993 & ~n33994 ;
  assign n33996 = n33992 & n33995 ;
  assign n33997 = \wishbone_rx_fifo_fifo_reg[15][31]/P0001  & n33172 ;
  assign n33998 = \wishbone_rx_fifo_fifo_reg[13][31]/P0001  & n33201 ;
  assign n33999 = ~n33997 & ~n33998 ;
  assign n34000 = \wishbone_rx_fifo_fifo_reg[7][31]/P0001  & n33192 ;
  assign n34001 = \wishbone_rx_fifo_fifo_reg[14][31]/P0001  & n33212 ;
  assign n34002 = ~n34000 & ~n34001 ;
  assign n34003 = n33999 & n34002 ;
  assign n34004 = n33996 & n34003 ;
  assign n34005 = n33989 & n34004 ;
  assign n34006 = ~\wishbone_rx_fifo_fifo_reg[0][31]/P0001  & n33164 ;
  assign n34007 = ~n34005 & ~n34006 ;
  assign n34008 = \wishbone_rx_fifo_fifo_reg[0][31]/P0001  & n33167 ;
  assign n34009 = ~n34007 & ~n34008 ;
  assign n34010 = \wishbone_rx_fifo_fifo_reg[0][3]/P0001  & ~n33168 ;
  assign n34011 = \wishbone_rx_fifo_fifo_reg[5][3]/P0001  & n33209 ;
  assign n34012 = \wishbone_rx_fifo_fifo_reg[1][3]/P0001  & n33181 ;
  assign n34013 = ~n34011 & ~n34012 ;
  assign n34014 = \wishbone_rx_fifo_fifo_reg[11][3]/P0001  & n33203 ;
  assign n34015 = \wishbone_rx_fifo_fifo_reg[4][3]/P0001  & n33194 ;
  assign n34016 = ~n34014 & ~n34015 ;
  assign n34017 = n34013 & n34016 ;
  assign n34018 = \wishbone_rx_fifo_fifo_reg[8][3]/P0001  & n33179 ;
  assign n34019 = \wishbone_rx_fifo_fifo_reg[7][3]/P0001  & n33192 ;
  assign n34020 = ~n34018 & ~n34019 ;
  assign n34021 = \wishbone_rx_fifo_fifo_reg[10][3]/P0001  & n33189 ;
  assign n34022 = \wishbone_rx_fifo_fifo_reg[12][3]/P0001  & n33214 ;
  assign n34023 = ~n34021 & ~n34022 ;
  assign n34024 = n34020 & n34023 ;
  assign n34025 = n34017 & n34024 ;
  assign n34026 = \wishbone_rx_fifo_fifo_reg[3][3]/P0001  & n33199 ;
  assign n34027 = \wishbone_rx_fifo_fifo_reg[9][3]/P0001  & n33176 ;
  assign n34028 = \wishbone_rx_fifo_fifo_reg[2][3]/P0001  & n33207 ;
  assign n34029 = ~n34027 & ~n34028 ;
  assign n34030 = ~n34026 & n34029 ;
  assign n34031 = \wishbone_rx_fifo_fifo_reg[13][3]/P0001  & n33201 ;
  assign n34032 = \wishbone_rx_fifo_fifo_reg[6][3]/P0001  & n33187 ;
  assign n34033 = ~n34031 & ~n34032 ;
  assign n34034 = \wishbone_rx_fifo_fifo_reg[14][3]/P0001  & n33212 ;
  assign n34035 = \wishbone_rx_fifo_fifo_reg[15][3]/P0001  & n33172 ;
  assign n34036 = ~n34034 & ~n34035 ;
  assign n34037 = n34033 & n34036 ;
  assign n34038 = n34030 & n34037 ;
  assign n34039 = n34025 & n34038 ;
  assign n34040 = ~n33164 & ~n34039 ;
  assign n34041 = ~n34010 & ~n34040 ;
  assign n34042 = \wishbone_rx_fifo_fifo_reg[11][4]/P0001  & n33203 ;
  assign n34043 = \wishbone_rx_fifo_fifo_reg[3][4]/P0001  & n33199 ;
  assign n34044 = ~n34042 & ~n34043 ;
  assign n34045 = \wishbone_rx_fifo_fifo_reg[9][4]/P0001  & n33176 ;
  assign n34046 = \wishbone_rx_fifo_fifo_reg[8][4]/P0001  & n33179 ;
  assign n34047 = ~n34045 & ~n34046 ;
  assign n34048 = n34044 & n34047 ;
  assign n34049 = \wishbone_rx_fifo_fifo_reg[12][4]/P0001  & n33214 ;
  assign n34050 = ~n33164 & ~n34049 ;
  assign n34051 = \wishbone_rx_fifo_fifo_reg[5][4]/P0001  & n33209 ;
  assign n34052 = \wishbone_rx_fifo_fifo_reg[2][4]/P0001  & n33207 ;
  assign n34053 = ~n34051 & ~n34052 ;
  assign n34054 = n34050 & n34053 ;
  assign n34055 = n34048 & n34054 ;
  assign n34056 = \wishbone_rx_fifo_fifo_reg[1][4]/P0001  & n33181 ;
  assign n34057 = \wishbone_rx_fifo_fifo_reg[10][4]/P0001  & n33189 ;
  assign n34058 = ~n34056 & ~n34057 ;
  assign n34059 = \wishbone_rx_fifo_fifo_reg[6][4]/P0001  & n33187 ;
  assign n34060 = \wishbone_rx_fifo_fifo_reg[4][4]/P0001  & n33194 ;
  assign n34061 = ~n34059 & ~n34060 ;
  assign n34062 = n34058 & n34061 ;
  assign n34063 = \wishbone_rx_fifo_fifo_reg[15][4]/P0001  & n33172 ;
  assign n34064 = \wishbone_rx_fifo_fifo_reg[13][4]/P0001  & n33201 ;
  assign n34065 = ~n34063 & ~n34064 ;
  assign n34066 = \wishbone_rx_fifo_fifo_reg[7][4]/P0001  & n33192 ;
  assign n34067 = \wishbone_rx_fifo_fifo_reg[14][4]/P0001  & n33212 ;
  assign n34068 = ~n34066 & ~n34067 ;
  assign n34069 = n34065 & n34068 ;
  assign n34070 = n34062 & n34069 ;
  assign n34071 = n34055 & n34070 ;
  assign n34072 = ~\wishbone_rx_fifo_fifo_reg[0][4]/P0001  & n33164 ;
  assign n34073 = ~n34071 & ~n34072 ;
  assign n34074 = \wishbone_rx_fifo_fifo_reg[0][4]/P0001  & n33167 ;
  assign n34075 = ~n34073 & ~n34074 ;
  assign n34076 = \wishbone_rx_fifo_fifo_reg[4][5]/P0001  & n33194 ;
  assign n34077 = \wishbone_rx_fifo_fifo_reg[13][5]/P0001  & n33201 ;
  assign n34078 = ~n34076 & ~n34077 ;
  assign n34079 = \wishbone_rx_fifo_fifo_reg[2][5]/P0001  & n33207 ;
  assign n34080 = \wishbone_rx_fifo_fifo_reg[12][5]/P0001  & n33214 ;
  assign n34081 = ~n34079 & ~n34080 ;
  assign n34082 = n34078 & n34081 ;
  assign n34083 = \wishbone_rx_fifo_fifo_reg[10][5]/P0001  & n33189 ;
  assign n34084 = ~n33164 & ~n34083 ;
  assign n34085 = \wishbone_rx_fifo_fifo_reg[1][5]/P0001  & n33181 ;
  assign n34086 = \wishbone_rx_fifo_fifo_reg[8][5]/P0001  & n33179 ;
  assign n34087 = ~n34085 & ~n34086 ;
  assign n34088 = n34084 & n34087 ;
  assign n34089 = n34082 & n34088 ;
  assign n34090 = \wishbone_rx_fifo_fifo_reg[6][5]/P0001  & n33187 ;
  assign n34091 = \wishbone_rx_fifo_fifo_reg[7][5]/P0001  & n33192 ;
  assign n34092 = ~n34090 & ~n34091 ;
  assign n34093 = \wishbone_rx_fifo_fifo_reg[9][5]/P0001  & n33176 ;
  assign n34094 = \wishbone_rx_fifo_fifo_reg[5][5]/P0001  & n33209 ;
  assign n34095 = ~n34093 & ~n34094 ;
  assign n34096 = n34092 & n34095 ;
  assign n34097 = \wishbone_rx_fifo_fifo_reg[15][5]/P0001  & n33172 ;
  assign n34098 = \wishbone_rx_fifo_fifo_reg[3][5]/P0001  & n33199 ;
  assign n34099 = ~n34097 & ~n34098 ;
  assign n34100 = \wishbone_rx_fifo_fifo_reg[14][5]/P0001  & n33212 ;
  assign n34101 = \wishbone_rx_fifo_fifo_reg[11][5]/P0001  & n33203 ;
  assign n34102 = ~n34100 & ~n34101 ;
  assign n34103 = n34099 & n34102 ;
  assign n34104 = n34096 & n34103 ;
  assign n34105 = n34089 & n34104 ;
  assign n34106 = ~n33167 & n34105 ;
  assign n34107 = \wishbone_rx_fifo_fifo_reg[0][5]/P0001  & ~n34106 ;
  assign n34108 = ~n33164 & ~n34105 ;
  assign n34109 = ~n34107 & ~n34108 ;
  assign n34110 = \wishbone_rx_fifo_fifo_reg[0][6]/P0001  & ~n33168 ;
  assign n34111 = \wishbone_rx_fifo_fifo_reg[9][6]/P0001  & n33176 ;
  assign n34112 = \wishbone_rx_fifo_fifo_reg[6][6]/P0001  & n33187 ;
  assign n34113 = ~n34111 & ~n34112 ;
  assign n34114 = \wishbone_rx_fifo_fifo_reg[2][6]/P0001  & n33207 ;
  assign n34115 = \wishbone_rx_fifo_fifo_reg[1][6]/P0001  & n33181 ;
  assign n34116 = ~n34114 & ~n34115 ;
  assign n34117 = n34113 & n34116 ;
  assign n34118 = \wishbone_rx_fifo_fifo_reg[5][6]/P0001  & n33209 ;
  assign n34119 = \wishbone_rx_fifo_fifo_reg[14][6]/P0001  & n33212 ;
  assign n34120 = ~n34118 & ~n34119 ;
  assign n34121 = \wishbone_rx_fifo_fifo_reg[12][6]/P0001  & n33214 ;
  assign n34122 = \wishbone_rx_fifo_fifo_reg[3][6]/P0001  & n33199 ;
  assign n34123 = ~n34121 & ~n34122 ;
  assign n34124 = n34120 & n34123 ;
  assign n34125 = n34117 & n34124 ;
  assign n34126 = \wishbone_rx_fifo_fifo_reg[7][6]/P0001  & n33192 ;
  assign n34127 = \wishbone_rx_fifo_fifo_reg[10][6]/P0001  & n33189 ;
  assign n34128 = \wishbone_rx_fifo_fifo_reg[8][6]/P0001  & n33179 ;
  assign n34129 = ~n34127 & ~n34128 ;
  assign n34130 = ~n34126 & n34129 ;
  assign n34131 = \wishbone_rx_fifo_fifo_reg[4][6]/P0001  & n33194 ;
  assign n34132 = \wishbone_rx_fifo_fifo_reg[11][6]/P0001  & n33203 ;
  assign n34133 = ~n34131 & ~n34132 ;
  assign n34134 = \wishbone_rx_fifo_fifo_reg[15][6]/P0001  & n33172 ;
  assign n34135 = \wishbone_rx_fifo_fifo_reg[13][6]/P0001  & n33201 ;
  assign n34136 = ~n34134 & ~n34135 ;
  assign n34137 = n34133 & n34136 ;
  assign n34138 = n34130 & n34137 ;
  assign n34139 = n34125 & n34138 ;
  assign n34140 = ~n33164 & ~n34139 ;
  assign n34141 = ~n34110 & ~n34140 ;
  assign n34142 = \wishbone_rx_fifo_fifo_reg[13][7]/P0001  & n33201 ;
  assign n34143 = \wishbone_rx_fifo_fifo_reg[9][7]/P0001  & n33176 ;
  assign n34144 = ~n34142 & ~n34143 ;
  assign n34145 = \wishbone_rx_fifo_fifo_reg[6][7]/P0001  & n33187 ;
  assign n34146 = \wishbone_rx_fifo_fifo_reg[12][7]/P0001  & n33214 ;
  assign n34147 = ~n34145 & ~n34146 ;
  assign n34148 = n34144 & n34147 ;
  assign n34149 = \wishbone_rx_fifo_fifo_reg[3][7]/P0001  & n33199 ;
  assign n34150 = ~n33164 & ~n34149 ;
  assign n34151 = \wishbone_rx_fifo_fifo_reg[2][7]/P0001  & n33207 ;
  assign n34152 = \wishbone_rx_fifo_fifo_reg[15][7]/P0001  & n33172 ;
  assign n34153 = ~n34151 & ~n34152 ;
  assign n34154 = n34150 & n34153 ;
  assign n34155 = n34148 & n34154 ;
  assign n34156 = \wishbone_rx_fifo_fifo_reg[8][7]/P0001  & n33179 ;
  assign n34157 = \wishbone_rx_fifo_fifo_reg[5][7]/P0001  & n33209 ;
  assign n34158 = ~n34156 & ~n34157 ;
  assign n34159 = \wishbone_rx_fifo_fifo_reg[11][7]/P0001  & n33203 ;
  assign n34160 = \wishbone_rx_fifo_fifo_reg[7][7]/P0001  & n33192 ;
  assign n34161 = ~n34159 & ~n34160 ;
  assign n34162 = n34158 & n34161 ;
  assign n34163 = \wishbone_rx_fifo_fifo_reg[14][7]/P0001  & n33212 ;
  assign n34164 = \wishbone_rx_fifo_fifo_reg[10][7]/P0001  & n33189 ;
  assign n34165 = ~n34163 & ~n34164 ;
  assign n34166 = \wishbone_rx_fifo_fifo_reg[1][7]/P0001  & n33181 ;
  assign n34167 = \wishbone_rx_fifo_fifo_reg[4][7]/P0001  & n33194 ;
  assign n34168 = ~n34166 & ~n34167 ;
  assign n34169 = n34165 & n34168 ;
  assign n34170 = n34162 & n34169 ;
  assign n34171 = n34155 & n34170 ;
  assign n34172 = ~\wishbone_rx_fifo_fifo_reg[0][7]/P0001  & n33164 ;
  assign n34173 = ~n34171 & ~n34172 ;
  assign n34174 = \wishbone_rx_fifo_fifo_reg[0][7]/P0001  & n33167 ;
  assign n34175 = ~n34173 & ~n34174 ;
  assign n34176 = \wishbone_rx_fifo_fifo_reg[0][8]/P0001  & ~n33168 ;
  assign n34177 = \wishbone_rx_fifo_fifo_reg[13][8]/P0001  & n33201 ;
  assign n34178 = \wishbone_rx_fifo_fifo_reg[5][8]/P0001  & n33209 ;
  assign n34179 = ~n34177 & ~n34178 ;
  assign n34180 = \wishbone_rx_fifo_fifo_reg[9][8]/P0001  & n33176 ;
  assign n34181 = \wishbone_rx_fifo_fifo_reg[7][8]/P0001  & n33192 ;
  assign n34182 = ~n34180 & ~n34181 ;
  assign n34183 = n34179 & n34182 ;
  assign n34184 = \wishbone_rx_fifo_fifo_reg[3][8]/P0001  & n33199 ;
  assign n34185 = \wishbone_rx_fifo_fifo_reg[6][8]/P0001  & n33187 ;
  assign n34186 = ~n34184 & ~n34185 ;
  assign n34187 = \wishbone_rx_fifo_fifo_reg[12][8]/P0001  & n33214 ;
  assign n34188 = \wishbone_rx_fifo_fifo_reg[2][8]/P0001  & n33207 ;
  assign n34189 = ~n34187 & ~n34188 ;
  assign n34190 = n34186 & n34189 ;
  assign n34191 = n34183 & n34190 ;
  assign n34192 = \wishbone_rx_fifo_fifo_reg[1][8]/P0001  & n33181 ;
  assign n34193 = \wishbone_rx_fifo_fifo_reg[4][8]/P0001  & n33194 ;
  assign n34194 = \wishbone_rx_fifo_fifo_reg[8][8]/P0001  & n33179 ;
  assign n34195 = ~n34193 & ~n34194 ;
  assign n34196 = ~n34192 & n34195 ;
  assign n34197 = \wishbone_rx_fifo_fifo_reg[14][8]/P0001  & n33212 ;
  assign n34198 = \wishbone_rx_fifo_fifo_reg[10][8]/P0001  & n33189 ;
  assign n34199 = ~n34197 & ~n34198 ;
  assign n34200 = \wishbone_rx_fifo_fifo_reg[11][8]/P0001  & n33203 ;
  assign n34201 = \wishbone_rx_fifo_fifo_reg[15][8]/P0001  & n33172 ;
  assign n34202 = ~n34200 & ~n34201 ;
  assign n34203 = n34199 & n34202 ;
  assign n34204 = n34196 & n34203 ;
  assign n34205 = n34191 & n34204 ;
  assign n34206 = ~n33164 & ~n34205 ;
  assign n34207 = ~n34176 & ~n34206 ;
  assign n34208 = \wishbone_rx_fifo_fifo_reg[14][9]/P0001  & n33212 ;
  assign n34209 = \wishbone_rx_fifo_fifo_reg[9][9]/P0001  & n33176 ;
  assign n34210 = ~n34208 & ~n34209 ;
  assign n34211 = \wishbone_rx_fifo_fifo_reg[6][9]/P0001  & n33187 ;
  assign n34212 = \wishbone_rx_fifo_fifo_reg[15][9]/P0001  & n33172 ;
  assign n34213 = ~n34211 & ~n34212 ;
  assign n34214 = n34210 & n34213 ;
  assign n34215 = \wishbone_rx_fifo_fifo_reg[3][9]/P0001  & n33199 ;
  assign n34216 = ~n33164 & ~n34215 ;
  assign n34217 = \wishbone_rx_fifo_fifo_reg[12][9]/P0001  & n33214 ;
  assign n34218 = \wishbone_rx_fifo_fifo_reg[5][9]/P0001  & n33209 ;
  assign n34219 = ~n34217 & ~n34218 ;
  assign n34220 = n34216 & n34219 ;
  assign n34221 = n34214 & n34220 ;
  assign n34222 = \wishbone_rx_fifo_fifo_reg[1][9]/P0001  & n33181 ;
  assign n34223 = \wishbone_rx_fifo_fifo_reg[10][9]/P0001  & n33189 ;
  assign n34224 = ~n34222 & ~n34223 ;
  assign n34225 = \wishbone_rx_fifo_fifo_reg[8][9]/P0001  & n33179 ;
  assign n34226 = \wishbone_rx_fifo_fifo_reg[4][9]/P0001  & n33194 ;
  assign n34227 = ~n34225 & ~n34226 ;
  assign n34228 = n34224 & n34227 ;
  assign n34229 = \wishbone_rx_fifo_fifo_reg[7][9]/P0001  & n33192 ;
  assign n34230 = \wishbone_rx_fifo_fifo_reg[2][9]/P0001  & n33207 ;
  assign n34231 = ~n34229 & ~n34230 ;
  assign n34232 = \wishbone_rx_fifo_fifo_reg[13][9]/P0001  & n33201 ;
  assign n34233 = \wishbone_rx_fifo_fifo_reg[11][9]/P0001  & n33203 ;
  assign n34234 = ~n34232 & ~n34233 ;
  assign n34235 = n34231 & n34234 ;
  assign n34236 = n34228 & n34235 ;
  assign n34237 = n34221 & n34236 ;
  assign n34238 = ~\wishbone_rx_fifo_fifo_reg[0][9]/P0001  & n33164 ;
  assign n34239 = ~n34237 & ~n34238 ;
  assign n34240 = \wishbone_rx_fifo_fifo_reg[0][9]/P0001  & n33167 ;
  assign n34241 = ~n34239 & ~n34240 ;
  assign n34242 = ~\wishbone_TxAbortPacket_reg/NET0131  & ~\wishbone_TxRetryPacket_reg/NET0131  ;
  assign n34243 = ~\wishbone_tx_fifo_read_pointer_reg[0]/NET0131  & ~\wishbone_tx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n34244 = ~\wishbone_tx_fifo_read_pointer_reg[2]/NET0131  & ~\wishbone_tx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n34245 = n34243 & n34244 ;
  assign n34246 = n34242 & ~n34245 ;
  assign n34247 = \wishbone_tx_fifo_fifo_reg[0][0]/P0001  & ~n34246 ;
  assign n34248 = \wishbone_tx_fifo_read_pointer_reg[0]/NET0131  & ~\wishbone_tx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n34249 = \wishbone_tx_fifo_read_pointer_reg[2]/NET0131  & \wishbone_tx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n34250 = n34248 & n34249 ;
  assign n34251 = \wishbone_tx_fifo_fifo_reg[13][0]/P0001  & n34250 ;
  assign n34252 = ~\wishbone_tx_fifo_read_pointer_reg[0]/NET0131  & \wishbone_tx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n34253 = n34249 & n34252 ;
  assign n34254 = \wishbone_tx_fifo_fifo_reg[14][0]/P0001  & n34253 ;
  assign n34255 = ~n34251 & ~n34254 ;
  assign n34256 = ~\wishbone_tx_fifo_read_pointer_reg[2]/NET0131  & \wishbone_tx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n34257 = n34248 & n34256 ;
  assign n34258 = \wishbone_tx_fifo_fifo_reg[9][0]/P0001  & n34257 ;
  assign n34259 = \wishbone_tx_fifo_read_pointer_reg[0]/NET0131  & \wishbone_tx_fifo_read_pointer_reg[1]/NET0131  ;
  assign n34260 = \wishbone_tx_fifo_read_pointer_reg[2]/NET0131  & ~\wishbone_tx_fifo_read_pointer_reg[3]/NET0131  ;
  assign n34261 = n34259 & n34260 ;
  assign n34262 = \wishbone_tx_fifo_fifo_reg[7][0]/P0001  & n34261 ;
  assign n34263 = ~n34258 & ~n34262 ;
  assign n34264 = n34255 & n34263 ;
  assign n34265 = n34256 & n34259 ;
  assign n34266 = \wishbone_tx_fifo_fifo_reg[11][0]/P0001  & n34265 ;
  assign n34267 = n34248 & n34260 ;
  assign n34268 = \wishbone_tx_fifo_fifo_reg[5][0]/P0001  & n34267 ;
  assign n34269 = ~n34266 & ~n34268 ;
  assign n34270 = n34243 & n34256 ;
  assign n34271 = \wishbone_tx_fifo_fifo_reg[8][0]/P0001  & n34270 ;
  assign n34272 = n34249 & n34259 ;
  assign n34273 = \wishbone_tx_fifo_fifo_reg[15][0]/P0001  & n34272 ;
  assign n34274 = ~n34271 & ~n34273 ;
  assign n34275 = n34269 & n34274 ;
  assign n34276 = n34264 & n34275 ;
  assign n34277 = n34244 & n34252 ;
  assign n34278 = \wishbone_tx_fifo_fifo_reg[2][0]/P0001  & n34277 ;
  assign n34279 = n34243 & n34260 ;
  assign n34280 = \wishbone_tx_fifo_fifo_reg[4][0]/P0001  & n34279 ;
  assign n34281 = n34252 & n34256 ;
  assign n34282 = \wishbone_tx_fifo_fifo_reg[10][0]/P0001  & n34281 ;
  assign n34283 = ~n34280 & ~n34282 ;
  assign n34284 = ~n34278 & n34283 ;
  assign n34285 = n34252 & n34260 ;
  assign n34286 = \wishbone_tx_fifo_fifo_reg[6][0]/P0001  & n34285 ;
  assign n34287 = n34243 & n34249 ;
  assign n34288 = \wishbone_tx_fifo_fifo_reg[12][0]/P0001  & n34287 ;
  assign n34289 = ~n34286 & ~n34288 ;
  assign n34290 = n34244 & n34248 ;
  assign n34291 = \wishbone_tx_fifo_fifo_reg[1][0]/P0001  & n34290 ;
  assign n34292 = n34244 & n34259 ;
  assign n34293 = \wishbone_tx_fifo_fifo_reg[3][0]/P0001  & n34292 ;
  assign n34294 = ~n34291 & ~n34293 ;
  assign n34295 = n34289 & n34294 ;
  assign n34296 = n34284 & n34295 ;
  assign n34297 = n34276 & n34296 ;
  assign n34298 = n34242 & ~n34297 ;
  assign n34299 = ~n34247 & ~n34298 ;
  assign n34300 = \wishbone_tx_fifo_fifo_reg[0][10]/P0001  & ~n34246 ;
  assign n34301 = \wishbone_tx_fifo_fifo_reg[3][10]/P0001  & n34292 ;
  assign n34302 = \wishbone_tx_fifo_fifo_reg[7][10]/P0001  & n34261 ;
  assign n34303 = ~n34301 & ~n34302 ;
  assign n34304 = \wishbone_tx_fifo_fifo_reg[15][10]/P0001  & n34272 ;
  assign n34305 = \wishbone_tx_fifo_fifo_reg[14][10]/P0001  & n34253 ;
  assign n34306 = ~n34304 & ~n34305 ;
  assign n34307 = n34303 & n34306 ;
  assign n34308 = \wishbone_tx_fifo_fifo_reg[2][10]/P0001  & n34277 ;
  assign n34309 = \wishbone_tx_fifo_fifo_reg[13][10]/P0001  & n34250 ;
  assign n34310 = ~n34308 & ~n34309 ;
  assign n34311 = \wishbone_tx_fifo_fifo_reg[5][10]/P0001  & n34267 ;
  assign n34312 = \wishbone_tx_fifo_fifo_reg[11][10]/P0001  & n34265 ;
  assign n34313 = ~n34311 & ~n34312 ;
  assign n34314 = n34310 & n34313 ;
  assign n34315 = n34307 & n34314 ;
  assign n34316 = \wishbone_tx_fifo_fifo_reg[8][10]/P0001  & n34270 ;
  assign n34317 = \wishbone_tx_fifo_fifo_reg[10][10]/P0001  & n34281 ;
  assign n34318 = \wishbone_tx_fifo_fifo_reg[6][10]/P0001  & n34285 ;
  assign n34319 = ~n34317 & ~n34318 ;
  assign n34320 = ~n34316 & n34319 ;
  assign n34321 = \wishbone_tx_fifo_fifo_reg[12][10]/P0001  & n34287 ;
  assign n34322 = \wishbone_tx_fifo_fifo_reg[4][10]/P0001  & n34279 ;
  assign n34323 = ~n34321 & ~n34322 ;
  assign n34324 = \wishbone_tx_fifo_fifo_reg[1][10]/P0001  & n34290 ;
  assign n34325 = \wishbone_tx_fifo_fifo_reg[9][10]/P0001  & n34257 ;
  assign n34326 = ~n34324 & ~n34325 ;
  assign n34327 = n34323 & n34326 ;
  assign n34328 = n34320 & n34327 ;
  assign n34329 = n34315 & n34328 ;
  assign n34330 = n34242 & ~n34329 ;
  assign n34331 = ~n34300 & ~n34330 ;
  assign n34332 = \wishbone_tx_fifo_fifo_reg[0][11]/P0001  & ~n34246 ;
  assign n34333 = \wishbone_tx_fifo_fifo_reg[10][11]/P0001  & n34281 ;
  assign n34334 = \wishbone_tx_fifo_fifo_reg[5][11]/P0001  & n34267 ;
  assign n34335 = ~n34333 & ~n34334 ;
  assign n34336 = \wishbone_tx_fifo_fifo_reg[14][11]/P0001  & n34253 ;
  assign n34337 = \wishbone_tx_fifo_fifo_reg[4][11]/P0001  & n34279 ;
  assign n34338 = ~n34336 & ~n34337 ;
  assign n34339 = n34335 & n34338 ;
  assign n34340 = \wishbone_tx_fifo_fifo_reg[3][11]/P0001  & n34292 ;
  assign n34341 = \wishbone_tx_fifo_fifo_reg[6][11]/P0001  & n34285 ;
  assign n34342 = ~n34340 & ~n34341 ;
  assign n34343 = \wishbone_tx_fifo_fifo_reg[8][11]/P0001  & n34270 ;
  assign n34344 = \wishbone_tx_fifo_fifo_reg[7][11]/P0001  & n34261 ;
  assign n34345 = ~n34343 & ~n34344 ;
  assign n34346 = n34342 & n34345 ;
  assign n34347 = n34339 & n34346 ;
  assign n34348 = \wishbone_tx_fifo_fifo_reg[9][11]/P0001  & n34257 ;
  assign n34349 = \wishbone_tx_fifo_fifo_reg[15][11]/P0001  & n34272 ;
  assign n34350 = \wishbone_tx_fifo_fifo_reg[11][11]/P0001  & n34265 ;
  assign n34351 = ~n34349 & ~n34350 ;
  assign n34352 = ~n34348 & n34351 ;
  assign n34353 = \wishbone_tx_fifo_fifo_reg[1][11]/P0001  & n34290 ;
  assign n34354 = \wishbone_tx_fifo_fifo_reg[13][11]/P0001  & n34250 ;
  assign n34355 = ~n34353 & ~n34354 ;
  assign n34356 = \wishbone_tx_fifo_fifo_reg[2][11]/P0001  & n34277 ;
  assign n34357 = \wishbone_tx_fifo_fifo_reg[12][11]/P0001  & n34287 ;
  assign n34358 = ~n34356 & ~n34357 ;
  assign n34359 = n34355 & n34358 ;
  assign n34360 = n34352 & n34359 ;
  assign n34361 = n34347 & n34360 ;
  assign n34362 = n34242 & ~n34361 ;
  assign n34363 = ~n34332 & ~n34362 ;
  assign n34364 = \wishbone_tx_fifo_fifo_reg[0][12]/P0001  & ~n34246 ;
  assign n34365 = \wishbone_tx_fifo_fifo_reg[5][12]/P0001  & n34267 ;
  assign n34366 = \wishbone_tx_fifo_fifo_reg[9][12]/P0001  & n34257 ;
  assign n34367 = ~n34365 & ~n34366 ;
  assign n34368 = \wishbone_tx_fifo_fifo_reg[10][12]/P0001  & n34281 ;
  assign n34369 = \wishbone_tx_fifo_fifo_reg[13][12]/P0001  & n34250 ;
  assign n34370 = ~n34368 & ~n34369 ;
  assign n34371 = n34367 & n34370 ;
  assign n34372 = \wishbone_tx_fifo_fifo_reg[6][12]/P0001  & n34285 ;
  assign n34373 = \wishbone_tx_fifo_fifo_reg[12][12]/P0001  & n34287 ;
  assign n34374 = ~n34372 & ~n34373 ;
  assign n34375 = \wishbone_tx_fifo_fifo_reg[8][12]/P0001  & n34270 ;
  assign n34376 = \wishbone_tx_fifo_fifo_reg[11][12]/P0001  & n34265 ;
  assign n34377 = ~n34375 & ~n34376 ;
  assign n34378 = n34374 & n34377 ;
  assign n34379 = n34371 & n34378 ;
  assign n34380 = \wishbone_tx_fifo_fifo_reg[2][12]/P0001  & n34277 ;
  assign n34381 = \wishbone_tx_fifo_fifo_reg[7][12]/P0001  & n34261 ;
  assign n34382 = \wishbone_tx_fifo_fifo_reg[14][12]/P0001  & n34253 ;
  assign n34383 = ~n34381 & ~n34382 ;
  assign n34384 = ~n34380 & n34383 ;
  assign n34385 = \wishbone_tx_fifo_fifo_reg[1][12]/P0001  & n34290 ;
  assign n34386 = \wishbone_tx_fifo_fifo_reg[15][12]/P0001  & n34272 ;
  assign n34387 = ~n34385 & ~n34386 ;
  assign n34388 = \wishbone_tx_fifo_fifo_reg[4][12]/P0001  & n34279 ;
  assign n34389 = \wishbone_tx_fifo_fifo_reg[3][12]/P0001  & n34292 ;
  assign n34390 = ~n34388 & ~n34389 ;
  assign n34391 = n34387 & n34390 ;
  assign n34392 = n34384 & n34391 ;
  assign n34393 = n34379 & n34392 ;
  assign n34394 = n34242 & ~n34393 ;
  assign n34395 = ~n34364 & ~n34394 ;
  assign n34396 = \wishbone_tx_fifo_fifo_reg[0][13]/P0001  & ~n34246 ;
  assign n34397 = \wishbone_tx_fifo_fifo_reg[13][13]/P0001  & n34250 ;
  assign n34398 = \wishbone_tx_fifo_fifo_reg[9][13]/P0001  & n34257 ;
  assign n34399 = ~n34397 & ~n34398 ;
  assign n34400 = \wishbone_tx_fifo_fifo_reg[8][13]/P0001  & n34270 ;
  assign n34401 = \wishbone_tx_fifo_fifo_reg[14][13]/P0001  & n34253 ;
  assign n34402 = ~n34400 & ~n34401 ;
  assign n34403 = n34399 & n34402 ;
  assign n34404 = \wishbone_tx_fifo_fifo_reg[3][13]/P0001  & n34292 ;
  assign n34405 = \wishbone_tx_fifo_fifo_reg[5][13]/P0001  & n34267 ;
  assign n34406 = ~n34404 & ~n34405 ;
  assign n34407 = \wishbone_tx_fifo_fifo_reg[15][13]/P0001  & n34272 ;
  assign n34408 = \wishbone_tx_fifo_fifo_reg[2][13]/P0001  & n34277 ;
  assign n34409 = ~n34407 & ~n34408 ;
  assign n34410 = n34406 & n34409 ;
  assign n34411 = n34403 & n34410 ;
  assign n34412 = \wishbone_tx_fifo_fifo_reg[1][13]/P0001  & n34290 ;
  assign n34413 = \wishbone_tx_fifo_fifo_reg[4][13]/P0001  & n34279 ;
  assign n34414 = \wishbone_tx_fifo_fifo_reg[6][13]/P0001  & n34285 ;
  assign n34415 = ~n34413 & ~n34414 ;
  assign n34416 = ~n34412 & n34415 ;
  assign n34417 = \wishbone_tx_fifo_fifo_reg[7][13]/P0001  & n34261 ;
  assign n34418 = \wishbone_tx_fifo_fifo_reg[10][13]/P0001  & n34281 ;
  assign n34419 = ~n34417 & ~n34418 ;
  assign n34420 = \wishbone_tx_fifo_fifo_reg[11][13]/P0001  & n34265 ;
  assign n34421 = \wishbone_tx_fifo_fifo_reg[12][13]/P0001  & n34287 ;
  assign n34422 = ~n34420 & ~n34421 ;
  assign n34423 = n34419 & n34422 ;
  assign n34424 = n34416 & n34423 ;
  assign n34425 = n34411 & n34424 ;
  assign n34426 = n34242 & ~n34425 ;
  assign n34427 = ~n34396 & ~n34426 ;
  assign n34428 = \wishbone_tx_fifo_fifo_reg[0][14]/P0001  & ~n34246 ;
  assign n34429 = \wishbone_tx_fifo_fifo_reg[15][14]/P0001  & n34272 ;
  assign n34430 = \wishbone_tx_fifo_fifo_reg[6][14]/P0001  & n34285 ;
  assign n34431 = ~n34429 & ~n34430 ;
  assign n34432 = \wishbone_tx_fifo_fifo_reg[3][14]/P0001  & n34292 ;
  assign n34433 = \wishbone_tx_fifo_fifo_reg[11][14]/P0001  & n34265 ;
  assign n34434 = ~n34432 & ~n34433 ;
  assign n34435 = n34431 & n34434 ;
  assign n34436 = \wishbone_tx_fifo_fifo_reg[10][14]/P0001  & n34281 ;
  assign n34437 = \wishbone_tx_fifo_fifo_reg[9][14]/P0001  & n34257 ;
  assign n34438 = ~n34436 & ~n34437 ;
  assign n34439 = \wishbone_tx_fifo_fifo_reg[12][14]/P0001  & n34287 ;
  assign n34440 = \wishbone_tx_fifo_fifo_reg[8][14]/P0001  & n34270 ;
  assign n34441 = ~n34439 & ~n34440 ;
  assign n34442 = n34438 & n34441 ;
  assign n34443 = n34435 & n34442 ;
  assign n34444 = \wishbone_tx_fifo_fifo_reg[2][14]/P0001  & n34277 ;
  assign n34445 = \wishbone_tx_fifo_fifo_reg[4][14]/P0001  & n34279 ;
  assign n34446 = \wishbone_tx_fifo_fifo_reg[1][14]/P0001  & n34290 ;
  assign n34447 = ~n34445 & ~n34446 ;
  assign n34448 = ~n34444 & n34447 ;
  assign n34449 = \wishbone_tx_fifo_fifo_reg[5][14]/P0001  & n34267 ;
  assign n34450 = \wishbone_tx_fifo_fifo_reg[14][14]/P0001  & n34253 ;
  assign n34451 = ~n34449 & ~n34450 ;
  assign n34452 = \wishbone_tx_fifo_fifo_reg[7][14]/P0001  & n34261 ;
  assign n34453 = \wishbone_tx_fifo_fifo_reg[13][14]/P0001  & n34250 ;
  assign n34454 = ~n34452 & ~n34453 ;
  assign n34455 = n34451 & n34454 ;
  assign n34456 = n34448 & n34455 ;
  assign n34457 = n34443 & n34456 ;
  assign n34458 = n34242 & ~n34457 ;
  assign n34459 = ~n34428 & ~n34458 ;
  assign n34460 = \wishbone_tx_fifo_fifo_reg[0][15]/P0001  & ~n34246 ;
  assign n34461 = \wishbone_tx_fifo_fifo_reg[2][15]/P0001  & n34277 ;
  assign n34462 = \wishbone_tx_fifo_fifo_reg[7][15]/P0001  & n34261 ;
  assign n34463 = ~n34461 & ~n34462 ;
  assign n34464 = \wishbone_tx_fifo_fifo_reg[15][15]/P0001  & n34272 ;
  assign n34465 = \wishbone_tx_fifo_fifo_reg[14][15]/P0001  & n34253 ;
  assign n34466 = ~n34464 & ~n34465 ;
  assign n34467 = n34463 & n34466 ;
  assign n34468 = \wishbone_tx_fifo_fifo_reg[1][15]/P0001  & n34290 ;
  assign n34469 = \wishbone_tx_fifo_fifo_reg[13][15]/P0001  & n34250 ;
  assign n34470 = ~n34468 & ~n34469 ;
  assign n34471 = \wishbone_tx_fifo_fifo_reg[5][15]/P0001  & n34267 ;
  assign n34472 = \wishbone_tx_fifo_fifo_reg[3][15]/P0001  & n34292 ;
  assign n34473 = ~n34471 & ~n34472 ;
  assign n34474 = n34470 & n34473 ;
  assign n34475 = n34467 & n34474 ;
  assign n34476 = \wishbone_tx_fifo_fifo_reg[8][15]/P0001  & n34270 ;
  assign n34477 = \wishbone_tx_fifo_fifo_reg[10][15]/P0001  & n34281 ;
  assign n34478 = \wishbone_tx_fifo_fifo_reg[6][15]/P0001  & n34285 ;
  assign n34479 = ~n34477 & ~n34478 ;
  assign n34480 = ~n34476 & n34479 ;
  assign n34481 = \wishbone_tx_fifo_fifo_reg[12][15]/P0001  & n34287 ;
  assign n34482 = \wishbone_tx_fifo_fifo_reg[4][15]/P0001  & n34279 ;
  assign n34483 = ~n34481 & ~n34482 ;
  assign n34484 = \wishbone_tx_fifo_fifo_reg[11][15]/P0001  & n34265 ;
  assign n34485 = \wishbone_tx_fifo_fifo_reg[9][15]/P0001  & n34257 ;
  assign n34486 = ~n34484 & ~n34485 ;
  assign n34487 = n34483 & n34486 ;
  assign n34488 = n34480 & n34487 ;
  assign n34489 = n34475 & n34488 ;
  assign n34490 = n34242 & ~n34489 ;
  assign n34491 = ~n34460 & ~n34490 ;
  assign n34492 = \wishbone_tx_fifo_fifo_reg[0][16]/P0001  & ~n34246 ;
  assign n34493 = \wishbone_tx_fifo_fifo_reg[13][16]/P0001  & n34250 ;
  assign n34494 = \wishbone_tx_fifo_fifo_reg[6][16]/P0001  & n34285 ;
  assign n34495 = ~n34493 & ~n34494 ;
  assign n34496 = \wishbone_tx_fifo_fifo_reg[8][16]/P0001  & n34270 ;
  assign n34497 = \wishbone_tx_fifo_fifo_reg[14][16]/P0001  & n34253 ;
  assign n34498 = ~n34496 & ~n34497 ;
  assign n34499 = n34495 & n34498 ;
  assign n34500 = \wishbone_tx_fifo_fifo_reg[2][16]/P0001  & n34277 ;
  assign n34501 = \wishbone_tx_fifo_fifo_reg[5][16]/P0001  & n34267 ;
  assign n34502 = ~n34500 & ~n34501 ;
  assign n34503 = \wishbone_tx_fifo_fifo_reg[15][16]/P0001  & n34272 ;
  assign n34504 = \wishbone_tx_fifo_fifo_reg[1][16]/P0001  & n34290 ;
  assign n34505 = ~n34503 & ~n34504 ;
  assign n34506 = n34502 & n34505 ;
  assign n34507 = n34499 & n34506 ;
  assign n34508 = \wishbone_tx_fifo_fifo_reg[11][16]/P0001  & n34265 ;
  assign n34509 = \wishbone_tx_fifo_fifo_reg[4][16]/P0001  & n34279 ;
  assign n34510 = \wishbone_tx_fifo_fifo_reg[9][16]/P0001  & n34257 ;
  assign n34511 = ~n34509 & ~n34510 ;
  assign n34512 = ~n34508 & n34511 ;
  assign n34513 = \wishbone_tx_fifo_fifo_reg[7][16]/P0001  & n34261 ;
  assign n34514 = \wishbone_tx_fifo_fifo_reg[10][16]/P0001  & n34281 ;
  assign n34515 = ~n34513 & ~n34514 ;
  assign n34516 = \wishbone_tx_fifo_fifo_reg[3][16]/P0001  & n34292 ;
  assign n34517 = \wishbone_tx_fifo_fifo_reg[12][16]/P0001  & n34287 ;
  assign n34518 = ~n34516 & ~n34517 ;
  assign n34519 = n34515 & n34518 ;
  assign n34520 = n34512 & n34519 ;
  assign n34521 = n34507 & n34520 ;
  assign n34522 = n34242 & ~n34521 ;
  assign n34523 = ~n34492 & ~n34522 ;
  assign n34524 = \wishbone_tx_fifo_fifo_reg[0][17]/P0001  & ~n34246 ;
  assign n34525 = \wishbone_tx_fifo_fifo_reg[2][17]/P0001  & n34277 ;
  assign n34526 = \wishbone_tx_fifo_fifo_reg[7][17]/P0001  & n34261 ;
  assign n34527 = ~n34525 & ~n34526 ;
  assign n34528 = \wishbone_tx_fifo_fifo_reg[15][17]/P0001  & n34272 ;
  assign n34529 = \wishbone_tx_fifo_fifo_reg[14][17]/P0001  & n34253 ;
  assign n34530 = ~n34528 & ~n34529 ;
  assign n34531 = n34527 & n34530 ;
  assign n34532 = \wishbone_tx_fifo_fifo_reg[1][17]/P0001  & n34290 ;
  assign n34533 = \wishbone_tx_fifo_fifo_reg[13][17]/P0001  & n34250 ;
  assign n34534 = ~n34532 & ~n34533 ;
  assign n34535 = \wishbone_tx_fifo_fifo_reg[5][17]/P0001  & n34267 ;
  assign n34536 = \wishbone_tx_fifo_fifo_reg[3][17]/P0001  & n34292 ;
  assign n34537 = ~n34535 & ~n34536 ;
  assign n34538 = n34534 & n34537 ;
  assign n34539 = n34531 & n34538 ;
  assign n34540 = \wishbone_tx_fifo_fifo_reg[8][17]/P0001  & n34270 ;
  assign n34541 = \wishbone_tx_fifo_fifo_reg[10][17]/P0001  & n34281 ;
  assign n34542 = \wishbone_tx_fifo_fifo_reg[6][17]/P0001  & n34285 ;
  assign n34543 = ~n34541 & ~n34542 ;
  assign n34544 = ~n34540 & n34543 ;
  assign n34545 = \wishbone_tx_fifo_fifo_reg[12][17]/P0001  & n34287 ;
  assign n34546 = \wishbone_tx_fifo_fifo_reg[4][17]/P0001  & n34279 ;
  assign n34547 = ~n34545 & ~n34546 ;
  assign n34548 = \wishbone_tx_fifo_fifo_reg[11][17]/P0001  & n34265 ;
  assign n34549 = \wishbone_tx_fifo_fifo_reg[9][17]/P0001  & n34257 ;
  assign n34550 = ~n34548 & ~n34549 ;
  assign n34551 = n34547 & n34550 ;
  assign n34552 = n34544 & n34551 ;
  assign n34553 = n34539 & n34552 ;
  assign n34554 = n34242 & ~n34553 ;
  assign n34555 = ~n34524 & ~n34554 ;
  assign n34556 = \wishbone_tx_fifo_fifo_reg[0][18]/P0001  & ~n34246 ;
  assign n34557 = \wishbone_tx_fifo_fifo_reg[2][18]/P0001  & n34277 ;
  assign n34558 = \wishbone_tx_fifo_fifo_reg[5][18]/P0001  & n34267 ;
  assign n34559 = ~n34557 & ~n34558 ;
  assign n34560 = \wishbone_tx_fifo_fifo_reg[14][18]/P0001  & n34253 ;
  assign n34561 = \wishbone_tx_fifo_fifo_reg[12][18]/P0001  & n34287 ;
  assign n34562 = ~n34560 & ~n34561 ;
  assign n34563 = n34559 & n34562 ;
  assign n34564 = \wishbone_tx_fifo_fifo_reg[10][18]/P0001  & n34281 ;
  assign n34565 = \wishbone_tx_fifo_fifo_reg[4][18]/P0001  & n34279 ;
  assign n34566 = ~n34564 & ~n34565 ;
  assign n34567 = \wishbone_tx_fifo_fifo_reg[3][18]/P0001  & n34292 ;
  assign n34568 = \wishbone_tx_fifo_fifo_reg[11][18]/P0001  & n34265 ;
  assign n34569 = ~n34567 & ~n34568 ;
  assign n34570 = n34566 & n34569 ;
  assign n34571 = n34563 & n34570 ;
  assign n34572 = \wishbone_tx_fifo_fifo_reg[8][18]/P0001  & n34270 ;
  assign n34573 = \wishbone_tx_fifo_fifo_reg[6][18]/P0001  & n34285 ;
  assign n34574 = \wishbone_tx_fifo_fifo_reg[7][18]/P0001  & n34261 ;
  assign n34575 = ~n34573 & ~n34574 ;
  assign n34576 = ~n34572 & n34575 ;
  assign n34577 = \wishbone_tx_fifo_fifo_reg[15][18]/P0001  & n34272 ;
  assign n34578 = \wishbone_tx_fifo_fifo_reg[1][18]/P0001  & n34290 ;
  assign n34579 = ~n34577 & ~n34578 ;
  assign n34580 = \wishbone_tx_fifo_fifo_reg[13][18]/P0001  & n34250 ;
  assign n34581 = \wishbone_tx_fifo_fifo_reg[9][18]/P0001  & n34257 ;
  assign n34582 = ~n34580 & ~n34581 ;
  assign n34583 = n34579 & n34582 ;
  assign n34584 = n34576 & n34583 ;
  assign n34585 = n34571 & n34584 ;
  assign n34586 = n34242 & ~n34585 ;
  assign n34587 = ~n34556 & ~n34586 ;
  assign n34588 = \wishbone_tx_fifo_fifo_reg[0][19]/P0001  & ~n34246 ;
  assign n34589 = \wishbone_tx_fifo_fifo_reg[13][19]/P0001  & n34250 ;
  assign n34590 = \wishbone_tx_fifo_fifo_reg[5][19]/P0001  & n34267 ;
  assign n34591 = ~n34589 & ~n34590 ;
  assign n34592 = \wishbone_tx_fifo_fifo_reg[9][19]/P0001  & n34257 ;
  assign n34593 = \wishbone_tx_fifo_fifo_reg[7][19]/P0001  & n34261 ;
  assign n34594 = ~n34592 & ~n34593 ;
  assign n34595 = n34591 & n34594 ;
  assign n34596 = \wishbone_tx_fifo_fifo_reg[3][19]/P0001  & n34292 ;
  assign n34597 = \wishbone_tx_fifo_fifo_reg[6][19]/P0001  & n34285 ;
  assign n34598 = ~n34596 & ~n34597 ;
  assign n34599 = \wishbone_tx_fifo_fifo_reg[12][19]/P0001  & n34287 ;
  assign n34600 = \wishbone_tx_fifo_fifo_reg[2][19]/P0001  & n34277 ;
  assign n34601 = ~n34599 & ~n34600 ;
  assign n34602 = n34598 & n34601 ;
  assign n34603 = n34595 & n34602 ;
  assign n34604 = \wishbone_tx_fifo_fifo_reg[1][19]/P0001  & n34290 ;
  assign n34605 = \wishbone_tx_fifo_fifo_reg[4][19]/P0001  & n34279 ;
  assign n34606 = \wishbone_tx_fifo_fifo_reg[8][19]/P0001  & n34270 ;
  assign n34607 = ~n34605 & ~n34606 ;
  assign n34608 = ~n34604 & n34607 ;
  assign n34609 = \wishbone_tx_fifo_fifo_reg[14][19]/P0001  & n34253 ;
  assign n34610 = \wishbone_tx_fifo_fifo_reg[10][19]/P0001  & n34281 ;
  assign n34611 = ~n34609 & ~n34610 ;
  assign n34612 = \wishbone_tx_fifo_fifo_reg[11][19]/P0001  & n34265 ;
  assign n34613 = \wishbone_tx_fifo_fifo_reg[15][19]/P0001  & n34272 ;
  assign n34614 = ~n34612 & ~n34613 ;
  assign n34615 = n34611 & n34614 ;
  assign n34616 = n34608 & n34615 ;
  assign n34617 = n34603 & n34616 ;
  assign n34618 = n34242 & ~n34617 ;
  assign n34619 = ~n34588 & ~n34618 ;
  assign n34620 = \wishbone_tx_fifo_fifo_reg[0][1]/P0001  & ~n34246 ;
  assign n34621 = \wishbone_tx_fifo_fifo_reg[9][1]/P0001  & n34257 ;
  assign n34622 = \wishbone_tx_fifo_fifo_reg[6][1]/P0001  & n34285 ;
  assign n34623 = ~n34621 & ~n34622 ;
  assign n34624 = \wishbone_tx_fifo_fifo_reg[2][1]/P0001  & n34277 ;
  assign n34625 = \wishbone_tx_fifo_fifo_reg[1][1]/P0001  & n34290 ;
  assign n34626 = ~n34624 & ~n34625 ;
  assign n34627 = n34623 & n34626 ;
  assign n34628 = \wishbone_tx_fifo_fifo_reg[5][1]/P0001  & n34267 ;
  assign n34629 = \wishbone_tx_fifo_fifo_reg[14][1]/P0001  & n34253 ;
  assign n34630 = ~n34628 & ~n34629 ;
  assign n34631 = \wishbone_tx_fifo_fifo_reg[12][1]/P0001  & n34287 ;
  assign n34632 = \wishbone_tx_fifo_fifo_reg[3][1]/P0001  & n34292 ;
  assign n34633 = ~n34631 & ~n34632 ;
  assign n34634 = n34630 & n34633 ;
  assign n34635 = n34627 & n34634 ;
  assign n34636 = \wishbone_tx_fifo_fifo_reg[7][1]/P0001  & n34261 ;
  assign n34637 = \wishbone_tx_fifo_fifo_reg[10][1]/P0001  & n34281 ;
  assign n34638 = \wishbone_tx_fifo_fifo_reg[8][1]/P0001  & n34270 ;
  assign n34639 = ~n34637 & ~n34638 ;
  assign n34640 = ~n34636 & n34639 ;
  assign n34641 = \wishbone_tx_fifo_fifo_reg[4][1]/P0001  & n34279 ;
  assign n34642 = \wishbone_tx_fifo_fifo_reg[11][1]/P0001  & n34265 ;
  assign n34643 = ~n34641 & ~n34642 ;
  assign n34644 = \wishbone_tx_fifo_fifo_reg[15][1]/P0001  & n34272 ;
  assign n34645 = \wishbone_tx_fifo_fifo_reg[13][1]/P0001  & n34250 ;
  assign n34646 = ~n34644 & ~n34645 ;
  assign n34647 = n34643 & n34646 ;
  assign n34648 = n34640 & n34647 ;
  assign n34649 = n34635 & n34648 ;
  assign n34650 = n34242 & ~n34649 ;
  assign n34651 = ~n34620 & ~n34650 ;
  assign n34652 = \wishbone_tx_fifo_fifo_reg[0][20]/P0001  & ~n34246 ;
  assign n34653 = \wishbone_tx_fifo_fifo_reg[15][20]/P0001  & n34272 ;
  assign n34654 = \wishbone_tx_fifo_fifo_reg[9][20]/P0001  & n34257 ;
  assign n34655 = ~n34653 & ~n34654 ;
  assign n34656 = \wishbone_tx_fifo_fifo_reg[8][20]/P0001  & n34270 ;
  assign n34657 = \wishbone_tx_fifo_fifo_reg[3][20]/P0001  & n34292 ;
  assign n34658 = ~n34656 & ~n34657 ;
  assign n34659 = n34655 & n34658 ;
  assign n34660 = \wishbone_tx_fifo_fifo_reg[6][20]/P0001  & n34285 ;
  assign n34661 = \wishbone_tx_fifo_fifo_reg[10][20]/P0001  & n34281 ;
  assign n34662 = ~n34660 & ~n34661 ;
  assign n34663 = \wishbone_tx_fifo_fifo_reg[7][20]/P0001  & n34261 ;
  assign n34664 = \wishbone_tx_fifo_fifo_reg[4][20]/P0001  & n34279 ;
  assign n34665 = ~n34663 & ~n34664 ;
  assign n34666 = n34662 & n34665 ;
  assign n34667 = n34659 & n34666 ;
  assign n34668 = \wishbone_tx_fifo_fifo_reg[1][20]/P0001  & n34290 ;
  assign n34669 = \wishbone_tx_fifo_fifo_reg[13][20]/P0001  & n34250 ;
  assign n34670 = \wishbone_tx_fifo_fifo_reg[2][20]/P0001  & n34277 ;
  assign n34671 = ~n34669 & ~n34670 ;
  assign n34672 = ~n34668 & n34671 ;
  assign n34673 = \wishbone_tx_fifo_fifo_reg[11][20]/P0001  & n34265 ;
  assign n34674 = \wishbone_tx_fifo_fifo_reg[5][20]/P0001  & n34267 ;
  assign n34675 = ~n34673 & ~n34674 ;
  assign n34676 = \wishbone_tx_fifo_fifo_reg[14][20]/P0001  & n34253 ;
  assign n34677 = \wishbone_tx_fifo_fifo_reg[12][20]/P0001  & n34287 ;
  assign n34678 = ~n34676 & ~n34677 ;
  assign n34679 = n34675 & n34678 ;
  assign n34680 = n34672 & n34679 ;
  assign n34681 = n34667 & n34680 ;
  assign n34682 = n34242 & ~n34681 ;
  assign n34683 = ~n34652 & ~n34682 ;
  assign n34684 = \wishbone_tx_fifo_fifo_reg[0][21]/P0001  & ~n34246 ;
  assign n34685 = \wishbone_tx_fifo_fifo_reg[13][21]/P0001  & n34250 ;
  assign n34686 = \wishbone_tx_fifo_fifo_reg[14][21]/P0001  & n34253 ;
  assign n34687 = ~n34685 & ~n34686 ;
  assign n34688 = \wishbone_tx_fifo_fifo_reg[9][21]/P0001  & n34257 ;
  assign n34689 = \wishbone_tx_fifo_fifo_reg[7][21]/P0001  & n34261 ;
  assign n34690 = ~n34688 & ~n34689 ;
  assign n34691 = n34687 & n34690 ;
  assign n34692 = \wishbone_tx_fifo_fifo_reg[11][21]/P0001  & n34265 ;
  assign n34693 = \wishbone_tx_fifo_fifo_reg[5][21]/P0001  & n34267 ;
  assign n34694 = ~n34692 & ~n34693 ;
  assign n34695 = \wishbone_tx_fifo_fifo_reg[8][21]/P0001  & n34270 ;
  assign n34696 = \wishbone_tx_fifo_fifo_reg[15][21]/P0001  & n34272 ;
  assign n34697 = ~n34695 & ~n34696 ;
  assign n34698 = n34694 & n34697 ;
  assign n34699 = n34691 & n34698 ;
  assign n34700 = \wishbone_tx_fifo_fifo_reg[2][21]/P0001  & n34277 ;
  assign n34701 = \wishbone_tx_fifo_fifo_reg[4][21]/P0001  & n34279 ;
  assign n34702 = \wishbone_tx_fifo_fifo_reg[10][21]/P0001  & n34281 ;
  assign n34703 = ~n34701 & ~n34702 ;
  assign n34704 = ~n34700 & n34703 ;
  assign n34705 = \wishbone_tx_fifo_fifo_reg[6][21]/P0001  & n34285 ;
  assign n34706 = \wishbone_tx_fifo_fifo_reg[12][21]/P0001  & n34287 ;
  assign n34707 = ~n34705 & ~n34706 ;
  assign n34708 = \wishbone_tx_fifo_fifo_reg[1][21]/P0001  & n34290 ;
  assign n34709 = \wishbone_tx_fifo_fifo_reg[3][21]/P0001  & n34292 ;
  assign n34710 = ~n34708 & ~n34709 ;
  assign n34711 = n34707 & n34710 ;
  assign n34712 = n34704 & n34711 ;
  assign n34713 = n34699 & n34712 ;
  assign n34714 = n34242 & ~n34713 ;
  assign n34715 = ~n34684 & ~n34714 ;
  assign n34716 = \wishbone_tx_fifo_fifo_reg[0][22]/P0001  & ~n34246 ;
  assign n34717 = \wishbone_tx_fifo_fifo_reg[13][22]/P0001  & n34250 ;
  assign n34718 = \wishbone_tx_fifo_fifo_reg[12][22]/P0001  & n34287 ;
  assign n34719 = ~n34717 & ~n34718 ;
  assign n34720 = \wishbone_tx_fifo_fifo_reg[9][22]/P0001  & n34257 ;
  assign n34721 = \wishbone_tx_fifo_fifo_reg[7][22]/P0001  & n34261 ;
  assign n34722 = ~n34720 & ~n34721 ;
  assign n34723 = n34719 & n34722 ;
  assign n34724 = \wishbone_tx_fifo_fifo_reg[2][22]/P0001  & n34277 ;
  assign n34725 = \wishbone_tx_fifo_fifo_reg[6][22]/P0001  & n34285 ;
  assign n34726 = ~n34724 & ~n34725 ;
  assign n34727 = \wishbone_tx_fifo_fifo_reg[14][22]/P0001  & n34253 ;
  assign n34728 = \wishbone_tx_fifo_fifo_reg[1][22]/P0001  & n34290 ;
  assign n34729 = ~n34727 & ~n34728 ;
  assign n34730 = n34726 & n34729 ;
  assign n34731 = n34723 & n34730 ;
  assign n34732 = \wishbone_tx_fifo_fifo_reg[11][22]/P0001  & n34265 ;
  assign n34733 = \wishbone_tx_fifo_fifo_reg[4][22]/P0001  & n34279 ;
  assign n34734 = \wishbone_tx_fifo_fifo_reg[8][22]/P0001  & n34270 ;
  assign n34735 = ~n34733 & ~n34734 ;
  assign n34736 = ~n34732 & n34735 ;
  assign n34737 = \wishbone_tx_fifo_fifo_reg[5][22]/P0001  & n34267 ;
  assign n34738 = \wishbone_tx_fifo_fifo_reg[10][22]/P0001  & n34281 ;
  assign n34739 = ~n34737 & ~n34738 ;
  assign n34740 = \wishbone_tx_fifo_fifo_reg[3][22]/P0001  & n34292 ;
  assign n34741 = \wishbone_tx_fifo_fifo_reg[15][22]/P0001  & n34272 ;
  assign n34742 = ~n34740 & ~n34741 ;
  assign n34743 = n34739 & n34742 ;
  assign n34744 = n34736 & n34743 ;
  assign n34745 = n34731 & n34744 ;
  assign n34746 = n34242 & ~n34745 ;
  assign n34747 = ~n34716 & ~n34746 ;
  assign n34748 = \wishbone_tx_fifo_fifo_reg[0][23]/P0001  & ~n34246 ;
  assign n34749 = \wishbone_tx_fifo_fifo_reg[10][23]/P0001  & n34281 ;
  assign n34750 = \wishbone_tx_fifo_fifo_reg[5][23]/P0001  & n34267 ;
  assign n34751 = ~n34749 & ~n34750 ;
  assign n34752 = \wishbone_tx_fifo_fifo_reg[14][23]/P0001  & n34253 ;
  assign n34753 = \wishbone_tx_fifo_fifo_reg[4][23]/P0001  & n34279 ;
  assign n34754 = ~n34752 & ~n34753 ;
  assign n34755 = n34751 & n34754 ;
  assign n34756 = \wishbone_tx_fifo_fifo_reg[2][23]/P0001  & n34277 ;
  assign n34757 = \wishbone_tx_fifo_fifo_reg[6][23]/P0001  & n34285 ;
  assign n34758 = ~n34756 & ~n34757 ;
  assign n34759 = \wishbone_tx_fifo_fifo_reg[8][23]/P0001  & n34270 ;
  assign n34760 = \wishbone_tx_fifo_fifo_reg[7][23]/P0001  & n34261 ;
  assign n34761 = ~n34759 & ~n34760 ;
  assign n34762 = n34758 & n34761 ;
  assign n34763 = n34755 & n34762 ;
  assign n34764 = \wishbone_tx_fifo_fifo_reg[9][23]/P0001  & n34257 ;
  assign n34765 = \wishbone_tx_fifo_fifo_reg[15][23]/P0001  & n34272 ;
  assign n34766 = \wishbone_tx_fifo_fifo_reg[3][23]/P0001  & n34292 ;
  assign n34767 = ~n34765 & ~n34766 ;
  assign n34768 = ~n34764 & n34767 ;
  assign n34769 = \wishbone_tx_fifo_fifo_reg[11][23]/P0001  & n34265 ;
  assign n34770 = \wishbone_tx_fifo_fifo_reg[13][23]/P0001  & n34250 ;
  assign n34771 = ~n34769 & ~n34770 ;
  assign n34772 = \wishbone_tx_fifo_fifo_reg[1][23]/P0001  & n34290 ;
  assign n34773 = \wishbone_tx_fifo_fifo_reg[12][23]/P0001  & n34287 ;
  assign n34774 = ~n34772 & ~n34773 ;
  assign n34775 = n34771 & n34774 ;
  assign n34776 = n34768 & n34775 ;
  assign n34777 = n34763 & n34776 ;
  assign n34778 = n34242 & ~n34777 ;
  assign n34779 = ~n34748 & ~n34778 ;
  assign n34780 = \wishbone_tx_fifo_fifo_reg[0][24]/P0001  & ~n34246 ;
  assign n34781 = \wishbone_tx_fifo_fifo_reg[5][24]/P0001  & n34267 ;
  assign n34782 = \wishbone_tx_fifo_fifo_reg[3][24]/P0001  & n34292 ;
  assign n34783 = ~n34781 & ~n34782 ;
  assign n34784 = \wishbone_tx_fifo_fifo_reg[2][24]/P0001  & n34277 ;
  assign n34785 = \wishbone_tx_fifo_fifo_reg[4][24]/P0001  & n34279 ;
  assign n34786 = ~n34784 & ~n34785 ;
  assign n34787 = n34783 & n34786 ;
  assign n34788 = \wishbone_tx_fifo_fifo_reg[8][24]/P0001  & n34270 ;
  assign n34789 = \wishbone_tx_fifo_fifo_reg[7][24]/P0001  & n34261 ;
  assign n34790 = ~n34788 & ~n34789 ;
  assign n34791 = \wishbone_tx_fifo_fifo_reg[10][24]/P0001  & n34281 ;
  assign n34792 = \wishbone_tx_fifo_fifo_reg[12][24]/P0001  & n34287 ;
  assign n34793 = ~n34791 & ~n34792 ;
  assign n34794 = n34790 & n34793 ;
  assign n34795 = n34787 & n34794 ;
  assign n34796 = \wishbone_tx_fifo_fifo_reg[1][24]/P0001  & n34290 ;
  assign n34797 = \wishbone_tx_fifo_fifo_reg[9][24]/P0001  & n34257 ;
  assign n34798 = \wishbone_tx_fifo_fifo_reg[11][24]/P0001  & n34265 ;
  assign n34799 = ~n34797 & ~n34798 ;
  assign n34800 = ~n34796 & n34799 ;
  assign n34801 = \wishbone_tx_fifo_fifo_reg[13][24]/P0001  & n34250 ;
  assign n34802 = \wishbone_tx_fifo_fifo_reg[6][24]/P0001  & n34285 ;
  assign n34803 = ~n34801 & ~n34802 ;
  assign n34804 = \wishbone_tx_fifo_fifo_reg[14][24]/P0001  & n34253 ;
  assign n34805 = \wishbone_tx_fifo_fifo_reg[15][24]/P0001  & n34272 ;
  assign n34806 = ~n34804 & ~n34805 ;
  assign n34807 = n34803 & n34806 ;
  assign n34808 = n34800 & n34807 ;
  assign n34809 = n34795 & n34808 ;
  assign n34810 = n34242 & ~n34809 ;
  assign n34811 = ~n34780 & ~n34810 ;
  assign n34812 = \wishbone_tx_fifo_fifo_reg[0][25]/P0001  & ~n34246 ;
  assign n34813 = \wishbone_tx_fifo_fifo_reg[13][25]/P0001  & n34250 ;
  assign n34814 = \wishbone_tx_fifo_fifo_reg[3][25]/P0001  & n34292 ;
  assign n34815 = ~n34813 & ~n34814 ;
  assign n34816 = \wishbone_tx_fifo_fifo_reg[11][25]/P0001  & n34265 ;
  assign n34817 = \wishbone_tx_fifo_fifo_reg[5][25]/P0001  & n34267 ;
  assign n34818 = ~n34816 & ~n34817 ;
  assign n34819 = n34815 & n34818 ;
  assign n34820 = \wishbone_tx_fifo_fifo_reg[6][25]/P0001  & n34285 ;
  assign n34821 = \wishbone_tx_fifo_fifo_reg[10][25]/P0001  & n34281 ;
  assign n34822 = ~n34820 & ~n34821 ;
  assign n34823 = \wishbone_tx_fifo_fifo_reg[12][25]/P0001  & n34287 ;
  assign n34824 = \wishbone_tx_fifo_fifo_reg[14][25]/P0001  & n34253 ;
  assign n34825 = ~n34823 & ~n34824 ;
  assign n34826 = n34822 & n34825 ;
  assign n34827 = n34819 & n34826 ;
  assign n34828 = \wishbone_tx_fifo_fifo_reg[15][25]/P0001  & n34272 ;
  assign n34829 = \wishbone_tx_fifo_fifo_reg[2][25]/P0001  & n34277 ;
  assign n34830 = \wishbone_tx_fifo_fifo_reg[9][25]/P0001  & n34257 ;
  assign n34831 = ~n34829 & ~n34830 ;
  assign n34832 = ~n34828 & n34831 ;
  assign n34833 = \wishbone_tx_fifo_fifo_reg[1][25]/P0001  & n34290 ;
  assign n34834 = \wishbone_tx_fifo_fifo_reg[4][25]/P0001  & n34279 ;
  assign n34835 = ~n34833 & ~n34834 ;
  assign n34836 = \wishbone_tx_fifo_fifo_reg[8][25]/P0001  & n34270 ;
  assign n34837 = \wishbone_tx_fifo_fifo_reg[7][25]/P0001  & n34261 ;
  assign n34838 = ~n34836 & ~n34837 ;
  assign n34839 = n34835 & n34838 ;
  assign n34840 = n34832 & n34839 ;
  assign n34841 = n34827 & n34840 ;
  assign n34842 = n34242 & ~n34841 ;
  assign n34843 = ~n34812 & ~n34842 ;
  assign n34844 = \wishbone_tx_fifo_fifo_reg[0][26]/P0001  & ~n34246 ;
  assign n34845 = \wishbone_tx_fifo_fifo_reg[6][26]/P0001  & n34285 ;
  assign n34846 = \wishbone_tx_fifo_fifo_reg[9][26]/P0001  & n34257 ;
  assign n34847 = ~n34845 & ~n34846 ;
  assign n34848 = \wishbone_tx_fifo_fifo_reg[2][26]/P0001  & n34277 ;
  assign n34849 = \wishbone_tx_fifo_fifo_reg[1][26]/P0001  & n34290 ;
  assign n34850 = ~n34848 & ~n34849 ;
  assign n34851 = n34847 & n34850 ;
  assign n34852 = \wishbone_tx_fifo_fifo_reg[5][26]/P0001  & n34267 ;
  assign n34853 = \wishbone_tx_fifo_fifo_reg[14][26]/P0001  & n34253 ;
  assign n34854 = ~n34852 & ~n34853 ;
  assign n34855 = \wishbone_tx_fifo_fifo_reg[12][26]/P0001  & n34287 ;
  assign n34856 = \wishbone_tx_fifo_fifo_reg[3][26]/P0001  & n34292 ;
  assign n34857 = ~n34855 & ~n34856 ;
  assign n34858 = n34854 & n34857 ;
  assign n34859 = n34851 & n34858 ;
  assign n34860 = \wishbone_tx_fifo_fifo_reg[7][26]/P0001  & n34261 ;
  assign n34861 = \wishbone_tx_fifo_fifo_reg[10][26]/P0001  & n34281 ;
  assign n34862 = \wishbone_tx_fifo_fifo_reg[8][26]/P0001  & n34270 ;
  assign n34863 = ~n34861 & ~n34862 ;
  assign n34864 = ~n34860 & n34863 ;
  assign n34865 = \wishbone_tx_fifo_fifo_reg[4][26]/P0001  & n34279 ;
  assign n34866 = \wishbone_tx_fifo_fifo_reg[11][26]/P0001  & n34265 ;
  assign n34867 = ~n34865 & ~n34866 ;
  assign n34868 = \wishbone_tx_fifo_fifo_reg[15][26]/P0001  & n34272 ;
  assign n34869 = \wishbone_tx_fifo_fifo_reg[13][26]/P0001  & n34250 ;
  assign n34870 = ~n34868 & ~n34869 ;
  assign n34871 = n34867 & n34870 ;
  assign n34872 = n34864 & n34871 ;
  assign n34873 = n34859 & n34872 ;
  assign n34874 = n34242 & ~n34873 ;
  assign n34875 = ~n34844 & ~n34874 ;
  assign n34876 = \wishbone_tx_fifo_fifo_reg[0][27]/P0001  & ~n34246 ;
  assign n34877 = \wishbone_tx_fifo_fifo_reg[1][27]/P0001  & n34290 ;
  assign n34878 = \wishbone_tx_fifo_fifo_reg[12][27]/P0001  & n34287 ;
  assign n34879 = ~n34877 & ~n34878 ;
  assign n34880 = \wishbone_tx_fifo_fifo_reg[9][27]/P0001  & n34257 ;
  assign n34881 = \wishbone_tx_fifo_fifo_reg[11][27]/P0001  & n34265 ;
  assign n34882 = ~n34880 & ~n34881 ;
  assign n34883 = n34879 & n34882 ;
  assign n34884 = \wishbone_tx_fifo_fifo_reg[6][27]/P0001  & n34285 ;
  assign n34885 = \wishbone_tx_fifo_fifo_reg[10][27]/P0001  & n34281 ;
  assign n34886 = ~n34884 & ~n34885 ;
  assign n34887 = \wishbone_tx_fifo_fifo_reg[5][27]/P0001  & n34267 ;
  assign n34888 = \wishbone_tx_fifo_fifo_reg[7][27]/P0001  & n34261 ;
  assign n34889 = ~n34887 & ~n34888 ;
  assign n34890 = n34886 & n34889 ;
  assign n34891 = n34883 & n34890 ;
  assign n34892 = \wishbone_tx_fifo_fifo_reg[8][27]/P0001  & n34270 ;
  assign n34893 = \wishbone_tx_fifo_fifo_reg[15][27]/P0001  & n34272 ;
  assign n34894 = \wishbone_tx_fifo_fifo_reg[2][27]/P0001  & n34277 ;
  assign n34895 = ~n34893 & ~n34894 ;
  assign n34896 = ~n34892 & n34895 ;
  assign n34897 = \wishbone_tx_fifo_fifo_reg[4][27]/P0001  & n34279 ;
  assign n34898 = \wishbone_tx_fifo_fifo_reg[3][27]/P0001  & n34292 ;
  assign n34899 = ~n34897 & ~n34898 ;
  assign n34900 = \wishbone_tx_fifo_fifo_reg[13][27]/P0001  & n34250 ;
  assign n34901 = \wishbone_tx_fifo_fifo_reg[14][27]/P0001  & n34253 ;
  assign n34902 = ~n34900 & ~n34901 ;
  assign n34903 = n34899 & n34902 ;
  assign n34904 = n34896 & n34903 ;
  assign n34905 = n34891 & n34904 ;
  assign n34906 = n34242 & ~n34905 ;
  assign n34907 = ~n34876 & ~n34906 ;
  assign n34908 = \wishbone_tx_fifo_fifo_reg[0][28]/P0001  & ~n34246 ;
  assign n34909 = \wishbone_tx_fifo_fifo_reg[14][28]/P0001  & n34253 ;
  assign n34910 = \wishbone_tx_fifo_fifo_reg[6][28]/P0001  & n34285 ;
  assign n34911 = ~n34909 & ~n34910 ;
  assign n34912 = \wishbone_tx_fifo_fifo_reg[1][28]/P0001  & n34290 ;
  assign n34913 = \wishbone_tx_fifo_fifo_reg[10][28]/P0001  & n34281 ;
  assign n34914 = ~n34912 & ~n34913 ;
  assign n34915 = n34911 & n34914 ;
  assign n34916 = \wishbone_tx_fifo_fifo_reg[12][28]/P0001  & n34287 ;
  assign n34917 = \wishbone_tx_fifo_fifo_reg[5][28]/P0001  & n34267 ;
  assign n34918 = ~n34916 & ~n34917 ;
  assign n34919 = \wishbone_tx_fifo_fifo_reg[4][28]/P0001  & n34279 ;
  assign n34920 = \wishbone_tx_fifo_fifo_reg[8][28]/P0001  & n34270 ;
  assign n34921 = ~n34919 & ~n34920 ;
  assign n34922 = n34918 & n34921 ;
  assign n34923 = n34915 & n34922 ;
  assign n34924 = \wishbone_tx_fifo_fifo_reg[11][28]/P0001  & n34265 ;
  assign n34925 = \wishbone_tx_fifo_fifo_reg[15][28]/P0001  & n34272 ;
  assign n34926 = \wishbone_tx_fifo_fifo_reg[3][28]/P0001  & n34292 ;
  assign n34927 = ~n34925 & ~n34926 ;
  assign n34928 = ~n34924 & n34927 ;
  assign n34929 = \wishbone_tx_fifo_fifo_reg[7][28]/P0001  & n34261 ;
  assign n34930 = \wishbone_tx_fifo_fifo_reg[2][28]/P0001  & n34277 ;
  assign n34931 = ~n34929 & ~n34930 ;
  assign n34932 = \wishbone_tx_fifo_fifo_reg[13][28]/P0001  & n34250 ;
  assign n34933 = \wishbone_tx_fifo_fifo_reg[9][28]/P0001  & n34257 ;
  assign n34934 = ~n34932 & ~n34933 ;
  assign n34935 = n34931 & n34934 ;
  assign n34936 = n34928 & n34935 ;
  assign n34937 = n34923 & n34936 ;
  assign n34938 = n34242 & ~n34937 ;
  assign n34939 = ~n34908 & ~n34938 ;
  assign n34940 = \wishbone_tx_fifo_fifo_reg[0][29]/P0001  & ~n34246 ;
  assign n34941 = \wishbone_tx_fifo_fifo_reg[11][29]/P0001  & n34265 ;
  assign n34942 = \wishbone_tx_fifo_fifo_reg[10][29]/P0001  & n34281 ;
  assign n34943 = ~n34941 & ~n34942 ;
  assign n34944 = \wishbone_tx_fifo_fifo_reg[8][29]/P0001  & n34270 ;
  assign n34945 = \wishbone_tx_fifo_fifo_reg[4][29]/P0001  & n34279 ;
  assign n34946 = ~n34944 & ~n34945 ;
  assign n34947 = n34943 & n34946 ;
  assign n34948 = \wishbone_tx_fifo_fifo_reg[3][29]/P0001  & n34292 ;
  assign n34949 = \wishbone_tx_fifo_fifo_reg[13][29]/P0001  & n34250 ;
  assign n34950 = ~n34948 & ~n34949 ;
  assign n34951 = \wishbone_tx_fifo_fifo_reg[1][29]/P0001  & n34290 ;
  assign n34952 = \wishbone_tx_fifo_fifo_reg[12][29]/P0001  & n34287 ;
  assign n34953 = ~n34951 & ~n34952 ;
  assign n34954 = n34950 & n34953 ;
  assign n34955 = n34947 & n34954 ;
  assign n34956 = \wishbone_tx_fifo_fifo_reg[15][29]/P0001  & n34272 ;
  assign n34957 = \wishbone_tx_fifo_fifo_reg[9][29]/P0001  & n34257 ;
  assign n34958 = \wishbone_tx_fifo_fifo_reg[14][29]/P0001  & n34253 ;
  assign n34959 = ~n34957 & ~n34958 ;
  assign n34960 = ~n34956 & n34959 ;
  assign n34961 = \wishbone_tx_fifo_fifo_reg[6][29]/P0001  & n34285 ;
  assign n34962 = \wishbone_tx_fifo_fifo_reg[7][29]/P0001  & n34261 ;
  assign n34963 = ~n34961 & ~n34962 ;
  assign n34964 = \wishbone_tx_fifo_fifo_reg[5][29]/P0001  & n34267 ;
  assign n34965 = \wishbone_tx_fifo_fifo_reg[2][29]/P0001  & n34277 ;
  assign n34966 = ~n34964 & ~n34965 ;
  assign n34967 = n34963 & n34966 ;
  assign n34968 = n34960 & n34967 ;
  assign n34969 = n34955 & n34968 ;
  assign n34970 = n34242 & ~n34969 ;
  assign n34971 = ~n34940 & ~n34970 ;
  assign n34972 = \wishbone_tx_fifo_fifo_reg[0][2]/P0001  & ~n34246 ;
  assign n34973 = \wishbone_tx_fifo_fifo_reg[2][2]/P0001  & n34277 ;
  assign n34974 = \wishbone_tx_fifo_fifo_reg[7][2]/P0001  & n34261 ;
  assign n34975 = ~n34973 & ~n34974 ;
  assign n34976 = \wishbone_tx_fifo_fifo_reg[15][2]/P0001  & n34272 ;
  assign n34977 = \wishbone_tx_fifo_fifo_reg[14][2]/P0001  & n34253 ;
  assign n34978 = ~n34976 & ~n34977 ;
  assign n34979 = n34975 & n34978 ;
  assign n34980 = \wishbone_tx_fifo_fifo_reg[1][2]/P0001  & n34290 ;
  assign n34981 = \wishbone_tx_fifo_fifo_reg[13][2]/P0001  & n34250 ;
  assign n34982 = ~n34980 & ~n34981 ;
  assign n34983 = \wishbone_tx_fifo_fifo_reg[5][2]/P0001  & n34267 ;
  assign n34984 = \wishbone_tx_fifo_fifo_reg[3][2]/P0001  & n34292 ;
  assign n34985 = ~n34983 & ~n34984 ;
  assign n34986 = n34982 & n34985 ;
  assign n34987 = n34979 & n34986 ;
  assign n34988 = \wishbone_tx_fifo_fifo_reg[8][2]/P0001  & n34270 ;
  assign n34989 = \wishbone_tx_fifo_fifo_reg[10][2]/P0001  & n34281 ;
  assign n34990 = \wishbone_tx_fifo_fifo_reg[6][2]/P0001  & n34285 ;
  assign n34991 = ~n34989 & ~n34990 ;
  assign n34992 = ~n34988 & n34991 ;
  assign n34993 = \wishbone_tx_fifo_fifo_reg[12][2]/P0001  & n34287 ;
  assign n34994 = \wishbone_tx_fifo_fifo_reg[4][2]/P0001  & n34279 ;
  assign n34995 = ~n34993 & ~n34994 ;
  assign n34996 = \wishbone_tx_fifo_fifo_reg[11][2]/P0001  & n34265 ;
  assign n34997 = \wishbone_tx_fifo_fifo_reg[9][2]/P0001  & n34257 ;
  assign n34998 = ~n34996 & ~n34997 ;
  assign n34999 = n34995 & n34998 ;
  assign n35000 = n34992 & n34999 ;
  assign n35001 = n34987 & n35000 ;
  assign n35002 = n34242 & ~n35001 ;
  assign n35003 = ~n34972 & ~n35002 ;
  assign n35004 = \wishbone_tx_fifo_fifo_reg[0][30]/P0001  & ~n34246 ;
  assign n35005 = \wishbone_tx_fifo_fifo_reg[5][30]/P0001  & n34267 ;
  assign n35006 = \wishbone_tx_fifo_fifo_reg[9][30]/P0001  & n34257 ;
  assign n35007 = ~n35005 & ~n35006 ;
  assign n35008 = \wishbone_tx_fifo_fifo_reg[10][30]/P0001  & n34281 ;
  assign n35009 = \wishbone_tx_fifo_fifo_reg[13][30]/P0001  & n34250 ;
  assign n35010 = ~n35008 & ~n35009 ;
  assign n35011 = n35007 & n35010 ;
  assign n35012 = \wishbone_tx_fifo_fifo_reg[6][30]/P0001  & n34285 ;
  assign n35013 = \wishbone_tx_fifo_fifo_reg[12][30]/P0001  & n34287 ;
  assign n35014 = ~n35012 & ~n35013 ;
  assign n35015 = \wishbone_tx_fifo_fifo_reg[8][30]/P0001  & n34270 ;
  assign n35016 = \wishbone_tx_fifo_fifo_reg[11][30]/P0001  & n34265 ;
  assign n35017 = ~n35015 & ~n35016 ;
  assign n35018 = n35014 & n35017 ;
  assign n35019 = n35011 & n35018 ;
  assign n35020 = \wishbone_tx_fifo_fifo_reg[2][30]/P0001  & n34277 ;
  assign n35021 = \wishbone_tx_fifo_fifo_reg[7][30]/P0001  & n34261 ;
  assign n35022 = \wishbone_tx_fifo_fifo_reg[14][30]/P0001  & n34253 ;
  assign n35023 = ~n35021 & ~n35022 ;
  assign n35024 = ~n35020 & n35023 ;
  assign n35025 = \wishbone_tx_fifo_fifo_reg[1][30]/P0001  & n34290 ;
  assign n35026 = \wishbone_tx_fifo_fifo_reg[15][30]/P0001  & n34272 ;
  assign n35027 = ~n35025 & ~n35026 ;
  assign n35028 = \wishbone_tx_fifo_fifo_reg[4][30]/P0001  & n34279 ;
  assign n35029 = \wishbone_tx_fifo_fifo_reg[3][30]/P0001  & n34292 ;
  assign n35030 = ~n35028 & ~n35029 ;
  assign n35031 = n35027 & n35030 ;
  assign n35032 = n35024 & n35031 ;
  assign n35033 = n35019 & n35032 ;
  assign n35034 = n34242 & ~n35033 ;
  assign n35035 = ~n35004 & ~n35034 ;
  assign n35036 = \wishbone_tx_fifo_fifo_reg[0][31]/P0001  & ~n34246 ;
  assign n35037 = \wishbone_tx_fifo_fifo_reg[3][31]/P0001  & n34292 ;
  assign n35038 = \wishbone_tx_fifo_fifo_reg[7][31]/P0001  & n34261 ;
  assign n35039 = ~n35037 & ~n35038 ;
  assign n35040 = \wishbone_tx_fifo_fifo_reg[15][31]/P0001  & n34272 ;
  assign n35041 = \wishbone_tx_fifo_fifo_reg[14][31]/P0001  & n34253 ;
  assign n35042 = ~n35040 & ~n35041 ;
  assign n35043 = n35039 & n35042 ;
  assign n35044 = \wishbone_tx_fifo_fifo_reg[2][31]/P0001  & n34277 ;
  assign n35045 = \wishbone_tx_fifo_fifo_reg[13][31]/P0001  & n34250 ;
  assign n35046 = ~n35044 & ~n35045 ;
  assign n35047 = \wishbone_tx_fifo_fifo_reg[5][31]/P0001  & n34267 ;
  assign n35048 = \wishbone_tx_fifo_fifo_reg[11][31]/P0001  & n34265 ;
  assign n35049 = ~n35047 & ~n35048 ;
  assign n35050 = n35046 & n35049 ;
  assign n35051 = n35043 & n35050 ;
  assign n35052 = \wishbone_tx_fifo_fifo_reg[8][31]/P0001  & n34270 ;
  assign n35053 = \wishbone_tx_fifo_fifo_reg[10][31]/P0001  & n34281 ;
  assign n35054 = \wishbone_tx_fifo_fifo_reg[6][31]/P0001  & n34285 ;
  assign n35055 = ~n35053 & ~n35054 ;
  assign n35056 = ~n35052 & n35055 ;
  assign n35057 = \wishbone_tx_fifo_fifo_reg[12][31]/P0001  & n34287 ;
  assign n35058 = \wishbone_tx_fifo_fifo_reg[4][31]/P0001  & n34279 ;
  assign n35059 = ~n35057 & ~n35058 ;
  assign n35060 = \wishbone_tx_fifo_fifo_reg[1][31]/P0001  & n34290 ;
  assign n35061 = \wishbone_tx_fifo_fifo_reg[9][31]/P0001  & n34257 ;
  assign n35062 = ~n35060 & ~n35061 ;
  assign n35063 = n35059 & n35062 ;
  assign n35064 = n35056 & n35063 ;
  assign n35065 = n35051 & n35064 ;
  assign n35066 = n34242 & ~n35065 ;
  assign n35067 = ~n35036 & ~n35066 ;
  assign n35068 = \wishbone_tx_fifo_fifo_reg[0][3]/P0001  & ~n34246 ;
  assign n35069 = \wishbone_tx_fifo_fifo_reg[15][3]/P0001  & n34272 ;
  assign n35070 = \wishbone_tx_fifo_fifo_reg[6][3]/P0001  & n34285 ;
  assign n35071 = ~n35069 & ~n35070 ;
  assign n35072 = \wishbone_tx_fifo_fifo_reg[3][3]/P0001  & n34292 ;
  assign n35073 = \wishbone_tx_fifo_fifo_reg[11][3]/P0001  & n34265 ;
  assign n35074 = ~n35072 & ~n35073 ;
  assign n35075 = n35071 & n35074 ;
  assign n35076 = \wishbone_tx_fifo_fifo_reg[12][3]/P0001  & n34287 ;
  assign n35077 = \wishbone_tx_fifo_fifo_reg[10][3]/P0001  & n34281 ;
  assign n35078 = ~n35076 & ~n35077 ;
  assign n35079 = \wishbone_tx_fifo_fifo_reg[5][3]/P0001  & n34267 ;
  assign n35080 = \wishbone_tx_fifo_fifo_reg[8][3]/P0001  & n34270 ;
  assign n35081 = ~n35079 & ~n35080 ;
  assign n35082 = n35078 & n35081 ;
  assign n35083 = n35075 & n35082 ;
  assign n35084 = \wishbone_tx_fifo_fifo_reg[2][3]/P0001  & n34277 ;
  assign n35085 = \wishbone_tx_fifo_fifo_reg[14][3]/P0001  & n34253 ;
  assign n35086 = \wishbone_tx_fifo_fifo_reg[1][3]/P0001  & n34290 ;
  assign n35087 = ~n35085 & ~n35086 ;
  assign n35088 = ~n35084 & n35087 ;
  assign n35089 = \wishbone_tx_fifo_fifo_reg[13][3]/P0001  & n34250 ;
  assign n35090 = \wishbone_tx_fifo_fifo_reg[9][3]/P0001  & n34257 ;
  assign n35091 = ~n35089 & ~n35090 ;
  assign n35092 = \wishbone_tx_fifo_fifo_reg[7][3]/P0001  & n34261 ;
  assign n35093 = \wishbone_tx_fifo_fifo_reg[4][3]/P0001  & n34279 ;
  assign n35094 = ~n35092 & ~n35093 ;
  assign n35095 = n35091 & n35094 ;
  assign n35096 = n35088 & n35095 ;
  assign n35097 = n35083 & n35096 ;
  assign n35098 = n34242 & ~n35097 ;
  assign n35099 = ~n35068 & ~n35098 ;
  assign n35100 = \wishbone_tx_fifo_fifo_reg[0][4]/P0001  & ~n34246 ;
  assign n35101 = \wishbone_tx_fifo_fifo_reg[13][4]/P0001  & n34250 ;
  assign n35102 = \wishbone_tx_fifo_fifo_reg[6][4]/P0001  & n34285 ;
  assign n35103 = ~n35101 & ~n35102 ;
  assign n35104 = \wishbone_tx_fifo_fifo_reg[8][4]/P0001  & n34270 ;
  assign n35105 = \wishbone_tx_fifo_fifo_reg[14][4]/P0001  & n34253 ;
  assign n35106 = ~n35104 & ~n35105 ;
  assign n35107 = n35103 & n35106 ;
  assign n35108 = \wishbone_tx_fifo_fifo_reg[3][4]/P0001  & n34292 ;
  assign n35109 = \wishbone_tx_fifo_fifo_reg[5][4]/P0001  & n34267 ;
  assign n35110 = ~n35108 & ~n35109 ;
  assign n35111 = \wishbone_tx_fifo_fifo_reg[15][4]/P0001  & n34272 ;
  assign n35112 = \wishbone_tx_fifo_fifo_reg[2][4]/P0001  & n34277 ;
  assign n35113 = ~n35111 & ~n35112 ;
  assign n35114 = n35110 & n35113 ;
  assign n35115 = n35107 & n35114 ;
  assign n35116 = \wishbone_tx_fifo_fifo_reg[1][4]/P0001  & n34290 ;
  assign n35117 = \wishbone_tx_fifo_fifo_reg[4][4]/P0001  & n34279 ;
  assign n35118 = \wishbone_tx_fifo_fifo_reg[9][4]/P0001  & n34257 ;
  assign n35119 = ~n35117 & ~n35118 ;
  assign n35120 = ~n35116 & n35119 ;
  assign n35121 = \wishbone_tx_fifo_fifo_reg[7][4]/P0001  & n34261 ;
  assign n35122 = \wishbone_tx_fifo_fifo_reg[10][4]/P0001  & n34281 ;
  assign n35123 = ~n35121 & ~n35122 ;
  assign n35124 = \wishbone_tx_fifo_fifo_reg[11][4]/P0001  & n34265 ;
  assign n35125 = \wishbone_tx_fifo_fifo_reg[12][4]/P0001  & n34287 ;
  assign n35126 = ~n35124 & ~n35125 ;
  assign n35127 = n35123 & n35126 ;
  assign n35128 = n35120 & n35127 ;
  assign n35129 = n35115 & n35128 ;
  assign n35130 = n34242 & ~n35129 ;
  assign n35131 = ~n35100 & ~n35130 ;
  assign n35132 = \wishbone_tx_fifo_fifo_reg[0][5]/P0001  & ~n34246 ;
  assign n35133 = \wishbone_tx_fifo_fifo_reg[10][5]/P0001  & n34281 ;
  assign n35134 = \wishbone_tx_fifo_fifo_reg[6][5]/P0001  & n34285 ;
  assign n35135 = ~n35133 & ~n35134 ;
  assign n35136 = \wishbone_tx_fifo_fifo_reg[12][5]/P0001  & n34287 ;
  assign n35137 = \wishbone_tx_fifo_fifo_reg[4][5]/P0001  & n34279 ;
  assign n35138 = ~n35136 & ~n35137 ;
  assign n35139 = n35135 & n35138 ;
  assign n35140 = \wishbone_tx_fifo_fifo_reg[3][5]/P0001  & n34292 ;
  assign n35141 = \wishbone_tx_fifo_fifo_reg[9][5]/P0001  & n34257 ;
  assign n35142 = ~n35140 & ~n35141 ;
  assign n35143 = \wishbone_tx_fifo_fifo_reg[5][5]/P0001  & n34267 ;
  assign n35144 = \wishbone_tx_fifo_fifo_reg[7][5]/P0001  & n34261 ;
  assign n35145 = ~n35143 & ~n35144 ;
  assign n35146 = n35142 & n35145 ;
  assign n35147 = n35139 & n35146 ;
  assign n35148 = \wishbone_tx_fifo_fifo_reg[15][5]/P0001  & n34272 ;
  assign n35149 = \wishbone_tx_fifo_fifo_reg[8][5]/P0001  & n34270 ;
  assign n35150 = \wishbone_tx_fifo_fifo_reg[11][5]/P0001  & n34265 ;
  assign n35151 = ~n35149 & ~n35150 ;
  assign n35152 = ~n35148 & n35151 ;
  assign n35153 = \wishbone_tx_fifo_fifo_reg[1][5]/P0001  & n34290 ;
  assign n35154 = \wishbone_tx_fifo_fifo_reg[13][5]/P0001  & n34250 ;
  assign n35155 = ~n35153 & ~n35154 ;
  assign n35156 = \wishbone_tx_fifo_fifo_reg[2][5]/P0001  & n34277 ;
  assign n35157 = \wishbone_tx_fifo_fifo_reg[14][5]/P0001  & n34253 ;
  assign n35158 = ~n35156 & ~n35157 ;
  assign n35159 = n35155 & n35158 ;
  assign n35160 = n35152 & n35159 ;
  assign n35161 = n35147 & n35160 ;
  assign n35162 = n34242 & ~n35161 ;
  assign n35163 = ~n35132 & ~n35162 ;
  assign n35164 = \wishbone_tx_fifo_fifo_reg[0][6]/P0001  & ~n34246 ;
  assign n35165 = \wishbone_tx_fifo_fifo_reg[9][6]/P0001  & n34257 ;
  assign n35166 = \wishbone_tx_fifo_fifo_reg[6][6]/P0001  & n34285 ;
  assign n35167 = ~n35165 & ~n35166 ;
  assign n35168 = \wishbone_tx_fifo_fifo_reg[2][6]/P0001  & n34277 ;
  assign n35169 = \wishbone_tx_fifo_fifo_reg[1][6]/P0001  & n34290 ;
  assign n35170 = ~n35168 & ~n35169 ;
  assign n35171 = n35167 & n35170 ;
  assign n35172 = \wishbone_tx_fifo_fifo_reg[12][6]/P0001  & n34287 ;
  assign n35173 = \wishbone_tx_fifo_fifo_reg[5][6]/P0001  & n34267 ;
  assign n35174 = ~n35172 & ~n35173 ;
  assign n35175 = \wishbone_tx_fifo_fifo_reg[14][6]/P0001  & n34253 ;
  assign n35176 = \wishbone_tx_fifo_fifo_reg[3][6]/P0001  & n34292 ;
  assign n35177 = ~n35175 & ~n35176 ;
  assign n35178 = n35174 & n35177 ;
  assign n35179 = n35171 & n35178 ;
  assign n35180 = \wishbone_tx_fifo_fifo_reg[7][6]/P0001  & n34261 ;
  assign n35181 = \wishbone_tx_fifo_fifo_reg[10][6]/P0001  & n34281 ;
  assign n35182 = \wishbone_tx_fifo_fifo_reg[8][6]/P0001  & n34270 ;
  assign n35183 = ~n35181 & ~n35182 ;
  assign n35184 = ~n35180 & n35183 ;
  assign n35185 = \wishbone_tx_fifo_fifo_reg[4][6]/P0001  & n34279 ;
  assign n35186 = \wishbone_tx_fifo_fifo_reg[11][6]/P0001  & n34265 ;
  assign n35187 = ~n35185 & ~n35186 ;
  assign n35188 = \wishbone_tx_fifo_fifo_reg[15][6]/P0001  & n34272 ;
  assign n35189 = \wishbone_tx_fifo_fifo_reg[13][6]/P0001  & n34250 ;
  assign n35190 = ~n35188 & ~n35189 ;
  assign n35191 = n35187 & n35190 ;
  assign n35192 = n35184 & n35191 ;
  assign n35193 = n35179 & n35192 ;
  assign n35194 = n34242 & ~n35193 ;
  assign n35195 = ~n35164 & ~n35194 ;
  assign n35196 = \wishbone_tx_fifo_fifo_reg[0][7]/P0001  & ~n34246 ;
  assign n35197 = \wishbone_tx_fifo_fifo_reg[6][7]/P0001  & n34285 ;
  assign n35198 = \wishbone_tx_fifo_fifo_reg[1][7]/P0001  & n34290 ;
  assign n35199 = ~n35197 & ~n35198 ;
  assign n35200 = \wishbone_tx_fifo_fifo_reg[11][7]/P0001  & n34265 ;
  assign n35201 = \wishbone_tx_fifo_fifo_reg[4][7]/P0001  & n34279 ;
  assign n35202 = ~n35200 & ~n35201 ;
  assign n35203 = n35199 & n35202 ;
  assign n35204 = \wishbone_tx_fifo_fifo_reg[9][7]/P0001  & n34257 ;
  assign n35205 = \wishbone_tx_fifo_fifo_reg[14][7]/P0001  & n34253 ;
  assign n35206 = ~n35204 & ~n35205 ;
  assign n35207 = \wishbone_tx_fifo_fifo_reg[10][7]/P0001  & n34281 ;
  assign n35208 = \wishbone_tx_fifo_fifo_reg[15][7]/P0001  & n34272 ;
  assign n35209 = ~n35207 & ~n35208 ;
  assign n35210 = n35206 & n35209 ;
  assign n35211 = n35203 & n35210 ;
  assign n35212 = \wishbone_tx_fifo_fifo_reg[3][7]/P0001  & n34292 ;
  assign n35213 = \wishbone_tx_fifo_fifo_reg[8][7]/P0001  & n34270 ;
  assign n35214 = \wishbone_tx_fifo_fifo_reg[2][7]/P0001  & n34277 ;
  assign n35215 = ~n35213 & ~n35214 ;
  assign n35216 = ~n35212 & n35215 ;
  assign n35217 = \wishbone_tx_fifo_fifo_reg[13][7]/P0001  & n34250 ;
  assign n35218 = \wishbone_tx_fifo_fifo_reg[5][7]/P0001  & n34267 ;
  assign n35219 = ~n35217 & ~n35218 ;
  assign n35220 = \wishbone_tx_fifo_fifo_reg[7][7]/P0001  & n34261 ;
  assign n35221 = \wishbone_tx_fifo_fifo_reg[12][7]/P0001  & n34287 ;
  assign n35222 = ~n35220 & ~n35221 ;
  assign n35223 = n35219 & n35222 ;
  assign n35224 = n35216 & n35223 ;
  assign n35225 = n35211 & n35224 ;
  assign n35226 = n34242 & ~n35225 ;
  assign n35227 = ~n35196 & ~n35226 ;
  assign n35228 = \wishbone_tx_fifo_fifo_reg[0][8]/P0001  & ~n34246 ;
  assign n35229 = \wishbone_tx_fifo_fifo_reg[8][8]/P0001  & n34270 ;
  assign n35230 = \wishbone_tx_fifo_fifo_reg[5][8]/P0001  & n34267 ;
  assign n35231 = ~n35229 & ~n35230 ;
  assign n35232 = \wishbone_tx_fifo_fifo_reg[13][8]/P0001  & n34250 ;
  assign n35233 = \wishbone_tx_fifo_fifo_reg[4][8]/P0001  & n34279 ;
  assign n35234 = ~n35232 & ~n35233 ;
  assign n35235 = n35231 & n35234 ;
  assign n35236 = \wishbone_tx_fifo_fifo_reg[9][8]/P0001  & n34257 ;
  assign n35237 = \wishbone_tx_fifo_fifo_reg[3][8]/P0001  & n34292 ;
  assign n35238 = ~n35236 & ~n35237 ;
  assign n35239 = \wishbone_tx_fifo_fifo_reg[6][8]/P0001  & n34285 ;
  assign n35240 = \wishbone_tx_fifo_fifo_reg[15][8]/P0001  & n34272 ;
  assign n35241 = ~n35239 & ~n35240 ;
  assign n35242 = n35238 & n35241 ;
  assign n35243 = n35235 & n35242 ;
  assign n35244 = \wishbone_tx_fifo_fifo_reg[11][8]/P0001  & n34265 ;
  assign n35245 = \wishbone_tx_fifo_fifo_reg[1][8]/P0001  & n34290 ;
  assign n35246 = \wishbone_tx_fifo_fifo_reg[10][8]/P0001  & n34281 ;
  assign n35247 = ~n35245 & ~n35246 ;
  assign n35248 = ~n35244 & n35247 ;
  assign n35249 = \wishbone_tx_fifo_fifo_reg[14][8]/P0001  & n34253 ;
  assign n35250 = \wishbone_tx_fifo_fifo_reg[12][8]/P0001  & n34287 ;
  assign n35251 = ~n35249 & ~n35250 ;
  assign n35252 = \wishbone_tx_fifo_fifo_reg[7][8]/P0001  & n34261 ;
  assign n35253 = \wishbone_tx_fifo_fifo_reg[2][8]/P0001  & n34277 ;
  assign n35254 = ~n35252 & ~n35253 ;
  assign n35255 = n35251 & n35254 ;
  assign n35256 = n35248 & n35255 ;
  assign n35257 = n35243 & n35256 ;
  assign n35258 = n34242 & ~n35257 ;
  assign n35259 = ~n35228 & ~n35258 ;
  assign n35260 = \wishbone_tx_fifo_fifo_reg[0][9]/P0001  & ~n34246 ;
  assign n35261 = \wishbone_tx_fifo_fifo_reg[13][9]/P0001  & n34250 ;
  assign n35262 = \wishbone_tx_fifo_fifo_reg[14][9]/P0001  & n34253 ;
  assign n35263 = ~n35261 & ~n35262 ;
  assign n35264 = \wishbone_tx_fifo_fifo_reg[9][9]/P0001  & n34257 ;
  assign n35265 = \wishbone_tx_fifo_fifo_reg[7][9]/P0001  & n34261 ;
  assign n35266 = ~n35264 & ~n35265 ;
  assign n35267 = n35263 & n35266 ;
  assign n35268 = \wishbone_tx_fifo_fifo_reg[11][9]/P0001  & n34265 ;
  assign n35269 = \wishbone_tx_fifo_fifo_reg[5][9]/P0001  & n34267 ;
  assign n35270 = ~n35268 & ~n35269 ;
  assign n35271 = \wishbone_tx_fifo_fifo_reg[8][9]/P0001  & n34270 ;
  assign n35272 = \wishbone_tx_fifo_fifo_reg[15][9]/P0001  & n34272 ;
  assign n35273 = ~n35271 & ~n35272 ;
  assign n35274 = n35270 & n35273 ;
  assign n35275 = n35267 & n35274 ;
  assign n35276 = \wishbone_tx_fifo_fifo_reg[2][9]/P0001  & n34277 ;
  assign n35277 = \wishbone_tx_fifo_fifo_reg[4][9]/P0001  & n34279 ;
  assign n35278 = \wishbone_tx_fifo_fifo_reg[10][9]/P0001  & n34281 ;
  assign n35279 = ~n35277 & ~n35278 ;
  assign n35280 = ~n35276 & n35279 ;
  assign n35281 = \wishbone_tx_fifo_fifo_reg[6][9]/P0001  & n34285 ;
  assign n35282 = \wishbone_tx_fifo_fifo_reg[12][9]/P0001  & n34287 ;
  assign n35283 = ~n35281 & ~n35282 ;
  assign n35284 = \wishbone_tx_fifo_fifo_reg[1][9]/P0001  & n34290 ;
  assign n35285 = \wishbone_tx_fifo_fifo_reg[3][9]/P0001  & n34292 ;
  assign n35286 = ~n35284 & ~n35285 ;
  assign n35287 = n35283 & n35286 ;
  assign n35288 = n35280 & n35287 ;
  assign n35289 = n35275 & n35288 ;
  assign n35290 = n34242 & ~n35289 ;
  assign n35291 = ~n35260 & ~n35290 ;
  assign n35292 = \wishbone_tx_burst_cnt_reg[1]/NET0131  & ~n13174 ;
  assign n35293 = n32466 & n35292 ;
  assign n35294 = ~n13167 & ~n32461 ;
  assign n35295 = ~n13166 & n35294 ;
  assign n35296 = ~n13164 & n35295 ;
  assign n35297 = ~n35293 & ~n35296 ;
  assign n35298 = \wishbone_ReadTxDataFromFifo_sync2_reg/NET0131  & ~\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131  ;
  assign n35299 = n14049 & ~n35298 ;
  assign n35300 = ~\wishbone_tx_fifo_cnt_reg[0]/NET0131  & ~\wishbone_tx_fifo_cnt_reg[1]/NET0131  ;
  assign n35301 = ~\wishbone_tx_fifo_cnt_reg[2]/NET0131  & n35300 ;
  assign n35302 = ~\wishbone_tx_fifo_cnt_reg[3]/NET0131  & ~\wishbone_tx_fifo_cnt_reg[4]/NET0131  ;
  assign n35303 = n14049 & n35302 ;
  assign n35304 = n35301 & n35303 ;
  assign n35305 = ~n35299 & ~n35304 ;
  assign n35306 = n35301 & n35302 ;
  assign n35307 = ~n14049 & n35298 ;
  assign n35308 = ~n35306 & n35307 ;
  assign n35309 = n35305 & ~n35308 ;
  assign n35310 = \wishbone_tx_fifo_cnt_reg[0]/NET0131  & \wishbone_tx_fifo_cnt_reg[1]/NET0131  ;
  assign n35311 = n32477 & n35310 ;
  assign n35312 = n14049 & ~n35311 ;
  assign n35313 = ~\wishbone_tx_fifo_cnt_reg[2]/NET0131  & ~\wishbone_tx_fifo_cnt_reg[3]/NET0131  ;
  assign n35314 = n35300 & n35313 ;
  assign n35315 = n35298 & ~n35314 ;
  assign n35316 = ~n35312 & ~n35315 ;
  assign n35317 = ~n35309 & n35316 ;
  assign n35318 = ~\wishbone_tx_fifo_cnt_reg[4]/NET0131  & ~n35317 ;
  assign n35319 = \wishbone_tx_fifo_cnt_reg[4]/NET0131  & n35316 ;
  assign n35320 = ~n35309 & n35319 ;
  assign n35321 = n34242 & ~n35320 ;
  assign n35322 = ~n35318 & n35321 ;
  assign n35323 = ~\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131  & ~n32871 ;
  assign n35324 = \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  & \wishbone_RxStatusWriteLatched_sync2_reg/NET0131  ;
  assign n35325 = ~n13087 & ~n35324 ;
  assign n35326 = ~n35323 & n35325 ;
  assign n35327 = ~mdc_pad_o_pad & \miim1_InProgress_reg/NET0131  ;
  assign n35328 = n32264 & n35327 ;
  assign n35329 = \miim1_BitCounter_reg[0]/NET0131  & \miim1_BitCounter_reg[1]/NET0131  ;
  assign n35330 = \miim1_BitCounter_reg[2]/NET0131  & \miim1_BitCounter_reg[3]/NET0131  ;
  assign n35331 = n35329 & n35330 ;
  assign n35332 = \miim1_BitCounter_reg[4]/NET0131  & n35331 ;
  assign n35333 = ~\miim1_BitCounter_reg[5]/NET0131  & ~n35332 ;
  assign n35334 = \miim1_BitCounter_reg[4]/NET0131  & \miim1_BitCounter_reg[5]/NET0131  ;
  assign n35335 = n35331 & n35334 ;
  assign n35336 = ~n35333 & ~n35335 ;
  assign n35337 = n35328 & n35336 ;
  assign n35338 = ~mdc_pad_o_pad & n32264 ;
  assign n35339 = \miim1_BitCounter_reg[5]/NET0131  & ~n35338 ;
  assign n35340 = n32523 & n35338 ;
  assign n35341 = ~n35339 & ~n35340 ;
  assign n35342 = ~n35337 & n35341 ;
  assign n35343 = \wishbone_rx_burst_en_reg/NET0131  & ~n13191 ;
  assign n35344 = n32430 & n35343 ;
  assign n35345 = \wishbone_rx_burst_cnt_reg[0]/NET0131  & \wishbone_rx_burst_cnt_reg[1]/NET0131  ;
  assign n35346 = ~\wishbone_rx_burst_cnt_reg[2]/NET0131  & n35345 ;
  assign n35347 = ~n13149 & ~n35346 ;
  assign n35348 = n13143 & n35347 ;
  assign n35349 = n13137 & n35348 ;
  assign n35350 = \wishbone_MasterWbRX_reg/NET0131  & n13126 ;
  assign n35351 = \wishbone_rx_fifo_cnt_reg[2]/NET0131  & ~n35350 ;
  assign n35352 = n13128 & ~n35351 ;
  assign n35353 = n32415 & ~n35352 ;
  assign n35354 = ~n32423 & ~n35352 ;
  assign n35355 = n32428 & n35354 ;
  assign n35356 = ~n35353 & ~n35355 ;
  assign n35357 = ~n35349 & n35356 ;
  assign n35358 = ~n35344 & n35357 ;
  assign n35359 = \wishbone_WriteRxDataToFifoSync2_reg/NET0131  & ~\wishbone_WriteRxDataToFifoSync3_reg/NET0131  ;
  assign n35360 = n16307 & ~n35359 ;
  assign n35361 = ~\wishbone_rx_fifo_cnt_reg[3]/NET0131  & \wishbone_rx_fifo_cnt_reg[4]/NET0131  ;
  assign n35362 = n16307 & n35361 ;
  assign n35363 = n13127 & n35362 ;
  assign n35364 = ~n35360 & ~n35363 ;
  assign n35365 = n13127 & n35361 ;
  assign n35366 = ~n16307 & n35359 ;
  assign n35367 = ~n35365 & n35366 ;
  assign n35368 = n35364 & ~n35367 ;
  assign n35369 = n13127 & n16307 ;
  assign n35370 = ~\wishbone_rx_fifo_cnt_reg[3]/NET0131  & ~n35369 ;
  assign n35371 = \wishbone_rx_fifo_cnt_reg[0]/NET0131  & \wishbone_rx_fifo_cnt_reg[1]/NET0131  ;
  assign n35372 = \wishbone_rx_fifo_cnt_reg[2]/NET0131  & ~n16307 ;
  assign n35373 = n35371 & n35372 ;
  assign n35374 = \wishbone_rx_fifo_cnt_reg[3]/NET0131  & ~n35373 ;
  assign n35375 = ~n35370 & ~n35374 ;
  assign n35376 = ~n35368 & n35375 ;
  assign n35377 = \wishbone_rx_fifo_cnt_reg[4]/NET0131  & ~n33164 ;
  assign n35378 = ~n35376 & n35377 ;
  assign n35379 = ~\wishbone_rx_fifo_cnt_reg[4]/NET0131  & ~n33164 ;
  assign n35380 = n35376 & n35379 ;
  assign n35381 = ~n35378 & ~n35380 ;
  assign n35382 = ~\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131  & ~\rxethmac1_RxEndFrm_reg/NET0131  ;
  assign n35383 = \maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131  & \rxethmac1_RxValid_reg/NET0131  ;
  assign n35384 = n35382 & n35383 ;
  assign n35385 = \maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131  & ~n32446 ;
  assign n35386 = ~n35384 & n35385 ;
  assign n35387 = ~\maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131  & ~n32446 ;
  assign n35388 = n35384 & n35387 ;
  assign n35389 = ~n35386 & ~n35388 ;
  assign n35390 = \rxethmac1_RxValid_reg/NET0131  & n35382 ;
  assign n35391 = ~\maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131  & ~n35390 ;
  assign n35392 = ~n32446 & ~n35384 ;
  assign n35393 = ~n35391 & n35392 ;
  assign n35394 = \maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131  & ~n32446 ;
  assign n35395 = n35384 & n35385 ;
  assign n35396 = ~n35394 & ~n35395 ;
  assign n35397 = ~\txethmac1_txstatem1_StateData_reg[1]/NET0131  & \txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n35398 = ~\txethmac1_txcrc_Crc_reg[28]/NET0131  & n35397 ;
  assign n35399 = ~\txethmac1_txstatem1_StateData_reg[1]/NET0131  & ~\txethmac1_txstatem1_StateFCS_reg/NET0131  ;
  assign n35400 = \txethmac1_txstatem1_StateJam_reg/NET0131  & n35399 ;
  assign n35401 = \txethmac1_txstatem1_StatePreamble_reg/NET0131  & n35399 ;
  assign n35402 = n11124 & n35401 ;
  assign n35403 = ~n35400 & ~n35402 ;
  assign n35404 = ~n35398 & n35403 ;
  assign n35405 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n35404 ;
  assign n35406 = n11443 & ~n35405 ;
  assign n35407 = ~\txethmac1_txcrc_Crc_reg[1]/NET0131  & n13011 ;
  assign n35408 = n12998 & n35407 ;
  assign n35409 = ~\txethmac1_txcrc_Crc_reg[1]/NET0131  & n11464 ;
  assign n35410 = n11464 & n13011 ;
  assign n35411 = n12998 & n35410 ;
  assign n35412 = ~n35409 & ~n35411 ;
  assign n35413 = ~n35408 & ~n35412 ;
  assign n35414 = \wishbone_ShiftWillEnd_reg/NET0131  & n15732 ;
  assign n35415 = \wishbone_LastByteIn_reg/NET0131  & ~n35414 ;
  assign n35416 = \rxethmac1_RxEndFrm_reg/NET0131  & ~n15732 ;
  assign n35417 = n32274 & n35416 ;
  assign n35418 = ~n35415 & ~n35417 ;
  assign n35419 = ~\RxAbort_wb_reg/NET0131  & ~n35418 ;
  assign n35420 = \rxethmac1_LatchedByte_reg[4]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n35421 = ~n33020 & n35420 ;
  assign n35422 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[4]/NET0131  ;
  assign n35423 = ~n33021 & n35422 ;
  assign n35424 = ~n35421 & ~n35423 ;
  assign n35425 = \miim1_BitCounter_reg[4]/NET0131  & ~\miim1_BitCounter_reg[6]/NET0131  ;
  assign n35426 = \miim1_BitCounter_reg[5]/NET0131  & n35425 ;
  assign n35427 = n35331 & n35426 ;
  assign n35428 = ~\miim1_InProgress_q1_reg/NET0131  & ~\miim1_InProgress_q2_reg/NET0131  ;
  assign n35429 = ~\miim1_InProgress_reg/NET0131  & \miim1_SyncStatMdcEn_reg/NET0131  ;
  assign n35430 = n35428 & n35429 ;
  assign n35431 = \miim1_WCtrlDataStart_q1_reg/NET0131  & ~\miim1_WCtrlDataStart_q2_reg/NET0131  ;
  assign n35432 = \miim1_RStatStart_q1_reg/NET0131  & ~\miim1_RStatStart_q2_reg/NET0131  ;
  assign n35433 = ~n35431 & ~n35432 ;
  assign n35434 = ~n35430 & n35433 ;
  assign n35435 = ~n35427 & n35434 ;
  assign n35436 = n35338 & ~n35435 ;
  assign n35437 = \miim1_WriteOp_reg/NET0131  & ~n35436 ;
  assign n35438 = \miim1_InProgress_reg/NET0131  & ~\miim1_WriteOp_reg/NET0131  ;
  assign n35439 = ~\miim1_InProgress_reg/NET0131  & ~n35431 ;
  assign n35440 = ~n35438 & ~n35439 ;
  assign n35441 = ~n35434 & n35440 ;
  assign n35442 = n35338 & n35441 ;
  assign n35443 = ~n35437 & ~n35442 ;
  assign n35444 = \ethreg1_MODER_0_DataOut_reg[0]/NET0131  & ~\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131  ;
  assign n35445 = ~\wishbone_r_RxEn_q_reg/NET0131  & n35444 ;
  assign n35446 = \wishbone_RxStatus_reg[13]/NET0131  & \wishbone_ShiftEnded_reg/NET0131  ;
  assign n35447 = n15779 & n35446 ;
  assign n35448 = ~n35445 & ~n35447 ;
  assign n35449 = \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131  & ~n35448 ;
  assign n35450 = \wishbone_ShiftEnded_reg/NET0131  & n15779 ;
  assign n35451 = \wishbone_RxBDAddress_reg[1]/NET0131  & \wishbone_RxBDAddress_reg[2]/NET0131  ;
  assign n35452 = \wishbone_RxBDAddress_reg[3]/NET0131  & n35451 ;
  assign n35453 = n35450 & n35452 ;
  assign n35454 = ~\wishbone_RxBDAddress_reg[4]/NET0131  & ~n35453 ;
  assign n35455 = \wishbone_RxBDAddress_reg[4]/NET0131  & \wishbone_ShiftEnded_reg/NET0131  ;
  assign n35456 = n15779 & n35455 ;
  assign n35457 = n35452 & n35456 ;
  assign n35458 = n35448 & ~n35457 ;
  assign n35459 = ~n35454 & n35458 ;
  assign n35460 = ~n35449 & ~n35459 ;
  assign n35461 = ~\wishbone_LastByteIn_reg/NET0131  & ~\wishbone_ShiftWillEnd_reg/NET0131  ;
  assign n35462 = ~n32449 & n35461 ;
  assign n35463 = n32279 & ~n35462 ;
  assign n35464 = \miim1_BitCounter_reg[1]/NET0131  & ~n35338 ;
  assign n35465 = ~n32519 & ~n35329 ;
  assign n35466 = ~n32522 & n35465 ;
  assign n35467 = n35328 & n35466 ;
  assign n35468 = ~n35464 & ~n35467 ;
  assign n35469 = \miim1_BitCounter_reg[2]/NET0131  & ~n35338 ;
  assign n35470 = \miim1_BitCounter_reg[2]/NET0131  & n35329 ;
  assign n35471 = ~\miim1_BitCounter_reg[2]/NET0131  & ~n35329 ;
  assign n35472 = ~n35470 & ~n35471 ;
  assign n35473 = ~n32522 & n35472 ;
  assign n35474 = n35328 & n35473 ;
  assign n35475 = ~n35469 & ~n35474 ;
  assign n35476 = \miim1_BitCounter_reg[3]/NET0131  & ~n35338 ;
  assign n35477 = ~n32522 & n35328 ;
  assign n35478 = ~\miim1_BitCounter_reg[3]/NET0131  & ~n35470 ;
  assign n35479 = ~n35331 & ~n35478 ;
  assign n35480 = n35477 & n35479 ;
  assign n35481 = ~n35476 & ~n35480 ;
  assign n35482 = \miim1_BitCounter_reg[4]/NET0131  & ~n35338 ;
  assign n35483 = ~\miim1_BitCounter_reg[4]/NET0131  & ~n35331 ;
  assign n35484 = ~n35332 & ~n35483 ;
  assign n35485 = n35477 & n35484 ;
  assign n35486 = ~n35482 & ~n35485 ;
  assign n35487 = \miim1_BitCounter_reg[6]/NET0131  & ~n35338 ;
  assign n35488 = \miim1_BitCounter_reg[6]/NET0131  & ~n35335 ;
  assign n35489 = ~n35427 & ~n35488 ;
  assign n35490 = n35477 & ~n35489 ;
  assign n35491 = ~n35487 & ~n35490 ;
  assign n35492 = ~\miim1_clkgen_Counter_reg[4]/NET0131  & ~\miim1_clkgen_Counter_reg[5]/NET0131  ;
  assign n35493 = n32249 & n35492 ;
  assign n35494 = \miim1_clkgen_Counter_reg[6]/NET0131  & ~n35493 ;
  assign n35495 = ~\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  & ~\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  ;
  assign n35496 = ~\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  & n35495 ;
  assign n35497 = n32258 & n35496 ;
  assign n35498 = \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  & n32264 ;
  assign n35499 = ~n35497 & n35498 ;
  assign n35500 = ~\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  & n32264 ;
  assign n35501 = n35497 & n35500 ;
  assign n35502 = ~n35499 & ~n35501 ;
  assign n35503 = ~n35494 & n35502 ;
  assign n35504 = \rxethmac1_Multicast_reg/NET0131  & n13019 ;
  assign n35505 = \rxethmac1_LatchedByte_reg[0]/NET0131  & n13027 ;
  assign n35506 = n13022 & n35505 ;
  assign n35507 = ~n35504 & ~n35506 ;
  assign n35508 = ~\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131  & ~\macstatus1_ReceiveEnd_reg/NET0131  ;
  assign n35509 = ~n32311 & ~n35508 ;
  assign n35510 = ~\rxethmac1_crcrx_Crc_reg[13]/NET0131  & n10663 ;
  assign n35511 = ~n10662 & n35510 ;
  assign n35512 = \rxethmac1_crcrx_Crc_reg[13]/NET0131  & n10663 ;
  assign n35513 = n10662 & n35512 ;
  assign n35514 = ~n35511 & ~n35513 ;
  assign n35515 = ~\maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001  & \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  ;
  assign n35516 = ~\txethmac1_TxUsedData_reg/NET0131  & ~n35515 ;
  assign n35517 = \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131  & \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131  ;
  assign n35518 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & ~n35517 ;
  assign n35519 = \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~n35518 ;
  assign n35520 = ~n35516 & n35519 ;
  assign n35521 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  ;
  assign n35522 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  & n35521 ;
  assign n35523 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  ;
  assign n35524 = \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & \txethmac1_TxUsedData_reg/NET0131  ;
  assign n35525 = n35523 & n35524 ;
  assign n35526 = n35522 & n35525 ;
  assign n35527 = \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  & ~n35526 ;
  assign n35528 = n35520 & n35527 ;
  assign n35529 = \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & \txethmac1_TxUsedData_reg/NET0131  ;
  assign n35530 = n35515 & n35529 ;
  assign n35531 = ~n35518 & n35530 ;
  assign n35532 = ~n35528 & ~n35531 ;
  assign n35533 = \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n35534 = ~n35532 & n35533 ;
  assign n35535 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  & ~n35534 ;
  assign n35536 = ~\txethmac1_TxAbort_reg/NET0131  & ~\txethmac1_TxDone_reg/NET0131  ;
  assign n35537 = ~\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  & ~n35536 ;
  assign n35538 = ~wb_rst_i_pad & ~n35537 ;
  assign n35539 = \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n35540 = \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  & n35539 ;
  assign n35541 = ~n35532 & n35540 ;
  assign n35542 = n35538 & ~n35541 ;
  assign n35543 = ~n35535 & n35542 ;
  assign n35544 = ~\wishbone_LatchValidBytes_q_reg/NET0131  & \wishbone_LatchValidBytes_reg/NET0131  ;
  assign n35545 = \wishbone_TxLength_reg[0]/NET0131  & n35544 ;
  assign n35546 = n14063 & n35545 ;
  assign n35547 = n14058 & n35546 ;
  assign n35548 = ~\wishbone_TxAbort_wb_q_reg/NET0131  & \wishbone_TxAbort_wb_reg/NET0131  ;
  assign n35549 = ~\wishbone_TxRetry_wb_q_reg/NET0131  & \wishbone_TxRetry_wb_reg/NET0131  ;
  assign n35550 = ~n35548 & ~n35549 ;
  assign n35551 = ~\wishbone_TxDone_wb_q_reg/NET0131  & \wishbone_TxDone_wb_reg/NET0131  ;
  assign n35552 = ~n35544 & ~n35551 ;
  assign n35553 = n35550 & n35552 ;
  assign n35554 = \wishbone_TxValidBytesLatched_reg[0]/NET0131  & n35553 ;
  assign n35555 = ~n35547 & ~n35554 ;
  assign n35556 = \wishbone_TxLength_reg[1]/NET0131  & n35544 ;
  assign n35557 = n14063 & n35556 ;
  assign n35558 = n14058 & n35557 ;
  assign n35559 = \wishbone_TxValidBytesLatched_reg[1]/NET0131  & n35553 ;
  assign n35560 = ~n35558 & ~n35559 ;
  assign n35561 = n11464 & n12554 ;
  assign n35562 = n11464 & n12676 ;
  assign n35563 = ~\miim1_BitCounter_reg[0]/NET0131  & n35327 ;
  assign n35564 = n32264 & n35563 ;
  assign n35565 = \miim1_BitCounter_reg[0]/NET0131  & ~n35338 ;
  assign n35566 = ~n35340 & ~n35565 ;
  assign n35567 = ~n35564 & n35566 ;
  assign n35568 = \txethmac1_txstatem1_StateData_reg[1]/NET0131  & n10693 ;
  assign n35569 = ~n11166 & ~n35568 ;
  assign n35570 = ~n10694 & ~n35569 ;
  assign n35571 = ~\txethmac1_txstatem1_StatePreamble_reg/NET0131  & ~n11348 ;
  assign n35572 = ~n11171 & ~n35571 ;
  assign n35573 = ~n35570 & n35572 ;
  assign n35574 = n35338 & ~n35434 ;
  assign n35575 = n35338 & n35427 ;
  assign n35576 = \miim1_InProgress_reg/NET0131  & ~n35575 ;
  assign n35577 = ~n35574 & ~n35576 ;
  assign n35578 = \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  & \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  ;
  assign n35579 = \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  & \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  ;
  assign n35580 = ~n35578 & ~n35579 ;
  assign n35581 = ~n32258 & n32264 ;
  assign n35582 = n35580 & n35581 ;
  assign n35583 = \miim1_clkgen_Counter_reg[2]/NET0131  & ~n32247 ;
  assign n35584 = ~n32508 & ~n35583 ;
  assign n35585 = ~n32264 & n35584 ;
  assign n35586 = ~n35582 & ~n35585 ;
  assign n35587 = \miim1_LatchByte1_d_reg/NET0131  & ~n35338 ;
  assign n35588 = \miim1_BitCounter_reg[4]/NET0131  & n32526 ;
  assign n35589 = \miim1_BitCounter_reg[1]/NET0131  & \miim1_BitCounter_reg[2]/NET0131  ;
  assign n35590 = \miim1_BitCounter_reg[0]/NET0131  & ~\miim1_BitCounter_reg[3]/NET0131  ;
  assign n35591 = \miim1_BitCounter_reg[5]/NET0131  & ~\miim1_WriteOp_reg/NET0131  ;
  assign n35592 = n35590 & n35591 ;
  assign n35593 = n35589 & n35592 ;
  assign n35594 = n35588 & n35593 ;
  assign n35595 = n35338 & n35594 ;
  assign n35596 = ~n35587 & ~n35595 ;
  assign n35597 = \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131  & ~n35448 ;
  assign n35598 = \wishbone_RxBDAddress_reg[4]/NET0131  & \wishbone_RxBDAddress_reg[5]/NET0131  ;
  assign n35599 = \wishbone_RxBDAddress_reg[6]/NET0131  & n35598 ;
  assign n35600 = n35453 & n35599 ;
  assign n35601 = ~\wishbone_RxBDAddress_reg[7]/NET0131  & ~n35600 ;
  assign n35602 = \wishbone_RxBDAddress_reg[7]/NET0131  & n35599 ;
  assign n35603 = n35453 & n35602 ;
  assign n35604 = n35448 & ~n35603 ;
  assign n35605 = ~n35601 & n35604 ;
  assign n35606 = ~n35597 & ~n35605 ;
  assign n35607 = ~\wishbone_LastByteIn_reg/NET0131  & n32270 ;
  assign n35608 = \rxethmac1_RxStartFrm_reg/NET0131  & n32304 ;
  assign n35609 = ~\rxethmac1_RxStartFrm_reg/NET0131  & ~\wishbone_RxByteCnt_reg[0]/NET0131  ;
  assign n35610 = n32447 & n35609 ;
  assign n35611 = ~n35608 & ~n35610 ;
  assign n35612 = n35607 & ~n35611 ;
  assign n35613 = ~\wishbone_RxDataLatched1_reg[10]/NET0131  & ~n35612 ;
  assign n35614 = ~\rxethmac1_RxData_reg[2]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35615 = n32270 & n35614 ;
  assign n35616 = ~n35611 & n35615 ;
  assign n35617 = ~n35613 & ~n35616 ;
  assign n35618 = ~\wishbone_RxDataLatched1_reg[11]/NET0131  & ~n35612 ;
  assign n35619 = ~\rxethmac1_RxData_reg[3]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35620 = n32270 & n35619 ;
  assign n35621 = ~n35611 & n35620 ;
  assign n35622 = ~n35618 & ~n35621 ;
  assign n35623 = ~\wishbone_RxDataLatched1_reg[12]/NET0131  & ~n35612 ;
  assign n35624 = ~\rxethmac1_RxData_reg[4]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35625 = n32270 & n35624 ;
  assign n35626 = ~n35611 & n35625 ;
  assign n35627 = ~n35623 & ~n35626 ;
  assign n35628 = ~\wishbone_RxDataLatched1_reg[13]/NET0131  & ~n35612 ;
  assign n35629 = ~\rxethmac1_RxData_reg[5]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35630 = n32270 & n35629 ;
  assign n35631 = ~n35611 & n35630 ;
  assign n35632 = ~n35628 & ~n35631 ;
  assign n35633 = ~\wishbone_RxDataLatched1_reg[14]/NET0131  & ~n35612 ;
  assign n35634 = ~\rxethmac1_RxData_reg[6]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35635 = n32270 & n35634 ;
  assign n35636 = ~n35611 & n35635 ;
  assign n35637 = ~n35633 & ~n35636 ;
  assign n35638 = ~\wishbone_RxDataLatched1_reg[15]/NET0131  & ~n35612 ;
  assign n35639 = ~\rxethmac1_RxData_reg[7]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35640 = n32270 & n35639 ;
  assign n35641 = ~n35611 & n35640 ;
  assign n35642 = ~n35638 & ~n35641 ;
  assign n35643 = \rxethmac1_RxStartFrm_reg/NET0131  & n32303 ;
  assign n35644 = ~\wishbone_RxByteCnt_reg[1]/NET0131  & \wishbone_RxEnableWindow_reg/NET0131  ;
  assign n35645 = ~\rxethmac1_RxStartFrm_reg/NET0131  & \wishbone_RxByteCnt_reg[0]/NET0131  ;
  assign n35646 = n35644 & n35645 ;
  assign n35647 = ~n35643 & ~n35646 ;
  assign n35648 = n35607 & ~n35647 ;
  assign n35649 = ~\wishbone_RxDataLatched1_reg[16]/NET0131  & ~n35648 ;
  assign n35650 = ~\rxethmac1_RxData_reg[0]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35651 = n32270 & n35650 ;
  assign n35652 = ~n35647 & n35651 ;
  assign n35653 = ~n35649 & ~n35652 ;
  assign n35654 = ~\wishbone_RxDataLatched1_reg[17]/NET0131  & ~n35648 ;
  assign n35655 = ~\rxethmac1_RxData_reg[1]/NET0131  & ~\wishbone_LastByteIn_reg/NET0131  ;
  assign n35656 = n32270 & n35655 ;
  assign n35657 = ~n35647 & n35656 ;
  assign n35658 = ~n35654 & ~n35657 ;
  assign n35659 = ~\wishbone_RxDataLatched1_reg[18]/NET0131  & ~n35648 ;
  assign n35660 = n35615 & ~n35647 ;
  assign n35661 = ~n35659 & ~n35660 ;
  assign n35662 = ~\wishbone_RxDataLatched1_reg[19]/NET0131  & ~n35648 ;
  assign n35663 = n35620 & ~n35647 ;
  assign n35664 = ~n35662 & ~n35663 ;
  assign n35665 = ~\wishbone_RxDataLatched1_reg[20]/NET0131  & ~n35648 ;
  assign n35666 = n35625 & ~n35647 ;
  assign n35667 = ~n35665 & ~n35666 ;
  assign n35668 = ~\wishbone_RxDataLatched1_reg[21]/NET0131  & ~n35648 ;
  assign n35669 = n35630 & ~n35647 ;
  assign n35670 = ~n35668 & ~n35669 ;
  assign n35671 = ~\wishbone_RxDataLatched1_reg[22]/NET0131  & ~n35648 ;
  assign n35672 = n35635 & ~n35647 ;
  assign n35673 = ~n35671 & ~n35672 ;
  assign n35674 = ~\wishbone_RxDataLatched1_reg[23]/NET0131  & ~n35648 ;
  assign n35675 = n35640 & ~n35647 ;
  assign n35676 = ~n35674 & ~n35675 ;
  assign n35677 = n35609 & n35644 ;
  assign n35678 = \rxethmac1_RxStartFrm_reg/NET0131  & n32967 ;
  assign n35679 = ~n35677 & ~n35678 ;
  assign n35680 = n35607 & ~n35679 ;
  assign n35681 = ~\wishbone_RxDataLatched1_reg[24]/NET0131  & ~n35680 ;
  assign n35682 = n35651 & ~n35679 ;
  assign n35683 = ~n35681 & ~n35682 ;
  assign n35684 = ~\wishbone_RxDataLatched1_reg[25]/NET0131  & ~n35680 ;
  assign n35685 = n35656 & ~n35679 ;
  assign n35686 = ~n35684 & ~n35685 ;
  assign n35687 = ~\wishbone_RxDataLatched1_reg[26]/NET0131  & ~n35680 ;
  assign n35688 = n35615 & ~n35679 ;
  assign n35689 = ~n35687 & ~n35688 ;
  assign n35690 = ~\wishbone_RxDataLatched1_reg[27]/NET0131  & ~n35680 ;
  assign n35691 = n35620 & ~n35679 ;
  assign n35692 = ~n35690 & ~n35691 ;
  assign n35693 = ~\wishbone_RxDataLatched1_reg[28]/NET0131  & ~n35680 ;
  assign n35694 = n35625 & ~n35679 ;
  assign n35695 = ~n35693 & ~n35694 ;
  assign n35696 = ~\wishbone_RxDataLatched1_reg[29]/NET0131  & ~n35680 ;
  assign n35697 = n35630 & ~n35679 ;
  assign n35698 = ~n35696 & ~n35697 ;
  assign n35699 = ~\wishbone_RxDataLatched1_reg[30]/NET0131  & ~n35680 ;
  assign n35700 = n35635 & ~n35679 ;
  assign n35701 = ~n35699 & ~n35700 ;
  assign n35702 = ~\wishbone_RxDataLatched1_reg[31]/NET0131  & ~n35680 ;
  assign n35703 = n35640 & ~n35679 ;
  assign n35704 = ~n35702 & ~n35703 ;
  assign n35705 = ~\wishbone_RxDataLatched1_reg[8]/NET0131  & ~n35612 ;
  assign n35706 = ~n35611 & n35651 ;
  assign n35707 = ~n35705 & ~n35706 ;
  assign n35708 = ~\wishbone_RxDataLatched1_reg[9]/NET0131  & ~n35612 ;
  assign n35709 = ~n35611 & n35656 ;
  assign n35710 = ~n35708 & ~n35709 ;
  assign n35711 = \miim1_LatchByte0_d_reg/NET0131  & ~n35338 ;
  assign n35712 = n35427 & n35438 ;
  assign n35713 = n35338 & n35712 ;
  assign n35714 = ~n35711 & ~n35713 ;
  assign n35715 = \wishbone_rx_burst_cnt_reg[1]/NET0131  & ~n13191 ;
  assign n35716 = n32430 & n35715 ;
  assign n35717 = ~n13144 & ~n35345 ;
  assign n35718 = ~n13149 & n35717 ;
  assign n35719 = n13143 & n35718 ;
  assign n35720 = n13137 & n35719 ;
  assign n35721 = ~n35716 & ~n35720 ;
  assign n35722 = \wishbone_rx_burst_cnt_reg[2]/NET0131  & ~n13191 ;
  assign n35723 = n32430 & n35722 ;
  assign n35724 = \wishbone_rx_burst_cnt_reg[2]/NET0131  & ~n35345 ;
  assign n35725 = ~n35346 & ~n35724 ;
  assign n35726 = ~n13149 & ~n35725 ;
  assign n35727 = n13143 & n35726 ;
  assign n35728 = n13137 & n35727 ;
  assign n35729 = ~n35723 & ~n35728 ;
  assign n35730 = ~\wishbone_tx_fifo_write_pointer_reg[0]/NET0131  & \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n35731 = \wishbone_tx_fifo_cnt_reg[4]/NET0131  & n35314 ;
  assign n35732 = \wishbone_tx_fifo_write_pointer_reg[1]/NET0131  & ~\wishbone_tx_fifo_write_pointer_reg[2]/NET0131  ;
  assign n35733 = n14049 & n34242 ;
  assign n35734 = n35732 & n35733 ;
  assign n35735 = ~n35731 & n35734 ;
  assign n35736 = n35730 & n35735 ;
  assign n35737 = ~\wishbone_tx_fifo_write_pointer_reg[1]/NET0131  & \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  ;
  assign n35738 = n35733 & n35737 ;
  assign n35739 = ~n35731 & n35738 ;
  assign n35740 = n35730 & n35739 ;
  assign n35741 = \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  & \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n35742 = n35739 & n35741 ;
  assign n35743 = \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  & n14049 ;
  assign n35744 = ~\wishbone_tx_fifo_write_pointer_reg[1]/NET0131  & ~\wishbone_tx_fifo_write_pointer_reg[2]/NET0131  ;
  assign n35745 = n35743 & n35744 ;
  assign n35746 = ~n35731 & n35745 ;
  assign n35747 = ~\wishbone_tx_fifo_write_pointer_reg[3]/NET0131  & n34242 ;
  assign n35748 = n35746 & n35747 ;
  assign n35749 = ~\wishbone_tx_fifo_write_pointer_reg[0]/NET0131  & ~\wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n35750 = n35735 & n35749 ;
  assign n35751 = \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  & ~\wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n35752 = n35735 & n35751 ;
  assign n35753 = n35739 & n35749 ;
  assign n35754 = n35739 & n35751 ;
  assign n35755 = n14049 & n35749 ;
  assign n35756 = \wishbone_tx_fifo_write_pointer_reg[1]/NET0131  & \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  ;
  assign n35757 = n34242 & n35756 ;
  assign n35758 = n35755 & n35757 ;
  assign n35759 = ~n35731 & n35758 ;
  assign n35760 = \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  & \wishbone_tx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n35761 = n14049 & n35760 ;
  assign n35762 = ~n35731 & n35761 ;
  assign n35763 = \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  & ~\wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n35764 = n34242 & n35763 ;
  assign n35765 = n35762 & n35764 ;
  assign n35766 = n34242 & n35744 ;
  assign n35767 = n14049 & n35741 ;
  assign n35768 = n35766 & n35767 ;
  assign n35769 = ~n35731 & n35768 ;
  assign n35770 = ~\wishbone_rx_burst_cnt_reg[0]/NET0131  & n13191 ;
  assign n35771 = \wishbone_rx_burst_cnt_reg[0]/NET0131  & ~n13191 ;
  assign n35772 = n32430 & n35771 ;
  assign n35773 = ~n35770 & ~n35772 ;
  assign n35774 = n35298 & ~n35302 ;
  assign n35775 = n35301 & n35774 ;
  assign n35776 = \wishbone_tx_fifo_cnt_reg[2]/NET0131  & n35310 ;
  assign n35777 = ~n35298 & n35776 ;
  assign n35778 = ~n35775 & ~n35777 ;
  assign n35779 = \wishbone_tx_fifo_cnt_reg[3]/NET0131  & ~n35778 ;
  assign n35780 = ~n35309 & n35779 ;
  assign n35781 = \wishbone_tx_fifo_cnt_reg[3]/NET0131  & n34242 ;
  assign n35782 = n34242 & ~n35778 ;
  assign n35783 = ~n35309 & n35782 ;
  assign n35784 = ~n35781 & ~n35783 ;
  assign n35785 = ~n35780 & ~n35784 ;
  assign n35786 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  & ~n35531 ;
  assign n35787 = ~n35528 & n35786 ;
  assign n35788 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  & n35538 ;
  assign n35789 = ~n35531 & n35538 ;
  assign n35790 = ~n35528 & n35789 ;
  assign n35791 = ~n35788 & ~n35790 ;
  assign n35792 = ~n35787 & ~n35791 ;
  assign n35793 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n35794 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  & ~n35531 ;
  assign n35795 = ~n35528 & n35794 ;
  assign n35796 = ~n35793 & ~n35795 ;
  assign n35797 = ~n35534 & n35538 ;
  assign n35798 = n35796 & n35797 ;
  assign n35799 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  & ~n35541 ;
  assign n35800 = \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  ;
  assign n35801 = n35533 & n35800 ;
  assign n35802 = ~n35532 & n35801 ;
  assign n35803 = n35538 & ~n35802 ;
  assign n35804 = ~n35799 & n35803 ;
  assign n35805 = \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  & \txethmac1_txstatem1_StateData_reg[1]/NET0131  ;
  assign n35806 = n11296 & n35805 ;
  assign n35807 = ~\txethmac1_PacketFinished_q_reg/NET0131  & ~n35806 ;
  assign n35808 = ~n11171 & n35807 ;
  assign n35809 = \txethmac1_txstatem1_StateData_reg[1]/NET0131  & ~n11297 ;
  assign n35810 = ~n11166 & ~n35809 ;
  assign n35811 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  ;
  assign n35812 = ~n35810 & n35811 ;
  assign n35813 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & ~n35810 ;
  assign n35814 = ~\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  & ~n35813 ;
  assign n35815 = ~n35812 & ~n35814 ;
  assign n35816 = n35808 & n35815 ;
  assign n35817 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131  ;
  assign n35818 = \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  & n35817 ;
  assign n35819 = ~n35810 & n35818 ;
  assign n35820 = \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  & n35819 ;
  assign n35821 = ~\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  & ~n35819 ;
  assign n35822 = n35808 & ~n35821 ;
  assign n35823 = ~n35820 & n35822 ;
  assign n35824 = ~n35369 & ~n35373 ;
  assign n35825 = \wishbone_rx_fifo_cnt_reg[3]/NET0131  & ~n35824 ;
  assign n35826 = ~n35368 & n35825 ;
  assign n35827 = \wishbone_rx_fifo_cnt_reg[3]/NET0131  & ~n33164 ;
  assign n35828 = ~n33164 & ~n35824 ;
  assign n35829 = ~n35368 & n35828 ;
  assign n35830 = ~n35827 & ~n35829 ;
  assign n35831 = ~n35826 & ~n35830 ;
  assign n35832 = n32819 & n32821 ;
  assign n35833 = n23733 & n35832 ;
  assign n35834 = n32818 & n35833 ;
  assign n35835 = ~\wb_dat_i[1]_pad  & n25057 ;
  assign n35836 = n35834 & n35835 ;
  assign n35837 = \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131  & ~\miim1_RStatStart_reg/NET0131  ;
  assign n35838 = ~\miim1_RStatStart_reg/NET0131  & n25057 ;
  assign n35839 = n35834 & n35838 ;
  assign n35840 = ~n35837 & ~n35839 ;
  assign n35841 = ~n35836 & ~n35840 ;
  assign n35842 = ~\wb_dat_i[2]_pad  & n25057 ;
  assign n35843 = n35834 & n35842 ;
  assign n35844 = \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131  & ~\miim1_WCtrlDataStart_reg/NET0131  ;
  assign n35845 = ~\miim1_WCtrlDataStart_reg/NET0131  & n25057 ;
  assign n35846 = n35834 & n35845 ;
  assign n35847 = ~n35844 & ~n35846 ;
  assign n35848 = ~n35843 & ~n35847 ;
  assign n35849 = ~n35526 & ~n35531 ;
  assign n35850 = n35520 & n35849 ;
  assign n35851 = \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  & n35538 ;
  assign n35852 = ~n35850 & n35851 ;
  assign n35853 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  & n35538 ;
  assign n35854 = n35850 & n35853 ;
  assign n35855 = ~n35852 & ~n35854 ;
  assign n35856 = \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & n35538 ;
  assign n35857 = ~n35802 & n35856 ;
  assign n35858 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & n35538 ;
  assign n35859 = n35802 & n35858 ;
  assign n35860 = ~n35857 & ~n35859 ;
  assign n35861 = ~n10986 & ~n35570 ;
  assign n35862 = n11008 & ~n35570 ;
  assign n35863 = n10984 & n35862 ;
  assign n35864 = ~n35861 & ~n35863 ;
  assign n35865 = ~\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131  & ~n35812 ;
  assign n35866 = n35808 & ~n35819 ;
  assign n35867 = ~n35865 & n35866 ;
  assign n35868 = \wishbone_MasterWbTX_reg/NET0131  & ~\wishbone_TxAbortPacket_NotCleared_reg/NET0131  ;
  assign n35869 = ~\wishbone_TxRetryPacket_NotCleared_reg/NET0131  & ~\wishbone_cyc_cleared_reg/NET0131  ;
  assign n35870 = n35868 & n35869 ;
  assign n35871 = n35311 & n35870 ;
  assign n35872 = \wishbone_TxLength_reg[2]/NET0131  & ~n17372 ;
  assign n35873 = ~\wishbone_TxLength_reg[3]/NET0131  & ~\wishbone_TxLength_reg[4]/NET0131  ;
  assign n35874 = ~n35872 & n35873 ;
  assign n35875 = n35870 & n35874 ;
  assign n35876 = n32475 & n35875 ;
  assign n35877 = ~n35871 & ~n35876 ;
  assign n35878 = \wishbone_BlockReadTxDataFromMemory_reg/NET0131  & ~\wishbone_TxDonePacket_reg/NET0131  ;
  assign n35879 = n34242 & n35878 ;
  assign n35880 = ~n35298 & n35879 ;
  assign n35881 = n35877 & ~n35880 ;
  assign n35882 = \miim1_InProgress_q1_reg/NET0131  & ~n35338 ;
  assign n35883 = ~n35328 & ~n35882 ;
  assign n35884 = ~\rxethmac1_RxEndFrm_d_reg/NET0131  & ~n12164 ;
  assign n35885 = ~\rxethmac1_RxEndFrm_d_reg/NET0131  & ~n12580 ;
  assign n35886 = n10525 & n35885 ;
  assign n35887 = ~n35884 & ~n35886 ;
  assign n35888 = \wb_adr_i[2]_pad  & n32819 ;
  assign n35889 = n23733 & n35888 ;
  assign n35890 = n32818 & n35889 ;
  assign n35891 = \wb_dat_i[2]_pad  & n23751 ;
  assign n35892 = n35890 & n35891 ;
  assign n35893 = \ethreg1_irq_rxb_reg/NET0131  & ~n35892 ;
  assign n35894 = ~\wishbone_RxB_IRQ_reg/NET0131  & ~n35893 ;
  assign n35895 = \wb_dat_i[6]_pad  & n23751 ;
  assign n35896 = n35890 & n35895 ;
  assign n35897 = \ethreg1_irq_rxc_reg/NET0131  & ~n35896 ;
  assign n35898 = ~\ethreg1_SetRxCIrq_reg/NET0131  & ~n35897 ;
  assign n35899 = \wb_dat_i[3]_pad  & n23751 ;
  assign n35900 = n35890 & n35899 ;
  assign n35901 = \ethreg1_irq_rxe_reg/NET0131  & ~n35900 ;
  assign n35902 = ~\wishbone_RxE_IRQ_reg/NET0131  & ~n35901 ;
  assign n35903 = \wb_dat_i[0]_pad  & n23751 ;
  assign n35904 = n35890 & n35903 ;
  assign n35905 = \ethreg1_irq_txb_reg/NET0131  & ~n35904 ;
  assign n35906 = ~\wishbone_TxB_IRQ_reg/NET0131  & ~n35905 ;
  assign n35907 = \wb_dat_i[5]_pad  & n23751 ;
  assign n35908 = n35890 & n35907 ;
  assign n35909 = \ethreg1_irq_txc_reg/NET0131  & ~n35908 ;
  assign n35910 = ~\ethreg1_SetTxCIrq_reg/NET0131  & ~n35909 ;
  assign n35911 = \wb_dat_i[1]_pad  & n23751 ;
  assign n35912 = n35890 & n35911 ;
  assign n35913 = \ethreg1_irq_txe_reg/NET0131  & ~n35912 ;
  assign n35914 = ~\wishbone_TxE_IRQ_reg/NET0131  & ~n35913 ;
  assign n35915 = \txethmac1_ColWindow_reg/NET0131  & ~n11164 ;
  assign n35916 = ~n11086 & n35915 ;
  assign n35917 = n11171 & n35916 ;
  assign n35918 = ~\txethmac1_TxRetry_reg/NET0131  & ~n35917 ;
  assign n35919 = n11567 & ~n35918 ;
  assign n35920 = ~\wishbone_RxReady_reg/NET0131  & n15726 ;
  assign n35921 = \wishbone_Busy_IRQ_rck_reg/NET0131  & ~\wishbone_Busy_IRQ_syncb2_reg/P0001  ;
  assign n35922 = ~n35920 & ~n35921 ;
  assign n35923 = \wishbone_RxBDAddress_reg[1]/NET0131  & \wishbone_ShiftEnded_reg/NET0131  ;
  assign n35924 = n15779 & n35923 ;
  assign n35925 = \wishbone_RxBDAddress_reg[2]/NET0131  & n35924 ;
  assign n35926 = ~\wishbone_RxBDAddress_reg[3]/NET0131  & ~n35925 ;
  assign n35927 = n35448 & ~n35453 ;
  assign n35928 = ~n35926 & n35927 ;
  assign n35929 = \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131  & ~n35448 ;
  assign n35930 = ~n35928 & ~n35929 ;
  assign n35931 = ~\wishbone_RxBDAddress_reg[5]/NET0131  & ~n35457 ;
  assign n35932 = \wishbone_RxBDAddress_reg[5]/NET0131  & n35457 ;
  assign n35933 = n35448 & ~n35932 ;
  assign n35934 = ~n35931 & n35933 ;
  assign n35935 = \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131  & ~n35448 ;
  assign n35936 = ~n35934 & ~n35935 ;
  assign n35937 = \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131  & ~n35448 ;
  assign n35938 = \wishbone_RxBDAddress_reg[6]/NET0131  & ~n35450 ;
  assign n35939 = n35452 & n35599 ;
  assign n35940 = ~\wishbone_RxStatus_reg[13]/NET0131  & ~n35939 ;
  assign n35941 = ~n35938 & ~n35940 ;
  assign n35942 = ~\wishbone_RxBDAddress_reg[6]/NET0131  & ~n35938 ;
  assign n35943 = ~n35932 & n35942 ;
  assign n35944 = ~n35941 & ~n35943 ;
  assign n35945 = ~n35445 & n35944 ;
  assign n35946 = ~n35937 & ~n35945 ;
  assign n35947 = \miim1_clkgen_Counter_reg[5]/NET0131  & ~n32250 ;
  assign n35948 = ~n35493 & ~n35947 ;
  assign n35949 = \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  & ~n32261 ;
  assign n35950 = n32264 & ~n35497 ;
  assign n35951 = ~n35949 & n35950 ;
  assign n35952 = ~n35948 & ~n35951 ;
  assign n35953 = n14049 & n35732 ;
  assign n35954 = ~n35731 & n35953 ;
  assign n35955 = n14049 & ~n34242 ;
  assign n35956 = n35730 & ~n35955 ;
  assign n35957 = n35954 & n35956 ;
  assign n35958 = \wishbone_tx_fifo_fifo_reg[10][14]/P0001  & ~n35957 ;
  assign n35959 = \m_wb_dat_i[14]_pad  & n35956 ;
  assign n35960 = n35954 & n35959 ;
  assign n35961 = ~n35958 & ~n35960 ;
  assign n35962 = \wishbone_tx_fifo_fifo_reg[10][18]/P0001  & ~n35957 ;
  assign n35963 = \m_wb_dat_i[18]_pad  & n35956 ;
  assign n35964 = n35954 & n35963 ;
  assign n35965 = ~n35962 & ~n35964 ;
  assign n35966 = \wishbone_tx_fifo_fifo_reg[10][27]/P0001  & ~n35957 ;
  assign n35967 = \m_wb_dat_i[27]_pad  & n35956 ;
  assign n35968 = n35954 & n35967 ;
  assign n35969 = ~n35966 & ~n35968 ;
  assign n35970 = \wishbone_tx_fifo_fifo_reg[10][29]/P0001  & ~n35957 ;
  assign n35971 = \m_wb_dat_i[29]_pad  & n35956 ;
  assign n35972 = n35954 & n35971 ;
  assign n35973 = ~n35970 & ~n35972 ;
  assign n35974 = \wishbone_tx_fifo_fifo_reg[10][3]/P0001  & ~n35957 ;
  assign n35975 = \m_wb_dat_i[3]_pad  & n35956 ;
  assign n35976 = n35954 & n35975 ;
  assign n35977 = ~n35974 & ~n35976 ;
  assign n35978 = n14049 & n35737 ;
  assign n35979 = ~n35731 & n35978 ;
  assign n35980 = n35956 & n35979 ;
  assign n35981 = \wishbone_tx_fifo_fifo_reg[12][12]/P0001  & ~n35980 ;
  assign n35982 = \m_wb_dat_i[12]_pad  & n35956 ;
  assign n35983 = n35979 & n35982 ;
  assign n35984 = ~n35981 & ~n35983 ;
  assign n35985 = \wishbone_tx_fifo_fifo_reg[12][14]/P0001  & ~n35980 ;
  assign n35986 = n35959 & n35979 ;
  assign n35987 = ~n35985 & ~n35986 ;
  assign n35988 = \wishbone_tx_fifo_fifo_reg[12][18]/P0001  & ~n35980 ;
  assign n35989 = n35963 & n35979 ;
  assign n35990 = ~n35988 & ~n35989 ;
  assign n35991 = \wishbone_tx_fifo_fifo_reg[12][22]/P0001  & ~n35980 ;
  assign n35992 = \m_wb_dat_i[22]_pad  & n35956 ;
  assign n35993 = n35979 & n35992 ;
  assign n35994 = ~n35991 & ~n35993 ;
  assign n35995 = \wishbone_tx_fifo_fifo_reg[12][25]/P0001  & ~n35980 ;
  assign n35996 = \m_wb_dat_i[25]_pad  & n35956 ;
  assign n35997 = n35979 & n35996 ;
  assign n35998 = ~n35995 & ~n35997 ;
  assign n35999 = \wishbone_tx_fifo_fifo_reg[12][27]/P0001  & ~n35980 ;
  assign n36000 = n35967 & n35979 ;
  assign n36001 = ~n35999 & ~n36000 ;
  assign n36002 = \wishbone_tx_fifo_fifo_reg[12][28]/P0001  & ~n35980 ;
  assign n36003 = \m_wb_dat_i[28]_pad  & n35956 ;
  assign n36004 = n35979 & n36003 ;
  assign n36005 = ~n36002 & ~n36004 ;
  assign n36006 = \wishbone_tx_fifo_fifo_reg[12][30]/P0001  & ~n35980 ;
  assign n36007 = \m_wb_dat_i[30]_pad  & n35956 ;
  assign n36008 = n35979 & n36007 ;
  assign n36009 = ~n36006 & ~n36008 ;
  assign n36010 = \wishbone_tx_fifo_fifo_reg[12][3]/P0001  & ~n35980 ;
  assign n36011 = n35975 & n35979 ;
  assign n36012 = ~n36010 & ~n36011 ;
  assign n36013 = \wishbone_tx_fifo_fifo_reg[12][6]/P0001  & ~n35980 ;
  assign n36014 = \m_wb_dat_i[6]_pad  & n35956 ;
  assign n36015 = n35979 & n36014 ;
  assign n36016 = ~n36013 & ~n36015 ;
  assign n36017 = n35751 & ~n35955 ;
  assign n36018 = n35954 & n36017 ;
  assign n36019 = \wishbone_tx_fifo_fifo_reg[3][10]/P0001  & ~n36018 ;
  assign n36020 = \m_wb_dat_i[10]_pad  & n36017 ;
  assign n36021 = n35954 & n36020 ;
  assign n36022 = ~n36019 & ~n36021 ;
  assign n36023 = \wishbone_tx_fifo_fifo_reg[3][11]/P0001  & ~n36018 ;
  assign n36024 = \m_wb_dat_i[11]_pad  & n36017 ;
  assign n36025 = n35954 & n36024 ;
  assign n36026 = ~n36023 & ~n36025 ;
  assign n36027 = \wishbone_tx_fifo_fifo_reg[3][13]/P0001  & ~n36018 ;
  assign n36028 = \m_wb_dat_i[13]_pad  & n36017 ;
  assign n36029 = n35954 & n36028 ;
  assign n36030 = ~n36027 & ~n36029 ;
  assign n36031 = \wishbone_tx_fifo_fifo_reg[3][18]/P0001  & ~n36018 ;
  assign n36032 = \m_wb_dat_i[18]_pad  & n36017 ;
  assign n36033 = n35954 & n36032 ;
  assign n36034 = ~n36031 & ~n36033 ;
  assign n36035 = \wishbone_tx_fifo_fifo_reg[3][19]/P0001  & ~n36018 ;
  assign n36036 = \m_wb_dat_i[19]_pad  & n36017 ;
  assign n36037 = n35954 & n36036 ;
  assign n36038 = ~n36035 & ~n36037 ;
  assign n36039 = \wishbone_tx_fifo_fifo_reg[3][25]/P0001  & ~n36018 ;
  assign n36040 = \m_wb_dat_i[25]_pad  & n36017 ;
  assign n36041 = n35954 & n36040 ;
  assign n36042 = ~n36039 & ~n36041 ;
  assign n36043 = \wishbone_tx_fifo_fifo_reg[3][29]/P0001  & ~n36018 ;
  assign n36044 = \m_wb_dat_i[29]_pad  & n36017 ;
  assign n36045 = n35954 & n36044 ;
  assign n36046 = ~n36043 & ~n36045 ;
  assign n36047 = \wishbone_tx_fifo_fifo_reg[3][31]/P0001  & ~n36018 ;
  assign n36048 = \m_wb_dat_i[31]_pad  & n36017 ;
  assign n36049 = n35954 & n36048 ;
  assign n36050 = ~n36047 & ~n36049 ;
  assign n36051 = \wishbone_tx_fifo_fifo_reg[3][4]/P0001  & ~n36018 ;
  assign n36052 = \m_wb_dat_i[4]_pad  & n36017 ;
  assign n36053 = n35954 & n36052 ;
  assign n36054 = ~n36051 & ~n36053 ;
  assign n36055 = \wishbone_tx_fifo_fifo_reg[3][5]/P0001  & ~n36018 ;
  assign n36056 = \m_wb_dat_i[5]_pad  & n36017 ;
  assign n36057 = n35954 & n36056 ;
  assign n36058 = ~n36055 & ~n36057 ;
  assign n36059 = \wishbone_tx_fifo_fifo_reg[3][8]/P0001  & ~n36018 ;
  assign n36060 = \m_wb_dat_i[8]_pad  & n36017 ;
  assign n36061 = n35954 & n36060 ;
  assign n36062 = ~n36059 & ~n36061 ;
  assign n36063 = n35979 & n36017 ;
  assign n36064 = \wishbone_tx_fifo_fifo_reg[5][11]/P0001  & ~n36063 ;
  assign n36065 = n35979 & n36024 ;
  assign n36066 = ~n36064 & ~n36065 ;
  assign n36067 = \wishbone_tx_fifo_fifo_reg[5][18]/P0001  & ~n36063 ;
  assign n36068 = n35979 & n36032 ;
  assign n36069 = ~n36067 & ~n36068 ;
  assign n36070 = \wishbone_tx_fifo_fifo_reg[5][19]/P0001  & ~n36063 ;
  assign n36071 = n35979 & n36036 ;
  assign n36072 = ~n36070 & ~n36071 ;
  assign n36073 = \wishbone_tx_fifo_fifo_reg[5][1]/P0001  & ~n36063 ;
  assign n36074 = \m_wb_dat_i[1]_pad  & n36017 ;
  assign n36075 = n35979 & n36074 ;
  assign n36076 = ~n36073 & ~n36075 ;
  assign n36077 = \wishbone_tx_fifo_fifo_reg[5][23]/P0001  & ~n36063 ;
  assign n36078 = \m_wb_dat_i[23]_pad  & n36017 ;
  assign n36079 = n35979 & n36078 ;
  assign n36080 = ~n36077 & ~n36079 ;
  assign n36081 = \wishbone_tx_fifo_fifo_reg[5][24]/P0001  & ~n36063 ;
  assign n36082 = \m_wb_dat_i[24]_pad  & n36017 ;
  assign n36083 = n35979 & n36082 ;
  assign n36084 = ~n36081 & ~n36083 ;
  assign n36085 = \wishbone_tx_fifo_fifo_reg[5][25]/P0001  & ~n36063 ;
  assign n36086 = n35979 & n36040 ;
  assign n36087 = ~n36085 & ~n36086 ;
  assign n36088 = \wishbone_tx_fifo_fifo_reg[5][26]/P0001  & ~n36063 ;
  assign n36089 = \m_wb_dat_i[26]_pad  & n36017 ;
  assign n36090 = n35979 & n36089 ;
  assign n36091 = ~n36088 & ~n36090 ;
  assign n36092 = \wishbone_tx_fifo_fifo_reg[5][28]/P0001  & ~n36063 ;
  assign n36093 = \m_wb_dat_i[28]_pad  & n36017 ;
  assign n36094 = n35979 & n36093 ;
  assign n36095 = ~n36092 & ~n36094 ;
  assign n36096 = \wishbone_tx_fifo_fifo_reg[5][3]/P0001  & ~n36063 ;
  assign n36097 = \m_wb_dat_i[3]_pad  & n36017 ;
  assign n36098 = n35979 & n36097 ;
  assign n36099 = ~n36096 & ~n36098 ;
  assign n36100 = \wishbone_tx_fifo_fifo_reg[5][8]/P0001  & ~n36063 ;
  assign n36101 = n35979 & n36060 ;
  assign n36102 = ~n36100 & ~n36101 ;
  assign n36103 = ~n35731 & n35755 ;
  assign n36104 = n35756 & ~n35955 ;
  assign n36105 = n36103 & n36104 ;
  assign n36106 = \wishbone_tx_fifo_fifo_reg[6][11]/P0001  & ~n36105 ;
  assign n36107 = \m_wb_dat_i[11]_pad  & n36104 ;
  assign n36108 = n36103 & n36107 ;
  assign n36109 = ~n36106 & ~n36108 ;
  assign n36110 = \wishbone_tx_fifo_fifo_reg[6][12]/P0001  & ~n36105 ;
  assign n36111 = \m_wb_dat_i[12]_pad  & n36104 ;
  assign n36112 = n36103 & n36111 ;
  assign n36113 = ~n36110 & ~n36112 ;
  assign n36114 = \wishbone_tx_fifo_fifo_reg[6][14]/P0001  & ~n36105 ;
  assign n36115 = \m_wb_dat_i[14]_pad  & n36104 ;
  assign n36116 = n36103 & n36115 ;
  assign n36117 = ~n36114 & ~n36116 ;
  assign n36118 = \wishbone_tx_fifo_fifo_reg[6][16]/P0001  & ~n36105 ;
  assign n36119 = \m_wb_dat_i[16]_pad  & n36104 ;
  assign n36120 = n36103 & n36119 ;
  assign n36121 = ~n36118 & ~n36120 ;
  assign n36122 = \wishbone_tx_fifo_fifo_reg[6][18]/P0001  & ~n36105 ;
  assign n36123 = \m_wb_dat_i[18]_pad  & n36104 ;
  assign n36124 = n36103 & n36123 ;
  assign n36125 = ~n36122 & ~n36124 ;
  assign n36126 = \wishbone_tx_fifo_fifo_reg[6][1]/P0001  & ~n36105 ;
  assign n36127 = \m_wb_dat_i[1]_pad  & n36104 ;
  assign n36128 = n36103 & n36127 ;
  assign n36129 = ~n36126 & ~n36128 ;
  assign n36130 = \wishbone_tx_fifo_fifo_reg[6][20]/P0001  & ~n36105 ;
  assign n36131 = \m_wb_dat_i[20]_pad  & n36104 ;
  assign n36132 = n36103 & n36131 ;
  assign n36133 = ~n36130 & ~n36132 ;
  assign n36134 = \wishbone_tx_fifo_fifo_reg[6][25]/P0001  & ~n36105 ;
  assign n36135 = \m_wb_dat_i[25]_pad  & n36104 ;
  assign n36136 = n36103 & n36135 ;
  assign n36137 = ~n36134 & ~n36136 ;
  assign n36138 = \wishbone_tx_fifo_fifo_reg[6][27]/P0001  & ~n36105 ;
  assign n36139 = \m_wb_dat_i[27]_pad  & n36104 ;
  assign n36140 = n36103 & n36139 ;
  assign n36141 = ~n36138 & ~n36140 ;
  assign n36142 = \wishbone_tx_fifo_fifo_reg[6][28]/P0001  & ~n36105 ;
  assign n36143 = \m_wb_dat_i[28]_pad  & n36104 ;
  assign n36144 = n36103 & n36143 ;
  assign n36145 = ~n36142 & ~n36144 ;
  assign n36146 = \wishbone_tx_fifo_fifo_reg[6][30]/P0001  & ~n36105 ;
  assign n36147 = \m_wb_dat_i[30]_pad  & n36104 ;
  assign n36148 = n36103 & n36147 ;
  assign n36149 = ~n36146 & ~n36148 ;
  assign n36150 = \wishbone_tx_fifo_fifo_reg[6][3]/P0001  & ~n36105 ;
  assign n36151 = \m_wb_dat_i[3]_pad  & n36104 ;
  assign n36152 = n36103 & n36151 ;
  assign n36153 = ~n36150 & ~n36152 ;
  assign n36154 = \wishbone_tx_fifo_fifo_reg[6][4]/P0001  & ~n36105 ;
  assign n36155 = \m_wb_dat_i[4]_pad  & n36104 ;
  assign n36156 = n36103 & n36155 ;
  assign n36157 = ~n36154 & ~n36156 ;
  assign n36158 = \wishbone_tx_fifo_fifo_reg[6][5]/P0001  & ~n36105 ;
  assign n36159 = \m_wb_dat_i[5]_pad  & n36104 ;
  assign n36160 = n36103 & n36159 ;
  assign n36161 = ~n36158 & ~n36160 ;
  assign n36162 = \wishbone_tx_fifo_fifo_reg[6][6]/P0001  & ~n36105 ;
  assign n36163 = \m_wb_dat_i[6]_pad  & n36104 ;
  assign n36164 = n36103 & n36163 ;
  assign n36165 = ~n36162 & ~n36164 ;
  assign n36166 = \wishbone_tx_fifo_fifo_reg[6][7]/P0001  & ~n36105 ;
  assign n36167 = \m_wb_dat_i[7]_pad  & n36104 ;
  assign n36168 = n36103 & n36167 ;
  assign n36169 = ~n36166 & ~n36168 ;
  assign n36170 = \wishbone_tx_fifo_fifo_reg[6][8]/P0001  & ~n36105 ;
  assign n36171 = \m_wb_dat_i[8]_pad  & n36104 ;
  assign n36172 = n36103 & n36171 ;
  assign n36173 = ~n36170 & ~n36172 ;
  assign n36174 = \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  & ~n35955 ;
  assign n36175 = n35746 & n36174 ;
  assign n36176 = \wishbone_tx_fifo_fifo_reg[9][12]/P0001  & ~n36175 ;
  assign n36177 = \m_wb_dat_i[12]_pad  & n36174 ;
  assign n36178 = n35746 & n36177 ;
  assign n36179 = ~n36176 & ~n36178 ;
  assign n36180 = \wishbone_tx_fifo_fifo_reg[9][13]/P0001  & ~n36175 ;
  assign n36181 = \m_wb_dat_i[13]_pad  & n36174 ;
  assign n36182 = n35746 & n36181 ;
  assign n36183 = ~n36180 & ~n36182 ;
  assign n36184 = \wishbone_tx_fifo_fifo_reg[9][14]/P0001  & ~n36175 ;
  assign n36185 = \m_wb_dat_i[14]_pad  & n36174 ;
  assign n36186 = n35746 & n36185 ;
  assign n36187 = ~n36184 & ~n36186 ;
  assign n36188 = \wishbone_tx_fifo_fifo_reg[9][20]/P0001  & ~n36175 ;
  assign n36189 = \m_wb_dat_i[20]_pad  & n36174 ;
  assign n36190 = n35746 & n36189 ;
  assign n36191 = ~n36188 & ~n36190 ;
  assign n36192 = \wishbone_tx_fifo_fifo_reg[9][25]/P0001  & ~n36175 ;
  assign n36193 = \m_wb_dat_i[25]_pad  & n36174 ;
  assign n36194 = n35746 & n36193 ;
  assign n36195 = ~n36192 & ~n36194 ;
  assign n36196 = \wishbone_tx_fifo_fifo_reg[9][26]/P0001  & ~n36175 ;
  assign n36197 = \m_wb_dat_i[26]_pad  & n36174 ;
  assign n36198 = n35746 & n36197 ;
  assign n36199 = ~n36196 & ~n36198 ;
  assign n36200 = \wishbone_tx_fifo_fifo_reg[9][30]/P0001  & ~n36175 ;
  assign n36201 = \m_wb_dat_i[30]_pad  & n36174 ;
  assign n36202 = n35746 & n36201 ;
  assign n36203 = ~n36200 & ~n36202 ;
  assign n36204 = \wishbone_tx_fifo_fifo_reg[9][5]/P0001  & ~n36175 ;
  assign n36205 = \m_wb_dat_i[5]_pad  & n36174 ;
  assign n36206 = n35746 & n36205 ;
  assign n36207 = ~n36204 & ~n36206 ;
  assign n36208 = \wishbone_tx_fifo_fifo_reg[9][8]/P0001  & ~n36175 ;
  assign n36209 = \m_wb_dat_i[8]_pad  & n36174 ;
  assign n36210 = n35746 & n36209 ;
  assign n36211 = ~n36208 & ~n36210 ;
  assign n36212 = \wishbone_tx_fifo_fifo_reg[6][23]/P0001  & ~n36105 ;
  assign n36213 = \m_wb_dat_i[23]_pad  & n36104 ;
  assign n36214 = n36103 & n36213 ;
  assign n36215 = ~n36212 & ~n36214 ;
  assign n36216 = n14049 & n35744 ;
  assign n36217 = n35749 & n36216 ;
  assign n36218 = ~n35731 & n36217 ;
  assign n36219 = ~n35955 & ~n36218 ;
  assign n36220 = n35735 & n35741 ;
  assign n36221 = n14049 & n35730 ;
  assign n36222 = n35757 & n36221 ;
  assign n36223 = ~n35731 & n36222 ;
  assign n36224 = n35757 & n35767 ;
  assign n36225 = ~n35731 & n36224 ;
  assign n36226 = n35766 & n36221 ;
  assign n36227 = ~n35731 & n36226 ;
  assign n36228 = \wishbone_Busy_IRQ_sync2_reg/P0001  & ~\wishbone_Busy_IRQ_sync3_reg/P0001  ;
  assign n36229 = \wb_dat_i[4]_pad  & n23751 ;
  assign n36230 = n35890 & n36229 ;
  assign n36231 = \ethreg1_irq_busy_reg/NET0131  & ~n36230 ;
  assign n36232 = ~n36228 & ~n36231 ;
  assign n36233 = ~\miim1_LatchByte_reg[0]/NET0131  & \miim1_LatchByte_reg[1]/NET0131  ;
  assign n36234 = n32545 & n36233 ;
  assign n36235 = n32531 & n36234 ;
  assign n36236 = n32513 & n36235 ;
  assign n36237 = \wishbone_rx_fifo_cnt_reg[0]/NET0131  & ~n33164 ;
  assign n36238 = n35368 & ~n36237 ;
  assign n36239 = ~n35368 & n36237 ;
  assign n36240 = ~n36238 & ~n36239 ;
  assign n36241 = \macstatus1_LoadRxStatus_reg/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n36242 = ~n11693 & n36241 ;
  assign n36243 = \macstatus1_LoadRxStatus_reg/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
  assign n36244 = n11693 & n36243 ;
  assign n36245 = ~n36242 & ~n36244 ;
  assign n36246 = ~\macstatus1_LoadRxStatus_reg/NET0131  & ~\wishbone_LatchedRxLength_reg[13]/NET0131  ;
  assign n36247 = n36245 & ~n36246 ;
  assign n36248 = ~\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  & ~n11674 ;
  assign n36249 = ~n11675 & ~n36248 ;
  assign n36250 = ~n11671 & ~n11723 ;
  assign n36251 = n10663 & ~n12178 ;
  assign n36252 = n10663 & ~n11635 ;
  assign n36253 = n11353 & n11362 ;
  assign n36254 = n10663 & ~n36253 ;
  assign n36255 = n35364 & ~n35371 ;
  assign n36256 = ~n13126 & ~n35367 ;
  assign n36257 = ~n36255 & ~n36256 ;
  assign n36258 = \wishbone_rx_fifo_cnt_reg[2]/NET0131  & ~n33164 ;
  assign n36259 = ~n36257 & n36258 ;
  assign n36260 = ~\wishbone_rx_fifo_cnt_reg[2]/NET0131  & ~n33164 ;
  assign n36261 = n36257 & n36260 ;
  assign n36262 = ~n36259 & ~n36261 ;
  assign n36263 = ~\rxethmac1_RxStartFrm_reg/NET0131  & ~\wishbone_LatchedRxStartFrm_reg/NET0131  ;
  assign n36264 = ~\wishbone_SyncRxStartFrm_q_reg/NET0131  & ~n36263 ;
  assign n36265 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  ;
  assign n36266 = \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  & \rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  ;
  assign n36267 = n36265 & n36266 ;
  assign n36268 = \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  & n36267 ;
  assign n36269 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & \rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
  assign n36270 = \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  & ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  ;
  assign n36271 = ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  & \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  ;
  assign n36272 = n36270 & n36271 ;
  assign n36273 = ~n36269 & ~n36272 ;
  assign n36274 = ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  & ~n36267 ;
  assign n36275 = n36273 & ~n36274 ;
  assign n36276 = ~n36268 & n36275 ;
  assign n36277 = \wishbone_rx_fifo_cnt_reg[1]/NET0131  & n35368 ;
  assign n36278 = ~n13126 & ~n35371 ;
  assign n36279 = ~n35364 & ~n36278 ;
  assign n36280 = n35366 & n36278 ;
  assign n36281 = ~n35365 & n36280 ;
  assign n36282 = ~n36279 & ~n36281 ;
  assign n36283 = ~n36277 & n36282 ;
  assign n36284 = ~n33164 & ~n36283 ;
  assign n36285 = \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  & \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131  ;
  assign n36286 = n11980 & n36285 ;
  assign n36287 = ~\maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131  & ~n36286 ;
  assign n36288 = ~wb_rst_i_pad & ~n11983 ;
  assign n36289 = ~n36287 & n36288 ;
  assign n36290 = \wishbone_StartOccured_reg/NET0131  & ~n35551 ;
  assign n36291 = n35550 & n36290 ;
  assign n36292 = ~\wishbone_TxStartFrm_wb_reg/NET0131  & ~n36291 ;
  assign n36293 = ~\ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131  & ~\ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131  ;
  assign n36294 = ~\ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131  & ~\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131  ;
  assign n36295 = n36293 & n36294 ;
  assign n36296 = ~\ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131  & ~\ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131  ;
  assign n36297 = ~\ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131  & ~\ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131  ;
  assign n36298 = n36296 & n36297 ;
  assign n36299 = n36295 & n36298 ;
  assign n36300 = \ethreg1_MODER_0_DataOut_reg[1]/NET0131  & ~\wishbone_r_TxEn_q_reg/NET0131  ;
  assign n36301 = ~n36299 & n36300 ;
  assign n36302 = ~\wishbone_TxAbortPacket_NotCleared_reg/NET0131  & ~\wishbone_TxDonePacket_NotCleared_reg/NET0131  ;
  assign n36303 = n14045 & ~n36302 ;
  assign n36304 = ~\wishbone_BlockingTxStatusWrite_reg/NET0131  & n36303 ;
  assign n36305 = \wishbone_TxBDAddress_reg[4]/NET0131  & ~n36304 ;
  assign n36306 = ~n36301 & n36305 ;
  assign n36307 = ~\wishbone_BlockingTxStatusWrite_reg/NET0131  & ~\wishbone_TxStatus_reg[13]/NET0131  ;
  assign n36308 = n36303 & n36307 ;
  assign n36309 = ~n36301 & n36308 ;
  assign n36310 = \wishbone_TxBDAddress_reg[1]/NET0131  & \wishbone_TxBDAddress_reg[2]/NET0131  ;
  assign n36311 = \wishbone_TxBDAddress_reg[3]/NET0131  & n36310 ;
  assign n36312 = ~\wishbone_TxBDAddress_reg[4]/NET0131  & ~n36311 ;
  assign n36313 = \wishbone_TxBDAddress_reg[3]/NET0131  & \wishbone_TxBDAddress_reg[4]/NET0131  ;
  assign n36314 = n36310 & n36313 ;
  assign n36315 = ~n36312 & ~n36314 ;
  assign n36316 = n36309 & n36315 ;
  assign n36317 = ~n36306 & ~n36316 ;
  assign n36318 = ~n36301 & ~n36304 ;
  assign n36319 = \wishbone_TxBDAddress_reg[5]/NET0131  & \wishbone_TxBDAddress_reg[6]/NET0131  ;
  assign n36320 = n36314 & n36319 ;
  assign n36321 = n36308 & ~n36320 ;
  assign n36322 = ~n36301 & n36321 ;
  assign n36323 = ~n36318 & ~n36322 ;
  assign n36324 = \wishbone_TxBDAddress_reg[6]/NET0131  & ~n36323 ;
  assign n36325 = \wishbone_TxBDAddress_reg[5]/NET0131  & n36314 ;
  assign n36326 = n36322 & n36325 ;
  assign n36327 = ~n36324 & ~n36326 ;
  assign n36328 = \wishbone_TxBDAddress_reg[7]/NET0131  & ~n36323 ;
  assign n36329 = \wishbone_TxBDAddress_reg[5]/NET0131  & ~\wishbone_TxBDAddress_reg[7]/NET0131  ;
  assign n36330 = \wishbone_TxBDAddress_reg[6]/NET0131  & n36329 ;
  assign n36331 = n36314 & n36330 ;
  assign n36332 = n36308 & n36331 ;
  assign n36333 = ~n36301 & n36332 ;
  assign n36334 = ~n36328 & ~n36333 ;
  assign n36335 = \wishbone_TxEndFrm_wb_reg/NET0131  & ~n35551 ;
  assign n36336 = n35550 & n36335 ;
  assign n36337 = n14063 & n17372 ;
  assign n36338 = n14058 & n36337 ;
  assign n36339 = \wishbone_tx_fifo_cnt_reg[0]/NET0131  & ~\wishbone_tx_fifo_cnt_reg[1]/NET0131  ;
  assign n36340 = ~\wishbone_tx_fifo_cnt_reg[2]/NET0131  & n36339 ;
  assign n36341 = n12725 & n35302 ;
  assign n36342 = n36340 & n36341 ;
  assign n36343 = n36338 & n36342 ;
  assign n36344 = ~n36336 & ~n36343 ;
  assign n36345 = \miim1_outctrl_Mdo_2d_reg/NET0131  & ~n32513 ;
  assign n36346 = ~\miim1_BitCounter_reg[4]/NET0131  & ~\miim1_BitCounter_reg[6]/NET0131  ;
  assign n36347 = ~\miim1_WriteOp_reg/NET0131  & ~n36346 ;
  assign n36348 = \miim1_BitCounter_reg[3]/NET0131  & ~\miim1_WriteOp_reg/NET0131  ;
  assign n36349 = n35589 & n36348 ;
  assign n36350 = ~n36347 & ~n36349 ;
  assign n36351 = \miim1_InProgress_reg/NET0131  & ~n32520 ;
  assign n36352 = n36350 & n36351 ;
  assign n36353 = ~n32523 & ~n36352 ;
  assign n36354 = mdc_pad_o_pad & n32520 ;
  assign n36355 = n32264 & n36354 ;
  assign n36356 = n36353 & n36355 ;
  assign n36357 = ~n36345 & ~n36356 ;
  assign n36358 = \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n36359 = n35523 & n36358 ;
  assign n36360 = \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  ;
  assign n36361 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & n36360 ;
  assign n36362 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  ;
  assign n36363 = \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n36364 = n36362 & n36363 ;
  assign n36365 = ~n36361 & ~n36364 ;
  assign n36366 = ~n36359 & n36365 ;
  assign n36367 = n35522 & ~n36366 ;
  assign n36368 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  ;
  assign n36369 = \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  & n36368 ;
  assign n36370 = \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n36371 = n36360 & n36370 ;
  assign n36372 = n36369 & n36371 ;
  assign n36373 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & n36362 ;
  assign n36374 = \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n36375 = n36368 & n36374 ;
  assign n36376 = n36373 & n36375 ;
  assign n36377 = ~n36372 & ~n36376 ;
  assign n36378 = ~n36367 & n36377 ;
  assign n36379 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  & n36368 ;
  assign n36380 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & n35523 ;
  assign n36381 = ~n35518 & n36380 ;
  assign n36382 = \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n36383 = n35523 & n36382 ;
  assign n36384 = \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n36385 = n36362 & n36384 ;
  assign n36386 = ~n36383 & ~n36385 ;
  assign n36387 = ~n36381 & n36386 ;
  assign n36388 = n36379 & ~n36387 ;
  assign n36389 = \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  & n35521 ;
  assign n36390 = \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n36391 = n36360 & n36390 ;
  assign n36392 = ~\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n36393 = \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n36394 = ~n36392 & n36393 ;
  assign n36395 = ~n36391 & ~n36394 ;
  assign n36396 = n36389 & ~n36395 ;
  assign n36397 = ~n36388 & ~n36396 ;
  assign n36398 = n36378 & n36397 ;
  assign n36399 = \txethmac1_txstatem1_StateJam_q_reg/NET0131  & \txethmac1_txstatem1_StateJam_reg/NET0131  ;
  assign n36400 = \txethmac1_random1_RandomLatched_reg[9]/NET0131  & ~n36399 ;
  assign n36401 = ~\txethmac1_RetryCnt_reg[1]/NET0131  & ~\txethmac1_RetryCnt_reg[2]/NET0131  ;
  assign n36402 = \txethmac1_RetryCnt_reg[3]/NET0131  & \txethmac1_random1_x_reg[9]/NET0131  ;
  assign n36403 = n36399 & n36402 ;
  assign n36404 = ~n36401 & n36403 ;
  assign n36405 = ~n36400 & ~n36404 ;
  assign n36406 = ~\wishbone_TxEn_q_reg/NET0131  & \wishbone_WbEn_q_reg/NET0131  ;
  assign n36407 = ~\wishbone_RxEn_needed_reg/NET0131  & ~\wishbone_RxEn_q_reg/NET0131  ;
  assign n36408 = n36406 & n36407 ;
  assign n36409 = \wishbone_RxEn_q_reg/NET0131  & ~\wishbone_TxEn_q_reg/NET0131  ;
  assign n36410 = ~\wishbone_WbEn_q_reg/NET0131  & n36409 ;
  assign n36411 = ~n36408 & ~n36410 ;
  assign n36412 = \wishbone_TxEn_needed_reg/NET0131  & ~n36411 ;
  assign n36413 = \wishbone_RxEn_needed_reg/NET0131  & ~\wishbone_RxEn_q_reg/NET0131  ;
  assign n36414 = ~\wishbone_TxEn_needed_reg/NET0131  & ~n36413 ;
  assign n36415 = ~\wishbone_TxEn_q_reg/NET0131  & ~n36414 ;
  assign n36416 = \wishbone_RxEn_q_reg/NET0131  & \wishbone_TxEn_q_reg/NET0131  ;
  assign n36417 = ~\wishbone_WbEn_q_reg/NET0131  & ~n36416 ;
  assign n36418 = ~n36415 & n36417 ;
  assign n36419 = ~n36412 & ~n36418 ;
  assign n36420 = n36406 & n36413 ;
  assign n36421 = \wishbone_ram_addr_reg[0]/NET0131  & ~n36420 ;
  assign n36422 = n36419 & n36421 ;
  assign n36423 = \wb_adr_i[2]_pad  & n36417 ;
  assign n36424 = ~n36415 & n36423 ;
  assign n36425 = \wishbone_TxEn_needed_reg/NET0131  & \wishbone_TxPointerRead_reg/NET0131  ;
  assign n36426 = ~n36411 & n36425 ;
  assign n36427 = \wishbone_RxPointerRead_reg/NET0131  & n36420 ;
  assign n36428 = ~n36426 & ~n36427 ;
  assign n36429 = ~n36424 & n36428 ;
  assign n36430 = ~n36422 & n36429 ;
  assign n36431 = \wishbone_ram_addr_reg[1]/NET0131  & ~n36420 ;
  assign n36432 = n36419 & n36431 ;
  assign n36433 = \wb_adr_i[3]_pad  & n36417 ;
  assign n36434 = ~n36415 & n36433 ;
  assign n36435 = \wishbone_TxBDAddress_reg[1]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36436 = ~n36411 & n36435 ;
  assign n36437 = \wishbone_RxBDAddress_reg[1]/NET0131  & n36420 ;
  assign n36438 = ~n36436 & ~n36437 ;
  assign n36439 = ~n36434 & n36438 ;
  assign n36440 = ~n36432 & n36439 ;
  assign n36441 = \wishbone_ram_addr_reg[2]/NET0131  & ~n36420 ;
  assign n36442 = n36419 & n36441 ;
  assign n36443 = \wb_adr_i[4]_pad  & n36417 ;
  assign n36444 = ~n36415 & n36443 ;
  assign n36445 = \wishbone_TxBDAddress_reg[2]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36446 = ~n36411 & n36445 ;
  assign n36447 = \wishbone_RxBDAddress_reg[2]/NET0131  & n36420 ;
  assign n36448 = ~n36446 & ~n36447 ;
  assign n36449 = ~n36444 & n36448 ;
  assign n36450 = ~n36442 & n36449 ;
  assign n36451 = \wishbone_ram_addr_reg[3]/NET0131  & ~n36420 ;
  assign n36452 = n36419 & n36451 ;
  assign n36453 = \wb_adr_i[5]_pad  & n36417 ;
  assign n36454 = ~n36415 & n36453 ;
  assign n36455 = \wishbone_TxBDAddress_reg[3]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36456 = ~n36411 & n36455 ;
  assign n36457 = \wishbone_RxBDAddress_reg[3]/NET0131  & n36420 ;
  assign n36458 = ~n36456 & ~n36457 ;
  assign n36459 = ~n36454 & n36458 ;
  assign n36460 = ~n36452 & n36459 ;
  assign n36461 = \wishbone_ram_addr_reg[4]/NET0131  & ~n36420 ;
  assign n36462 = n36419 & n36461 ;
  assign n36463 = \wb_adr_i[6]_pad  & n36417 ;
  assign n36464 = ~n36415 & n36463 ;
  assign n36465 = \wishbone_TxBDAddress_reg[4]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36466 = ~n36411 & n36465 ;
  assign n36467 = \wishbone_RxBDAddress_reg[4]/NET0131  & n36420 ;
  assign n36468 = ~n36466 & ~n36467 ;
  assign n36469 = ~n36464 & n36468 ;
  assign n36470 = ~n36462 & n36469 ;
  assign n36471 = \wishbone_ram_addr_reg[5]/NET0131  & ~n36420 ;
  assign n36472 = n36419 & n36471 ;
  assign n36473 = \wb_adr_i[7]_pad  & n36417 ;
  assign n36474 = ~n36415 & n36473 ;
  assign n36475 = \wishbone_TxBDAddress_reg[5]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36476 = ~n36411 & n36475 ;
  assign n36477 = \wishbone_RxBDAddress_reg[5]/NET0131  & n36420 ;
  assign n36478 = ~n36476 & ~n36477 ;
  assign n36479 = ~n36474 & n36478 ;
  assign n36480 = ~n36472 & n36479 ;
  assign n36481 = \wishbone_ram_addr_reg[6]/NET0131  & ~n36420 ;
  assign n36482 = n36419 & n36481 ;
  assign n36483 = \wb_adr_i[8]_pad  & n36417 ;
  assign n36484 = ~n36415 & n36483 ;
  assign n36485 = \wishbone_TxBDAddress_reg[6]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36486 = ~n36411 & n36485 ;
  assign n36487 = \wishbone_RxBDAddress_reg[6]/NET0131  & n36420 ;
  assign n36488 = ~n36486 & ~n36487 ;
  assign n36489 = ~n36484 & n36488 ;
  assign n36490 = ~n36482 & n36489 ;
  assign n36491 = \wishbone_ram_addr_reg[7]/NET0131  & ~n36420 ;
  assign n36492 = n36419 & n36491 ;
  assign n36493 = \wb_adr_i[9]_pad  & n36417 ;
  assign n36494 = ~n36415 & n36493 ;
  assign n36495 = \wishbone_TxBDAddress_reg[7]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36496 = ~n36411 & n36495 ;
  assign n36497 = \wishbone_RxBDAddress_reg[7]/NET0131  & n36420 ;
  assign n36498 = ~n36496 & ~n36497 ;
  assign n36499 = ~n36494 & n36498 ;
  assign n36500 = ~n36492 & n36499 ;
  assign n36501 = \wishbone_ram_di_reg[0]/NET0131  & ~n36420 ;
  assign n36502 = n36419 & n36501 ;
  assign n36503 = \wb_dat_i[0]_pad  & n36417 ;
  assign n36504 = ~n36415 & n36503 ;
  assign n36505 = \macstatus1_CarrierSenseLost_reg/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36506 = ~n36411 & n36505 ;
  assign n36507 = \wishbone_RxStatusInLatched_reg[0]/NET0131  & n36420 ;
  assign n36508 = ~n36506 & ~n36507 ;
  assign n36509 = ~n36504 & n36508 ;
  assign n36510 = ~n36502 & n36509 ;
  assign n36511 = \wishbone_ram_di_reg[13]/NET0131  & ~n36420 ;
  assign n36512 = n36419 & n36511 ;
  assign n36513 = \wb_dat_i[13]_pad  & n36417 ;
  assign n36514 = ~n36415 & n36513 ;
  assign n36515 = \wishbone_TxEn_needed_reg/NET0131  & \wishbone_TxStatus_reg[13]/NET0131  ;
  assign n36516 = ~n36411 & n36515 ;
  assign n36517 = \wishbone_RxStatus_reg[13]/NET0131  & n36420 ;
  assign n36518 = ~n36516 & ~n36517 ;
  assign n36519 = ~n36514 & n36518 ;
  assign n36520 = ~n36512 & n36519 ;
  assign n36521 = \wishbone_ram_di_reg[14]/NET0131  & ~n36420 ;
  assign n36522 = n36419 & n36521 ;
  assign n36523 = \wb_dat_i[14]_pad  & n36417 ;
  assign n36524 = ~n36415 & n36523 ;
  assign n36525 = \wishbone_TxEn_needed_reg/NET0131  & \wishbone_TxStatus_reg[14]/NET0131  ;
  assign n36526 = ~n36411 & n36525 ;
  assign n36527 = \wishbone_RxStatus_reg[14]/NET0131  & n36420 ;
  assign n36528 = ~n36526 & ~n36527 ;
  assign n36529 = ~n36524 & n36528 ;
  assign n36530 = ~n36522 & n36529 ;
  assign n36531 = \wishbone_ram_di_reg[16]/NET0131  & ~n36420 ;
  assign n36532 = n36419 & n36531 ;
  assign n36533 = \wishbone_LatchedTxLength_reg[0]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36534 = ~n36411 & n36533 ;
  assign n36535 = \wb_dat_i[16]_pad  & n36417 ;
  assign n36536 = ~n36415 & n36535 ;
  assign n36537 = \wishbone_LatchedRxLength_reg[0]/NET0131  & n36420 ;
  assign n36538 = ~n36536 & ~n36537 ;
  assign n36539 = ~n36534 & n36538 ;
  assign n36540 = ~n36532 & n36539 ;
  assign n36541 = \wishbone_ram_di_reg[17]/NET0131  & ~n36420 ;
  assign n36542 = n36419 & n36541 ;
  assign n36543 = \wishbone_LatchedTxLength_reg[1]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36544 = ~n36411 & n36543 ;
  assign n36545 = \wb_dat_i[17]_pad  & n36417 ;
  assign n36546 = ~n36415 & n36545 ;
  assign n36547 = \wishbone_LatchedRxLength_reg[1]/NET0131  & n36420 ;
  assign n36548 = ~n36546 & ~n36547 ;
  assign n36549 = ~n36544 & n36548 ;
  assign n36550 = ~n36542 & n36549 ;
  assign n36551 = \wishbone_ram_di_reg[18]/NET0131  & ~n36420 ;
  assign n36552 = n36419 & n36551 ;
  assign n36553 = \wishbone_LatchedTxLength_reg[2]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36554 = ~n36411 & n36553 ;
  assign n36555 = \wb_dat_i[18]_pad  & n36417 ;
  assign n36556 = ~n36415 & n36555 ;
  assign n36557 = \wishbone_LatchedRxLength_reg[2]/NET0131  & n36420 ;
  assign n36558 = ~n36556 & ~n36557 ;
  assign n36559 = ~n36554 & n36558 ;
  assign n36560 = ~n36552 & n36559 ;
  assign n36561 = \wishbone_ram_di_reg[19]/NET0131  & ~n36420 ;
  assign n36562 = n36419 & n36561 ;
  assign n36563 = \wishbone_LatchedTxLength_reg[3]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36564 = ~n36411 & n36563 ;
  assign n36565 = \wb_dat_i[19]_pad  & n36417 ;
  assign n36566 = ~n36415 & n36565 ;
  assign n36567 = \wishbone_LatchedRxLength_reg[3]/NET0131  & n36420 ;
  assign n36568 = ~n36566 & ~n36567 ;
  assign n36569 = ~n36564 & n36568 ;
  assign n36570 = ~n36562 & n36569 ;
  assign n36571 = \wishbone_ram_di_reg[1]/NET0131  & ~n36420 ;
  assign n36572 = n36419 & n36571 ;
  assign n36573 = \wb_dat_i[1]_pad  & n36417 ;
  assign n36574 = ~n36415 & n36573 ;
  assign n36575 = \macstatus1_DeferLatched_reg/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36576 = ~n36411 & n36575 ;
  assign n36577 = \wishbone_RxStatusInLatched_reg[1]/NET0131  & n36420 ;
  assign n36578 = ~n36576 & ~n36577 ;
  assign n36579 = ~n36574 & n36578 ;
  assign n36580 = ~n36572 & n36579 ;
  assign n36581 = \wishbone_ram_di_reg[20]/NET0131  & ~n36420 ;
  assign n36582 = n36419 & n36581 ;
  assign n36583 = \wishbone_LatchedTxLength_reg[4]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36584 = ~n36411 & n36583 ;
  assign n36585 = \wb_dat_i[20]_pad  & n36417 ;
  assign n36586 = ~n36415 & n36585 ;
  assign n36587 = \wishbone_LatchedRxLength_reg[4]/NET0131  & n36420 ;
  assign n36588 = ~n36586 & ~n36587 ;
  assign n36589 = ~n36584 & n36588 ;
  assign n36590 = ~n36582 & n36589 ;
  assign n36591 = \wishbone_ram_di_reg[21]/NET0131  & ~n36420 ;
  assign n36592 = n36419 & n36591 ;
  assign n36593 = \wishbone_LatchedTxLength_reg[5]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36594 = ~n36411 & n36593 ;
  assign n36595 = \wb_dat_i[21]_pad  & n36417 ;
  assign n36596 = ~n36415 & n36595 ;
  assign n36597 = \wishbone_LatchedRxLength_reg[5]/NET0131  & n36420 ;
  assign n36598 = ~n36596 & ~n36597 ;
  assign n36599 = ~n36594 & n36598 ;
  assign n36600 = ~n36592 & n36599 ;
  assign n36601 = \wishbone_ram_di_reg[22]/NET0131  & ~n36420 ;
  assign n36602 = n36419 & n36601 ;
  assign n36603 = \wishbone_LatchedTxLength_reg[6]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36604 = ~n36411 & n36603 ;
  assign n36605 = \wb_dat_i[22]_pad  & n36417 ;
  assign n36606 = ~n36415 & n36605 ;
  assign n36607 = \wishbone_LatchedRxLength_reg[6]/NET0131  & n36420 ;
  assign n36608 = ~n36606 & ~n36607 ;
  assign n36609 = ~n36604 & n36608 ;
  assign n36610 = ~n36602 & n36609 ;
  assign n36611 = \wishbone_ram_di_reg[23]/NET0131  & ~n36420 ;
  assign n36612 = n36419 & n36611 ;
  assign n36613 = \wb_dat_i[23]_pad  & n36417 ;
  assign n36614 = ~n36415 & n36613 ;
  assign n36615 = \wishbone_LatchedTxLength_reg[7]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36616 = ~n36411 & n36615 ;
  assign n36617 = \wishbone_LatchedRxLength_reg[7]/NET0131  & n36420 ;
  assign n36618 = ~n36616 & ~n36617 ;
  assign n36619 = ~n36614 & n36618 ;
  assign n36620 = ~n36612 & n36619 ;
  assign n36621 = \wishbone_ram_di_reg[24]/NET0131  & ~n36420 ;
  assign n36622 = n36419 & n36621 ;
  assign n36623 = \wb_dat_i[24]_pad  & n36417 ;
  assign n36624 = ~n36415 & n36623 ;
  assign n36625 = \wishbone_LatchedTxLength_reg[8]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36626 = ~n36411 & n36625 ;
  assign n36627 = \wishbone_LatchedRxLength_reg[8]/NET0131  & n36420 ;
  assign n36628 = ~n36626 & ~n36627 ;
  assign n36629 = ~n36624 & n36628 ;
  assign n36630 = ~n36622 & n36629 ;
  assign n36631 = \wishbone_ram_di_reg[25]/NET0131  & ~n36420 ;
  assign n36632 = n36419 & n36631 ;
  assign n36633 = \wishbone_LatchedTxLength_reg[9]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36634 = ~n36411 & n36633 ;
  assign n36635 = \wb_dat_i[25]_pad  & n36417 ;
  assign n36636 = ~n36415 & n36635 ;
  assign n36637 = \wishbone_LatchedRxLength_reg[9]/NET0131  & n36420 ;
  assign n36638 = ~n36636 & ~n36637 ;
  assign n36639 = ~n36634 & n36638 ;
  assign n36640 = ~n36632 & n36639 ;
  assign n36641 = \wishbone_ram_di_reg[26]/NET0131  & ~n36420 ;
  assign n36642 = n36419 & n36641 ;
  assign n36643 = \wishbone_LatchedTxLength_reg[10]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36644 = ~n36411 & n36643 ;
  assign n36645 = \wb_dat_i[26]_pad  & n36417 ;
  assign n36646 = ~n36415 & n36645 ;
  assign n36647 = \wishbone_LatchedRxLength_reg[10]/NET0131  & n36420 ;
  assign n36648 = ~n36646 & ~n36647 ;
  assign n36649 = ~n36644 & n36648 ;
  assign n36650 = ~n36642 & n36649 ;
  assign n36651 = \wishbone_ram_di_reg[27]/NET0131  & ~n36420 ;
  assign n36652 = n36419 & n36651 ;
  assign n36653 = \wb_dat_i[27]_pad  & n36417 ;
  assign n36654 = ~n36415 & n36653 ;
  assign n36655 = \wishbone_LatchedTxLength_reg[11]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36656 = ~n36411 & n36655 ;
  assign n36657 = \wishbone_LatchedRxLength_reg[11]/NET0131  & n36420 ;
  assign n36658 = ~n36656 & ~n36657 ;
  assign n36659 = ~n36654 & n36658 ;
  assign n36660 = ~n36652 & n36659 ;
  assign n36661 = \wishbone_ram_di_reg[28]/NET0131  & ~n36420 ;
  assign n36662 = n36419 & n36661 ;
  assign n36663 = \wishbone_LatchedTxLength_reg[12]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36664 = ~n36411 & n36663 ;
  assign n36665 = \wb_dat_i[28]_pad  & n36417 ;
  assign n36666 = ~n36415 & n36665 ;
  assign n36667 = \wishbone_LatchedRxLength_reg[12]/NET0131  & n36420 ;
  assign n36668 = ~n36666 & ~n36667 ;
  assign n36669 = ~n36664 & n36668 ;
  assign n36670 = ~n36662 & n36669 ;
  assign n36671 = \wishbone_ram_di_reg[29]/NET0131  & ~n36420 ;
  assign n36672 = n36419 & n36671 ;
  assign n36673 = \wb_dat_i[29]_pad  & n36417 ;
  assign n36674 = ~n36415 & n36673 ;
  assign n36675 = \wishbone_LatchedTxLength_reg[13]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36676 = ~n36411 & n36675 ;
  assign n36677 = \wishbone_LatchedRxLength_reg[13]/NET0131  & n36420 ;
  assign n36678 = ~n36676 & ~n36677 ;
  assign n36679 = ~n36674 & n36678 ;
  assign n36680 = ~n36672 & n36679 ;
  assign n36681 = \wishbone_ram_di_reg[2]/NET0131  & ~n36420 ;
  assign n36682 = n36419 & n36681 ;
  assign n36683 = \macstatus1_LateCollLatched_reg/P0002  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36684 = ~n36411 & n36683 ;
  assign n36685 = \wb_dat_i[2]_pad  & n36417 ;
  assign n36686 = ~n36415 & n36685 ;
  assign n36687 = \wishbone_RxStatusInLatched_reg[2]/NET0131  & n36420 ;
  assign n36688 = ~n36686 & ~n36687 ;
  assign n36689 = ~n36684 & n36688 ;
  assign n36690 = ~n36682 & n36689 ;
  assign n36691 = \wishbone_ram_di_reg[30]/NET0131  & ~n36420 ;
  assign n36692 = n36419 & n36691 ;
  assign n36693 = \wishbone_LatchedTxLength_reg[14]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36694 = ~n36411 & n36693 ;
  assign n36695 = \wb_dat_i[30]_pad  & n36417 ;
  assign n36696 = ~n36415 & n36695 ;
  assign n36697 = \wishbone_LatchedRxLength_reg[14]/NET0131  & n36420 ;
  assign n36698 = ~n36696 & ~n36697 ;
  assign n36699 = ~n36694 & n36698 ;
  assign n36700 = ~n36692 & n36699 ;
  assign n36701 = \wishbone_ram_di_reg[31]/NET0131  & ~n36420 ;
  assign n36702 = n36419 & n36701 ;
  assign n36703 = \wishbone_LatchedTxLength_reg[15]/NET0131  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36704 = ~n36411 & n36703 ;
  assign n36705 = \wb_dat_i[31]_pad  & n36417 ;
  assign n36706 = ~n36415 & n36705 ;
  assign n36707 = \wishbone_LatchedRxLength_reg[15]/NET0131  & n36420 ;
  assign n36708 = ~n36706 & ~n36707 ;
  assign n36709 = ~n36704 & n36708 ;
  assign n36710 = ~n36702 & n36709 ;
  assign n36711 = \wishbone_ram_di_reg[3]/NET0131  & ~n36420 ;
  assign n36712 = n36419 & n36711 ;
  assign n36713 = \wb_dat_i[3]_pad  & n36417 ;
  assign n36714 = ~n36415 & n36713 ;
  assign n36715 = \macstatus1_RetryLimit_reg/P0002  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36716 = ~n36411 & n36715 ;
  assign n36717 = \wishbone_RxStatusInLatched_reg[3]/NET0131  & n36420 ;
  assign n36718 = ~n36716 & ~n36717 ;
  assign n36719 = ~n36714 & n36718 ;
  assign n36720 = ~n36712 & n36719 ;
  assign n36721 = \wishbone_ram_di_reg[4]/NET0131  & ~n36420 ;
  assign n36722 = n36419 & n36721 ;
  assign n36723 = \macstatus1_RetryCntLatched_reg[0]/P0002  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36724 = ~n36411 & n36723 ;
  assign n36725 = \wb_dat_i[4]_pad  & n36417 ;
  assign n36726 = ~n36415 & n36725 ;
  assign n36727 = \wishbone_RxStatusInLatched_reg[4]/NET0131  & n36420 ;
  assign n36728 = ~n36726 & ~n36727 ;
  assign n36729 = ~n36724 & n36728 ;
  assign n36730 = ~n36722 & n36729 ;
  assign n36731 = \wishbone_ram_di_reg[5]/NET0131  & ~n36420 ;
  assign n36732 = n36419 & n36731 ;
  assign n36733 = \macstatus1_RetryCntLatched_reg[1]/P0002  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36734 = ~n36411 & n36733 ;
  assign n36735 = \wb_dat_i[5]_pad  & n36417 ;
  assign n36736 = ~n36415 & n36735 ;
  assign n36737 = \wishbone_RxStatusInLatched_reg[5]/NET0131  & n36420 ;
  assign n36738 = ~n36736 & ~n36737 ;
  assign n36739 = ~n36734 & n36738 ;
  assign n36740 = ~n36732 & n36739 ;
  assign n36741 = \wishbone_ram_di_reg[6]/NET0131  & ~n36420 ;
  assign n36742 = n36419 & n36741 ;
  assign n36743 = \macstatus1_RetryCntLatched_reg[2]/P0002  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36744 = ~n36411 & n36743 ;
  assign n36745 = \wb_dat_i[6]_pad  & n36417 ;
  assign n36746 = ~n36415 & n36745 ;
  assign n36747 = \wishbone_RxStatusInLatched_reg[6]/NET0131  & n36420 ;
  assign n36748 = ~n36746 & ~n36747 ;
  assign n36749 = ~n36744 & n36748 ;
  assign n36750 = ~n36742 & n36749 ;
  assign n36751 = \wishbone_ram_di_reg[7]/NET0131  & ~n36420 ;
  assign n36752 = n36419 & n36751 ;
  assign n36753 = \macstatus1_RetryCntLatched_reg[3]/P0002  & \wishbone_TxEn_needed_reg/NET0131  ;
  assign n36754 = ~n36411 & n36753 ;
  assign n36755 = \wb_dat_i[7]_pad  & n36417 ;
  assign n36756 = ~n36415 & n36755 ;
  assign n36757 = \wishbone_RxStatusInLatched_reg[7]/NET0131  & n36420 ;
  assign n36758 = ~n36756 & ~n36757 ;
  assign n36759 = ~n36754 & n36758 ;
  assign n36760 = ~n36752 & n36759 ;
  assign n36761 = \wishbone_ram_di_reg[8]/NET0131  & ~n36420 ;
  assign n36762 = n36419 & n36761 ;
  assign n36763 = \wishbone_TxEn_needed_reg/NET0131  & \wishbone_TxUnderRun_reg/NET0131  ;
  assign n36764 = ~n36411 & n36763 ;
  assign n36765 = \wb_dat_i[8]_pad  & n36417 ;
  assign n36766 = ~n36415 & n36765 ;
  assign n36767 = \wishbone_RxStatusInLatched_reg[8]/NET0131  & n36420 ;
  assign n36768 = ~n36766 & ~n36767 ;
  assign n36769 = ~n36764 & n36768 ;
  assign n36770 = ~n36762 & n36769 ;
  assign n36771 = n35359 & ~n35365 ;
  assign n36772 = \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  & ~n33164 ;
  assign n36773 = ~n36771 & n36772 ;
  assign n36774 = n35359 & ~n36772 ;
  assign n36775 = ~n35365 & n36774 ;
  assign n36776 = ~n36773 & ~n36775 ;
  assign n36777 = ~\wishbone_tx_fifo_write_pointer_reg[0]/NET0131  & ~n14049 ;
  assign n36778 = \wishbone_tx_fifo_cnt_reg[4]/NET0131  & ~\wishbone_tx_fifo_write_pointer_reg[0]/NET0131  ;
  assign n36779 = n35314 & n36778 ;
  assign n36780 = ~n36777 & ~n36779 ;
  assign n36781 = ~n35731 & n35743 ;
  assign n36782 = n34242 & ~n36781 ;
  assign n36783 = n36780 & n36782 ;
  assign n36784 = ~n35955 & ~n36783 ;
  assign n36785 = ~\wishbone_rx_fifo_write_pointer_reg[0]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n36786 = ~n33164 & n35359 ;
  assign n36787 = \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[2]/NET0131  ;
  assign n36788 = n36786 & n36787 ;
  assign n36789 = ~n35365 & n36788 ;
  assign n36790 = n36785 & n36789 ;
  assign n36791 = \wishbone_rx_fifo_fifo_reg[10][10]/P0001  & ~n36790 ;
  assign n36792 = \wishbone_RxDataLatched2_reg[10]/NET0131  & n36785 ;
  assign n36793 = n36789 & n36792 ;
  assign n36794 = ~n36791 & ~n36793 ;
  assign n36795 = \wishbone_rx_fifo_fifo_reg[10][12]/P0001  & ~n36790 ;
  assign n36796 = \wishbone_RxDataLatched2_reg[12]/NET0131  & n36785 ;
  assign n36797 = n36789 & n36796 ;
  assign n36798 = ~n36795 & ~n36797 ;
  assign n36799 = \wishbone_rx_fifo_fifo_reg[10][14]/P0001  & ~n36790 ;
  assign n36800 = \wishbone_RxDataLatched2_reg[14]/NET0131  & n36785 ;
  assign n36801 = n36789 & n36800 ;
  assign n36802 = ~n36799 & ~n36801 ;
  assign n36803 = \wishbone_rx_fifo_fifo_reg[10][16]/P0001  & ~n36790 ;
  assign n36804 = \wishbone_RxDataLatched2_reg[16]/NET0131  & n36785 ;
  assign n36805 = n36789 & n36804 ;
  assign n36806 = ~n36803 & ~n36805 ;
  assign n36807 = \wishbone_rx_fifo_fifo_reg[10][1]/P0001  & ~n36790 ;
  assign n36808 = \wishbone_RxDataLatched2_reg[1]/NET0131  & n36785 ;
  assign n36809 = n36789 & n36808 ;
  assign n36810 = ~n36807 & ~n36809 ;
  assign n36811 = \wishbone_rx_fifo_fifo_reg[10][20]/P0001  & ~n36790 ;
  assign n36812 = \wishbone_RxDataLatched2_reg[20]/NET0131  & n36785 ;
  assign n36813 = n36789 & n36812 ;
  assign n36814 = ~n36811 & ~n36813 ;
  assign n36815 = \wishbone_rx_fifo_fifo_reg[10][27]/P0001  & ~n36790 ;
  assign n36816 = \wishbone_RxDataLatched2_reg[27]/NET0131  & n36785 ;
  assign n36817 = n36789 & n36816 ;
  assign n36818 = ~n36815 & ~n36817 ;
  assign n36819 = \wishbone_rx_fifo_fifo_reg[10][28]/P0001  & ~n36790 ;
  assign n36820 = \wishbone_RxDataLatched2_reg[28]/NET0131  & n36785 ;
  assign n36821 = n36789 & n36820 ;
  assign n36822 = ~n36819 & ~n36821 ;
  assign n36823 = \wishbone_rx_fifo_fifo_reg[10][29]/P0001  & ~n36790 ;
  assign n36824 = \wishbone_RxDataLatched2_reg[29]/NET0131  & n36785 ;
  assign n36825 = n36789 & n36824 ;
  assign n36826 = ~n36823 & ~n36825 ;
  assign n36827 = \wishbone_rx_fifo_fifo_reg[10][31]/P0001  & ~n36790 ;
  assign n36828 = \wishbone_RxDataLatched2_reg[31]/NET0131  & n36785 ;
  assign n36829 = n36789 & n36828 ;
  assign n36830 = ~n36827 & ~n36829 ;
  assign n36831 = \wishbone_rx_fifo_fifo_reg[10][4]/P0001  & ~n36790 ;
  assign n36832 = \wishbone_RxDataLatched2_reg[4]/NET0131  & n36785 ;
  assign n36833 = n36789 & n36832 ;
  assign n36834 = ~n36831 & ~n36833 ;
  assign n36835 = \wishbone_rx_fifo_fifo_reg[10][5]/P0001  & ~n36790 ;
  assign n36836 = \wishbone_RxDataLatched2_reg[5]/NET0131  & n36785 ;
  assign n36837 = n36789 & n36836 ;
  assign n36838 = ~n36835 & ~n36837 ;
  assign n36839 = \wishbone_rx_fifo_fifo_reg[10][7]/P0001  & ~n36790 ;
  assign n36840 = \wishbone_RxDataLatched2_reg[7]/NET0131  & n36785 ;
  assign n36841 = n36789 & n36840 ;
  assign n36842 = ~n36839 & ~n36841 ;
  assign n36843 = \wishbone_rx_fifo_fifo_reg[10][9]/P0001  & ~n36790 ;
  assign n36844 = \wishbone_RxDataLatched2_reg[9]/NET0131  & n36785 ;
  assign n36845 = n36789 & n36844 ;
  assign n36846 = ~n36843 & ~n36845 ;
  assign n36847 = \wishbone_rx_fifo_write_pointer_reg[2]/NET0131  & n35359 ;
  assign n36848 = ~n33164 & n36847 ;
  assign n36849 = ~n35365 & n36848 ;
  assign n36850 = ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n36785 ;
  assign n36851 = n36849 & n36850 ;
  assign n36852 = \wishbone_rx_fifo_fifo_reg[12][11]/P0001  & ~n36851 ;
  assign n36853 = \wishbone_RxDataLatched2_reg[11]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36854 = n36785 & n36853 ;
  assign n36855 = n36849 & n36854 ;
  assign n36856 = ~n36852 & ~n36855 ;
  assign n36857 = \wishbone_rx_fifo_fifo_reg[12][12]/P0001  & ~n36851 ;
  assign n36858 = \wishbone_RxDataLatched2_reg[12]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36859 = n36785 & n36858 ;
  assign n36860 = n36849 & n36859 ;
  assign n36861 = ~n36857 & ~n36860 ;
  assign n36862 = \wishbone_rx_fifo_fifo_reg[12][14]/P0001  & ~n36851 ;
  assign n36863 = \wishbone_RxDataLatched2_reg[14]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36864 = n36785 & n36863 ;
  assign n36865 = n36849 & n36864 ;
  assign n36866 = ~n36862 & ~n36865 ;
  assign n36867 = \wishbone_rx_fifo_fifo_reg[12][15]/P0001  & ~n36851 ;
  assign n36868 = \wishbone_RxDataLatched2_reg[15]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36869 = n36785 & n36868 ;
  assign n36870 = n36849 & n36869 ;
  assign n36871 = ~n36867 & ~n36870 ;
  assign n36872 = \wishbone_rx_fifo_fifo_reg[12][16]/P0001  & ~n36851 ;
  assign n36873 = \wishbone_RxDataLatched2_reg[16]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36874 = n36785 & n36873 ;
  assign n36875 = n36849 & n36874 ;
  assign n36876 = ~n36872 & ~n36875 ;
  assign n36877 = \wishbone_rx_fifo_fifo_reg[12][17]/P0001  & ~n36851 ;
  assign n36878 = \wishbone_RxDataLatched2_reg[17]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36879 = n36785 & n36878 ;
  assign n36880 = n36849 & n36879 ;
  assign n36881 = ~n36877 & ~n36880 ;
  assign n36882 = \wishbone_rx_fifo_fifo_reg[12][19]/P0001  & ~n36851 ;
  assign n36883 = \wishbone_RxDataLatched2_reg[19]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36884 = n36785 & n36883 ;
  assign n36885 = n36849 & n36884 ;
  assign n36886 = ~n36882 & ~n36885 ;
  assign n36887 = \wishbone_rx_fifo_fifo_reg[12][21]/P0001  & ~n36851 ;
  assign n36888 = \wishbone_RxDataLatched2_reg[21]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36889 = n36785 & n36888 ;
  assign n36890 = n36849 & n36889 ;
  assign n36891 = ~n36887 & ~n36890 ;
  assign n36892 = \wishbone_rx_fifo_fifo_reg[12][22]/P0001  & ~n36851 ;
  assign n36893 = \wishbone_RxDataLatched2_reg[22]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36894 = n36785 & n36893 ;
  assign n36895 = n36849 & n36894 ;
  assign n36896 = ~n36892 & ~n36895 ;
  assign n36897 = \wishbone_rx_fifo_fifo_reg[12][23]/P0001  & ~n36851 ;
  assign n36898 = \wishbone_RxDataLatched2_reg[23]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36899 = n36785 & n36898 ;
  assign n36900 = n36849 & n36899 ;
  assign n36901 = ~n36897 & ~n36900 ;
  assign n36902 = \wishbone_rx_fifo_fifo_reg[12][24]/P0001  & ~n36851 ;
  assign n36903 = \wishbone_RxDataLatched2_reg[24]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36904 = n36785 & n36903 ;
  assign n36905 = n36849 & n36904 ;
  assign n36906 = ~n36902 & ~n36905 ;
  assign n36907 = \wishbone_rx_fifo_fifo_reg[12][27]/P0001  & ~n36851 ;
  assign n36908 = \wishbone_RxDataLatched2_reg[27]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36909 = n36785 & n36908 ;
  assign n36910 = n36849 & n36909 ;
  assign n36911 = ~n36907 & ~n36910 ;
  assign n36912 = \wishbone_rx_fifo_fifo_reg[12][28]/P0001  & ~n36851 ;
  assign n36913 = \wishbone_RxDataLatched2_reg[28]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36914 = n36785 & n36913 ;
  assign n36915 = n36849 & n36914 ;
  assign n36916 = ~n36912 & ~n36915 ;
  assign n36917 = \wishbone_rx_fifo_fifo_reg[12][31]/P0001  & ~n36851 ;
  assign n36918 = \wishbone_RxDataLatched2_reg[31]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36919 = n36785 & n36918 ;
  assign n36920 = n36849 & n36919 ;
  assign n36921 = ~n36917 & ~n36920 ;
  assign n36922 = \wishbone_rx_fifo_fifo_reg[12][4]/P0001  & ~n36851 ;
  assign n36923 = \wishbone_RxDataLatched2_reg[4]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36924 = n36785 & n36923 ;
  assign n36925 = n36849 & n36924 ;
  assign n36926 = ~n36922 & ~n36925 ;
  assign n36927 = \wishbone_rx_fifo_fifo_reg[12][7]/P0001  & ~n36851 ;
  assign n36928 = \wishbone_RxDataLatched2_reg[7]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n36929 = n36785 & n36928 ;
  assign n36930 = n36849 & n36929 ;
  assign n36931 = ~n36927 & ~n36930 ;
  assign n36932 = \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n36933 = n36789 & n36932 ;
  assign n36934 = \wishbone_rx_fifo_fifo_reg[3][10]/P0001  & ~n36933 ;
  assign n36935 = \wishbone_RxDataLatched2_reg[10]/NET0131  & n36932 ;
  assign n36936 = n36789 & n36935 ;
  assign n36937 = ~n36934 & ~n36936 ;
  assign n36938 = \wishbone_rx_fifo_fifo_reg[3][12]/P0001  & ~n36933 ;
  assign n36939 = \wishbone_RxDataLatched2_reg[12]/NET0131  & n36932 ;
  assign n36940 = n36789 & n36939 ;
  assign n36941 = ~n36938 & ~n36940 ;
  assign n36942 = \wishbone_rx_fifo_fifo_reg[3][13]/P0001  & ~n36933 ;
  assign n36943 = \wishbone_RxDataLatched2_reg[13]/NET0131  & n36932 ;
  assign n36944 = n36789 & n36943 ;
  assign n36945 = ~n36942 & ~n36944 ;
  assign n36946 = \wishbone_rx_fifo_fifo_reg[3][14]/P0001  & ~n36933 ;
  assign n36947 = \wishbone_RxDataLatched2_reg[14]/NET0131  & n36932 ;
  assign n36948 = n36789 & n36947 ;
  assign n36949 = ~n36946 & ~n36948 ;
  assign n36950 = \wishbone_rx_fifo_fifo_reg[3][18]/P0001  & ~n36933 ;
  assign n36951 = \wishbone_RxDataLatched2_reg[18]/NET0131  & n36932 ;
  assign n36952 = n36789 & n36951 ;
  assign n36953 = ~n36950 & ~n36952 ;
  assign n36954 = \wishbone_rx_fifo_fifo_reg[3][19]/P0001  & ~n36933 ;
  assign n36955 = \wishbone_RxDataLatched2_reg[19]/NET0131  & n36932 ;
  assign n36956 = n36789 & n36955 ;
  assign n36957 = ~n36954 & ~n36956 ;
  assign n36958 = \wishbone_rx_fifo_fifo_reg[3][24]/P0001  & ~n36933 ;
  assign n36959 = \wishbone_RxDataLatched2_reg[24]/NET0131  & n36932 ;
  assign n36960 = n36789 & n36959 ;
  assign n36961 = ~n36958 & ~n36960 ;
  assign n36962 = \wishbone_rx_fifo_fifo_reg[3][26]/P0001  & ~n36933 ;
  assign n36963 = \wishbone_RxDataLatched2_reg[26]/NET0131  & n36932 ;
  assign n36964 = n36789 & n36963 ;
  assign n36965 = ~n36962 & ~n36964 ;
  assign n36966 = \wishbone_rx_fifo_fifo_reg[3][29]/P0001  & ~n36933 ;
  assign n36967 = \wishbone_RxDataLatched2_reg[29]/NET0131  & n36932 ;
  assign n36968 = n36789 & n36967 ;
  assign n36969 = ~n36966 & ~n36968 ;
  assign n36970 = \wishbone_rx_fifo_fifo_reg[3][28]/P0001  & ~n36933 ;
  assign n36971 = \wishbone_RxDataLatched2_reg[28]/NET0131  & n36932 ;
  assign n36972 = n36789 & n36971 ;
  assign n36973 = ~n36970 & ~n36972 ;
  assign n36974 = \wishbone_rx_fifo_fifo_reg[3][2]/P0001  & ~n36933 ;
  assign n36975 = \wishbone_RxDataLatched2_reg[2]/NET0131  & n36932 ;
  assign n36976 = n36789 & n36975 ;
  assign n36977 = ~n36974 & ~n36976 ;
  assign n36978 = \wishbone_rx_fifo_fifo_reg[3][30]/P0001  & ~n36933 ;
  assign n36979 = \wishbone_RxDataLatched2_reg[30]/NET0131  & n36932 ;
  assign n36980 = n36789 & n36979 ;
  assign n36981 = ~n36978 & ~n36980 ;
  assign n36982 = \wishbone_rx_fifo_fifo_reg[3][31]/P0001  & ~n36933 ;
  assign n36983 = \wishbone_RxDataLatched2_reg[31]/NET0131  & n36932 ;
  assign n36984 = n36789 & n36983 ;
  assign n36985 = ~n36982 & ~n36984 ;
  assign n36986 = \wishbone_rx_fifo_fifo_reg[3][4]/P0001  & ~n36933 ;
  assign n36987 = \wishbone_RxDataLatched2_reg[4]/NET0131  & n36932 ;
  assign n36988 = n36789 & n36987 ;
  assign n36989 = ~n36986 & ~n36988 ;
  assign n36990 = \wishbone_rx_fifo_fifo_reg[3][7]/P0001  & ~n36933 ;
  assign n36991 = \wishbone_RxDataLatched2_reg[7]/NET0131  & n36932 ;
  assign n36992 = n36789 & n36991 ;
  assign n36993 = ~n36990 & ~n36992 ;
  assign n36994 = \wishbone_rx_fifo_fifo_reg[3][8]/P0001  & ~n36933 ;
  assign n36995 = \wishbone_RxDataLatched2_reg[8]/NET0131  & n36932 ;
  assign n36996 = n36789 & n36995 ;
  assign n36997 = ~n36994 & ~n36996 ;
  assign n36998 = \wishbone_rx_fifo_fifo_reg[3][9]/P0001  & ~n36933 ;
  assign n36999 = \wishbone_RxDataLatched2_reg[9]/NET0131  & n36932 ;
  assign n37000 = n36789 & n36999 ;
  assign n37001 = ~n36998 & ~n37000 ;
  assign n37002 = ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n36932 ;
  assign n37003 = n36849 & n37002 ;
  assign n37004 = \wishbone_rx_fifo_fifo_reg[5][10]/P0001  & ~n37003 ;
  assign n37005 = \wishbone_RxDataLatched2_reg[10]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37006 = n36932 & n37005 ;
  assign n37007 = n36849 & n37006 ;
  assign n37008 = ~n37004 & ~n37007 ;
  assign n37009 = \wishbone_rx_fifo_fifo_reg[5][13]/P0001  & ~n37003 ;
  assign n37010 = \wishbone_RxDataLatched2_reg[13]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37011 = n36932 & n37010 ;
  assign n37012 = n36849 & n37011 ;
  assign n37013 = ~n37009 & ~n37012 ;
  assign n37014 = \wishbone_rx_fifo_fifo_reg[5][15]/P0001  & ~n37003 ;
  assign n37015 = n36868 & n36932 ;
  assign n37016 = n36849 & n37015 ;
  assign n37017 = ~n37014 & ~n37016 ;
  assign n37018 = \wishbone_rx_fifo_fifo_reg[5][17]/P0001  & ~n37003 ;
  assign n37019 = n36878 & n36932 ;
  assign n37020 = n36849 & n37019 ;
  assign n37021 = ~n37018 & ~n37020 ;
  assign n37022 = \wishbone_rx_fifo_fifo_reg[5][19]/P0001  & ~n37003 ;
  assign n37023 = n36883 & n36932 ;
  assign n37024 = n36849 & n37023 ;
  assign n37025 = ~n37022 & ~n37024 ;
  assign n37026 = \wishbone_rx_fifo_fifo_reg[5][1]/P0001  & ~n37003 ;
  assign n37027 = \wishbone_RxDataLatched2_reg[1]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37028 = n36932 & n37027 ;
  assign n37029 = n36849 & n37028 ;
  assign n37030 = ~n37026 & ~n37029 ;
  assign n37031 = \wishbone_rx_fifo_fifo_reg[5][21]/P0001  & ~n37003 ;
  assign n37032 = n36888 & n36932 ;
  assign n37033 = n36849 & n37032 ;
  assign n37034 = ~n37031 & ~n37033 ;
  assign n37035 = \wishbone_rx_fifo_fifo_reg[5][22]/P0001  & ~n37003 ;
  assign n37036 = n36893 & n36932 ;
  assign n37037 = n36849 & n37036 ;
  assign n37038 = ~n37035 & ~n37037 ;
  assign n37039 = \wishbone_rx_fifo_fifo_reg[5][20]/P0001  & ~n37003 ;
  assign n37040 = \wishbone_RxDataLatched2_reg[20]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37041 = n36932 & n37040 ;
  assign n37042 = n36849 & n37041 ;
  assign n37043 = ~n37039 & ~n37042 ;
  assign n37044 = \wishbone_rx_fifo_fifo_reg[5][23]/P0001  & ~n37003 ;
  assign n37045 = n36898 & n36932 ;
  assign n37046 = n36849 & n37045 ;
  assign n37047 = ~n37044 & ~n37046 ;
  assign n37048 = \wishbone_rx_fifo_fifo_reg[5][24]/P0001  & ~n37003 ;
  assign n37049 = n36903 & n36932 ;
  assign n37050 = n36849 & n37049 ;
  assign n37051 = ~n37048 & ~n37050 ;
  assign n37052 = \wishbone_rx_fifo_fifo_reg[5][26]/P0001  & ~n37003 ;
  assign n37053 = \wishbone_RxDataLatched2_reg[26]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37054 = n36932 & n37053 ;
  assign n37055 = n36849 & n37054 ;
  assign n37056 = ~n37052 & ~n37055 ;
  assign n37057 = \wishbone_rx_fifo_fifo_reg[5][28]/P0001  & ~n37003 ;
  assign n37058 = n36913 & n36932 ;
  assign n37059 = n36849 & n37058 ;
  assign n37060 = ~n37057 & ~n37059 ;
  assign n37061 = \wishbone_rx_fifo_fifo_reg[5][3]/P0001  & ~n37003 ;
  assign n37062 = \wishbone_RxDataLatched2_reg[3]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37063 = n36932 & n37062 ;
  assign n37064 = n36849 & n37063 ;
  assign n37065 = ~n37061 & ~n37064 ;
  assign n37066 = \wishbone_rx_fifo_fifo_reg[5][6]/P0001  & ~n37003 ;
  assign n37067 = \wishbone_RxDataLatched2_reg[6]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37068 = n36932 & n37067 ;
  assign n37069 = n36849 & n37068 ;
  assign n37070 = ~n37066 & ~n37069 ;
  assign n37071 = \wishbone_rx_fifo_fifo_reg[5][8]/P0001  & ~n37003 ;
  assign n37072 = \wishbone_RxDataLatched2_reg[8]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37073 = n36932 & n37072 ;
  assign n37074 = n36849 & n37073 ;
  assign n37075 = ~n37071 & ~n37074 ;
  assign n37076 = ~\wishbone_rx_fifo_write_pointer_reg[0]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n37077 = \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n37076 ;
  assign n37078 = n36849 & n37077 ;
  assign n37079 = \wishbone_rx_fifo_fifo_reg[6][0]/P0001  & ~n37078 ;
  assign n37080 = \wishbone_RxDataLatched2_reg[0]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37081 = n37076 & n37080 ;
  assign n37082 = n36849 & n37081 ;
  assign n37083 = ~n37079 & ~n37082 ;
  assign n37084 = \wishbone_rx_fifo_fifo_reg[6][10]/P0001  & ~n37078 ;
  assign n37085 = \wishbone_RxDataLatched2_reg[10]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37086 = n37076 & n37085 ;
  assign n37087 = n36849 & n37086 ;
  assign n37088 = ~n37084 & ~n37087 ;
  assign n37089 = \wishbone_rx_fifo_fifo_reg[6][11]/P0001  & ~n37078 ;
  assign n37090 = \wishbone_RxDataLatched2_reg[11]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37091 = n37076 & n37090 ;
  assign n37092 = n36849 & n37091 ;
  assign n37093 = ~n37089 & ~n37092 ;
  assign n37094 = \wishbone_rx_fifo_fifo_reg[6][14]/P0001  & ~n37078 ;
  assign n37095 = \wishbone_RxDataLatched2_reg[14]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37096 = n37076 & n37095 ;
  assign n37097 = n36849 & n37096 ;
  assign n37098 = ~n37094 & ~n37097 ;
  assign n37099 = \wishbone_rx_fifo_fifo_reg[6][15]/P0001  & ~n37078 ;
  assign n37100 = \wishbone_RxDataLatched2_reg[15]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37101 = n37076 & n37100 ;
  assign n37102 = n36849 & n37101 ;
  assign n37103 = ~n37099 & ~n37102 ;
  assign n37104 = \wishbone_rx_fifo_fifo_reg[6][16]/P0001  & ~n37078 ;
  assign n37105 = \wishbone_RxDataLatched2_reg[16]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37106 = n37076 & n37105 ;
  assign n37107 = n36849 & n37106 ;
  assign n37108 = ~n37104 & ~n37107 ;
  assign n37109 = \wishbone_rx_fifo_fifo_reg[6][18]/P0001  & ~n37078 ;
  assign n37110 = \wishbone_RxDataLatched2_reg[18]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37111 = n37076 & n37110 ;
  assign n37112 = n36849 & n37111 ;
  assign n37113 = ~n37109 & ~n37112 ;
  assign n37114 = \wishbone_rx_fifo_fifo_reg[6][19]/P0001  & ~n37078 ;
  assign n37115 = \wishbone_RxDataLatched2_reg[19]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37116 = n37076 & n37115 ;
  assign n37117 = n36849 & n37116 ;
  assign n37118 = ~n37114 & ~n37117 ;
  assign n37119 = \wishbone_rx_fifo_fifo_reg[6][1]/P0001  & ~n37078 ;
  assign n37120 = \wishbone_RxDataLatched2_reg[1]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37121 = n37076 & n37120 ;
  assign n37122 = n36849 & n37121 ;
  assign n37123 = ~n37119 & ~n37122 ;
  assign n37124 = \wishbone_rx_fifo_fifo_reg[6][21]/P0001  & ~n37078 ;
  assign n37125 = \wishbone_RxDataLatched2_reg[21]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37126 = n37076 & n37125 ;
  assign n37127 = n36849 & n37126 ;
  assign n37128 = ~n37124 & ~n37127 ;
  assign n37129 = \wishbone_rx_fifo_fifo_reg[6][22]/P0001  & ~n37078 ;
  assign n37130 = \wishbone_RxDataLatched2_reg[22]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37131 = n37076 & n37130 ;
  assign n37132 = n36849 & n37131 ;
  assign n37133 = ~n37129 & ~n37132 ;
  assign n37134 = \wishbone_rx_fifo_fifo_reg[6][23]/P0001  & ~n37078 ;
  assign n37135 = \wishbone_RxDataLatched2_reg[23]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37136 = n37076 & n37135 ;
  assign n37137 = n36849 & n37136 ;
  assign n37138 = ~n37134 & ~n37137 ;
  assign n37139 = \wishbone_rx_fifo_fifo_reg[6][25]/P0001  & ~n37078 ;
  assign n37140 = \wishbone_RxDataLatched2_reg[25]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37141 = n37076 & n37140 ;
  assign n37142 = n36849 & n37141 ;
  assign n37143 = ~n37139 & ~n37142 ;
  assign n37144 = \wishbone_rx_fifo_fifo_reg[6][26]/P0001  & ~n37078 ;
  assign n37145 = \wishbone_RxDataLatched2_reg[26]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37146 = n37076 & n37145 ;
  assign n37147 = n36849 & n37146 ;
  assign n37148 = ~n37144 & ~n37147 ;
  assign n37149 = \wishbone_rx_fifo_fifo_reg[6][24]/P0001  & ~n37078 ;
  assign n37150 = \wishbone_RxDataLatched2_reg[24]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37151 = n37076 & n37150 ;
  assign n37152 = n36849 & n37151 ;
  assign n37153 = ~n37149 & ~n37152 ;
  assign n37154 = \wishbone_rx_fifo_fifo_reg[6][27]/P0001  & ~n37078 ;
  assign n37155 = \wishbone_RxDataLatched2_reg[27]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37156 = n37076 & n37155 ;
  assign n37157 = n36849 & n37156 ;
  assign n37158 = ~n37154 & ~n37157 ;
  assign n37159 = \wishbone_rx_fifo_fifo_reg[6][28]/P0001  & ~n37078 ;
  assign n37160 = \wishbone_RxDataLatched2_reg[28]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37161 = n37076 & n37160 ;
  assign n37162 = n36849 & n37161 ;
  assign n37163 = ~n37159 & ~n37162 ;
  assign n37164 = \wishbone_rx_fifo_fifo_reg[6][2]/P0001  & ~n37078 ;
  assign n37165 = \wishbone_RxDataLatched2_reg[2]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37166 = n37076 & n37165 ;
  assign n37167 = n36849 & n37166 ;
  assign n37168 = ~n37164 & ~n37167 ;
  assign n37169 = \wishbone_rx_fifo_fifo_reg[6][31]/P0001  & ~n37078 ;
  assign n37170 = \wishbone_RxDataLatched2_reg[31]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37171 = n37076 & n37170 ;
  assign n37172 = n36849 & n37171 ;
  assign n37173 = ~n37169 & ~n37172 ;
  assign n37174 = \wishbone_rx_fifo_fifo_reg[6][5]/P0001  & ~n37078 ;
  assign n37175 = \wishbone_RxDataLatched2_reg[5]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37176 = n37076 & n37175 ;
  assign n37177 = n36849 & n37176 ;
  assign n37178 = ~n37174 & ~n37177 ;
  assign n37179 = \wishbone_rx_fifo_fifo_reg[6][6]/P0001  & ~n37078 ;
  assign n37180 = \wishbone_RxDataLatched2_reg[6]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37181 = n37076 & n37180 ;
  assign n37182 = n36849 & n37181 ;
  assign n37183 = ~n37179 & ~n37182 ;
  assign n37184 = \wishbone_rx_fifo_fifo_reg[6][7]/P0001  & ~n37078 ;
  assign n37185 = \wishbone_RxDataLatched2_reg[7]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37186 = n37076 & n37185 ;
  assign n37187 = n36849 & n37186 ;
  assign n37188 = ~n37184 & ~n37187 ;
  assign n37189 = \wishbone_rx_fifo_fifo_reg[6][9]/P0001  & ~n37078 ;
  assign n37190 = \wishbone_RxDataLatched2_reg[9]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37191 = n37076 & n37190 ;
  assign n37192 = n36849 & n37191 ;
  assign n37193 = ~n37189 & ~n37192 ;
  assign n37194 = ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & ~\wishbone_rx_fifo_write_pointer_reg[2]/NET0131  ;
  assign n37195 = n35359 & n37194 ;
  assign n37196 = \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n37197 = ~n33164 & n37196 ;
  assign n37198 = n37195 & n37197 ;
  assign n37199 = ~n35365 & n37198 ;
  assign n37200 = \wishbone_rx_fifo_fifo_reg[9][0]/P0001  & ~n37199 ;
  assign n37201 = \wishbone_RxDataLatched2_reg[0]/NET0131  & n37199 ;
  assign n37202 = ~n37200 & ~n37201 ;
  assign n37203 = \wishbone_rx_fifo_fifo_reg[9][10]/P0001  & ~n37199 ;
  assign n37204 = \wishbone_RxDataLatched2_reg[10]/NET0131  & n37199 ;
  assign n37205 = ~n37203 & ~n37204 ;
  assign n37206 = \wishbone_rx_fifo_fifo_reg[9][11]/P0001  & ~n37199 ;
  assign n37207 = \wishbone_RxDataLatched2_reg[11]/NET0131  & n37199 ;
  assign n37208 = ~n37206 & ~n37207 ;
  assign n37209 = \wishbone_rx_fifo_fifo_reg[9][13]/P0001  & ~n37199 ;
  assign n37210 = \wishbone_RxDataLatched2_reg[13]/NET0131  & n37199 ;
  assign n37211 = ~n37209 & ~n37210 ;
  assign n37212 = \wishbone_rx_fifo_fifo_reg[9][16]/P0001  & ~n37199 ;
  assign n37213 = \wishbone_RxDataLatched2_reg[16]/NET0131  & n37199 ;
  assign n37214 = ~n37212 & ~n37213 ;
  assign n37215 = \wishbone_rx_fifo_fifo_reg[9][17]/P0001  & ~n37199 ;
  assign n37216 = \wishbone_RxDataLatched2_reg[17]/NET0131  & n37199 ;
  assign n37217 = ~n37215 & ~n37216 ;
  assign n37218 = \wishbone_rx_fifo_fifo_reg[9][18]/P0001  & ~n37199 ;
  assign n37219 = \wishbone_RxDataLatched2_reg[18]/NET0131  & n37199 ;
  assign n37220 = ~n37218 & ~n37219 ;
  assign n37221 = \wishbone_rx_fifo_fifo_reg[9][19]/P0001  & ~n37199 ;
  assign n37222 = \wishbone_RxDataLatched2_reg[19]/NET0131  & n37199 ;
  assign n37223 = ~n37221 & ~n37222 ;
  assign n37224 = \wishbone_rx_fifo_fifo_reg[9][1]/P0001  & ~n37199 ;
  assign n37225 = \wishbone_RxDataLatched2_reg[1]/NET0131  & n37199 ;
  assign n37226 = ~n37224 & ~n37225 ;
  assign n37227 = \wishbone_rx_fifo_fifo_reg[9][20]/P0001  & ~n37199 ;
  assign n37228 = \wishbone_RxDataLatched2_reg[20]/NET0131  & n37199 ;
  assign n37229 = ~n37227 & ~n37228 ;
  assign n37230 = \wishbone_rx_fifo_fifo_reg[9][21]/P0001  & ~n37199 ;
  assign n37231 = \wishbone_RxDataLatched2_reg[21]/NET0131  & n37199 ;
  assign n37232 = ~n37230 & ~n37231 ;
  assign n37233 = \wishbone_rx_fifo_fifo_reg[9][22]/P0001  & ~n37199 ;
  assign n37234 = \wishbone_RxDataLatched2_reg[22]/NET0131  & n37199 ;
  assign n37235 = ~n37233 & ~n37234 ;
  assign n37236 = \wishbone_rx_fifo_fifo_reg[9][23]/P0001  & ~n37199 ;
  assign n37237 = \wishbone_RxDataLatched2_reg[23]/NET0131  & n37199 ;
  assign n37238 = ~n37236 & ~n37237 ;
  assign n37239 = \wishbone_rx_fifo_fifo_reg[9][24]/P0001  & ~n37199 ;
  assign n37240 = \wishbone_RxDataLatched2_reg[24]/NET0131  & n37199 ;
  assign n37241 = ~n37239 & ~n37240 ;
  assign n37242 = \wishbone_rx_fifo_fifo_reg[9][25]/P0001  & ~n37199 ;
  assign n37243 = \wishbone_RxDataLatched2_reg[25]/NET0131  & n37199 ;
  assign n37244 = ~n37242 & ~n37243 ;
  assign n37245 = \wishbone_rx_fifo_fifo_reg[9][26]/P0001  & ~n37199 ;
  assign n37246 = \wishbone_RxDataLatched2_reg[26]/NET0131  & n37199 ;
  assign n37247 = ~n37245 & ~n37246 ;
  assign n37248 = \wishbone_rx_fifo_fifo_reg[9][27]/P0001  & ~n37199 ;
  assign n37249 = \wishbone_RxDataLatched2_reg[27]/NET0131  & n37199 ;
  assign n37250 = ~n37248 & ~n37249 ;
  assign n37251 = \wishbone_rx_fifo_fifo_reg[9][29]/P0001  & ~n37199 ;
  assign n37252 = \wishbone_RxDataLatched2_reg[29]/NET0131  & n37199 ;
  assign n37253 = ~n37251 & ~n37252 ;
  assign n37254 = \wishbone_rx_fifo_fifo_reg[9][2]/P0001  & ~n37199 ;
  assign n37255 = \wishbone_RxDataLatched2_reg[2]/NET0131  & n37199 ;
  assign n37256 = ~n37254 & ~n37255 ;
  assign n37257 = \wishbone_rx_fifo_fifo_reg[9][30]/P0001  & ~n37199 ;
  assign n37258 = \wishbone_RxDataLatched2_reg[30]/NET0131  & n37199 ;
  assign n37259 = ~n37257 & ~n37258 ;
  assign n37260 = \wishbone_rx_fifo_fifo_reg[9][4]/P0001  & ~n37199 ;
  assign n37261 = \wishbone_RxDataLatched2_reg[4]/NET0131  & n37199 ;
  assign n37262 = ~n37260 & ~n37261 ;
  assign n37263 = \wishbone_rx_fifo_fifo_reg[9][5]/P0001  & ~n37199 ;
  assign n37264 = \wishbone_RxDataLatched2_reg[5]/NET0131  & n37199 ;
  assign n37265 = ~n37263 & ~n37264 ;
  assign n37266 = \wishbone_rx_fifo_fifo_reg[9][7]/P0001  & ~n37199 ;
  assign n37267 = \wishbone_RxDataLatched2_reg[7]/NET0131  & n37199 ;
  assign n37268 = ~n37266 & ~n37267 ;
  assign n37269 = \wishbone_rx_fifo_fifo_reg[9][9]/P0001  & ~n37199 ;
  assign n37270 = \wishbone_RxDataLatched2_reg[9]/NET0131  & n37199 ;
  assign n37271 = ~n37269 & ~n37270 ;
  assign n37272 = \wishbone_tx_fifo_cnt_reg[0]/NET0131  & n34242 ;
  assign n37273 = n35309 & n37272 ;
  assign n37274 = ~n35309 & ~n37272 ;
  assign n37275 = ~n37273 & ~n37274 ;
  assign n37276 = n37076 & n37194 ;
  assign n37277 = ~n33164 & ~n37276 ;
  assign n37278 = n36771 & ~n37277 ;
  assign n37279 = n36789 & n37196 ;
  assign n37280 = ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n37196 ;
  assign n37281 = n36849 & n37280 ;
  assign n37282 = \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n36785 ;
  assign n37283 = n36849 & n37282 ;
  assign n37284 = \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n37196 ;
  assign n37285 = n36849 & n37284 ;
  assign n37286 = ~n33164 & n36932 ;
  assign n37287 = n37195 & n37286 ;
  assign n37288 = ~n35365 & n37287 ;
  assign n37289 = n36789 & n37076 ;
  assign n37290 = ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n37076 ;
  assign n37291 = n36849 & n37290 ;
  assign n37292 = \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & n36932 ;
  assign n37293 = n36849 & n37292 ;
  assign n37294 = n36785 & n37194 ;
  assign n37295 = n36786 & n37294 ;
  assign n37296 = ~n35365 & n37295 ;
  assign n37297 = \miim1_LatchByte_reg[0]/NET0131  & n32545 ;
  assign n37298 = n32531 & n37297 ;
  assign n37299 = n32513 & n37298 ;
  assign n37300 = n35298 & ~n35306 ;
  assign n37301 = \wishbone_tx_fifo_read_pointer_reg[0]/NET0131  & n34242 ;
  assign n37302 = ~n37300 & n37301 ;
  assign n37303 = n35298 & ~n37301 ;
  assign n37304 = ~n35306 & n37303 ;
  assign n37305 = ~n37302 & ~n37304 ;
  assign n37306 = ~n11732 & ~n11734 ;
  assign n37307 = \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37308 = n35523 & n37307 ;
  assign n37309 = ~\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  ;
  assign n37310 = n36393 & ~n37309 ;
  assign n37311 = ~n37308 & ~n37310 ;
  assign n37312 = n36379 & ~n37311 ;
  assign n37313 = ~n35522 & ~n36369 ;
  assign n37314 = n36380 & ~n37313 ;
  assign n37315 = \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37316 = n35523 & n37315 ;
  assign n37317 = n35522 & n37316 ;
  assign n37318 = \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37319 = n36360 & n37318 ;
  assign n37320 = n36369 & n37319 ;
  assign n37321 = ~n37317 & ~n37320 ;
  assign n37322 = ~n37314 & n37321 ;
  assign n37323 = \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37324 = n36360 & n37323 ;
  assign n37325 = n36389 & n37324 ;
  assign n37326 = \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37327 = n36368 & n37326 ;
  assign n37328 = n36373 & n37327 ;
  assign n37329 = ~n37325 & ~n37328 ;
  assign n37330 = \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37331 = n35521 & n37330 ;
  assign n37332 = n36373 & n37331 ;
  assign n37333 = \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37334 = n36362 & n37333 ;
  assign n37335 = n36389 & n37334 ;
  assign n37336 = ~n37332 & ~n37335 ;
  assign n37337 = n37329 & n37336 ;
  assign n37338 = n37322 & n37337 ;
  assign n37339 = ~n37312 & n37338 ;
  assign n37340 = n16307 & n33170 ;
  assign n37341 = ~n13129 & n37340 ;
  assign n37342 = \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  & n37341 ;
  assign n37343 = \wishbone_rx_fifo_read_pointer_reg[3]/NET0131  & ~n33164 ;
  assign n37344 = ~n37342 & n37343 ;
  assign n37345 = ~\wishbone_rx_fifo_read_pointer_reg[3]/NET0131  & ~n33164 ;
  assign n37346 = n37342 & n37345 ;
  assign n37347 = ~n37344 & ~n37346 ;
  assign n37348 = ~n35308 & ~n35310 ;
  assign n37349 = ~n35300 & n35305 ;
  assign n37350 = ~n37348 & ~n37349 ;
  assign n37351 = \wishbone_tx_fifo_cnt_reg[2]/NET0131  & n34242 ;
  assign n37352 = ~n37350 & n37351 ;
  assign n37353 = ~\wishbone_tx_fifo_cnt_reg[2]/NET0131  & n34242 ;
  assign n37354 = n37350 & n37353 ;
  assign n37355 = ~n37352 & ~n37354 ;
  assign n37356 = ~\wishbone_tx_fifo_read_pointer_reg[1]/NET0131  & ~n35298 ;
  assign n37357 = ~\wishbone_tx_fifo_read_pointer_reg[1]/NET0131  & n35302 ;
  assign n37358 = n35301 & n37357 ;
  assign n37359 = ~n37356 & ~n37358 ;
  assign n37360 = ~n34248 & ~n34252 ;
  assign n37361 = n35298 & n37360 ;
  assign n37362 = ~n35306 & n37361 ;
  assign n37363 = n34242 & ~n37362 ;
  assign n37364 = n37359 & n37363 ;
  assign n37365 = \wishbone_tx_fifo_read_pointer_reg[2]/NET0131  & n35298 ;
  assign n37366 = n34259 & n37365 ;
  assign n37367 = ~n35306 & n37366 ;
  assign n37368 = ~\wishbone_tx_fifo_read_pointer_reg[3]/NET0131  & ~n37367 ;
  assign n37369 = n34272 & n35298 ;
  assign n37370 = ~n35306 & n37369 ;
  assign n37371 = n34242 & ~n37370 ;
  assign n37372 = ~n37368 & n37371 ;
  assign n37373 = \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
  assign n37374 = n35359 & n37373 ;
  assign n37375 = ~n35365 & n37374 ;
  assign n37376 = \wishbone_rx_fifo_write_pointer_reg[2]/NET0131  & ~n33164 ;
  assign n37377 = ~n37375 & n37376 ;
  assign n37378 = ~\wishbone_rx_fifo_write_pointer_reg[2]/NET0131  & ~n33164 ;
  assign n37379 = n37375 & n37378 ;
  assign n37380 = ~n37377 & ~n37379 ;
  assign n37381 = \wishbone_rx_fifo_write_pointer_reg[2]/NET0131  & \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
  assign n37382 = n37375 & n37381 ;
  assign n37383 = \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  & ~n33164 ;
  assign n37384 = n37375 & n37376 ;
  assign n37385 = ~n37383 & ~n37384 ;
  assign n37386 = ~n37382 & ~n37385 ;
  assign n37387 = \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  & n34242 ;
  assign n37388 = ~n35762 & n37387 ;
  assign n37389 = ~\wishbone_tx_fifo_write_pointer_reg[2]/NET0131  & n34242 ;
  assign n37390 = n35762 & n37389 ;
  assign n37391 = ~n37388 & ~n37390 ;
  assign n37392 = \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  & n35762 ;
  assign n37393 = n35747 & n37392 ;
  assign n37394 = \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  & n34242 ;
  assign n37395 = ~n37392 & n37394 ;
  assign n37396 = ~n37393 & ~n37395 ;
  assign n37397 = \wishbone_TxEn_reg/NET0131  & ~n36420 ;
  assign n37398 = n36419 & n37397 ;
  assign n37399 = ~n36412 & ~n37398 ;
  assign n37400 = n10525 & ~n12580 ;
  assign n37401 = ~n10648 & n37400 ;
  assign n37402 = ~n12168 & ~n37401 ;
  assign n37403 = \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  & n35359 ;
  assign n37404 = ~n35365 & n37403 ;
  assign n37405 = ~\wishbone_rx_fifo_write_pointer_reg[1]/NET0131  & ~n37404 ;
  assign n37406 = ~n33164 & ~n37375 ;
  assign n37407 = ~n37405 & n37406 ;
  assign n37408 = \wishbone_tx_fifo_cnt_reg[1]/NET0131  & n35309 ;
  assign n37409 = ~n35300 & ~n35310 ;
  assign n37410 = n35307 & ~n37409 ;
  assign n37411 = ~n35306 & n37410 ;
  assign n37412 = ~n35305 & n37409 ;
  assign n37413 = ~n37411 & ~n37412 ;
  assign n37414 = ~n37408 & n37413 ;
  assign n37415 = n34242 & ~n37414 ;
  assign n37416 = n34259 & n35298 ;
  assign n37417 = ~n35306 & n37416 ;
  assign n37418 = ~\wishbone_tx_fifo_read_pointer_reg[2]/NET0131  & ~n37417 ;
  assign n37419 = n34242 & ~n37367 ;
  assign n37420 = ~n37418 & n37419 ;
  assign n37421 = ~\wishbone_tx_fifo_write_pointer_reg[1]/NET0131  & ~n36781 ;
  assign n37422 = n34242 & ~n35762 ;
  assign n37423 = ~n37421 & n37422 ;
  assign n37424 = \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  & ~\maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131  ;
  assign n37425 = n11464 & n11608 ;
  assign n37426 = n23741 & n23794 ;
  assign n37427 = ~\wb_adr_i[11]_pad  & \wb_sel_i[2]_pad  ;
  assign n37428 = n23726 & n37427 ;
  assign n37429 = ~n23725 & n37428 ;
  assign n37430 = n32819 & n37429 ;
  assign n37431 = n37426 & n37430 ;
  assign n37432 = ~\ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131  & ~n37431 ;
  assign n37433 = ~\wb_dat_i[16]_pad  & n23794 ;
  assign n37434 = n23741 & n37433 ;
  assign n37435 = n37430 & n37434 ;
  assign n37436 = ~\RstTxPauseRq_reg/NET0131  & ~n37435 ;
  assign n37437 = ~n37432 & n37436 ;
  assign n37438 = ~\RxAbort_wb_reg/NET0131  & ~\rxethmac1_RxEndFrm_reg/NET0131  ;
  assign n37439 = \wishbone_RxEnableWindow_reg/NET0131  & n37438 ;
  assign n37440 = ~\rxethmac1_RxStartFrm_reg/NET0131  & ~n37439 ;
  assign n37441 = \miim1_clkgen_Counter_reg[0]/NET0131  & \miim1_clkgen_Counter_reg[1]/NET0131  ;
  assign n37442 = ~n32247 & ~n37441 ;
  assign n37443 = ~n32264 & n37442 ;
  assign n37444 = \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  & ~\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  ;
  assign n37445 = ~\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  & \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  ;
  assign n37446 = ~n37444 & ~n37445 ;
  assign n37447 = ~\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  & ~\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  ;
  assign n37448 = ~\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  & n37447 ;
  assign n37449 = n32255 & n37448 ;
  assign n37450 = n37446 & ~n37449 ;
  assign n37451 = n32264 & ~n37450 ;
  assign n37452 = ~n37443 & ~n37451 ;
  assign n37453 = \rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131  & ~n13066 ;
  assign n37454 = ~\ethreg1_MODER_0_DataOut_reg[3]/NET0131  & \rxethmac1_Broadcast_reg/NET0131  ;
  assign n37455 = ~\rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131  & ~\rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131  ;
  assign n37456 = ~n37454 & n37455 ;
  assign n37457 = \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  & \maccontrol1_receivecontrol1_AddressOK_reg/NET0131  ;
  assign n37458 = n37456 & ~n37457 ;
  assign n37459 = n12580 & n13051 ;
  assign n37460 = n37458 & n37459 ;
  assign n37461 = n10564 & n37460 ;
  assign n37462 = ~n37453 & ~n37461 ;
  assign n37463 = \wishbone_ram_di_reg[11]/NET0131  & ~n36420 ;
  assign n37464 = n36419 & n37463 ;
  assign n37465 = \wb_dat_i[11]_pad  & n36417 ;
  assign n37466 = ~n36415 & n37465 ;
  assign n37467 = \wishbone_TxEn_needed_reg/NET0131  & \wishbone_TxStatus_reg[11]/NET0131  ;
  assign n37468 = ~n36411 & n37467 ;
  assign n37469 = ~n37466 & ~n37468 ;
  assign n37470 = ~n37464 & n37469 ;
  assign n37471 = \wishbone_ram_di_reg[12]/NET0131  & ~n36420 ;
  assign n37472 = n36419 & n37471 ;
  assign n37473 = \wb_dat_i[12]_pad  & n36417 ;
  assign n37474 = ~n36415 & n37473 ;
  assign n37475 = \wishbone_TxEn_needed_reg/NET0131  & \wishbone_TxStatus_reg[12]/NET0131  ;
  assign n37476 = ~n36411 & n37475 ;
  assign n37477 = ~n37474 & ~n37476 ;
  assign n37478 = ~n37472 & n37477 ;
  assign n37479 = \txethmac1_random1_RandomLatched_reg[8]/NET0131  & ~n36399 ;
  assign n37480 = ~\txethmac1_RetryCnt_reg[0]/NET0131  & ~\txethmac1_RetryCnt_reg[1]/NET0131  ;
  assign n37481 = ~\txethmac1_RetryCnt_reg[2]/NET0131  & n37480 ;
  assign n37482 = \txethmac1_RetryCnt_reg[3]/NET0131  & \txethmac1_random1_x_reg[8]/NET0131  ;
  assign n37483 = n36399 & n37482 ;
  assign n37484 = ~n37481 & n37483 ;
  assign n37485 = ~n37479 & ~n37484 ;
  assign n37486 = \wishbone_BDRead_reg/NET0131  & ~n36417 ;
  assign n37487 = \wishbone_BDRead_reg/NET0131  & ~\wishbone_TxEn_q_reg/NET0131  ;
  assign n37488 = ~n36414 & n37487 ;
  assign n37489 = ~n37486 & ~n37488 ;
  assign n37490 = ~\wb_adr_i[11]_pad  & n23726 ;
  assign n37491 = ~n23725 & n37490 ;
  assign n37492 = \wb_adr_i[10]_pad  & ~wb_we_i_pad ;
  assign n37493 = n37491 & n37492 ;
  assign n37494 = n36418 & n37493 ;
  assign n37495 = n37489 & ~n37494 ;
  assign n37496 = \wishbone_TxAbort_wb_q_reg/NET0131  & ~\wishbone_TxAbort_wb_reg/NET0131  ;
  assign n37497 = ~\wishbone_TxAbortPacketBlocked_reg/NET0131  & ~\wishbone_TxAbortPacket_reg/NET0131  ;
  assign n37498 = ~n37496 & ~n37497 ;
  assign n37499 = \wishbone_TxDone_wb_q_reg/NET0131  & ~\wishbone_TxDone_wb_reg/NET0131  ;
  assign n37500 = ~\wishbone_TxDonePacketBlocked_reg/NET0131  & ~\wishbone_TxDonePacket_reg/NET0131  ;
  assign n37501 = ~n37499 & ~n37500 ;
  assign n37502 = ~\txethmac1_random1_x_reg[2]/NET0131  & ~\txethmac1_random1_x_reg[9]/NET0131  ;
  assign n37503 = \txethmac1_random1_x_reg[2]/NET0131  & \txethmac1_random1_x_reg[9]/NET0131  ;
  assign n37504 = ~n37502 & ~n37503 ;
  assign n37505 = \macstatus1_LoadRxStatus_reg/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n37506 = ~n11671 & n37505 ;
  assign n37507 = \macstatus1_LoadRxStatus_reg/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
  assign n37508 = n11671 & n37507 ;
  assign n37509 = ~n37506 & ~n37508 ;
  assign n37510 = ~\macstatus1_LoadRxStatus_reg/NET0131  & ~\wishbone_LatchedRxLength_reg[11]/NET0131  ;
  assign n37511 = n37509 & ~n37510 ;
  assign n37512 = \TPauseRq_reg/NET0131  & \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  ;
  assign n37513 = ~\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131  & ~n37512 ;
  assign n37514 = ~n10692 & ~n37513 ;
  assign n37515 = n10984 & n11008 ;
  assign n37516 = n10986 & ~n37515 ;
  assign n37517 = \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  & ~wb_rst_i_pad ;
  assign n37518 = ~n11983 & n37517 ;
  assign n37519 = ~\maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  & ~wb_rst_i_pad ;
  assign n37520 = n11983 & n37519 ;
  assign n37521 = ~n37518 & ~n37520 ;
  assign n37522 = ~\wishbone_TxBDAddress_reg[1]/NET0131  & ~n36308 ;
  assign n37523 = ~\wishbone_BlockingTxStatusWrite_reg/NET0131  & \wishbone_TxBDAddress_reg[1]/NET0131  ;
  assign n37524 = n36303 & n37523 ;
  assign n37525 = ~n36301 & ~n37524 ;
  assign n37526 = ~n37522 & n37525 ;
  assign n37527 = \wishbone_TxBDAddress_reg[2]/NET0131  & ~n36304 ;
  assign n37528 = ~\wishbone_TxBDAddress_reg[1]/NET0131  & ~\wishbone_TxBDAddress_reg[2]/NET0131  ;
  assign n37529 = ~n36310 & ~n37528 ;
  assign n37530 = n36308 & n37529 ;
  assign n37531 = ~n37527 & ~n37530 ;
  assign n37532 = ~n36301 & ~n37531 ;
  assign n37533 = \wishbone_TxBDAddress_reg[3]/NET0131  & ~n36304 ;
  assign n37534 = ~\wishbone_TxBDAddress_reg[3]/NET0131  & ~n36310 ;
  assign n37535 = ~n36311 & ~n37534 ;
  assign n37536 = n36308 & n37535 ;
  assign n37537 = ~n37533 & ~n37536 ;
  assign n37538 = ~n36301 & ~n37537 ;
  assign n37539 = \wishbone_TxBDAddress_reg[5]/NET0131  & ~n36304 ;
  assign n37540 = ~\wishbone_TxBDAddress_reg[5]/NET0131  & ~n36314 ;
  assign n37541 = n36308 & ~n36325 ;
  assign n37542 = ~n37540 & n37541 ;
  assign n37543 = ~n37539 & ~n37542 ;
  assign n37544 = ~n36301 & ~n37543 ;
  assign n37545 = \wishbone_Flop_reg/NET0131  & \wishbone_TxByteCnt_reg[0]/NET0131  ;
  assign n37546 = n12725 & n37545 ;
  assign n37547 = ~\wishbone_TxByteCnt_reg[0]/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n37548 = ~n12725 & n37547 ;
  assign n37549 = ~\wishbone_Flop_reg/NET0131  & ~\wishbone_TxByteCnt_reg[0]/NET0131  ;
  assign n37550 = n12725 & n37549 ;
  assign n37551 = ~n37548 & ~n37550 ;
  assign n37552 = ~n37546 & n37551 ;
  assign n37553 = \wishbone_TxPointerLSB_reg[0]/NET0131  & \wishbone_TxStartFrm_reg/NET0131  ;
  assign n37554 = ~n12725 & n37553 ;
  assign n37555 = ~\wishbone_TxAbort_q_reg/NET0131  & ~\wishbone_TxRetry_q_reg/NET0131  ;
  assign n37556 = ~n37554 & n37555 ;
  assign n37557 = n37552 & n37556 ;
  assign n37558 = \wishbone_TxStartFrm_reg/NET0131  & ~n12725 ;
  assign n37559 = ~n12753 & ~n12756 ;
  assign n37560 = n37558 & ~n37559 ;
  assign n37561 = n37555 & n37560 ;
  assign n37562 = ~\wishbone_TxByteCnt_reg[1]/NET0131  & ~n37546 ;
  assign n37563 = ~n37558 & ~n37562 ;
  assign n37564 = \wishbone_TxByteCnt_reg[1]/NET0131  & n37546 ;
  assign n37565 = n37555 & ~n37564 ;
  assign n37566 = n37563 & n37565 ;
  assign n37567 = ~n37561 & ~n37566 ;
  assign n37568 = ~\wishbone_TxEn_needed_reg/NET0131  & n36408 ;
  assign n37569 = \wishbone_WbEn_reg/NET0131  & ~n37568 ;
  assign n37570 = ~n36420 & n37569 ;
  assign n37571 = n36419 & n37570 ;
  assign n37572 = ~n36418 & ~n37571 ;
  assign n37573 = ~\miim1_BitCounter_reg[5]/NET0131  & n32526 ;
  assign n37574 = n36353 & ~n37573 ;
  assign n37575 = \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  & n36265 ;
  assign n37576 = ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  & ~n37575 ;
  assign n37577 = ~n36267 & n36273 ;
  assign n37578 = ~n37576 & n37577 ;
  assign n37579 = ~\wishbone_WB_ACK_O_reg/P0001  & ~n23729 ;
  assign n37580 = ~wb_ack_o_pad & ~n37579 ;
  assign n37581 = n25057 & n35834 ;
  assign n37582 = \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  & n11980 ;
  assign n37583 = ~\maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131  & ~n37582 ;
  assign n37584 = ~wb_rst_i_pad & ~n36286 ;
  assign n37585 = ~n37583 & n37584 ;
  assign n37586 = n23794 & n35890 ;
  assign n37587 = \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37588 = n35521 & n37587 ;
  assign n37589 = n36373 & n37588 ;
  assign n37590 = \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37591 = n36360 & n37590 ;
  assign n37592 = n36389 & n37591 ;
  assign n37593 = \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37594 = n35523 & n37593 ;
  assign n37595 = n36379 & n37594 ;
  assign n37596 = ~n37592 & ~n37595 ;
  assign n37597 = ~n37589 & n37596 ;
  assign n37598 = \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37599 = n36360 & n37598 ;
  assign n37600 = n36369 & n37599 ;
  assign n37601 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & n35800 ;
  assign n37602 = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37603 = n37601 & n37602 ;
  assign n37604 = ~n37600 & ~n37603 ;
  assign n37605 = \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37606 = n36362 & n37605 ;
  assign n37607 = n36389 & n37606 ;
  assign n37608 = \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37609 = n36368 & n37608 ;
  assign n37610 = n36373 & n37609 ;
  assign n37611 = ~n37607 & ~n37610 ;
  assign n37612 = \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37613 = n35523 & n37612 ;
  assign n37614 = n35522 & n37613 ;
  assign n37615 = \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37616 = n36362 & n37615 ;
  assign n37617 = n36379 & n37616 ;
  assign n37618 = ~n37614 & ~n37617 ;
  assign n37619 = n37611 & n37618 ;
  assign n37620 = n37604 & n37619 ;
  assign n37621 = n37597 & n37620 ;
  assign n37622 = ~\macstatus1_DribbleNibble_reg/NET0131  & ~n12164 ;
  assign n37623 = ~\rxethmac1_rxstatem1_StateSFD_reg/NET0131  & ~n37622 ;
  assign n37624 = ~\rxethmac1_crcrx_Crc_reg[28]/NET0131  & n10567 ;
  assign n37625 = n10564 & n37624 ;
  assign n37626 = \rxethmac1_CrcHash_reg[2]/P0001  & n10570 ;
  assign n37627 = n10567 & n10570 ;
  assign n37628 = n10564 & n37627 ;
  assign n37629 = ~n37626 & ~n37628 ;
  assign n37630 = ~n37625 & ~n37629 ;
  assign n37631 = ~\rxethmac1_crcrx_Crc_reg[29]/NET0131  & n10567 ;
  assign n37632 = n10564 & n37631 ;
  assign n37633 = \rxethmac1_CrcHash_reg[3]/P0001  & n10570 ;
  assign n37634 = ~n37628 & ~n37633 ;
  assign n37635 = ~n37632 & ~n37634 ;
  assign n37636 = ~\rxethmac1_crcrx_Crc_reg[30]/NET0131  & n10567 ;
  assign n37637 = n10564 & n37636 ;
  assign n37638 = \rxethmac1_CrcHash_reg[4]/P0001  & n10570 ;
  assign n37639 = ~n37628 & ~n37638 ;
  assign n37640 = ~n37637 & ~n37639 ;
  assign n37641 = ~\rxethmac1_crcrx_Crc_reg[31]/NET0131  & n10567 ;
  assign n37642 = n10564 & n37641 ;
  assign n37643 = \rxethmac1_CrcHash_reg[5]/P0001  & n10570 ;
  assign n37644 = ~n37628 & ~n37643 ;
  assign n37645 = ~n37642 & ~n37644 ;
  assign n37646 = ~\wishbone_ReadTxDataFromMemory_reg/NET0131  & ~n18545 ;
  assign n37647 = n35550 & ~n37646 ;
  assign n37648 = ~n36338 & n37647 ;
  assign n37649 = \wishbone_RxEn_reg/NET0131  & n36419 ;
  assign n37650 = ~n36420 & ~n37649 ;
  assign n37651 = mdc_pad_o_pad & ~n32264 ;
  assign n37652 = ~n35338 & ~n37651 ;
  assign n37653 = \rxethmac1_LatchedByte_reg[1]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n37654 = ~n33020 & n37653 ;
  assign n37655 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[1]/NET0131  ;
  assign n37656 = ~n33021 & n37655 ;
  assign n37657 = ~n37654 & ~n37656 ;
  assign n37658 = \rxethmac1_LatchedByte_reg[2]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n37659 = ~n33020 & n37658 ;
  assign n37660 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[2]/NET0131  ;
  assign n37661 = ~n33021 & n37660 ;
  assign n37662 = ~n37659 & ~n37661 ;
  assign n37663 = \rxethmac1_LatchedByte_reg[3]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n37664 = ~n33020 & n37663 ;
  assign n37665 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[3]/NET0131  ;
  assign n37666 = ~n33021 & n37665 ;
  assign n37667 = ~n37664 & ~n37666 ;
  assign n37668 = \rxethmac1_LatchedByte_reg[5]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n37669 = ~n33020 & n37668 ;
  assign n37670 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[5]/NET0131  ;
  assign n37671 = ~n33021 & n37670 ;
  assign n37672 = ~n37669 & ~n37671 ;
  assign n37673 = \rxethmac1_LatchedByte_reg[6]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n37674 = ~n33020 & n37673 ;
  assign n37675 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[6]/NET0131  ;
  assign n37676 = ~n33021 & n37675 ;
  assign n37677 = ~n37674 & ~n37676 ;
  assign n37678 = \rxethmac1_LatchedByte_reg[7]/NET0131  & \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
  assign n37679 = ~n33020 & n37678 ;
  assign n37680 = \rxethmac1_DelayData_reg/NET0131  & \rxethmac1_RxData_d_reg[7]/NET0131  ;
  assign n37681 = ~n33021 & n37680 ;
  assign n37682 = ~n37679 & ~n37681 ;
  assign n37683 = \ethreg1_MODER_1_DataOut_reg[4]/NET0131  & ~n36269 ;
  assign n37684 = n10580 & n37683 ;
  assign n37685 = n36265 & ~n36269 ;
  assign n37686 = ~\ethreg1_MODER_1_DataOut_reg[4]/NET0131  & ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  ;
  assign n37687 = ~n36269 & n37686 ;
  assign n37688 = ~n37685 & ~n37687 ;
  assign n37689 = ~n37684 & n37688 ;
  assign n37690 = ~n36272 & n37689 ;
  assign n37691 = \wb_adr_i[2]_pad  & ~\wb_adr_i[3]_pad  ;
  assign n37692 = n35834 & n37691 ;
  assign n37693 = ~\wb_adr_i[5]_pad  & n23734 ;
  assign n37694 = n23733 & n37693 ;
  assign n37695 = ~\wb_adr_i[4]_pad  & n32819 ;
  assign n37696 = n32818 & n37695 ;
  assign n37697 = n37694 & n37696 ;
  assign n37698 = \wishbone_TxByteCnt_reg[1]/NET0131  & ~\wishbone_TxEndFrm_wb_reg/NET0131  ;
  assign n37699 = n37546 & n37698 ;
  assign n37700 = ~\txethmac1_TxRetry_reg/NET0131  & ~\wishbone_TxEndFrm_reg/NET0131  ;
  assign n37701 = \wishbone_Flop_reg/NET0131  & ~n37700 ;
  assign n37702 = ~\maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n37703 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\txethmac1_TxAbort_reg/NET0131  ;
  assign n37704 = n37702 & ~n37703 ;
  assign n37705 = ~\maccontrol1_MuxedAbort_reg/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n37706 = \wishbone_Flop_reg/NET0131  & ~n37705 ;
  assign n37707 = n37704 & n37706 ;
  assign n37708 = ~n37701 & ~n37707 ;
  assign n37709 = ~\wishbone_LastWord_reg/NET0131  & ~n37564 ;
  assign n37710 = n37708 & ~n37709 ;
  assign n37711 = ~n37699 & n37710 ;
  assign n37712 = \wishbone_BDWrite_reg[0]/NET0131  & ~n36417 ;
  assign n37713 = \wishbone_BDWrite_reg[0]/NET0131  & ~\wishbone_TxEn_q_reg/NET0131  ;
  assign n37714 = ~n36414 & n37713 ;
  assign n37715 = ~n37712 & ~n37714 ;
  assign n37716 = \wb_adr_i[10]_pad  & wb_we_i_pad ;
  assign n37717 = n36417 & n37716 ;
  assign n37718 = ~n36415 & n37717 ;
  assign n37719 = n32818 & n37718 ;
  assign n37720 = n37715 & ~n37719 ;
  assign n37721 = \wishbone_BDWrite_reg[1]/NET0131  & ~n36417 ;
  assign n37722 = \wishbone_BDWrite_reg[1]/NET0131  & ~\wishbone_TxEn_q_reg/NET0131  ;
  assign n37723 = ~n36414 & n37722 ;
  assign n37724 = ~n37721 & ~n37723 ;
  assign n37725 = ~\wb_adr_i[11]_pad  & \wb_sel_i[1]_pad  ;
  assign n37726 = n23726 & n37725 ;
  assign n37727 = ~n23725 & n37726 ;
  assign n37728 = n37718 & n37727 ;
  assign n37729 = n37724 & ~n37728 ;
  assign n37730 = \wishbone_BDWrite_reg[2]/NET0131  & ~n36417 ;
  assign n37731 = \wishbone_BDWrite_reg[2]/NET0131  & ~\wishbone_TxEn_q_reg/NET0131  ;
  assign n37732 = ~n36414 & n37731 ;
  assign n37733 = ~n37730 & ~n37732 ;
  assign n37734 = n37429 & n37718 ;
  assign n37735 = n37733 & ~n37734 ;
  assign n37736 = ~\wishbone_LastWord_reg/NET0131  & \wishbone_TxByteCnt_reg[1]/NET0131  ;
  assign n37737 = n37546 & n37736 ;
  assign n37738 = \wishbone_TxStartFrm_reg/NET0131  & n12738 ;
  assign n37739 = n12728 & n37738 ;
  assign n37740 = \wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131  & ~\wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131  ;
  assign n37741 = \wishbone_ReadTxDataFromFifo_tck_reg/NET0131  & ~n37740 ;
  assign n37742 = ~n12747 & ~n37741 ;
  assign n37743 = ~n37739 & n37742 ;
  assign n37744 = ~n37737 & n37743 ;
  assign n37745 = n32255 & n37447 ;
  assign n37746 = ~\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  & ~n37745 ;
  assign n37747 = n32264 & ~n37746 ;
  assign n37748 = \miim1_clkgen_Counter_reg[0]/NET0131  & ~n32264 ;
  assign n37749 = ~n37747 & ~n37748 ;
  assign n37750 = \wishbone_TxAbortPacket_NotCleared_reg/NET0131  & ~n14045 ;
  assign n37751 = ~\wishbone_tx_burst_en_reg/NET0131  & ~n13131 ;
  assign n37752 = \wishbone_MasterWbTX_reg/NET0131  & ~n37751 ;
  assign n37753 = ~\wishbone_TxAbortPacketBlocked_reg/NET0131  & \wishbone_TxAbort_wb_reg/NET0131  ;
  assign n37754 = ~\wishbone_TxAbortPacket_NotCleared_reg/NET0131  & n37753 ;
  assign n37755 = ~n37752 & n37754 ;
  assign n37756 = ~n37750 & ~n37755 ;
  assign n37757 = \wishbone_TxDonePacket_NotCleared_reg/NET0131  & ~n14045 ;
  assign n37758 = ~\wishbone_TxDonePacketBlocked_reg/NET0131  & \wishbone_TxDone_wb_reg/NET0131  ;
  assign n37759 = ~\wishbone_TxDonePacket_NotCleared_reg/NET0131  & n37758 ;
  assign n37760 = ~n37752 & n37759 ;
  assign n37761 = ~n37757 & ~n37760 ;
  assign n37762 = n16307 & n33164 ;
  assign n37763 = ~\wishbone_rx_fifo_read_pointer_reg[0]/NET0131  & ~n16307 ;
  assign n37764 = ~\wishbone_rx_fifo_read_pointer_reg[0]/NET0131  & n13128 ;
  assign n37765 = n13127 & n37764 ;
  assign n37766 = ~n37763 & ~n37765 ;
  assign n37767 = \wishbone_rx_fifo_read_pointer_reg[0]/NET0131  & n16307 ;
  assign n37768 = ~n13129 & n37767 ;
  assign n37769 = ~n33164 & ~n37768 ;
  assign n37770 = n37766 & n37769 ;
  assign n37771 = ~n37762 & ~n37770 ;
  assign n37772 = \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131  & ~n35448 ;
  assign n37773 = ~\wishbone_RxBDAddress_reg[2]/NET0131  & ~n35924 ;
  assign n37774 = n35448 & ~n35925 ;
  assign n37775 = ~n37773 & n37774 ;
  assign n37776 = ~n37772 & ~n37775 ;
  assign n37777 = \wb_dat_i[10]_pad  & n36417 ;
  assign n37778 = ~n36415 & n37777 ;
  assign n37779 = \wishbone_ram_di_reg[10]/NET0131  & ~n36420 ;
  assign n37780 = n36419 & n37779 ;
  assign n37781 = ~n37778 & ~n37780 ;
  assign n37782 = \wb_dat_i[15]_pad  & n36417 ;
  assign n37783 = ~n36415 & n37782 ;
  assign n37784 = \wishbone_ram_di_reg[15]/NET0131  & ~n36420 ;
  assign n37785 = n36419 & n37784 ;
  assign n37786 = ~n37783 & ~n37785 ;
  assign n37787 = \wb_dat_i[9]_pad  & n36417 ;
  assign n37788 = ~n36415 & n37787 ;
  assign n37789 = \wishbone_ram_di_reg[9]/NET0131  & ~n36420 ;
  assign n37790 = n36419 & n37789 ;
  assign n37791 = ~n37788 & ~n37790 ;
  assign n37792 = \macstatus1_LoadRxStatus_reg/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n37793 = ~n11668 & n37792 ;
  assign n37794 = \macstatus1_LoadRxStatus_reg/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
  assign n37795 = n11668 & n37794 ;
  assign n37796 = ~n37793 & ~n37795 ;
  assign n37797 = ~\macstatus1_LoadRxStatus_reg/NET0131  & \wishbone_LatchedRxLength_reg[8]/NET0131  ;
  assign n37798 = n37796 & ~n37797 ;
  assign n37799 = \macstatus1_LoadRxStatus_reg/NET0131  & ~\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n37800 = ~n11734 & n37799 ;
  assign n37801 = \macstatus1_LoadRxStatus_reg/NET0131  & \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
  assign n37802 = n11734 & n37801 ;
  assign n37803 = ~n37800 & ~n37802 ;
  assign n37804 = ~\macstatus1_LoadRxStatus_reg/NET0131  & ~\wishbone_LatchedRxLength_reg[7]/NET0131  ;
  assign n37805 = n37803 & ~n37804 ;
  assign n37806 = ~n11680 & ~n11682 ;
  assign n37807 = ~n11722 & ~n11726 ;
  assign n37808 = ~\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  & ~n11665 ;
  assign n37809 = ~n11731 & ~n37808 ;
  assign n37810 = \txethmac1_TxRetry_reg/NET0131  & ~\wishbone_TxRetry_q_reg/NET0131  ;
  assign n37811 = \wishbone_TxStartFrm_reg/NET0131  & ~\wishbone_TxUsedData_q_reg/NET0131  ;
  assign n37812 = ~n37810 & n37811 ;
  assign n37813 = ~\wishbone_TxStartFrm_sync2_reg/NET0131  & ~n37812 ;
  assign n37814 = ~\wishbone_rx_fifo_read_pointer_reg[1]/NET0131  & ~n37768 ;
  assign n37815 = ~n33164 & ~n37341 ;
  assign n37816 = ~n37814 & n37815 ;
  assign n37817 = n23733 & n32819 ;
  assign n37818 = n32818 & n37817 ;
  assign n37819 = \wb_adr_i[4]_pad  & \wb_adr_i[5]_pad  ;
  assign n37820 = n37691 & n37819 ;
  assign n37821 = n37818 & n37820 ;
  assign n37822 = n37727 & n37817 ;
  assign n37823 = n37820 & n37822 ;
  assign n37824 = n35359 & n35361 ;
  assign n37825 = n13127 & n37824 ;
  assign n37826 = ~\wishbone_RxOverrun_reg/NET0131  & ~n37825 ;
  assign n37827 = ~n35450 & ~n37826 ;
  assign n37828 = n35298 & n35302 ;
  assign n37829 = n35301 & n37828 ;
  assign n37830 = ~\wishbone_TxUnderRun_wb_reg/NET0131  & ~n37829 ;
  assign n37831 = ~n35548 & ~n37830 ;
  assign n37832 = n25059 & n32820 ;
  assign n37833 = n25059 & n37430 ;
  assign n37834 = ~\ethreg1_MODER_0_DataOut_reg[5]/NET0131  & n37456 ;
  assign n37835 = n37459 & n37834 ;
  assign n37836 = n10564 & n37835 ;
  assign n37837 = n23747 & n23751 ;
  assign n37838 = n32820 & n37837 ;
  assign n37839 = ~\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  & ~n36265 ;
  assign n37840 = ~n37575 & ~n37839 ;
  assign n37841 = n36273 & n37840 ;
  assign n37842 = n32819 & n37727 ;
  assign n37843 = n37837 & n37842 ;
  assign n37844 = \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  & ~\maccontrol1_receivecontrol1_Divider2_reg/NET0131  ;
  assign n37845 = ~n11977 & n37844 ;
  assign n37846 = \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  & ~n33164 ;
  assign n37847 = ~n37341 & n37846 ;
  assign n37848 = ~\wishbone_rx_fifo_read_pointer_reg[2]/NET0131  & ~n33164 ;
  assign n37849 = n37341 & n37848 ;
  assign n37850 = ~n37847 & ~n37849 ;
  assign n37851 = ~\wb_adr_i[2]_pad  & ~\wb_adr_i[5]_pad  ;
  assign n37852 = n23793 & n37851 ;
  assign n37853 = n37818 & n37852 ;
  assign n37854 = \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  & n11983 ;
  assign n37855 = ~\maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131  & ~n37854 ;
  assign n37856 = ~wb_rst_i_pad & ~n11985 ;
  assign n37857 = ~n37855 & n37856 ;
  assign n37858 = ~\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  & ~n35517 ;
  assign n37859 = ~\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  & ~\txethmac1_TxUsedData_reg/NET0131  ;
  assign n37860 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  ;
  assign n37861 = ~n37859 & ~n37860 ;
  assign n37862 = ~n37858 & n37861 ;
  assign n37863 = n35538 & n37862 ;
  assign n37864 = n11203 & ~n11348 ;
  assign n37865 = \txethmac1_random1_RandomLatched_reg[5]/NET0131  & ~n36399 ;
  assign n37866 = \txethmac1_RetryCnt_reg[1]/NET0131  & \txethmac1_RetryCnt_reg[2]/NET0131  ;
  assign n37867 = ~\txethmac1_RetryCnt_reg[3]/NET0131  & ~n37866 ;
  assign n37868 = \txethmac1_random1_x_reg[5]/NET0131  & n36399 ;
  assign n37869 = ~n37867 & n37868 ;
  assign n37870 = ~n37865 & ~n37869 ;
  assign n37871 = ~\wb_adr_i[5]_pad  & n25057 ;
  assign n37872 = n23733 & n37871 ;
  assign n37873 = n37696 & n37872 ;
  assign n37874 = n11464 & n11588 ;
  assign n37875 = \wishbone_BDWrite_reg[3]/NET0131  & ~n36417 ;
  assign n37876 = \wishbone_BDWrite_reg[3]/NET0131  & ~\wishbone_TxEn_q_reg/NET0131  ;
  assign n37877 = ~n36414 & n37876 ;
  assign n37878 = ~n37875 & ~n37877 ;
  assign n37879 = ~\wb_adr_i[11]_pad  & \wb_sel_i[3]_pad  ;
  assign n37880 = n23726 & n37879 ;
  assign n37881 = ~n23725 & n37880 ;
  assign n37882 = n37718 & n37881 ;
  assign n37883 = n37878 & ~n37882 ;
  assign n37884 = \wishbone_BlockingTxBDRead_reg/NET0131  & ~\wishbone_TxBDReady_reg/NET0131  ;
  assign n37885 = ~\wishbone_BlockingTxBDRead_reg/NET0131  & \wishbone_TxBDReady_reg/NET0131  ;
  assign n37886 = ~n37884 & ~n37885 ;
  assign n37887 = ~\wishbone_BlockingTxBDRead_reg/NET0131  & ~\wishbone_TxRetryPacket_NotCleared_reg/NET0131  ;
  assign n37888 = ~n36304 & n37887 ;
  assign n37889 = n37886 & ~n37888 ;
  assign n37890 = ~\wishbone_TxStartFrm_syncb2_reg/NET0131  & \wishbone_TxStartFrm_wb_reg/NET0131  ;
  assign n37891 = ~\wishbone_StartOccured_reg/NET0131  & \wishbone_TxBDReady_reg/NET0131  ;
  assign n37892 = ~n37890 & ~n37891 ;
  assign n37893 = ~n35731 & ~n37890 ;
  assign n37894 = ~n36338 & n37893 ;
  assign n37895 = ~n37892 & ~n37894 ;
  assign n37896 = n32822 & n37819 ;
  assign n37897 = n37818 & n37896 ;
  assign n37898 = n37822 & n37896 ;
  assign n37899 = n23734 & n32821 ;
  assign n37900 = n37818 & n37899 ;
  assign n37901 = n37822 & n37899 ;
  assign n37902 = \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37903 = n36368 & n37902 ;
  assign n37904 = n36373 & n37903 ;
  assign n37905 = \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37906 = n35523 & n37905 ;
  assign n37907 = n36379 & n37906 ;
  assign n37908 = \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37909 = n36360 & n37908 ;
  assign n37910 = n36369 & n37909 ;
  assign n37911 = ~n37907 & ~n37910 ;
  assign n37912 = ~n37904 & n37911 ;
  assign n37913 = \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37914 = n36360 & n37913 ;
  assign n37915 = n36389 & n37914 ;
  assign n37916 = n36369 & n36380 ;
  assign n37917 = ~n37915 & ~n37916 ;
  assign n37918 = \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37919 = n36362 & n37918 ;
  assign n37920 = n36379 & n37919 ;
  assign n37921 = \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37922 = n35523 & n37921 ;
  assign n37923 = n35522 & n37922 ;
  assign n37924 = ~n37920 & ~n37923 ;
  assign n37925 = \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37926 = n35521 & n37925 ;
  assign n37927 = n36373 & n37926 ;
  assign n37928 = \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37929 = n36362 & n37928 ;
  assign n37930 = n36389 & n37929 ;
  assign n37931 = ~n37927 & ~n37930 ;
  assign n37932 = n37924 & n37931 ;
  assign n37933 = n37917 & n37932 ;
  assign n37934 = n37912 & n37933 ;
  assign n37935 = \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37936 = n36368 & n37935 ;
  assign n37937 = n36373 & n37936 ;
  assign n37938 = \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37939 = n35523 & n37938 ;
  assign n37940 = n36379 & n37939 ;
  assign n37941 = \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37942 = n36360 & n37941 ;
  assign n37943 = n36369 & n37942 ;
  assign n37944 = ~n37940 & ~n37943 ;
  assign n37945 = ~n37937 & n37944 ;
  assign n37946 = \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37947 = n36360 & n37946 ;
  assign n37948 = n36389 & n37947 ;
  assign n37949 = ~n37916 & ~n37948 ;
  assign n37950 = \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37951 = n36362 & n37950 ;
  assign n37952 = n36379 & n37951 ;
  assign n37953 = \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37954 = n35523 & n37953 ;
  assign n37955 = n35522 & n37954 ;
  assign n37956 = ~n37952 & ~n37955 ;
  assign n37957 = \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n37958 = n35521 & n37957 ;
  assign n37959 = n36373 & n37958 ;
  assign n37960 = \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n37961 = n36362 & n37960 ;
  assign n37962 = n36389 & n37961 ;
  assign n37963 = ~n37959 & ~n37962 ;
  assign n37964 = n37956 & n37963 ;
  assign n37965 = n37949 & n37964 ;
  assign n37966 = n37945 & n37965 ;
  assign n37967 = \txethmac1_RetryCnt_reg[3]/NET0131  & \txethmac1_random1_x_reg[6]/NET0131  ;
  assign n37968 = \txethmac1_RetryCnt_reg[2]/NET0131  & \txethmac1_random1_x_reg[6]/NET0131  ;
  assign n37969 = n11418 & n37968 ;
  assign n37970 = ~n37967 & ~n37969 ;
  assign n37971 = n36399 & n37970 ;
  assign n37972 = ~\txethmac1_random1_RandomLatched_reg[6]/NET0131  & ~n36399 ;
  assign n37973 = ~n37971 & ~n37972 ;
  assign n37974 = ~\wishbone_BlockingTxBDRead_reg/NET0131  & \wishbone_TxRetryPacket_NotCleared_reg/NET0131  ;
  assign n37975 = ~\wishbone_BlockingTxBDRead_reg/NET0131  & ~\wishbone_BlockingTxStatusWrite_reg/NET0131  ;
  assign n37976 = n36303 & n37975 ;
  assign n37977 = ~n37974 & ~n37976 ;
  assign n37978 = ~\wishbone_TxBDRead_reg/NET0131  & n37977 ;
  assign n37979 = ~\wishbone_TxBDReady_reg/NET0131  & ~n37978 ;
  assign n37980 = ~\wishbone_TxBDReady_reg/NET0131  & ~n37977 ;
  assign n37981 = ~\wishbone_TxRetryPacketBlocked_reg/NET0131  & \wishbone_TxRetry_wb_reg/NET0131  ;
  assign n37982 = ~\wishbone_TxRetryPacket_NotCleared_reg/NET0131  & ~n37981 ;
  assign n37983 = \wishbone_MasterWbTX_reg/NET0131  & ~\wishbone_TxRetryPacket_NotCleared_reg/NET0131  ;
  assign n37984 = ~n37751 & n37983 ;
  assign n37985 = ~n37982 & ~n37984 ;
  assign n37986 = ~n37980 & n37985 ;
  assign n37987 = \wishbone_TxByteCnt_reg[0]/NET0131  & ~\wishbone_TxValidBytesLatched_reg[0]/NET0131  ;
  assign n37988 = ~\wishbone_TxByteCnt_reg[0]/NET0131  & \wishbone_TxValidBytesLatched_reg[0]/NET0131  ;
  assign n37989 = ~n37987 & ~n37988 ;
  assign n37990 = \wishbone_LastWord_reg/NET0131  & ~\wishbone_TxEndFrm_reg/NET0131  ;
  assign n37991 = ~n37989 & n37990 ;
  assign n37992 = \wishbone_Flop_reg/NET0131  & ~n37991 ;
  assign n37993 = ~n12733 & ~n12736 ;
  assign n37994 = \wishbone_Flop_reg/NET0131  & ~\wishbone_TxValidBytesLatched_reg[1]/NET0131  ;
  assign n37995 = ~n37993 & n37994 ;
  assign n37996 = \wishbone_Flop_reg/NET0131  & \wishbone_TxValidBytesLatched_reg[1]/NET0131  ;
  assign n37997 = n37993 & n37996 ;
  assign n37998 = ~n37995 & ~n37997 ;
  assign n37999 = ~n37992 & n37998 ;
  assign n38000 = n37704 & ~n37705 ;
  assign n38001 = ~\wishbone_Flop_reg/NET0131  & ~\wishbone_TxEndFrm_reg/NET0131  ;
  assign n38002 = ~\wishbone_TxRetry_q_reg/NET0131  & ~n38001 ;
  assign n38003 = ~n38000 & n38002 ;
  assign n38004 = n37999 & n38003 ;
  assign n38005 = \wishbone_WbEn_q_reg/NET0131  & \wishbone_WbEn_reg/NET0131  ;
  assign n38006 = \wishbone_BDWrite_reg[1]/NET0131  & n38005 ;
  assign n38007 = ~n35450 & ~n38006 ;
  assign n38008 = ~n36304 & n38007 ;
  assign n38009 = ~\wishbone_ram_addr_reg[3]/NET0131  & ~\wishbone_ram_addr_reg[4]/NET0131  ;
  assign n38010 = \wishbone_ram_addr_reg[0]/NET0131  & \wishbone_ram_addr_reg[6]/NET0131  ;
  assign n38011 = n38009 & n38010 ;
  assign n38012 = \wishbone_ram_addr_reg[1]/NET0131  & ~\wishbone_ram_addr_reg[7]/NET0131  ;
  assign n38013 = ~\wishbone_ram_addr_reg[2]/NET0131  & \wishbone_ram_addr_reg[5]/NET0131  ;
  assign n38014 = n38012 & n38013 ;
  assign n38015 = n38011 & n38014 ;
  assign n38016 = ~n38008 & n38015 ;
  assign n38017 = \wishbone_BDWrite_reg[2]/NET0131  & n38005 ;
  assign n38018 = ~n35450 & ~n38017 ;
  assign n38019 = ~n36304 & n38018 ;
  assign n38020 = \wishbone_ram_addr_reg[2]/NET0131  & \wishbone_ram_addr_reg[5]/NET0131  ;
  assign n38021 = ~\wishbone_ram_addr_reg[1]/NET0131  & ~\wishbone_ram_addr_reg[7]/NET0131  ;
  assign n38022 = n38020 & n38021 ;
  assign n38023 = n38011 & n38022 ;
  assign n38024 = ~n38019 & n38023 ;
  assign n38025 = n38012 & n38020 ;
  assign n38026 = ~\wishbone_ram_addr_reg[0]/NET0131  & \wishbone_ram_addr_reg[6]/NET0131  ;
  assign n38027 = n38009 & n38026 ;
  assign n38028 = n38025 & n38027 ;
  assign n38029 = ~n38019 & n38028 ;
  assign n38030 = \wishbone_ram_addr_reg[3]/NET0131  & ~\wishbone_ram_addr_reg[4]/NET0131  ;
  assign n38031 = n38010 & n38030 ;
  assign n38032 = n38013 & n38021 ;
  assign n38033 = n38031 & n38032 ;
  assign n38034 = ~n38019 & n38033 ;
  assign n38035 = n38026 & n38030 ;
  assign n38036 = n38014 & n38035 ;
  assign n38037 = ~n38019 & n38036 ;
  assign n38038 = n38022 & n38035 ;
  assign n38039 = ~n38019 & n38038 ;
  assign n38040 = \wishbone_BDWrite_reg[0]/NET0131  & n38005 ;
  assign n38041 = ~n35450 & ~n38040 ;
  assign n38042 = ~n36304 & n38041 ;
  assign n38043 = ~\wishbone_ram_addr_reg[2]/NET0131  & ~\wishbone_ram_addr_reg[5]/NET0131  ;
  assign n38044 = n38012 & n38043 ;
  assign n38045 = \wishbone_ram_addr_reg[3]/NET0131  & \wishbone_ram_addr_reg[4]/NET0131  ;
  assign n38046 = n38010 & n38045 ;
  assign n38047 = n38044 & n38046 ;
  assign n38048 = ~n38042 & n38047 ;
  assign n38049 = ~\wishbone_ram_addr_reg[3]/NET0131  & \wishbone_ram_addr_reg[4]/NET0131  ;
  assign n38050 = n38010 & n38049 ;
  assign n38051 = n38032 & n38050 ;
  assign n38052 = ~n38019 & n38051 ;
  assign n38053 = n38026 & n38049 ;
  assign n38054 = n38014 & n38053 ;
  assign n38055 = ~n38019 & n38054 ;
  assign n38056 = n38022 & n38053 ;
  assign n38057 = ~n38019 & n38056 ;
  assign n38058 = n38026 & n38045 ;
  assign n38059 = n38032 & n38058 ;
  assign n38060 = ~n38019 & n38059 ;
  assign n38061 = n38032 & n38046 ;
  assign n38062 = ~n38019 & n38061 ;
  assign n38063 = \wishbone_ram_addr_reg[1]/NET0131  & \wishbone_ram_addr_reg[7]/NET0131  ;
  assign n38064 = \wishbone_ram_addr_reg[2]/NET0131  & ~\wishbone_ram_addr_reg[5]/NET0131  ;
  assign n38065 = n38063 & n38064 ;
  assign n38066 = ~\wishbone_ram_addr_reg[0]/NET0131  & ~\wishbone_ram_addr_reg[6]/NET0131  ;
  assign n38067 = n38009 & n38066 ;
  assign n38068 = n38065 & n38067 ;
  assign n38069 = ~n38019 & n38068 ;
  assign n38070 = \wishbone_ram_addr_reg[0]/NET0131  & ~\wishbone_ram_addr_reg[6]/NET0131  ;
  assign n38071 = n38009 & n38070 ;
  assign n38072 = n38065 & n38071 ;
  assign n38073 = ~n38019 & n38072 ;
  assign n38074 = n38043 & n38063 ;
  assign n38075 = n38030 & n38070 ;
  assign n38076 = n38074 & n38075 ;
  assign n38077 = ~n38019 & n38076 ;
  assign n38078 = ~\wishbone_ram_addr_reg[1]/NET0131  & \wishbone_ram_addr_reg[7]/NET0131  ;
  assign n38079 = n38064 & n38078 ;
  assign n38080 = n38075 & n38079 ;
  assign n38081 = ~n38019 & n38080 ;
  assign n38082 = n38030 & n38066 ;
  assign n38083 = n38065 & n38082 ;
  assign n38084 = ~n38019 & n38083 ;
  assign n38085 = n38049 & n38070 ;
  assign n38086 = n38074 & n38085 ;
  assign n38087 = ~n38019 & n38086 ;
  assign n38088 = n38079 & n38085 ;
  assign n38089 = ~n38019 & n38088 ;
  assign n38090 = n38049 & n38066 ;
  assign n38091 = n38065 & n38090 ;
  assign n38092 = ~n38019 & n38091 ;
  assign n38093 = ~n38008 & n38068 ;
  assign n38094 = n38043 & n38078 ;
  assign n38095 = n38045 & n38070 ;
  assign n38096 = n38094 & n38095 ;
  assign n38097 = ~n38019 & n38096 ;
  assign n38098 = n38045 & n38066 ;
  assign n38099 = n38074 & n38098 ;
  assign n38100 = ~n38019 & n38099 ;
  assign n38101 = n38079 & n38098 ;
  assign n38102 = ~n38019 & n38101 ;
  assign n38103 = n38012 & n38064 ;
  assign n38104 = n38075 & n38103 ;
  assign n38105 = ~n38019 & n38104 ;
  assign n38106 = n38013 & n38063 ;
  assign n38107 = n38067 & n38106 ;
  assign n38108 = ~n38019 & n38107 ;
  assign n38109 = n38071 & n38106 ;
  assign n38110 = ~n38019 & n38109 ;
  assign n38111 = n38020 & n38078 ;
  assign n38112 = n38067 & n38111 ;
  assign n38113 = ~n38019 & n38112 ;
  assign n38114 = n38071 & n38111 ;
  assign n38115 = ~n38019 & n38114 ;
  assign n38116 = n38020 & n38063 ;
  assign n38117 = n38067 & n38116 ;
  assign n38118 = ~n38019 & n38117 ;
  assign n38119 = n38071 & n38116 ;
  assign n38120 = ~n38019 & n38119 ;
  assign n38121 = n38013 & n38078 ;
  assign n38122 = n38075 & n38121 ;
  assign n38123 = ~n38019 & n38122 ;
  assign n38124 = n38082 & n38106 ;
  assign n38125 = ~n38019 & n38124 ;
  assign n38126 = n38082 & n38111 ;
  assign n38127 = ~n38019 & n38126 ;
  assign n38128 = n38082 & n38116 ;
  assign n38129 = ~n38019 & n38128 ;
  assign n38130 = n38085 & n38121 ;
  assign n38131 = ~n38019 & n38130 ;
  assign n38132 = n38090 & n38106 ;
  assign n38133 = ~n38019 & n38132 ;
  assign n38134 = n38090 & n38111 ;
  assign n38135 = ~n38019 & n38134 ;
  assign n38136 = n38090 & n38116 ;
  assign n38137 = ~n38019 & n38136 ;
  assign n38138 = n38098 & n38121 ;
  assign n38139 = ~n38019 & n38138 ;
  assign n38140 = n38011 & n38074 ;
  assign n38141 = ~n38019 & n38140 ;
  assign n38142 = n38011 & n38079 ;
  assign n38143 = ~n38019 & n38142 ;
  assign n38144 = n38027 & n38065 ;
  assign n38145 = ~n38019 & n38144 ;
  assign n38146 = n38031 & n38094 ;
  assign n38147 = ~n38019 & n38146 ;
  assign n38148 = n38035 & n38074 ;
  assign n38149 = ~n38019 & n38148 ;
  assign n38150 = n38035 & n38079 ;
  assign n38151 = ~n38019 & n38150 ;
  assign n38152 = n38050 & n38094 ;
  assign n38153 = ~n38019 & n38152 ;
  assign n38154 = n38053 & n38074 ;
  assign n38155 = ~n38019 & n38154 ;
  assign n38156 = n38053 & n38079 ;
  assign n38157 = ~n38019 & n38156 ;
  assign n38158 = n38058 & n38094 ;
  assign n38159 = ~n38019 & n38158 ;
  assign n38160 = n38046 & n38094 ;
  assign n38161 = ~n38019 & n38160 ;
  assign n38162 = ~n38008 & n38072 ;
  assign n38163 = n38011 & n38121 ;
  assign n38164 = ~n38019 & n38163 ;
  assign n38165 = n38027 & n38106 ;
  assign n38166 = ~n38019 & n38165 ;
  assign n38167 = n38023 & ~n38042 ;
  assign n38168 = n38027 & n38111 ;
  assign n38169 = ~n38019 & n38168 ;
  assign n38170 = n38028 & ~n38042 ;
  assign n38171 = n38027 & n38116 ;
  assign n38172 = ~n38019 & n38171 ;
  assign n38173 = n38035 & n38121 ;
  assign n38174 = ~n38019 & n38173 ;
  assign n38175 = n38033 & ~n38042 ;
  assign n38176 = n38036 & ~n38042 ;
  assign n38177 = n38085 & n38103 ;
  assign n38178 = ~n38019 & n38177 ;
  assign n38179 = n38038 & ~n38042 ;
  assign n38180 = n38053 & n38121 ;
  assign n38181 = ~n38019 & n38180 ;
  assign n38182 = ~n38042 & n38051 ;
  assign n38183 = n38021 & n38064 ;
  assign n38184 = n38031 & n38183 ;
  assign n38185 = ~n38042 & n38184 ;
  assign n38186 = ~n38042 & n38054 ;
  assign n38187 = n38021 & n38043 ;
  assign n38188 = n38095 & n38187 ;
  assign n38189 = ~n38019 & n38188 ;
  assign n38190 = ~n38042 & n38056 ;
  assign n38191 = n38044 & n38095 ;
  assign n38192 = ~n38019 & n38191 ;
  assign n38193 = n38095 & n38183 ;
  assign n38194 = ~n38019 & n38193 ;
  assign n38195 = n38098 & n38103 ;
  assign n38196 = ~n38019 & n38195 ;
  assign n38197 = ~n38042 & n38059 ;
  assign n38198 = ~n38042 & n38061 ;
  assign n38199 = n38025 & n38067 ;
  assign n38200 = ~n38019 & n38199 ;
  assign n38201 = n38025 & n38071 ;
  assign n38202 = ~n38019 & n38201 ;
  assign n38203 = n38014 & n38075 ;
  assign n38204 = ~n38019 & n38203 ;
  assign n38205 = n38022 & n38075 ;
  assign n38206 = ~n38019 & n38205 ;
  assign n38207 = n38025 & n38082 ;
  assign n38208 = ~n38019 & n38207 ;
  assign n38209 = n38014 & n38085 ;
  assign n38210 = ~n38019 & n38209 ;
  assign n38211 = n38022 & n38085 ;
  assign n38212 = ~n38019 & n38211 ;
  assign n38213 = n38025 & n38090 ;
  assign n38214 = ~n38019 & n38213 ;
  assign n38215 = n38032 & n38095 ;
  assign n38216 = ~n38019 & n38215 ;
  assign n38217 = n38014 & n38098 ;
  assign n38218 = ~n38019 & n38217 ;
  assign n38219 = n38022 & n38098 ;
  assign n38220 = ~n38019 & n38219 ;
  assign n38221 = ~n38042 & n38068 ;
  assign n38222 = ~n38042 & n38072 ;
  assign n38223 = n38011 & n38103 ;
  assign n38224 = ~n38019 & n38223 ;
  assign n38225 = ~n38042 & n38076 ;
  assign n38226 = n38031 & n38187 ;
  assign n38227 = ~n38019 & n38226 ;
  assign n38228 = n38031 & n38044 ;
  assign n38229 = ~n38019 & n38228 ;
  assign n38230 = ~n38019 & n38184 ;
  assign n38231 = n38035 & n38103 ;
  assign n38232 = ~n38019 & n38231 ;
  assign n38233 = ~n38042 & n38080 ;
  assign n38234 = ~n38042 & n38083 ;
  assign n38235 = n38050 & n38187 ;
  assign n38236 = ~n38019 & n38235 ;
  assign n38237 = n38044 & n38050 ;
  assign n38238 = ~n38019 & n38237 ;
  assign n38239 = n38050 & n38183 ;
  assign n38240 = ~n38019 & n38239 ;
  assign n38241 = n38053 & n38103 ;
  assign n38242 = ~n38019 & n38241 ;
  assign n38243 = n38058 & n38187 ;
  assign n38244 = ~n38019 & n38243 ;
  assign n38245 = n38046 & n38187 ;
  assign n38246 = ~n38019 & n38245 ;
  assign n38247 = ~n38042 & n38086 ;
  assign n38248 = n38044 & n38058 ;
  assign n38249 = ~n38019 & n38248 ;
  assign n38250 = ~n38019 & n38047 ;
  assign n38251 = n38058 & n38183 ;
  assign n38252 = ~n38019 & n38251 ;
  assign n38253 = ~n38042 & n38088 ;
  assign n38254 = n38046 & n38183 ;
  assign n38255 = ~n38019 & n38254 ;
  assign n38256 = ~n38042 & n38091 ;
  assign n38257 = n38015 & ~n38019 ;
  assign n38258 = ~n38042 & n38096 ;
  assign n38259 = \wishbone_BDWrite_reg[3]/NET0131  & n38005 ;
  assign n38260 = ~n35450 & ~n38259 ;
  assign n38261 = ~n36304 & n38260 ;
  assign n38262 = n38023 & ~n38261 ;
  assign n38263 = n38028 & ~n38261 ;
  assign n38264 = ~n38042 & n38099 ;
  assign n38265 = n38033 & ~n38261 ;
  assign n38266 = n38036 & ~n38261 ;
  assign n38267 = ~n38042 & n38101 ;
  assign n38268 = n38038 & ~n38261 ;
  assign n38269 = n38051 & ~n38261 ;
  assign n38270 = ~n38042 & n38104 ;
  assign n38271 = n38054 & ~n38261 ;
  assign n38272 = n38056 & ~n38261 ;
  assign n38273 = ~n38042 & n38107 ;
  assign n38274 = n38059 & ~n38261 ;
  assign n38275 = n38061 & ~n38261 ;
  assign n38276 = ~n38042 & n38109 ;
  assign n38277 = ~n38042 & n38112 ;
  assign n38278 = ~n38042 & n38114 ;
  assign n38279 = ~n38042 & n38117 ;
  assign n38280 = ~n38042 & n38119 ;
  assign n38281 = ~n38042 & n38122 ;
  assign n38282 = n38068 & ~n38261 ;
  assign n38283 = n38072 & ~n38261 ;
  assign n38284 = ~n38042 & n38124 ;
  assign n38285 = n38076 & ~n38261 ;
  assign n38286 = ~n38042 & n38126 ;
  assign n38287 = n38080 & ~n38261 ;
  assign n38288 = n38083 & ~n38261 ;
  assign n38289 = ~n38042 & n38128 ;
  assign n38290 = n38086 & ~n38261 ;
  assign n38291 = n38088 & ~n38261 ;
  assign n38292 = ~n38042 & n38130 ;
  assign n38293 = n38091 & ~n38261 ;
  assign n38294 = ~n38042 & n38132 ;
  assign n38295 = n38096 & ~n38261 ;
  assign n38296 = n38099 & ~n38261 ;
  assign n38297 = n38101 & ~n38261 ;
  assign n38298 = ~n38042 & n38134 ;
  assign n38299 = n38104 & ~n38261 ;
  assign n38300 = ~n38042 & n38136 ;
  assign n38301 = n38107 & ~n38261 ;
  assign n38302 = n38109 & ~n38261 ;
  assign n38303 = n38112 & ~n38261 ;
  assign n38304 = ~n38042 & n38138 ;
  assign n38305 = n38114 & ~n38261 ;
  assign n38306 = n38117 & ~n38261 ;
  assign n38307 = n38119 & ~n38261 ;
  assign n38308 = n38122 & ~n38261 ;
  assign n38309 = n38124 & ~n38261 ;
  assign n38310 = n38126 & ~n38261 ;
  assign n38311 = n38128 & ~n38261 ;
  assign n38312 = n38130 & ~n38261 ;
  assign n38313 = n38132 & ~n38261 ;
  assign n38314 = n38134 & ~n38261 ;
  assign n38315 = n38136 & ~n38261 ;
  assign n38316 = n38138 & ~n38261 ;
  assign n38317 = ~n38042 & n38140 ;
  assign n38318 = ~n38042 & n38142 ;
  assign n38319 = ~n38042 & n38144 ;
  assign n38320 = n38140 & ~n38261 ;
  assign n38321 = n38142 & ~n38261 ;
  assign n38322 = n38144 & ~n38261 ;
  assign n38323 = ~n38042 & n38146 ;
  assign n38324 = n38146 & ~n38261 ;
  assign n38325 = ~n38042 & n38148 ;
  assign n38326 = n38148 & ~n38261 ;
  assign n38327 = n38150 & ~n38261 ;
  assign n38328 = ~n38042 & n38150 ;
  assign n38329 = n38152 & ~n38261 ;
  assign n38330 = n38154 & ~n38261 ;
  assign n38331 = n38156 & ~n38261 ;
  assign n38332 = ~n38042 & n38152 ;
  assign n38333 = n38158 & ~n38261 ;
  assign n38334 = n38160 & ~n38261 ;
  assign n38335 = ~n38042 & n38154 ;
  assign n38336 = ~n38042 & n38156 ;
  assign n38337 = n38163 & ~n38261 ;
  assign n38338 = n38165 & ~n38261 ;
  assign n38339 = n38168 & ~n38261 ;
  assign n38340 = ~n38042 & n38158 ;
  assign n38341 = n38171 & ~n38261 ;
  assign n38342 = ~n38042 & n38160 ;
  assign n38343 = n38173 & ~n38261 ;
  assign n38344 = n38177 & ~n38261 ;
  assign n38345 = n38180 & ~n38261 ;
  assign n38346 = ~n38042 & n38163 ;
  assign n38347 = ~n38042 & n38165 ;
  assign n38348 = ~n38042 & n38168 ;
  assign n38349 = n38188 & ~n38261 ;
  assign n38350 = n38191 & ~n38261 ;
  assign n38351 = ~n38042 & n38171 ;
  assign n38352 = n38193 & ~n38261 ;
  assign n38353 = n38195 & ~n38261 ;
  assign n38354 = ~n38042 & n38173 ;
  assign n38355 = n38199 & ~n38261 ;
  assign n38356 = n38201 & ~n38261 ;
  assign n38357 = n38203 & ~n38261 ;
  assign n38358 = n38205 & ~n38261 ;
  assign n38359 = n38207 & ~n38261 ;
  assign n38360 = ~n38042 & n38177 ;
  assign n38361 = ~n38042 & n38180 ;
  assign n38362 = n38209 & ~n38261 ;
  assign n38363 = n38211 & ~n38261 ;
  assign n38364 = n38213 & ~n38261 ;
  assign n38365 = n38215 & ~n38261 ;
  assign n38366 = n38217 & ~n38261 ;
  assign n38367 = n38219 & ~n38261 ;
  assign n38368 = n38223 & ~n38261 ;
  assign n38369 = n38226 & ~n38261 ;
  assign n38370 = n38228 & ~n38261 ;
  assign n38371 = n38184 & ~n38261 ;
  assign n38372 = n38231 & ~n38261 ;
  assign n38373 = ~n38042 & n38188 ;
  assign n38374 = n38235 & ~n38261 ;
  assign n38375 = n38237 & ~n38261 ;
  assign n38376 = ~n38042 & n38191 ;
  assign n38377 = n38239 & ~n38261 ;
  assign n38378 = n38241 & ~n38261 ;
  assign n38379 = n38243 & ~n38261 ;
  assign n38380 = ~n38042 & n38193 ;
  assign n38381 = n38245 & ~n38261 ;
  assign n38382 = n38248 & ~n38261 ;
  assign n38383 = n38047 & ~n38261 ;
  assign n38384 = ~n38042 & n38195 ;
  assign n38385 = n38251 & ~n38261 ;
  assign n38386 = n38254 & ~n38261 ;
  assign n38387 = n38015 & ~n38261 ;
  assign n38388 = ~n38042 & n38199 ;
  assign n38389 = ~n38042 & n38201 ;
  assign n38390 = ~n38042 & n38239 ;
  assign n38391 = ~n38042 & n38203 ;
  assign n38392 = ~n38042 & n38205 ;
  assign n38393 = ~n38042 & n38207 ;
  assign n38394 = ~n38008 & n38061 ;
  assign n38395 = ~n38042 & n38209 ;
  assign n38396 = ~n38042 & n38211 ;
  assign n38397 = ~n38042 & n38213 ;
  assign n38398 = ~n38042 & n38215 ;
  assign n38399 = ~n38042 & n38217 ;
  assign n38400 = ~n38042 & n38219 ;
  assign n38401 = ~n38042 & n38223 ;
  assign n38402 = ~n38042 & n38226 ;
  assign n38403 = ~n38042 & n38251 ;
  assign n38404 = ~n38042 & n38228 ;
  assign n38405 = ~n38042 & n38231 ;
  assign n38406 = ~n38042 & n38235 ;
  assign n38407 = ~n38042 & n38237 ;
  assign n38408 = ~n38042 & n38241 ;
  assign n38409 = ~n38042 & n38243 ;
  assign n38410 = ~n38042 & n38245 ;
  assign n38411 = ~n38042 & n38248 ;
  assign n38412 = ~n38042 & n38254 ;
  assign n38413 = n38015 & ~n38042 ;
  assign n38414 = ~n38008 & n38023 ;
  assign n38415 = ~n38008 & n38028 ;
  assign n38416 = ~n38008 & n38033 ;
  assign n38417 = ~n38008 & n38036 ;
  assign n38418 = ~n38008 & n38038 ;
  assign n38419 = ~n38008 & n38059 ;
  assign n38420 = ~n38008 & n38051 ;
  assign n38421 = ~n38008 & n38054 ;
  assign n38422 = ~n38008 & n38056 ;
  assign n38423 = ~n38008 & n38076 ;
  assign n38424 = ~n38008 & n38080 ;
  assign n38425 = ~n38008 & n38083 ;
  assign n38426 = ~n38008 & n38086 ;
  assign n38427 = ~n38008 & n38088 ;
  assign n38428 = ~n38008 & n38091 ;
  assign n38429 = ~n38008 & n38096 ;
  assign n38430 = ~n38008 & n38099 ;
  assign n38431 = ~n38008 & n38101 ;
  assign n38432 = ~n38008 & n38104 ;
  assign n38433 = ~n38008 & n38107 ;
  assign n38434 = ~n38008 & n38109 ;
  assign n38435 = ~n38008 & n38112 ;
  assign n38436 = ~n38008 & n38114 ;
  assign n38437 = ~n38008 & n38117 ;
  assign n38438 = ~n38008 & n38119 ;
  assign n38439 = ~n38008 & n38122 ;
  assign n38440 = ~n38008 & n38124 ;
  assign n38441 = ~n38008 & n38126 ;
  assign n38442 = ~n38008 & n38128 ;
  assign n38443 = ~n38008 & n38130 ;
  assign n38444 = ~n38008 & n38132 ;
  assign n38445 = ~n38008 & n38134 ;
  assign n38446 = ~n38008 & n38136 ;
  assign n38447 = ~n38008 & n38138 ;
  assign n38448 = ~n38008 & n38140 ;
  assign n38449 = ~n38008 & n38142 ;
  assign n38450 = ~n38008 & n38144 ;
  assign n38451 = ~n38008 & n38146 ;
  assign n38452 = ~n38008 & n38148 ;
  assign n38453 = ~n38008 & n38150 ;
  assign n38454 = ~n38008 & n38152 ;
  assign n38455 = ~n38008 & n38154 ;
  assign n38456 = ~n38008 & n38156 ;
  assign n38457 = ~n38008 & n38158 ;
  assign n38458 = ~n38008 & n38160 ;
  assign n38459 = ~n38008 & n38163 ;
  assign n38460 = ~n38008 & n38165 ;
  assign n38461 = ~n38008 & n38168 ;
  assign n38462 = ~n38008 & n38171 ;
  assign n38463 = ~n38008 & n38173 ;
  assign n38464 = ~n38008 & n38177 ;
  assign n38465 = ~n38008 & n38180 ;
  assign n38466 = ~n38008 & n38188 ;
  assign n38467 = ~n38008 & n38191 ;
  assign n38468 = ~n38008 & n38193 ;
  assign n38469 = ~n38008 & n38195 ;
  assign n38470 = ~n38008 & n38199 ;
  assign n38471 = ~n38008 & n38201 ;
  assign n38472 = ~n38008 & n38203 ;
  assign n38473 = ~n38008 & n38205 ;
  assign n38474 = ~n38008 & n38207 ;
  assign n38475 = ~n38008 & n38209 ;
  assign n38476 = ~n38008 & n38211 ;
  assign n38477 = ~n38008 & n38213 ;
  assign n38478 = ~n38008 & n38215 ;
  assign n38479 = ~n38008 & n38217 ;
  assign n38480 = ~n38008 & n38219 ;
  assign n38481 = ~n38008 & n38223 ;
  assign n38482 = ~n38008 & n38226 ;
  assign n38483 = ~n38008 & n38228 ;
  assign n38484 = ~n38008 & n38184 ;
  assign n38485 = ~n38008 & n38231 ;
  assign n38486 = ~n38008 & n38235 ;
  assign n38487 = ~n38008 & n38237 ;
  assign n38488 = ~n38008 & n38239 ;
  assign n38489 = ~n38008 & n38241 ;
  assign n38490 = ~n38008 & n38243 ;
  assign n38491 = ~n38008 & n38245 ;
  assign n38492 = ~n38008 & n38248 ;
  assign n38493 = ~n38008 & n38047 ;
  assign n38494 = ~n38008 & n38251 ;
  assign n38495 = ~n38008 & n38254 ;
  assign n38496 = n38075 & n38187 ;
  assign n38497 = ~n38008 & n38496 ;
  assign n38498 = n38014 & n38050 ;
  assign n38499 = ~n38008 & n38498 ;
  assign n38500 = n38067 & n38187 ;
  assign n38501 = ~n38019 & n38500 ;
  assign n38502 = n38022 & n38027 ;
  assign n38503 = ~n38019 & n38502 ;
  assign n38504 = n38011 & n38025 ;
  assign n38505 = ~n38019 & n38504 ;
  assign n38506 = n38032 & n38035 ;
  assign n38507 = ~n38019 & n38506 ;
  assign n38508 = n38014 & n38031 ;
  assign n38509 = ~n38019 & n38508 ;
  assign n38510 = n38022 & n38031 ;
  assign n38511 = ~n38019 & n38510 ;
  assign n38512 = n38044 & n38082 ;
  assign n38513 = ~n38019 & n38512 ;
  assign n38514 = n38025 & n38035 ;
  assign n38515 = ~n38019 & n38514 ;
  assign n38516 = n38025 & n38031 ;
  assign n38517 = ~n38019 & n38516 ;
  assign n38518 = n38032 & n38053 ;
  assign n38519 = ~n38019 & n38518 ;
  assign n38520 = ~n38019 & n38498 ;
  assign n38521 = n38022 & n38050 ;
  assign n38522 = ~n38019 & n38521 ;
  assign n38523 = n38025 & n38053 ;
  assign n38524 = ~n38019 & n38523 ;
  assign n38525 = n38022 & n38082 ;
  assign n38526 = ~n38042 & n38525 ;
  assign n38527 = n38025 & n38050 ;
  assign n38528 = ~n38019 & n38527 ;
  assign n38529 = n38044 & n38075 ;
  assign n38530 = ~n38019 & n38529 ;
  assign n38531 = n38014 & n38058 ;
  assign n38532 = ~n38019 & n38531 ;
  assign n38533 = n38014 & n38046 ;
  assign n38534 = ~n38019 & n38533 ;
  assign n38535 = n38022 & n38058 ;
  assign n38536 = ~n38019 & n38535 ;
  assign n38537 = n38022 & n38046 ;
  assign n38538 = ~n38019 & n38537 ;
  assign n38539 = n38025 & n38058 ;
  assign n38540 = ~n38019 & n38539 ;
  assign n38541 = n38025 & n38046 ;
  assign n38542 = ~n38019 & n38541 ;
  assign n38543 = n38067 & n38094 ;
  assign n38544 = ~n38019 & n38543 ;
  assign n38545 = n38071 & n38094 ;
  assign n38546 = ~n38019 & n38545 ;
  assign n38547 = n38082 & n38183 ;
  assign n38548 = ~n38019 & n38547 ;
  assign n38549 = n38067 & n38074 ;
  assign n38550 = ~n38019 & n38549 ;
  assign n38551 = n38071 & n38074 ;
  assign n38552 = ~n38019 & n38551 ;
  assign n38553 = n38067 & n38079 ;
  assign n38554 = ~n38019 & n38553 ;
  assign n38555 = n38071 & n38079 ;
  assign n38556 = ~n38019 & n38555 ;
  assign n38557 = n38082 & n38094 ;
  assign n38558 = ~n38019 & n38557 ;
  assign n38559 = n38075 & n38094 ;
  assign n38560 = ~n38019 & n38559 ;
  assign n38561 = n38074 & n38082 ;
  assign n38562 = ~n38019 & n38561 ;
  assign n38563 = n38075 & n38183 ;
  assign n38564 = ~n38019 & n38563 ;
  assign n38565 = n38079 & n38082 ;
  assign n38566 = ~n38019 & n38565 ;
  assign n38567 = n38065 & n38075 ;
  assign n38568 = ~n38019 & n38567 ;
  assign n38569 = n38090 & n38094 ;
  assign n38570 = ~n38019 & n38569 ;
  assign n38571 = ~n38008 & n38545 ;
  assign n38572 = ~n38008 & n38555 ;
  assign n38573 = n38085 & n38094 ;
  assign n38574 = ~n38019 & n38573 ;
  assign n38575 = n38074 & n38090 ;
  assign n38576 = ~n38019 & n38575 ;
  assign n38577 = ~n38008 & n38541 ;
  assign n38578 = n38079 & n38090 ;
  assign n38579 = ~n38019 & n38578 ;
  assign n38580 = n38082 & n38103 ;
  assign n38581 = ~n38019 & n38580 ;
  assign n38582 = ~n38008 & n38557 ;
  assign n38583 = n38065 & n38085 ;
  assign n38584 = ~n38019 & n38583 ;
  assign n38585 = n38094 & n38098 ;
  assign n38586 = ~n38019 & n38585 ;
  assign n38587 = n38074 & n38095 ;
  assign n38588 = ~n38019 & n38587 ;
  assign n38589 = n38079 & n38095 ;
  assign n38590 = ~n38019 & n38589 ;
  assign n38591 = n38065 & n38098 ;
  assign n38592 = ~n38019 & n38591 ;
  assign n38593 = ~n38008 & n38549 ;
  assign n38594 = n38065 & n38095 ;
  assign n38595 = ~n38019 & n38594 ;
  assign n38596 = n38067 & n38121 ;
  assign n38597 = ~n38019 & n38596 ;
  assign n38598 = n38071 & n38121 ;
  assign n38599 = ~n38019 & n38598 ;
  assign n38600 = ~n38008 & n38547 ;
  assign n38601 = ~n38008 & n38563 ;
  assign n38602 = n38082 & n38121 ;
  assign n38603 = ~n38019 & n38602 ;
  assign n38604 = n38090 & n38187 ;
  assign n38605 = ~n38019 & n38604 ;
  assign n38606 = n38075 & n38106 ;
  assign n38607 = ~n38019 & n38606 ;
  assign n38608 = n38075 & n38111 ;
  assign n38609 = ~n38019 & n38608 ;
  assign n38610 = ~n38008 & n38561 ;
  assign n38611 = n38075 & n38116 ;
  assign n38612 = ~n38019 & n38611 ;
  assign n38613 = n38090 & n38121 ;
  assign n38614 = ~n38019 & n38613 ;
  assign n38615 = ~n38008 & n38553 ;
  assign n38616 = n38085 & n38106 ;
  assign n38617 = ~n38019 & n38616 ;
  assign n38618 = n38085 & n38187 ;
  assign n38619 = ~n38019 & n38618 ;
  assign n38620 = ~n38008 & n38539 ;
  assign n38621 = n38027 & n38187 ;
  assign n38622 = ~n38042 & n38621 ;
  assign n38623 = n38085 & n38111 ;
  assign n38624 = ~n38019 & n38623 ;
  assign n38625 = n38085 & n38116 ;
  assign n38626 = ~n38019 & n38625 ;
  assign n38627 = n38095 & n38121 ;
  assign n38628 = ~n38019 & n38627 ;
  assign n38629 = n38098 & n38106 ;
  assign n38630 = ~n38019 & n38629 ;
  assign n38631 = n38095 & n38106 ;
  assign n38632 = ~n38019 & n38631 ;
  assign n38633 = n38098 & n38111 ;
  assign n38634 = ~n38019 & n38633 ;
  assign n38635 = n38095 & n38111 ;
  assign n38636 = ~n38019 & n38635 ;
  assign n38637 = ~n38008 & n38502 ;
  assign n38638 = n38044 & n38090 ;
  assign n38639 = ~n38019 & n38638 ;
  assign n38640 = n38098 & n38116 ;
  assign n38641 = ~n38019 & n38640 ;
  assign n38642 = n38095 & n38116 ;
  assign n38643 = ~n38019 & n38642 ;
  assign n38644 = n38027 & n38094 ;
  assign n38645 = ~n38019 & n38644 ;
  assign n38646 = n38011 & n38094 ;
  assign n38647 = ~n38019 & n38646 ;
  assign n38648 = n38027 & n38074 ;
  assign n38649 = ~n38019 & n38648 ;
  assign n38650 = n38027 & n38079 ;
  assign n38651 = ~n38019 & n38650 ;
  assign n38652 = n38011 & n38065 ;
  assign n38653 = ~n38019 & n38652 ;
  assign n38654 = n38044 & n38085 ;
  assign n38655 = ~n38019 & n38654 ;
  assign n38656 = n38071 & n38187 ;
  assign n38657 = ~n38019 & n38656 ;
  assign n38658 = n38035 & n38094 ;
  assign n38659 = ~n38019 & n38658 ;
  assign n38660 = ~n38008 & n38537 ;
  assign n38661 = n38031 & n38074 ;
  assign n38662 = ~n38019 & n38661 ;
  assign n38663 = n38031 & n38079 ;
  assign n38664 = ~n38019 & n38663 ;
  assign n38665 = n38035 & n38065 ;
  assign n38666 = ~n38019 & n38665 ;
  assign n38667 = n38031 & n38065 ;
  assign n38668 = ~n38019 & n38667 ;
  assign n38669 = n38053 & n38094 ;
  assign n38670 = ~n38019 & n38669 ;
  assign n38671 = n38090 & n38183 ;
  assign n38672 = ~n38019 & n38671 ;
  assign n38673 = n38050 & n38074 ;
  assign n38674 = ~n38019 & n38673 ;
  assign n38675 = n38050 & n38079 ;
  assign n38676 = ~n38019 & n38675 ;
  assign n38677 = n38053 & n38065 ;
  assign n38678 = ~n38019 & n38677 ;
  assign n38679 = n38050 & n38065 ;
  assign n38680 = ~n38019 & n38679 ;
  assign n38681 = n38044 & n38053 ;
  assign n38682 = ~n38042 & n38681 ;
  assign n38683 = n38058 & n38074 ;
  assign n38684 = ~n38019 & n38683 ;
  assign n38685 = n38046 & n38074 ;
  assign n38686 = ~n38019 & n38685 ;
  assign n38687 = n38085 & n38183 ;
  assign n38688 = ~n38019 & n38687 ;
  assign n38689 = n38058 & n38079 ;
  assign n38690 = ~n38019 & n38689 ;
  assign n38691 = n38046 & n38079 ;
  assign n38692 = ~n38019 & n38691 ;
  assign n38693 = ~n38042 & n38500 ;
  assign n38694 = n38058 & n38065 ;
  assign n38695 = ~n38019 & n38694 ;
  assign n38696 = n38046 & n38065 ;
  assign n38697 = ~n38019 & n38696 ;
  assign n38698 = n38027 & n38121 ;
  assign n38699 = ~n38019 & n38698 ;
  assign n38700 = ~n38042 & n38502 ;
  assign n38701 = n38011 & n38106 ;
  assign n38702 = ~n38019 & n38701 ;
  assign n38703 = n38011 & n38111 ;
  assign n38704 = ~n38019 & n38703 ;
  assign n38705 = n38090 & n38103 ;
  assign n38706 = ~n38019 & n38705 ;
  assign n38707 = ~n38042 & n38504 ;
  assign n38708 = n38011 & n38116 ;
  assign n38709 = ~n38019 & n38708 ;
  assign n38710 = ~n38042 & n38506 ;
  assign n38711 = n38031 & n38121 ;
  assign n38712 = ~n38019 & n38711 ;
  assign n38713 = n38035 & n38106 ;
  assign n38714 = ~n38019 & n38713 ;
  assign n38715 = n38031 & n38106 ;
  assign n38716 = ~n38019 & n38715 ;
  assign n38717 = n38035 & n38111 ;
  assign n38718 = ~n38019 & n38717 ;
  assign n38719 = n38031 & n38111 ;
  assign n38720 = ~n38019 & n38719 ;
  assign n38721 = n38035 & n38116 ;
  assign n38722 = ~n38019 & n38721 ;
  assign n38723 = ~n38042 & n38508 ;
  assign n38724 = n38031 & n38116 ;
  assign n38725 = ~n38019 & n38724 ;
  assign n38726 = n38071 & n38103 ;
  assign n38727 = ~n38042 & n38726 ;
  assign n38728 = n38050 & n38121 ;
  assign n38729 = ~n38019 & n38728 ;
  assign n38730 = ~n38042 & n38510 ;
  assign n38731 = n38053 & n38106 ;
  assign n38732 = ~n38019 & n38731 ;
  assign n38733 = n38050 & n38106 ;
  assign n38734 = ~n38019 & n38733 ;
  assign n38735 = ~n38042 & n38512 ;
  assign n38736 = n38053 & n38111 ;
  assign n38737 = ~n38019 & n38736 ;
  assign n38738 = n38050 & n38111 ;
  assign n38739 = ~n38019 & n38738 ;
  assign n38740 = ~n38042 & n38514 ;
  assign n38741 = n38053 & n38116 ;
  assign n38742 = ~n38019 & n38741 ;
  assign n38743 = n38050 & n38116 ;
  assign n38744 = ~n38019 & n38743 ;
  assign n38745 = ~n38042 & n38516 ;
  assign n38746 = n38058 & n38121 ;
  assign n38747 = ~n38019 & n38746 ;
  assign n38748 = n38046 & n38121 ;
  assign n38749 = ~n38019 & n38748 ;
  assign n38750 = ~n38042 & n38518 ;
  assign n38751 = n38098 & n38187 ;
  assign n38752 = ~n38019 & n38751 ;
  assign n38753 = n38058 & n38106 ;
  assign n38754 = ~n38019 & n38753 ;
  assign n38755 = n38046 & n38106 ;
  assign n38756 = ~n38019 & n38755 ;
  assign n38757 = n38058 & n38111 ;
  assign n38758 = ~n38019 & n38757 ;
  assign n38759 = n38046 & n38111 ;
  assign n38760 = ~n38019 & n38759 ;
  assign n38761 = ~n38008 & n38535 ;
  assign n38762 = n38058 & n38116 ;
  assign n38763 = ~n38019 & n38762 ;
  assign n38764 = ~n38042 & n38498 ;
  assign n38765 = n38046 & n38116 ;
  assign n38766 = ~n38019 & n38765 ;
  assign n38767 = n38044 & n38098 ;
  assign n38768 = ~n38019 & n38767 ;
  assign n38769 = ~n38042 & n38521 ;
  assign n38770 = n38098 & n38183 ;
  assign n38771 = ~n38019 & n38770 ;
  assign n38772 = n38044 & n38067 ;
  assign n38773 = ~n38019 & n38772 ;
  assign n38774 = ~n38042 & n38523 ;
  assign n38775 = ~n38042 & n38527 ;
  assign n38776 = n38095 & n38103 ;
  assign n38777 = ~n38019 & n38776 ;
  assign n38778 = n38032 & n38067 ;
  assign n38779 = ~n38019 & n38778 ;
  assign n38780 = ~n38042 & n38529 ;
  assign n38781 = n38032 & n38071 ;
  assign n38782 = ~n38019 & n38781 ;
  assign n38783 = n38014 & n38067 ;
  assign n38784 = ~n38019 & n38783 ;
  assign n38785 = n38014 & n38071 ;
  assign n38786 = ~n38019 & n38785 ;
  assign n38787 = n38022 & n38067 ;
  assign n38788 = ~n38019 & n38787 ;
  assign n38789 = n38022 & n38071 ;
  assign n38790 = ~n38019 & n38789 ;
  assign n38791 = ~n38042 & n38531 ;
  assign n38792 = n38044 & n38071 ;
  assign n38793 = ~n38019 & n38792 ;
  assign n38794 = n38032 & n38082 ;
  assign n38795 = ~n38019 & n38794 ;
  assign n38796 = ~n38042 & n38533 ;
  assign n38797 = n38032 & n38075 ;
  assign n38798 = ~n38019 & n38797 ;
  assign n38799 = n38014 & n38082 ;
  assign n38800 = ~n38019 & n38799 ;
  assign n38801 = ~n38042 & n38535 ;
  assign n38802 = ~n38019 & n38525 ;
  assign n38803 = ~n38042 & n38537 ;
  assign n38804 = ~n38042 & n38539 ;
  assign n38805 = n38025 & n38075 ;
  assign n38806 = ~n38019 & n38805 ;
  assign n38807 = n38032 & n38090 ;
  assign n38808 = ~n38019 & n38807 ;
  assign n38809 = ~n38042 & n38541 ;
  assign n38810 = n38032 & n38085 ;
  assign n38811 = ~n38019 & n38810 ;
  assign n38812 = n38067 & n38183 ;
  assign n38813 = ~n38019 & n38812 ;
  assign n38814 = ~n38042 & n38543 ;
  assign n38815 = n38014 & n38090 ;
  assign n38816 = ~n38019 & n38815 ;
  assign n38817 = ~n38042 & n38545 ;
  assign n38818 = n38022 & n38090 ;
  assign n38819 = ~n38019 & n38818 ;
  assign n38820 = ~n38042 & n38547 ;
  assign n38821 = n38025 & n38085 ;
  assign n38822 = ~n38019 & n38821 ;
  assign n38823 = ~n38042 & n38549 ;
  assign n38824 = n38032 & n38098 ;
  assign n38825 = ~n38019 & n38824 ;
  assign n38826 = ~n38042 & n38551 ;
  assign n38827 = n38014 & n38095 ;
  assign n38828 = ~n38019 & n38827 ;
  assign n38829 = ~n38042 & n38553 ;
  assign n38830 = n38071 & n38183 ;
  assign n38831 = ~n38019 & n38830 ;
  assign n38832 = ~n38042 & n38555 ;
  assign n38833 = n38022 & n38095 ;
  assign n38834 = ~n38019 & n38833 ;
  assign n38835 = n38025 & n38098 ;
  assign n38836 = ~n38019 & n38835 ;
  assign n38837 = n38025 & n38095 ;
  assign n38838 = ~n38019 & n38837 ;
  assign n38839 = ~n38019 & n38621 ;
  assign n38840 = n38011 & n38187 ;
  assign n38841 = ~n38019 & n38840 ;
  assign n38842 = ~n38042 & n38833 ;
  assign n38843 = n38027 & n38044 ;
  assign n38844 = ~n38019 & n38843 ;
  assign n38845 = n38011 & n38044 ;
  assign n38846 = ~n38019 & n38845 ;
  assign n38847 = ~n38042 & n38557 ;
  assign n38848 = n38027 & n38183 ;
  assign n38849 = ~n38019 & n38848 ;
  assign n38850 = n38011 & n38183 ;
  assign n38851 = ~n38019 & n38850 ;
  assign n38852 = ~n38042 & n38559 ;
  assign n38853 = n38067 & n38103 ;
  assign n38854 = ~n38019 & n38853 ;
  assign n38855 = n38027 & n38103 ;
  assign n38856 = ~n38019 & n38855 ;
  assign n38857 = ~n38042 & n38561 ;
  assign n38858 = n38035 & n38187 ;
  assign n38859 = ~n38019 & n38858 ;
  assign n38860 = n38035 & n38044 ;
  assign n38861 = ~n38019 & n38860 ;
  assign n38862 = ~n38042 & n38563 ;
  assign n38863 = n38035 & n38183 ;
  assign n38864 = ~n38019 & n38863 ;
  assign n38865 = ~n38042 & n38565 ;
  assign n38866 = n38031 & n38103 ;
  assign n38867 = ~n38019 & n38866 ;
  assign n38868 = ~n38019 & n38726 ;
  assign n38869 = n38053 & n38187 ;
  assign n38870 = ~n38019 & n38869 ;
  assign n38871 = ~n38042 & n38567 ;
  assign n38872 = ~n38019 & n38681 ;
  assign n38873 = ~n38042 & n38569 ;
  assign n38874 = n38053 & n38183 ;
  assign n38875 = ~n38019 & n38874 ;
  assign n38876 = n38046 & n38103 ;
  assign n38877 = ~n38261 & n38876 ;
  assign n38878 = ~n38042 & n38573 ;
  assign n38879 = n38050 & n38103 ;
  assign n38880 = ~n38019 & n38879 ;
  assign n38881 = ~n38042 & n38575 ;
  assign n38882 = n38082 & n38187 ;
  assign n38883 = ~n38019 & n38882 ;
  assign n38884 = ~n38042 & n38578 ;
  assign n38885 = n38058 & n38103 ;
  assign n38886 = ~n38019 & n38885 ;
  assign n38887 = ~n38042 & n38580 ;
  assign n38888 = ~n38019 & n38876 ;
  assign n38889 = ~n38261 & n38885 ;
  assign n38890 = n38027 & n38032 ;
  assign n38891 = ~n38019 & n38890 ;
  assign n38892 = n38011 & n38032 ;
  assign n38893 = ~n38019 & n38892 ;
  assign n38894 = n38014 & n38027 ;
  assign n38895 = ~n38019 & n38894 ;
  assign n38896 = ~n38042 & n38583 ;
  assign n38897 = ~n38019 & n38496 ;
  assign n38898 = ~n38042 & n38585 ;
  assign n38899 = ~n38261 & n38500 ;
  assign n38900 = ~n38261 & n38502 ;
  assign n38901 = ~n38042 & n38830 ;
  assign n38902 = ~n38261 & n38504 ;
  assign n38903 = ~n38008 & n38543 ;
  assign n38904 = ~n38261 & n38506 ;
  assign n38905 = ~n38042 & n38587 ;
  assign n38906 = ~n38261 & n38508 ;
  assign n38907 = ~n38042 & n38589 ;
  assign n38908 = ~n38261 & n38510 ;
  assign n38909 = ~n38261 & n38512 ;
  assign n38910 = ~n38042 & n38591 ;
  assign n38911 = ~n38261 & n38514 ;
  assign n38912 = ~n38261 & n38516 ;
  assign n38913 = ~n38042 & n38594 ;
  assign n38914 = ~n38261 & n38518 ;
  assign n38915 = ~n38261 & n38498 ;
  assign n38916 = ~n38042 & n38596 ;
  assign n38917 = ~n38261 & n38521 ;
  assign n38918 = ~n38261 & n38523 ;
  assign n38919 = ~n38042 & n38598 ;
  assign n38920 = ~n38261 & n38527 ;
  assign n38921 = ~n38261 & n38529 ;
  assign n38922 = ~n38261 & n38531 ;
  assign n38923 = ~n38261 & n38533 ;
  assign n38924 = ~n38261 & n38535 ;
  assign n38925 = ~n38261 & n38537 ;
  assign n38926 = ~n38261 & n38539 ;
  assign n38927 = ~n38261 & n38541 ;
  assign n38928 = ~n38261 & n38543 ;
  assign n38929 = ~n38261 & n38545 ;
  assign n38930 = ~n38261 & n38547 ;
  assign n38931 = ~n38261 & n38549 ;
  assign n38932 = ~n38042 & n38602 ;
  assign n38933 = ~n38261 & n38551 ;
  assign n38934 = ~n38261 & n38553 ;
  assign n38935 = ~n38261 & n38555 ;
  assign n38936 = ~n38042 & n38604 ;
  assign n38937 = ~n38261 & n38557 ;
  assign n38938 = ~n38261 & n38559 ;
  assign n38939 = ~n38261 & n38561 ;
  assign n38940 = ~n38042 & n38827 ;
  assign n38941 = ~n38042 & n38606 ;
  assign n38942 = ~n38008 & n38518 ;
  assign n38943 = ~n38261 & n38563 ;
  assign n38944 = ~n38261 & n38565 ;
  assign n38945 = ~n38042 & n38608 ;
  assign n38946 = ~n38261 & n38567 ;
  assign n38947 = ~n38261 & n38569 ;
  assign n38948 = ~n38261 & n38573 ;
  assign n38949 = ~n38042 & n38611 ;
  assign n38950 = ~n38261 & n38575 ;
  assign n38951 = ~n38042 & n38613 ;
  assign n38952 = ~n38261 & n38578 ;
  assign n38953 = ~n38261 & n38580 ;
  assign n38954 = ~n38261 & n38583 ;
  assign n38955 = ~n38261 & n38585 ;
  assign n38956 = ~n38042 & n38616 ;
  assign n38957 = ~n38042 & n38618 ;
  assign n38958 = ~n38261 & n38587 ;
  assign n38959 = ~n38261 & n38589 ;
  assign n38960 = ~n38261 & n38591 ;
  assign n38961 = ~n38042 & n38623 ;
  assign n38962 = ~n38261 & n38594 ;
  assign n38963 = ~n38261 & n38596 ;
  assign n38964 = ~n38261 & n38598 ;
  assign n38965 = ~n38042 & n38625 ;
  assign n38966 = ~n38042 & n38627 ;
  assign n38967 = ~n38261 & n38602 ;
  assign n38968 = ~n38042 & n38629 ;
  assign n38969 = ~n38261 & n38604 ;
  assign n38970 = ~n38042 & n38631 ;
  assign n38971 = ~n38261 & n38606 ;
  assign n38972 = ~n38042 & n38633 ;
  assign n38973 = ~n38261 & n38608 ;
  assign n38974 = ~n38042 & n38635 ;
  assign n38975 = ~n38261 & n38611 ;
  assign n38976 = ~n38042 & n38638 ;
  assign n38977 = ~n38261 & n38613 ;
  assign n38978 = ~n38042 & n38640 ;
  assign n38979 = ~n38261 & n38616 ;
  assign n38980 = ~n38042 & n38642 ;
  assign n38981 = ~n38261 & n38618 ;
  assign n38982 = ~n38042 & n38644 ;
  assign n38983 = ~n38261 & n38623 ;
  assign n38984 = ~n38042 & n38646 ;
  assign n38985 = ~n38261 & n38625 ;
  assign n38986 = ~n38042 & n38648 ;
  assign n38987 = ~n38261 & n38627 ;
  assign n38988 = ~n38261 & n38629 ;
  assign n38989 = ~n38261 & n38631 ;
  assign n38990 = ~n38261 & n38633 ;
  assign n38991 = ~n38042 & n38650 ;
  assign n38992 = ~n38261 & n38635 ;
  assign n38993 = ~n38261 & n38638 ;
  assign n38994 = ~n38261 & n38640 ;
  assign n38995 = ~n38261 & n38642 ;
  assign n38996 = ~n38261 & n38644 ;
  assign n38997 = ~n38261 & n38646 ;
  assign n38998 = ~n38042 & n38652 ;
  assign n38999 = ~n38261 & n38648 ;
  assign n39000 = ~n38042 & n38654 ;
  assign n39001 = ~n38261 & n38650 ;
  assign n39002 = ~n38042 & n38656 ;
  assign n39003 = ~n38261 & n38652 ;
  assign n39004 = ~n38042 & n38658 ;
  assign n39005 = ~n38261 & n38654 ;
  assign n39006 = ~n38261 & n38656 ;
  assign n39007 = ~n38261 & n38658 ;
  assign n39008 = ~n38261 & n38661 ;
  assign n39009 = ~n38042 & n38661 ;
  assign n39010 = ~n38261 & n38663 ;
  assign n39011 = ~n38261 & n38665 ;
  assign n39012 = ~n38261 & n38667 ;
  assign n39013 = ~n38261 & n38669 ;
  assign n39014 = ~n38042 & n38663 ;
  assign n39015 = ~n38261 & n38866 ;
  assign n39016 = ~n38261 & n38671 ;
  assign n39017 = ~n38042 & n38665 ;
  assign n39018 = ~n38261 & n38673 ;
  assign n39019 = ~n38042 & n38667 ;
  assign n39020 = ~n38261 & n38675 ;
  assign n39021 = ~n38042 & n38669 ;
  assign n39022 = ~n38261 & n38677 ;
  assign n39023 = ~n38261 & n38679 ;
  assign n39024 = ~n38042 & n38821 ;
  assign n39025 = ~n38042 & n38671 ;
  assign n39026 = ~n38261 & n38683 ;
  assign n39027 = ~n38261 & n38685 ;
  assign n39028 = ~n38261 & n38687 ;
  assign n39029 = ~n38261 & n38689 ;
  assign n39030 = ~n38042 & n38673 ;
  assign n39031 = ~n38261 & n38691 ;
  assign n39032 = ~n38042 & n38762 ;
  assign n39033 = ~n38261 & n38694 ;
  assign n39034 = ~n38261 & n38696 ;
  assign n39035 = ~n38261 & n38698 ;
  assign n39036 = ~n38042 & n38675 ;
  assign n39037 = ~n38261 & n38863 ;
  assign n39038 = ~n38042 & n38677 ;
  assign n39039 = ~n38261 & n38701 ;
  assign n39040 = ~n38042 & n38679 ;
  assign n39041 = ~n38261 & n38703 ;
  assign n39042 = ~n38261 & n38705 ;
  assign n39043 = ~n38261 & n38708 ;
  assign n39044 = ~n38261 & n38711 ;
  assign n39045 = ~n38042 & n38683 ;
  assign n39046 = ~n38261 & n38713 ;
  assign n39047 = ~n38261 & n38715 ;
  assign n39048 = ~n38042 & n38685 ;
  assign n39049 = ~n38261 & n38717 ;
  assign n39050 = ~n38261 & n38719 ;
  assign n39051 = ~n38042 & n38687 ;
  assign n39052 = ~n38261 & n38721 ;
  assign n39053 = ~n38261 & n38724 ;
  assign n39054 = ~n38042 & n38689 ;
  assign n39055 = ~n38042 & n38691 ;
  assign n39056 = ~n38261 & n38728 ;
  assign n39057 = ~n38261 & n38731 ;
  assign n39058 = ~n38042 & n38863 ;
  assign n39059 = ~n38042 & n38694 ;
  assign n39060 = ~n38261 & n38733 ;
  assign n39061 = ~n38261 & n38736 ;
  assign n39062 = ~n38042 & n38696 ;
  assign n39063 = ~n38261 & n38738 ;
  assign n39064 = ~n38261 & n38741 ;
  assign n39065 = ~n38042 & n38698 ;
  assign n39066 = ~n38261 & n38743 ;
  assign n39067 = ~n38261 & n38746 ;
  assign n39068 = ~n38261 & n38748 ;
  assign n39069 = ~n38261 & n38751 ;
  assign n39070 = ~n38261 & n38753 ;
  assign n39071 = ~n38261 & n38755 ;
  assign n39072 = ~n38042 & n38701 ;
  assign n39073 = ~n38261 & n38757 ;
  assign n39074 = ~n38261 & n38759 ;
  assign n39075 = ~n38261 & n38762 ;
  assign n39076 = ~n38261 & n38765 ;
  assign n39077 = ~n38042 & n38703 ;
  assign n39078 = ~n38261 & n38767 ;
  assign n39079 = ~n38042 & n38705 ;
  assign n39080 = ~n38261 & n38770 ;
  assign n39081 = ~n38261 & n38772 ;
  assign n39082 = ~n38042 & n38708 ;
  assign n39083 = ~n38261 & n38776 ;
  assign n39084 = ~n38261 & n38778 ;
  assign n39085 = ~n38261 & n38781 ;
  assign n39086 = ~n38261 & n38783 ;
  assign n39087 = ~n38042 & n38711 ;
  assign n39088 = ~n38261 & n38785 ;
  assign n39089 = ~n38261 & n38787 ;
  assign n39090 = ~n38042 & n38713 ;
  assign n39091 = ~n38261 & n38789 ;
  assign n39092 = ~n38042 & n38715 ;
  assign n39093 = ~n38261 & n38792 ;
  assign n39094 = ~n38042 & n38717 ;
  assign n39095 = ~n38261 & n38794 ;
  assign n39096 = ~n38261 & n38797 ;
  assign n39097 = ~n38042 & n38719 ;
  assign n39098 = ~n38261 & n38799 ;
  assign n39099 = ~n38042 & n38721 ;
  assign n39100 = ~n38261 & n38850 ;
  assign n39101 = ~n38261 & n38525 ;
  assign n39102 = ~n38042 & n38724 ;
  assign n39103 = ~n38261 & n38805 ;
  assign n39104 = ~n38261 & n38807 ;
  assign n39105 = ~n38261 & n38848 ;
  assign n39106 = ~n38261 & n38810 ;
  assign n39107 = ~n38261 & n38812 ;
  assign n39108 = ~n38261 & n38815 ;
  assign n39109 = ~n38042 & n38728 ;
  assign n39110 = ~n38261 & n38818 ;
  assign n39111 = ~n38261 & n38845 ;
  assign n39112 = ~n38042 & n38731 ;
  assign n39113 = ~n38042 & n38733 ;
  assign n39114 = ~n38261 & n38821 ;
  assign n39115 = ~n38261 & n38824 ;
  assign n39116 = ~n38042 & n38736 ;
  assign n39117 = ~n38042 & n38738 ;
  assign n39118 = ~n38261 & n38827 ;
  assign n39119 = ~n38261 & n38830 ;
  assign n39120 = ~n38042 & n38741 ;
  assign n39121 = ~n38261 & n38833 ;
  assign n39122 = ~n38261 & n38843 ;
  assign n39123 = ~n38042 & n38743 ;
  assign n39124 = ~n38261 & n38835 ;
  assign n39125 = ~n38261 & n38837 ;
  assign n39126 = ~n38042 & n38746 ;
  assign n39127 = ~n38261 & n38621 ;
  assign n39128 = ~n38261 & n38840 ;
  assign n39129 = ~n38042 & n38748 ;
  assign n39130 = ~n38042 & n38751 ;
  assign n39131 = ~n38042 & n38753 ;
  assign n39132 = ~n38261 & n38853 ;
  assign n39133 = ~n38261 & n38855 ;
  assign n39134 = ~n38042 & n38755 ;
  assign n39135 = ~n38261 & n38858 ;
  assign n39136 = ~n38042 & n38757 ;
  assign n39137 = ~n38261 & n38860 ;
  assign n39138 = ~n38042 & n38759 ;
  assign n39139 = ~n38042 & n38765 ;
  assign n39140 = ~n38261 & n38726 ;
  assign n39141 = ~n38261 & n38869 ;
  assign n39142 = ~n38042 & n38767 ;
  assign n39143 = ~n38261 & n38681 ;
  assign n39144 = ~n38261 & n38874 ;
  assign n39145 = ~n38042 & n38770 ;
  assign n39146 = ~n38261 & n38879 ;
  assign n39147 = ~n38261 & n38882 ;
  assign n39148 = ~n38042 & n38772 ;
  assign n39149 = ~n38042 & n38776 ;
  assign n39150 = ~n38042 & n38778 ;
  assign n39151 = ~n38261 & n38890 ;
  assign n39152 = ~n38261 & n38892 ;
  assign n39153 = ~n38042 & n38781 ;
  assign n39154 = ~n38261 & n38894 ;
  assign n39155 = ~n38042 & n38783 ;
  assign n39156 = ~n38261 & n38496 ;
  assign n39157 = ~n38042 & n38785 ;
  assign n39158 = ~n38042 & n38787 ;
  assign n39159 = ~n38042 & n38882 ;
  assign n39160 = ~n38008 & n38514 ;
  assign n39161 = ~n38042 & n38789 ;
  assign n39162 = ~n38008 & n38512 ;
  assign n39163 = ~n38008 & n38531 ;
  assign n39164 = ~n38042 & n38792 ;
  assign n39165 = ~n38042 & n38794 ;
  assign n39166 = ~n38008 & n38559 ;
  assign n39167 = ~n38042 & n38797 ;
  assign n39168 = ~n38042 & n38799 ;
  assign n39169 = ~n38042 & n38805 ;
  assign n39170 = ~n38042 & n38807 ;
  assign n39171 = ~n38042 & n38810 ;
  assign n39172 = ~n38042 & n38812 ;
  assign n39173 = ~n38042 & n38815 ;
  assign n39174 = ~n38042 & n38818 ;
  assign n39175 = ~n38042 & n38824 ;
  assign n39176 = ~n38008 & n38504 ;
  assign n39177 = ~n38042 & n38835 ;
  assign n39178 = ~n38042 & n38837 ;
  assign n39179 = ~n38042 & n38840 ;
  assign n39180 = ~n38042 & n38843 ;
  assign n39181 = ~n38042 & n38845 ;
  assign n39182 = ~n38042 & n38848 ;
  assign n39183 = ~n38042 & n38850 ;
  assign n39184 = ~n38042 & n38853 ;
  assign n39185 = ~n38042 & n38855 ;
  assign n39186 = ~n38042 & n38858 ;
  assign n39187 = ~n38042 & n38860 ;
  assign n39188 = ~n38042 & n38866 ;
  assign n39189 = ~n38042 & n38869 ;
  assign n39190 = ~n38042 & n38874 ;
  assign n39191 = ~n38042 & n38879 ;
  assign n39192 = ~n38008 & n38523 ;
  assign n39193 = ~n38042 & n38885 ;
  assign n39194 = ~n38042 & n38876 ;
  assign n39195 = ~n38008 & n38521 ;
  assign n39196 = ~n38042 & n38890 ;
  assign n39197 = ~n38042 & n38892 ;
  assign n39198 = ~n38042 & n38894 ;
  assign n39199 = ~n38042 & n38496 ;
  assign n39200 = ~n38008 & n38500 ;
  assign n39201 = ~n38008 & n38506 ;
  assign n39202 = ~n38008 & n38508 ;
  assign n39203 = ~n38008 & n38510 ;
  assign n39204 = ~n38008 & n38516 ;
  assign n39205 = ~n38008 & n38527 ;
  assign n39206 = ~n38008 & n38529 ;
  assign n39207 = ~n38008 & n38533 ;
  assign n39208 = ~n38008 & n38551 ;
  assign n39209 = ~n38008 & n38565 ;
  assign n39210 = ~n38008 & n38567 ;
  assign n39211 = ~n38008 & n38569 ;
  assign n39212 = ~n38008 & n38573 ;
  assign n39213 = ~n38008 & n38575 ;
  assign n39214 = ~n38008 & n38578 ;
  assign n39215 = ~n38008 & n38580 ;
  assign n39216 = ~n38008 & n38583 ;
  assign n39217 = ~n38008 & n38585 ;
  assign n39218 = ~n38008 & n38587 ;
  assign n39219 = ~n38008 & n38589 ;
  assign n39220 = ~n38008 & n38591 ;
  assign n39221 = ~n38008 & n38594 ;
  assign n39222 = ~n38008 & n38596 ;
  assign n39223 = ~n38008 & n38598 ;
  assign n39224 = ~n38008 & n38602 ;
  assign n39225 = ~n38008 & n38604 ;
  assign n39226 = ~n38008 & n38606 ;
  assign n39227 = ~n38008 & n38608 ;
  assign n39228 = ~n38008 & n38611 ;
  assign n39229 = ~n38008 & n38613 ;
  assign n39230 = ~n38008 & n38616 ;
  assign n39231 = ~n38008 & n38618 ;
  assign n39232 = ~n38008 & n38623 ;
  assign n39233 = ~n38008 & n38625 ;
  assign n39234 = ~n38008 & n38627 ;
  assign n39235 = ~n38008 & n38629 ;
  assign n39236 = ~n38008 & n38631 ;
  assign n39237 = ~n38008 & n38633 ;
  assign n39238 = ~n38008 & n38635 ;
  assign n39239 = ~n38008 & n38638 ;
  assign n39240 = ~n38008 & n38640 ;
  assign n39241 = ~n38008 & n38642 ;
  assign n39242 = ~n38008 & n38644 ;
  assign n39243 = ~n38008 & n38646 ;
  assign n39244 = ~n38008 & n38648 ;
  assign n39245 = ~n38008 & n38650 ;
  assign n39246 = ~n38008 & n38652 ;
  assign n39247 = ~n38008 & n38654 ;
  assign n39248 = ~n38008 & n38656 ;
  assign n39249 = ~n38008 & n38658 ;
  assign n39250 = ~n38008 & n38661 ;
  assign n39251 = ~n38008 & n38663 ;
  assign n39252 = ~n38008 & n38665 ;
  assign n39253 = ~n38008 & n38667 ;
  assign n39254 = ~n38008 & n38669 ;
  assign n39255 = ~n38008 & n38671 ;
  assign n39256 = ~n38008 & n38673 ;
  assign n39257 = ~n38008 & n38675 ;
  assign n39258 = ~n38008 & n38677 ;
  assign n39259 = ~n38008 & n38679 ;
  assign n39260 = ~n38008 & n38683 ;
  assign n39261 = ~n38008 & n38685 ;
  assign n39262 = ~n38008 & n38687 ;
  assign n39263 = ~n38008 & n38689 ;
  assign n39264 = ~n38008 & n38691 ;
  assign n39265 = ~n38008 & n38694 ;
  assign n39266 = ~n38008 & n38696 ;
  assign n39267 = ~n38008 & n38698 ;
  assign n39268 = ~n38008 & n38701 ;
  assign n39269 = ~n38008 & n38703 ;
  assign n39270 = ~n38008 & n38705 ;
  assign n39271 = ~n38008 & n38708 ;
  assign n39272 = ~n38008 & n38711 ;
  assign n39273 = ~n38008 & n38713 ;
  assign n39274 = ~n38008 & n38715 ;
  assign n39275 = ~n38008 & n38717 ;
  assign n39276 = ~n38008 & n38719 ;
  assign n39277 = ~n38008 & n38721 ;
  assign n39278 = ~n38008 & n38724 ;
  assign n39279 = ~n38008 & n38728 ;
  assign n39280 = ~n38008 & n38731 ;
  assign n39281 = ~n38008 & n38733 ;
  assign n39282 = ~n38008 & n38736 ;
  assign n39283 = ~n38008 & n38738 ;
  assign n39284 = ~n38008 & n38741 ;
  assign n39285 = ~n38008 & n38743 ;
  assign n39286 = ~n38008 & n38746 ;
  assign n39287 = ~n38008 & n38748 ;
  assign n39288 = ~n38008 & n38751 ;
  assign n39289 = ~n38008 & n38753 ;
  assign n39290 = ~n38008 & n38755 ;
  assign n39291 = ~n38008 & n38757 ;
  assign n39292 = ~n38008 & n38759 ;
  assign n39293 = ~n38008 & n38762 ;
  assign n39294 = ~n38008 & n38765 ;
  assign n39295 = ~n38008 & n38767 ;
  assign n39296 = ~n38008 & n38770 ;
  assign n39297 = ~n38008 & n38772 ;
  assign n39298 = ~n38008 & n38776 ;
  assign n39299 = ~n38008 & n38778 ;
  assign n39300 = ~n38008 & n38781 ;
  assign n39301 = ~n38008 & n38783 ;
  assign n39302 = ~n38008 & n38785 ;
  assign n39303 = ~n38008 & n38787 ;
  assign n39304 = ~n38008 & n38789 ;
  assign n39305 = ~n38008 & n38792 ;
  assign n39306 = ~n38008 & n38794 ;
  assign n39307 = ~n38008 & n38797 ;
  assign n39308 = ~n38008 & n38799 ;
  assign n39309 = ~n38008 & n38525 ;
  assign n39310 = ~n38008 & n38805 ;
  assign n39311 = ~n38008 & n38807 ;
  assign n39312 = ~n38008 & n38810 ;
  assign n39313 = ~n38008 & n38812 ;
  assign n39314 = ~n38008 & n38815 ;
  assign n39315 = ~n38008 & n38818 ;
  assign n39316 = ~n38008 & n38821 ;
  assign n39317 = ~n38008 & n38824 ;
  assign n39318 = ~n38008 & n38827 ;
  assign n39319 = ~n38008 & n38830 ;
  assign n39320 = ~n38008 & n38833 ;
  assign n39321 = ~n38008 & n38835 ;
  assign n39322 = ~n38008 & n38837 ;
  assign n39323 = ~n38008 & n38621 ;
  assign n39324 = ~n38008 & n38840 ;
  assign n39325 = ~n38008 & n38843 ;
  assign n39326 = ~n38008 & n38845 ;
  assign n39327 = ~n38008 & n38848 ;
  assign n39328 = ~n38008 & n38850 ;
  assign n39329 = ~n38008 & n38853 ;
  assign n39330 = ~n38008 & n38855 ;
  assign n39331 = ~n38008 & n38858 ;
  assign n39332 = ~n38008 & n38860 ;
  assign n39333 = ~n38008 & n38863 ;
  assign n39334 = ~n38008 & n38866 ;
  assign n39335 = ~n38008 & n38726 ;
  assign n39336 = ~n38008 & n38869 ;
  assign n39337 = ~n38008 & n38681 ;
  assign n39338 = ~n38008 & n38874 ;
  assign n39339 = ~n38008 & n38879 ;
  assign n39340 = ~n38008 & n38882 ;
  assign n39341 = ~n38008 & n38885 ;
  assign n39342 = ~n38008 & n38876 ;
  assign n39343 = ~n38008 & n38890 ;
  assign n39344 = ~n38008 & n38892 ;
  assign n39345 = ~n38008 & n38894 ;
  assign n39346 = ~n11691 & ~n11693 ;
  assign n39347 = ~\ethreg1_MODER_1_DataOut_reg[4]/NET0131  & n13027 ;
  assign n39348 = n13022 & n39347 ;
  assign n39349 = \rxethmac1_rxstatem1_StateData0_reg/NET0131  & n10579 ;
  assign n39350 = n37575 & n39349 ;
  assign n39351 = ~n39348 & ~n39350 ;
  assign n39352 = \wishbone_TxBDReady_reg/NET0131  & n14063 ;
  assign n39353 = n14058 & n39352 ;
  assign n39354 = n23741 & n23751 ;
  assign n39355 = n32820 & n39354 ;
  assign n39356 = ~n37752 & n37753 ;
  assign n39357 = ~n12747 & ~n37739 ;
  assign n39358 = ~n37564 & n39357 ;
  assign n39359 = n23808 & n32820 ;
  assign n39360 = ~n37752 & n37758 ;
  assign n39361 = n23808 & n37842 ;
  assign n39362 = n37842 & n39354 ;
  assign n39363 = n23808 & n37430 ;
  assign n39364 = n23737 & n32820 ;
  assign n39365 = n32820 & n37426 ;
  assign n39366 = n23737 & n37842 ;
  assign n39367 = n37426 & n37842 ;
  assign n39368 = n37430 & n39354 ;
  assign n39369 = n23737 & n37430 ;
  assign n39370 = n32819 & n37881 ;
  assign n39371 = n23737 & n39370 ;
  assign n39372 = n39354 & n39370 ;
  assign n39373 = n23741 & n23743 ;
  assign n39374 = n37842 & n39373 ;
  assign n39375 = n37430 & n39373 ;
  assign n39376 = n39370 & n39373 ;
  assign n39377 = n32820 & n39373 ;
  assign n39378 = n23743 & n23747 ;
  assign n39379 = n32820 & n39378 ;
  assign n39380 = n37842 & n39378 ;
  assign n39381 = n37430 & n39378 ;
  assign n39382 = n39370 & n39378 ;
  assign n39383 = ~\txethmac1_txcrc_Crc_reg[31]/NET0131  & n35397 ;
  assign n39384 = ~\txethmac1_txstatem1_StateJam_reg/NET0131  & ~\txethmac1_txstatem1_StatePreamble_reg/NET0131  ;
  assign n39385 = n35399 & ~n39384 ;
  assign n39386 = ~n39383 & ~n39385 ;
  assign n39387 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n39386 ;
  assign n39388 = n11455 & ~n39387 ;
  assign n39389 = \txethmac1_RetryCnt_reg[3]/NET0131  & \txethmac1_random1_x_reg[7]/NET0131  ;
  assign n39390 = \wishbone_RxBDRead_reg/NET0131  & ~\wishbone_RxBDReady_reg/NET0131  ;
  assign n39391 = \wishbone_RxReady_reg/NET0131  & ~n39390 ;
  assign n39392 = ~n35445 & ~n35450 ;
  assign n39393 = \wishbone_RxAbortSync3_reg/NET0131  & ~\wishbone_RxAbortSync4_reg/NET0131  ;
  assign n39394 = ~n39390 & ~n39393 ;
  assign n39395 = n39392 & n39394 ;
  assign n39396 = ~n39391 & ~n39395 ;
  assign n39397 = \txethmac1_random1_RandomLatched_reg[2]/NET0131  & ~n36399 ;
  assign n39398 = ~\txethmac1_RetryCnt_reg[2]/NET0131  & ~\txethmac1_RetryCnt_reg[3]/NET0131  ;
  assign n39399 = ~n11418 & n39398 ;
  assign n39400 = \txethmac1_random1_x_reg[2]/NET0131  & n36399 ;
  assign n39401 = ~n39399 & n39400 ;
  assign n39402 = ~n39397 & ~n39401 ;
  assign n39403 = ~\wishbone_RxBDAddress_reg[1]/NET0131  & ~n35450 ;
  assign n39404 = ~n35924 & ~n39403 ;
  assign n39405 = n35448 & n39404 ;
  assign n39406 = \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131  & ~n35448 ;
  assign n39407 = ~n39405 & ~n39406 ;
  assign n39408 = \wishbone_TxEn_needed_reg/NET0131  & ~n18545 ;
  assign n39409 = ~\wishbone_WbEn_q_reg/NET0131  & \wishbone_WbEn_reg/NET0131  ;
  assign n39410 = ~\wishbone_TxBDReady_reg/NET0131  & n39409 ;
  assign n39411 = \ethreg1_MODER_0_DataOut_reg[1]/NET0131  & n39410 ;
  assign n39412 = ~n36299 & n39411 ;
  assign n39413 = ~n39408 & ~n39412 ;
  assign n39414 = \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39415 = n36360 & n39414 ;
  assign n39416 = n36369 & n39415 ;
  assign n39417 = \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39418 = n36360 & n39417 ;
  assign n39419 = n36389 & n39418 ;
  assign n39420 = ~n39416 & ~n39419 ;
  assign n39421 = \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n39422 = n36368 & n39421 ;
  assign n39423 = n36373 & n39422 ;
  assign n39424 = \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39425 = n35523 & n39424 ;
  assign n39426 = n35522 & n39425 ;
  assign n39427 = ~n39423 & ~n39426 ;
  assign n39428 = n39420 & n39427 ;
  assign n39429 = \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39430 = n36362 & n39429 ;
  assign n39431 = n36389 & n39430 ;
  assign n39432 = \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39433 = n35523 & n39432 ;
  assign n39434 = n36379 & n39433 ;
  assign n39435 = ~n39431 & ~n39434 ;
  assign n39436 = \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n39437 = n35521 & n39436 ;
  assign n39438 = n36373 & n39437 ;
  assign n39439 = \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39440 = n36362 & n39439 ;
  assign n39441 = n36379 & n39440 ;
  assign n39442 = ~n39438 & ~n39441 ;
  assign n39443 = n39435 & n39442 ;
  assign n39444 = n39428 & n39443 ;
  assign n39445 = \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39446 = n36360 & n39445 ;
  assign n39447 = n36369 & n39446 ;
  assign n39448 = \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39449 = n36360 & n39448 ;
  assign n39450 = n36389 & n39449 ;
  assign n39451 = ~n39447 & ~n39450 ;
  assign n39452 = \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n39453 = n36368 & n39452 ;
  assign n39454 = n36373 & n39453 ;
  assign n39455 = \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39456 = n35523 & n39455 ;
  assign n39457 = n35522 & n39456 ;
  assign n39458 = ~n39454 & ~n39457 ;
  assign n39459 = n39451 & n39458 ;
  assign n39460 = \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39461 = n36362 & n39460 ;
  assign n39462 = n36389 & n39461 ;
  assign n39463 = \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39464 = n35523 & n39463 ;
  assign n39465 = n36379 & n39464 ;
  assign n39466 = ~n39462 & ~n39465 ;
  assign n39467 = \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n39468 = n35521 & n39467 ;
  assign n39469 = n36373 & n39468 ;
  assign n39470 = \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39471 = n36362 & n39470 ;
  assign n39472 = n36379 & n39471 ;
  assign n39473 = ~n39469 & ~n39472 ;
  assign n39474 = n39466 & n39473 ;
  assign n39475 = n39459 & n39474 ;
  assign n39476 = \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39477 = n36360 & n39476 ;
  assign n39478 = n36369 & n39477 ;
  assign n39479 = \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39480 = n36360 & n39479 ;
  assign n39481 = n36389 & n39480 ;
  assign n39482 = ~n39478 & ~n39481 ;
  assign n39483 = \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n39484 = n36368 & n39483 ;
  assign n39485 = n36373 & n39484 ;
  assign n39486 = \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39487 = n35523 & n39486 ;
  assign n39488 = n35522 & n39487 ;
  assign n39489 = ~n39485 & ~n39488 ;
  assign n39490 = n39482 & n39489 ;
  assign n39491 = \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39492 = n36362 & n39491 ;
  assign n39493 = n36389 & n39492 ;
  assign n39494 = \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131  & \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39495 = n35523 & n39494 ;
  assign n39496 = n36379 & n39495 ;
  assign n39497 = ~n39493 & ~n39496 ;
  assign n39498 = \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
  assign n39499 = n35521 & n39498 ;
  assign n39500 = n36373 & n39499 ;
  assign n39501 = \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  & ~\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
  assign n39502 = n36362 & n39501 ;
  assign n39503 = n36379 & n39502 ;
  assign n39504 = ~n39500 & ~n39503 ;
  assign n39505 = n39497 & n39504 ;
  assign n39506 = n39490 & n39505 ;
  assign n39507 = ~\wishbone_TxAbort_wb_reg/NET0131  & ~\wishbone_TxDone_wb_reg/NET0131  ;
  assign n39508 = ~\wishbone_BlockingTxStatusWrite_reg/NET0131  & ~n36303 ;
  assign n39509 = ~n39507 & ~n39508 ;
  assign n39510 = \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n39511 = ~n10694 & ~n39510 ;
  assign n39512 = \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n39513 = \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n39514 = ~n39512 & ~n39513 ;
  assign n39515 = \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n39516 = ~\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
  assign n39517 = ~n39515 & ~n39516 ;
  assign n39518 = n39514 & n39517 ;
  assign n39519 = n39511 & n39518 ;
  assign n39520 = ~\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
  assign n39521 = ~\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n39522 = \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n39523 = ~n39521 & ~n39522 ;
  assign n39524 = ~n39520 & n39523 ;
  assign n39525 = ~\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
  assign n39526 = ~\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
  assign n39527 = ~n39525 & ~n39526 ;
  assign n39528 = ~\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  & \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
  assign n39529 = \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  & ~\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
  assign n39530 = ~n39528 & ~n39529 ;
  assign n39531 = n39527 & n39530 ;
  assign n39532 = n39524 & n39531 ;
  assign n39533 = ~n15133 & n39532 ;
  assign n39534 = n39519 & n39533 ;
  assign n39535 = ~\txethmac1_ColWindow_reg/NET0131  & ~\txethmac1_txstatem1_StateIPG_reg/NET0131  ;
  assign n39536 = ~\txethmac1_txstatem1_StateIdle_reg/NET0131  & n39535 ;
  assign n39537 = ~n39534 & ~n39536 ;
  assign n39538 = n10564 & n10567 ;
  assign n39539 = ~\txethmac1_txcrc_Crc_reg[30]/NET0131  & n35397 ;
  assign n39540 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & n39539 ;
  assign n39541 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n11495 ;
  assign n39542 = n11494 & n39541 ;
  assign n39543 = ~n39540 & ~n39542 ;
  assign n39544 = ~n11501 & n39543 ;
  assign n39545 = \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  & ~wb_rst_i_pad ;
  assign n39546 = ~n11980 & n39545 ;
  assign n39547 = ~\maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  & ~wb_rst_i_pad ;
  assign n39548 = n11980 & n39547 ;
  assign n39549 = ~n39546 & ~n39548 ;
  assign n39550 = \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  & ~\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  ;
  assign n39551 = \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131  & ~n39550 ;
  assign n39552 = \wishbone_RxStatus_reg[14]/NET0131  & \wishbone_ShiftEnded_reg/NET0131  ;
  assign n39553 = n15779 & n39552 ;
  assign n39554 = ~n39551 & n39553 ;
  assign n39555 = ~\wishbone_RxStatusInLatched_reg[3]/NET0131  & ~\wishbone_RxStatusInLatched_reg[4]/NET0131  ;
  assign n39556 = ~\wishbone_RxStatusInLatched_reg[5]/NET0131  & ~\wishbone_RxStatusInLatched_reg[6]/NET0131  ;
  assign n39557 = n39555 & n39556 ;
  assign n39558 = ~\wishbone_RxStatusInLatched_reg[0]/NET0131  & ~\wishbone_RxStatusInLatched_reg[1]/NET0131  ;
  assign n39559 = ~\macstatus1_LatchedCrcError_reg/NET0131  & n39558 ;
  assign n39560 = n39557 & n39559 ;
  assign n39561 = n39554 & n39560 ;
  assign n39562 = n39557 & n39558 ;
  assign n39563 = n39554 & ~n39562 ;
  assign n39564 = \miim1_RStat_q2_reg/NET0131  & ~\miim1_RStat_q3_reg/NET0131  ;
  assign n39565 = ~\miim1_RStatStart_reg/NET0131  & ~n39564 ;
  assign n39566 = ~\miim1_EndBusy_reg/NET0131  & ~n39565 ;
  assign n39567 = \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  ;
  assign n39568 = \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131  & \txethmac1_TxUsedData_reg/NET0131  ;
  assign n39569 = n39567 & n39568 ;
  assign n39570 = ~\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131  & ~n39569 ;
  assign n39571 = \txethmac1_TxUsedData_reg/NET0131  & n39567 ;
  assign n39572 = n35517 & n39571 ;
  assign n39573 = n35538 & ~n39572 ;
  assign n39574 = ~n39570 & n39573 ;
  assign n39575 = \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  & n35523 ;
  assign n39576 = n35522 & n39575 ;
  assign n39577 = ~\maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001  & ~n39576 ;
  assign n39578 = \wishbone_ShiftEnded_reg/NET0131  & ~n15779 ;
  assign n39579 = \wishbone_rx_fifo_cnt_reg[0]/NET0131  & ~\wishbone_rx_fifo_cnt_reg[1]/NET0131  ;
  assign n39580 = ~\wishbone_rx_fifo_cnt_reg[2]/NET0131  & n39579 ;
  assign n39581 = \wishbone_ShiftEndedSync3_reg/NET0131  & ~\wishbone_ShiftEnded_reg/NET0131  ;
  assign n39582 = n13128 & n16307 ;
  assign n39583 = n39581 & n39582 ;
  assign n39584 = n39580 & n39583 ;
  assign n39585 = ~n39578 & ~n39584 ;
  assign n39586 = \txethmac1_random1_RandomLatched_reg[4]/NET0131  & ~n36399 ;
  assign n39587 = \txethmac1_RetryCnt_reg[2]/NET0131  & ~n37480 ;
  assign n39588 = ~\txethmac1_RetryCnt_reg[3]/NET0131  & ~n39587 ;
  assign n39589 = \txethmac1_random1_x_reg[4]/NET0131  & n36399 ;
  assign n39590 = ~n39588 & n39589 ;
  assign n39591 = ~n39586 & ~n39590 ;
  assign n39592 = ~\wishbone_RxReady_reg/NET0131  & ~n16305 ;
  assign n39593 = \wishbone_r_RxEn_q_reg/NET0131  & ~n35444 ;
  assign n39594 = \wishbone_RxAbortSync2_reg/NET0131  & ~\wishbone_RxAbortSync3_reg/NET0131  ;
  assign n39595 = ~\wishbone_ShiftEnded_reg/NET0131  & ~n39594 ;
  assign n39596 = ~n39593 & n39595 ;
  assign n39597 = ~n39592 & n39596 ;
  assign n39598 = \macstatus1_CarrierSenseLost_reg/NET0131  & ~n11183 ;
  assign n39599 = ~n11185 & n39598 ;
  assign n39600 = ~\CarrierSense_Tx2_reg/NET0131  & ~\ethreg1_MODER_0_DataOut_reg[7]/NET0131  ;
  assign n39601 = ~\ethreg1_MODER_1_DataOut_reg[2]/NET0131  & ~mcoll_pad_i_pad ;
  assign n39602 = n39600 & n39601 ;
  assign n39603 = ~n11201 & n39602 ;
  assign n39604 = ~n39599 & ~n39603 ;
  assign n39605 = ~\wishbone_TxRetry_q_reg/NET0131  & ~n38000 ;
  assign n39606 = ~\maccontrol1_MuxedDone_reg/NET0131  & \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
  assign n39607 = ~\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\txethmac1_TxDone_reg/NET0131  ;
  assign n39608 = n37702 & ~n39607 ;
  assign n39609 = ~n39606 & n39608 ;
  assign n39610 = ~\wishbone_Flop_reg/NET0131  & ~n12725 ;
  assign n39611 = ~n12728 & ~n39610 ;
  assign n39612 = ~n39609 & n39611 ;
  assign n39613 = n39605 & n39612 ;
  assign n39614 = ~n11665 & ~n11766 ;
  assign n39615 = ~\txethmac1_txcrc_Crc_reg[29]/NET0131  & n35397 ;
  assign n39616 = ~\txethmac1_txstatem1_StateJam_reg/NET0131  & \txethmac1_txstatem1_StatePreamble_reg/NET0131  ;
  assign n39617 = n35399 & n39616 ;
  assign n39618 = ~n39615 & ~n39617 ;
  assign n39619 = ~\txethmac1_txstatem1_StateData_reg[0]/NET0131  & ~n39618 ;
  assign n39620 = n11478 & ~n39619 ;
  assign n39621 = \ethreg1_MODER_0_DataOut_reg[1]/NET0131  & ~n36299 ;
  assign n39622 = ~\wishbone_BlockingTxStatusWrite_reg/NET0131  & \wishbone_TxStatus_reg[14]/NET0131  ;
  assign n39623 = n36303 & n39622 ;
  assign n39624 = ~\macstatus1_CarrierSenseLost_reg/NET0131  & ~\macstatus1_LateCollLatched_reg/P0002  ;
  assign n39625 = ~\macstatus1_RetryLimit_reg/P0002  & ~\wishbone_TxUnderRun_reg/NET0131  ;
  assign n39626 = n39624 & n39625 ;
  assign n39627 = n39623 & n39626 ;
  assign n39628 = n39623 & ~n39626 ;
  assign n39629 = ~\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131  & ~n39571 ;
  assign n39630 = n35538 & ~n39569 ;
  assign n39631 = ~n39629 & n39630 ;
  assign n39632 = \maccontrol1_receivecontrol1_Pause_reg/NET0131  & n11978 ;
  assign n39633 = ~\maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131  & ~n39632 ;
  assign n39634 = ~wb_rst_i_pad & ~n11980 ;
  assign n39635 = ~n39633 & n39634 ;
  assign n39636 = \miim1_ScanStat_q2_reg/NET0131  & ~\miim1_SyncStatMdcEn_reg/NET0131  ;
  assign n39637 = ~\miim1_Nvalid_reg/NET0131  & ~n39636 ;
  assign n39638 = ~\miim1_InProgress_q2_reg/NET0131  & \miim1_InProgress_q3_reg/NET0131  ;
  assign n39639 = ~n39637 & ~n39638 ;
  assign n39640 = \TxPauseRq_sync2_reg/NET0131  & ~\TxPauseRq_sync3_reg/NET0131  ;
  assign n39641 = \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & \maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131  ;
  assign n39642 = \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131  & ~n12725 ;
  assign n39643 = \maccontrol1_TxUsedDataOutDetected_reg/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n39644 = n35536 & n39643 ;
  assign n39645 = n39642 & ~n39644 ;
  assign n39646 = ~\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  & ~n39645 ;
  assign n39647 = ~n39641 & ~n39646 ;
  assign n39648 = \wishbone_BlockingTxStatusWrite_sync2_reg/NET0131  & ~\wishbone_BlockingTxStatusWrite_sync3_reg/NET0131  ;
  assign n39649 = \macstatus1_DeferLatched_reg/NET0131  & ~n39648 ;
  assign n39650 = ~n11146 & ~n39649 ;
  assign n39651 = \txethmac1_random1_RandomLatched_reg[3]/NET0131  & ~n36399 ;
  assign n39652 = \txethmac1_random1_x_reg[3]/NET0131  & n36399 ;
  assign n39653 = ~n39398 & n39652 ;
  assign n39654 = ~n39651 & ~n39653 ;
  assign n39655 = \wishbone_RxStatusWriteLatched_reg/NET0131  & ~\wishbone_RxStatusWriteLatched_syncb2_reg/NET0131  ;
  assign n39656 = ~\wishbone_RxStatusWriteLatched_syncb2_reg/NET0131  & \wishbone_ShiftEnded_reg/NET0131  ;
  assign n39657 = n15779 & n39656 ;
  assign n39658 = ~n39655 & ~n39657 ;
  assign n39659 = \miim1_WCtrlData_q2_reg/NET0131  & ~\miim1_WCtrlData_q3_reg/NET0131  ;
  assign n39660 = ~\miim1_WCtrlDataStart_reg/NET0131  & ~n39659 ;
  assign n39661 = ~\miim1_EndBusy_reg/NET0131  & ~n39660 ;
  assign n39662 = ~\ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131  & ~\ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131  ;
  assign n39663 = ~\ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131  & n39662 ;
  assign n39664 = \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131  & ~\ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131  ;
  assign n39665 = ~\miim1_shftrg_ShiftReg_reg[1]/NET0131  & n39664 ;
  assign n39666 = n39663 & n39665 ;
  assign n39667 = n39663 & n39664 ;
  assign n39668 = \miim1_shftrg_LinkFail_reg/NET0131  & ~n39667 ;
  assign n39669 = ~n39666 & ~n39668 ;
  assign n39670 = \wishbone_RxEn_needed_reg/NET0131  & ~n16305 ;
  assign n39671 = ~\wishbone_RxReady_reg/NET0131  & n35444 ;
  assign n39672 = n39409 & n39671 ;
  assign n39673 = ~n39670 & ~n39672 ;
  assign n39674 = ~\wb_adr_i[11]_pad  & ~n23725 ;
  assign n39675 = ~wb_err_o_pad & n23726 ;
  assign n39676 = ~n39674 & n39675 ;
  assign n39677 = \maccontrol1_MuxedDone_reg/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n39678 = ~\maccontrol1_TxDoneInLatched_reg/NET0131  & \maccontrol1_TxUsedDataOutDetected_reg/NET0131  ;
  assign n39679 = \txethmac1_TxDone_reg/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n39680 = n39678 & n39679 ;
  assign n39681 = ~n39677 & ~n39680 ;
  assign n39682 = \maccontrol1_MuxedAbort_reg/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n39683 = ~\maccontrol1_TxAbortInLatched_reg/NET0131  & \maccontrol1_TxUsedDataOutDetected_reg/NET0131  ;
  assign n39684 = \txethmac1_TxAbort_reg/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n39685 = n39683 & n39684 ;
  assign n39686 = ~n39682 & ~n39685 ;
  assign n39687 = ~n37752 & n37981 ;
  assign n39688 = \ethreg1_SetTxCIrq_sync2_reg/NET0131  & ~\ethreg1_SetTxCIrq_sync3_reg/NET0131  ;
  assign n39689 = \ethreg1_SetRxCIrq_sync2_reg/NET0131  & ~\ethreg1_SetRxCIrq_sync3_reg/NET0131  ;
  assign n39690 = \wishbone_BDRead_reg/NET0131  & n39409 ;
  assign n39691 = ~\wishbone_BDWrite_reg[0]/NET0131  & ~\wishbone_BDWrite_reg[1]/NET0131  ;
  assign n39692 = ~\wishbone_BDWrite_reg[2]/NET0131  & ~\wishbone_BDWrite_reg[3]/NET0131  ;
  assign n39693 = n39691 & n39692 ;
  assign n39694 = n38005 & ~n39693 ;
  assign n39695 = ~n39690 & ~n39694 ;
  assign n39696 = \maccontrol1_TxUsedDataOutDetected_reg/NET0131  & n35536 ;
  assign n39697 = n11186 & ~n39696 ;
  assign n39698 = \WillSendControlFrame_sync2_reg/NET0131  & ~\WillSendControlFrame_sync3_reg/NET0131  ;
  assign n39699 = \txethmac1_random1_RandomLatched_reg[1]/NET0131  & ~n36399 ;
  assign n39700 = ~\txethmac1_RetryCnt_reg[1]/NET0131  & n39398 ;
  assign n39701 = \txethmac1_random1_x_reg[1]/NET0131  & n36399 ;
  assign n39702 = ~n39700 & n39701 ;
  assign n39703 = ~n39699 & ~n39702 ;
  assign n39704 = ~\ethreg1_MODER_2_DataOut_reg[0]/NET0131  & \macstatus1_RxColWindow_reg/NET0131  ;
  assign n39705 = ~\ethreg1_MODER_1_DataOut_reg[2]/NET0131  & mcoll_pad_i_pad ;
  assign n39706 = ~n39704 & n39705 ;
  assign n39707 = ~\macstatus1_RxLateCollision_reg/NET0131  & ~n39706 ;
  assign n39708 = ~\macstatus1_LoadRxStatus_reg/NET0131  & ~n39707 ;
  assign n39709 = n11167 & n11201 ;
  assign n39710 = ~\Collision_Tx1_reg/NET0131  & ~\Collision_Tx2_reg/NET0131  ;
  assign n39711 = ~n39709 & ~n39710 ;
  assign n39712 = \wishbone_RxPointerRead_reg/NET0131  & ~n15779 ;
  assign n39713 = \wishbone_RxBDRead_reg/NET0131  & \wishbone_RxBDReady_reg/NET0131  ;
  assign n39714 = ~n39712 & ~n39713 ;
  assign n39715 = ~\maccontrol1_TxUsedDataOutDetected_reg/NET0131  & ~n12725 ;
  assign n39716 = n35536 & ~n39715 ;
  assign n39717 = \wishbone_ShiftEndedSync1_reg/NET0131  & ~\wishbone_ShiftEndedSync2_reg/NET0131  ;
  assign n39718 = ~n39581 & ~n39717 ;
  assign n39719 = ~\ethreg1_MODER_1_DataOut_reg[2]/NET0131  & ~\txethmac1_txstatem1_Rule1_reg/NET0131  ;
  assign n39720 = ~\txethmac1_txstatem1_StatePreamble_reg/NET0131  & n39719 ;
  assign n39721 = ~\txethmac1_txstatem1_StateBackOff_reg/NET0131  & ~\txethmac1_txstatem1_StateIdle_reg/NET0131  ;
  assign n39722 = ~n39720 & n39721 ;
  assign n39723 = ~\wishbone_TxRetryPacketBlocked_reg/NET0131  & ~\wishbone_TxRetryPacket_reg/NET0131  ;
  assign n39724 = \wishbone_TxRetry_wb_q_reg/NET0131  & ~\wishbone_TxRetry_wb_reg/NET0131  ;
  assign n39725 = ~n39723 & ~n39724 ;
  assign n39726 = ~\RxAbort_wb_reg/NET0131  & ~\wishbone_RxAbortLatched_reg/NET0131  ;
  assign n39727 = ~\wishbone_RxAbortSyncb2_reg/NET0131  & ~n39726 ;
  assign n39728 = \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  & ~\txethmac1_TxDone_reg/NET0131  ;
  assign n39729 = ~n39642 & ~n39728 ;
  assign n39730 = ~\wishbone_TxEn_q_reg/NET0131  & \wishbone_TxPointerRead_reg/NET0131  ;
  assign n39731 = \wishbone_TxBDRead_reg/NET0131  & \wishbone_TxBDReady_reg/NET0131  ;
  assign n39732 = ~n39730 & ~n39731 ;
  assign n39733 = ~mrxdv_pad_i_pad & n35444 ;
  assign n39734 = ~n10651 & ~n39733 ;
  assign n39735 = ~\wishbone_BlockingIncrementTxPointer_reg/NET0131  & ~\wishbone_IncrTxPointer_reg/NET0131  ;
  assign n39736 = n13131 & ~n39735 ;
  assign n39737 = ~\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131  & \wishbone_TxUnderRun_sync1_reg/NET0131  ;
  assign n39738 = ~\wishbone_TxUnderRun_wb_reg/NET0131  & ~n39737 ;
  assign n39739 = \miim1_EndBusy_reg/NET0131  & ~\miim1_WCtrlDataStart_q_reg/NET0131  ;
  assign n39740 = ~n29536 & ~n39739 ;
  assign n39741 = \maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131  & ~\wishbone_TxStartFrm_reg/NET0131  ;
  assign n39742 = ~\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  & ~n39741 ;
  assign n39743 = ~\wishbone_TxUnderRun_reg/NET0131  & ~\wishbone_TxUnderRun_sync1_reg/NET0131  ;
  assign n39744 = ~\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131  & ~n39743 ;
  assign n39745 = \maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131  & ~\txethmac1_TxDone_reg/NET0131  ;
  assign n39746 = \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  & \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131  ;
  assign n39747 = ~n39745 & ~n39746 ;
  assign n39748 = ~\miim1_outctrl_Mdo_2d_reg/NET0131  & ~\miim1_shftrg_ShiftReg_reg[7]/NET0131  ;
  assign n39749 = \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  & \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131  ;
  assign n39750 = ~wb_rst_i_pad & ~n15114 ;
  assign n39751 = ~wb_rst_i_pad & ~n15695 ;
  assign n39752 = ~n39750 & ~n39751 ;
  assign n39753 = ~wb_rst_i_pad & ~n17358 ;
  assign n39754 = ~wb_rst_i_pad & ~n17905 ;
  assign n39755 = ~n39753 & ~n39754 ;
  assign n39756 = n39752 & n39755 ;
  assign n39757 = ~wb_rst_i_pad & ~n19273 ;
  assign n39758 = n19794 & n20833 ;
  assign n39759 = n39757 & ~n39758 ;
  assign n39760 = ~wb_rst_i_pad & ~n14044 ;
  assign n39761 = ~wb_rst_i_pad & ~n14593 ;
  assign n39762 = ~n39760 & ~n39761 ;
  assign n39763 = ~n39759 & n39762 ;
  assign n39764 = n39756 & n39763 ;
  assign n39765 = ~wb_rst_i_pad & ~n23718 ;
  assign n39766 = ~wb_rst_i_pad & ~n22688 ;
  assign n39767 = ~wb_rst_i_pad & ~n23202 ;
  assign n39768 = ~n39766 & ~n39767 ;
  assign n39769 = ~n39765 & n39768 ;
  assign n39770 = ~wb_rst_i_pad & ~n18434 ;
  assign n39771 = ~n20315 & ~n39770 ;
  assign n39772 = ~wb_rst_i_pad & ~n21643 ;
  assign n39773 = ~wb_rst_i_pad & ~n22172 ;
  assign n39774 = ~n39772 & ~n39773 ;
  assign n39775 = n39771 & n39774 ;
  assign n39776 = n39769 & n39775 ;
  assign n39777 = n39764 & n39776 ;
  assign n39778 = n14047 & ~n16296 ;
  assign n39779 = ~n39777 & n39778 ;
  assign n39780 = n35550 & ~n35551 ;
  assign n39781 = \wishbone_TxBDReady_reg/NET0131  & ~n14046 ;
  assign n39782 = n39780 & n39781 ;
  assign n39783 = ~n39779 & ~n39782 ;
  assign n39784 = ~wb_rst_i_pad & ~n31508 ;
  assign n39785 = ~wb_rst_i_pad & ~n30970 ;
  assign n39786 = ~wb_rst_i_pad & ~n28901 ;
  assign n39787 = ~\wishbone_RxPointerLSB_rst_reg[0]/NET0131  & ~n16305 ;
  assign n39788 = ~n16307 & ~n39787 ;
  assign n39789 = ~n16305 & n39788 ;
  assign n39790 = ~wb_rst_i_pad & n39788 ;
  assign n39791 = ~n24902 & n39790 ;
  assign n39792 = ~n39789 & ~n39791 ;
  assign n39793 = ~wb_rst_i_pad & ~n24329 ;
  assign n39794 = \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  & n23751 ;
  assign n39795 = n23747 & n39794 ;
  assign n39796 = \ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131  & n23782 ;
  assign n39797 = ~n39795 & ~n39796 ;
  assign n39798 = \ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131  & n23743 ;
  assign n39799 = n23741 & n39798 ;
  assign n39800 = \ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131  & n23743 ;
  assign n39801 = n23747 & n39800 ;
  assign n39802 = ~n39799 & ~n39801 ;
  assign n39803 = n39797 & n39802 ;
  assign n39804 = \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  & n23751 ;
  assign n39805 = n23741 & n39804 ;
  assign n39806 = \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131  & n23794 ;
  assign n39807 = n23741 & n39806 ;
  assign n39808 = ~n39805 & ~n39807 ;
  assign n39809 = n23730 & n39808 ;
  assign n39810 = n39803 & n39809 ;
  assign n39811 = \ethreg1_MODER_1_DataOut_reg[2]/NET0131  & n23808 ;
  assign n39812 = \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131  & n23802 ;
  assign n39813 = ~n39811 & ~n39812 ;
  assign n39814 = \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  & n23737 ;
  assign n39815 = \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131  & n23813 ;
  assign n39816 = ~n39814 & ~n39815 ;
  assign n39817 = n39813 & n39816 ;
  assign n39818 = n39810 & n39817 ;
  assign n39819 = n23730 & ~n39818 ;
  assign n39820 = ~wb_rst_i_pad & ~n39818 ;
  assign n39821 = ~n32189 & n39820 ;
  assign n39822 = ~n39819 & ~n39821 ;
  assign n39823 = ~\wishbone_RxPointerMSB_reg[10]/NET0131  & ~n30337 ;
  assign n39824 = ~n16305 & ~n18517 ;
  assign n39825 = ~n39823 & n39824 ;
  assign n39826 = n18507 & ~n32189 ;
  assign n39827 = ~n39825 & ~n39826 ;
  assign n39828 = \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131  & \ethreg1_irq_rxe_reg/NET0131  ;
  assign n39829 = \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131  & \ethreg1_irq_rxb_reg/NET0131  ;
  assign n39830 = \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131  & \ethreg1_irq_rxc_reg/NET0131  ;
  assign n39831 = ~n39829 & ~n39830 ;
  assign n39832 = ~n39828 & n39831 ;
  assign n39833 = \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131  & \ethreg1_irq_txc_reg/NET0131  ;
  assign n39834 = \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131  & \ethreg1_irq_busy_reg/NET0131  ;
  assign n39835 = ~n39833 & ~n39834 ;
  assign n39836 = \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131  & \ethreg1_irq_txe_reg/NET0131  ;
  assign n39837 = \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131  & \ethreg1_irq_txb_reg/NET0131  ;
  assign n39838 = ~n39836 & ~n39837 ;
  assign n39839 = n39835 & n39838 ;
  assign n39840 = n39832 & n39839 ;
  assign n39841 = \wishbone_tx_fifo_fifo_reg[2][15]/P0001  & ~n35750 ;
  assign n39842 = \m_wb_dat_i[15]_pad  & n35749 ;
  assign n39843 = n35735 & n39842 ;
  assign n39844 = ~n39841 & ~n39843 ;
  assign n39845 = \wishbone_tx_fifo_fifo_reg[2][16]/P0001  & ~n35750 ;
  assign n39846 = \m_wb_dat_i[16]_pad  & n35749 ;
  assign n39847 = n35735 & n39846 ;
  assign n39848 = ~n39845 & ~n39847 ;
  assign n39849 = \wishbone_tx_fifo_fifo_reg[2][17]/P0001  & ~n35750 ;
  assign n39850 = \m_wb_dat_i[17]_pad  & n35749 ;
  assign n39851 = n35735 & n39850 ;
  assign n39852 = ~n39849 & ~n39851 ;
  assign n39853 = \wishbone_tx_fifo_fifo_reg[2][22]/P0001  & ~n35750 ;
  assign n39854 = \m_wb_dat_i[22]_pad  & n35749 ;
  assign n39855 = n35735 & n39854 ;
  assign n39856 = ~n39853 & ~n39855 ;
  assign n39857 = \wishbone_tx_fifo_fifo_reg[2][23]/P0001  & ~n35750 ;
  assign n39858 = \m_wb_dat_i[23]_pad  & n35749 ;
  assign n39859 = n35735 & n39858 ;
  assign n39860 = ~n39857 & ~n39859 ;
  assign n39861 = \wishbone_tx_fifo_fifo_reg[2][25]/P0001  & ~n35750 ;
  assign n39862 = \m_wb_dat_i[25]_pad  & n35749 ;
  assign n39863 = n35735 & n39862 ;
  assign n39864 = ~n39861 & ~n39863 ;
  assign n39865 = \wishbone_tx_fifo_fifo_reg[2][2]/P0001  & ~n35750 ;
  assign n39866 = \m_wb_dat_i[2]_pad  & n35749 ;
  assign n39867 = n35735 & n39866 ;
  assign n39868 = ~n39865 & ~n39867 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g215539/_0_  = n10562 ;
  assign \g215543/_0_  = n10575 ;
  assign \g215547/_0_  = ~n10584 ;
  assign \g215551/_0_  = n10668 ;
  assign \g215552/_0_  = n10681 ;
  assign \g215578/_0_  = n10686 ;
  assign \g215587/_1_  = n11211 ;
  assign \g215589/_1_  = n11223 ;
  assign \g215591/_1_  = n11229 ;
  assign \g215593/_1_  = n11232 ;
  assign \g215595/_1_  = n11236 ;
  assign \g215597/_1_  = n11241 ;
  assign \g215599/_1_  = n11247 ;
  assign \g215601/_1_  = n11253 ;
  assign \g215603/_1_  = n11260 ;
  assign \g215605/_1_  = n11267 ;
  assign \g215607/_1_  = n11275 ;
  assign \g215609/_1_  = n11280 ;
  assign \g215611/_1_  = n11283 ;
  assign \g215613/_1_  = n11287 ;
  assign \g215615/_1_  = n11292 ;
  assign \g215617/_1_  = n11295 ;
  assign \g215618/_0_  = ~n11300 ;
  assign \g215619/_0_  = ~n11302 ;
  assign \g215620/_0_  = n11350 ;
  assign \g215632/_1_  = n11352 ;
  assign \g215634/_0_  = ~n11369 ;
  assign \g215635/_0_  = ~n11379 ;
  assign \g215636/_0_  = ~n11381 ;
  assign \g215637/_0_  = n11385 ;
  assign \g215638/_0_  = n11394 ;
  assign \g215639/_0_  = n11401 ;
  assign \g215655/_1_  = n11417 ;
  assign \g215657/_1_  = n11424 ;
  assign \g215659/_1_  = n11430 ;
  assign \g215661/_1_  = n11433 ;
  assign \g215662/_0_  = ~n11469 ;
  assign \g215663/_0_  = ~n11492 ;
  assign \g215664/_0_  = ~n11516 ;
  assign \g215665/_0_  = n11519 ;
  assign \g215668/_0_  = n11521 ;
  assign \g215674/_0_  = n11536 ;
  assign \g215677/_0_  = ~n11550 ;
  assign \g215686/_0_  = ~n11561 ;
  assign \g215695/_0_  = n11568 ;
  assign \g215696/_0_  = n11574 ;
  assign \g215702/_1__syn_2  = ~n11561 ;
  assign \g215705/_0_  = n11581 ;
  assign \g215706/_0_  = ~n11583 ;
  assign \g215716/_0_  = ~n11597 ;
  assign \g215717/_0_  = ~n11617 ;
  assign \g215718/_0_  = ~n11633 ;
  assign \g215726/_0_  = n11640 ;
  assign \g215727/_0_  = n11645 ;
  assign \g215728/_0_  = ~n11655 ;
  assign \g215760/_0_  = n11660 ;
  assign \g215764/_0_  = ~n11962 ;
  assign \g215765/_0_  = n11998 ;
  assign \g215766/_0_  = n12010 ;
  assign \g215767/_3_  = n12025 ;
  assign \g215768/_3_  = n12036 ;
  assign \g215769/_3_  = n12045 ;
  assign \g215770/_3_  = n12052 ;
  assign \g215771/_3_  = ~n12059 ;
  assign \g215772/_3_  = n12066 ;
  assign \g215773/_3_  = n12076 ;
  assign \g215774/_3_  = n12083 ;
  assign \g215775/_3_  = n12093 ;
  assign \g215776/_3_  = n12100 ;
  assign \g215777/_3_  = n12109 ;
  assign \g215778/_3_  = n12116 ;
  assign \g215779/_3_  = n12123 ;
  assign \g215780/_3_  = n12130 ;
  assign \g215790/_0_  = n12142 ;
  assign \g215791/_0_  = ~n12151 ;
  assign \g215792/_0_  = ~n12160 ;
  assign \g215793/_0_  = ~n12162 ;
  assign \g215801/_0_  = n12174 ;
  assign \g215802/_0_  = n12183 ;
  assign \g215803/_0_  = n12188 ;
  assign \g215804/_0_  = ~n12190 ;
  assign \g215812/_0_  = n12197 ;
  assign \g215813/_0_  = ~n12206 ;
  assign \g215821/_0_  = n12223 ;
  assign \g215823/_0_  = ~n12232 ;
  assign \g215831/_0_  = ~n12237 ;
  assign \g215832/_0_  = ~n12243 ;
  assign \g215833/_0_  = ~n12252 ;
  assign \g215845/_0_  = ~n12259 ;
  assign \g215846/_0_  = n12264 ;
  assign \g215847/_0_  = n12508 ;
  assign \g215872/_0_  = n12513 ;
  assign \g215873/_0_  = n12549 ;
  assign \g215874/_0_  = ~n12563 ;
  assign \g215904/_0_  = n12572 ;
  assign \g215905/_0_  = n12599 ;
  assign \g215906/_0_  = n12610 ;
  assign \g215907/_0_  = n12614 ;
  assign \g215908/_0_  = n12619 ;
  assign \g215909/_0_  = n12622 ;
  assign \g215910/_0_  = n12628 ;
  assign \g215911/_0_  = n12632 ;
  assign \g215912/_0_  = n12636 ;
  assign \g215913/_0_  = n12641 ;
  assign \g215914/_0_  = n12646 ;
  assign \g215915/_0_  = n12651 ;
  assign \g215916/_0_  = n12657 ;
  assign \g215917/_0_  = n12661 ;
  assign \g215918/_0_  = n12665 ;
  assign \g215919/_0_  = n12668 ;
  assign \g215920/_0_  = n12671 ;
  assign \g215923/_0_  = ~n12685 ;
  assign \g215926/_0_  = n12690 ;
  assign \g215941/_0_  = ~n12708 ;
  assign \g215942/_0_  = n12714 ;
  assign \g215943/_0_  = n12717 ;
  assign \g215944/_0_  = ~n12723 ;
  assign \g215945/_0_  = n12761 ;
  assign \g215946/_0_  = n12785 ;
  assign \g215947/_0_  = n12809 ;
  assign \g215948/_0_  = n12833 ;
  assign \g215949/_0_  = n12857 ;
  assign \g215950/_0_  = n12881 ;
  assign \g215951/_0_  = n12905 ;
  assign \g215952/_0_  = n12929 ;
  assign \g215953/_0_  = n12934 ;
  assign \g215954/_0_  = ~n12941 ;
  assign \g215955/_0_  = n12944 ;
  assign \g215956/_0_  = ~n12981 ;
  assign \g215957/_0_  = ~n13018 ;
  assign \g215959/_00_  = n13039 ;
  assign \g215960/_0_  = n13043 ;
  assign \g215962/_0_  = n13048 ;
  assign \g215964/_0_  = n13082 ;
  assign \g215966/_0_  = n13086 ;
  assign \g215972/_0_  = ~n13094 ;
  assign \g216035/_0_  = ~n13212 ;
  assign \g216037/_0_  = ~n13229 ;
  assign \g216038/_0_  = ~n14082 ;
  assign \g216039/_0_  = ~n14603 ;
  assign \g216040/_0_  = ~n15121 ;
  assign \g216041/_0_  = n15126 ;
  assign \g216042/_0_  = n15131 ;
  assign \g216046/_0_  = ~n15167 ;
  assign \g216048/_0_  = ~n15184 ;
  assign \g216057/_0_  = ~n15709 ;
  assign \g216263/_0_  = ~n15725 ;
  assign \g216264/_0_  = ~n15748 ;
  assign \g216265/_0_  = ~n15753 ;
  assign \g216266/_0_  = ~n15758 ;
  assign \g216267/_0_  = ~n15763 ;
  assign \g216268/_0_  = ~n15768 ;
  assign \g216269/_0_  = ~n15773 ;
  assign \g216270/_0_  = ~n15778 ;
  assign \g216271/_0_  = ~n16299 ;
  assign \g216272/_0_  = ~n16304 ;
  assign \g216273/_0_  = ~n16823 ;
  assign \g216284/_0_  = ~n16828 ;
  assign \g216289/_0_  = ~n16833 ;
  assign \g216290/_0_  = ~n16847 ;
  assign \g216292/_0_  = ~n17394 ;
  assign \g216296/_0_  = ~n17923 ;
  assign \g216297/_0_  = ~n18450 ;
  assign \g216300/_0_  = ~n18457 ;
  assign \g216301/_0_  = ~n18464 ;
  assign \g216302/_0_  = ~n18471 ;
  assign \g216303/_0_  = ~n18478 ;
  assign \g216304/_0_  = ~n18485 ;
  assign \g216305/_0_  = ~n18492 ;
  assign \g216306/_0_  = ~n18499 ;
  assign \g216307/_0_  = ~n18506 ;
  assign \g216310/_3_  = ~n18544 ;
  assign \g216311/_3_  = ~n18585 ;
  assign \g216314/u3_syn_7  = ~n15745 ;
  assign \g216322/_3_  = ~n18592 ;
  assign \g216323/_3_  = ~n18597 ;
  assign \g216324/_3_  = ~n18602 ;
  assign \g216325/_3_  = ~n18607 ;
  assign \g216326/_3_  = ~n18612 ;
  assign \g216327/_3_  = ~n18617 ;
  assign \g216328/_3_  = ~n18622 ;
  assign \g216329/_3_  = ~n18627 ;
  assign \g216369/_0_  = ~n18646 ;
  assign \g216370/_0_  = ~n18662 ;
  assign \g216371/_0_  = ~n18674 ;
  assign \g216372/_0_  = ~n18691 ;
  assign \g216373/_0_  = ~n18704 ;
  assign \g216374/_0_  = ~n18715 ;
  assign \g216375/_0_  = ~n18729 ;
  assign \g216376/_0_  = ~n18747 ;
  assign \g216379/_0_  = ~n18762 ;
  assign \g216380/_0_  = ~n19282 ;
  assign \g216381/_0_  = ~n19283 ;
  assign \g216385/_0_  = ~n19803 ;
  assign \g216389/_0_  = n20322 ;
  assign \g216390/_0_  = ~n20851 ;
  assign \g216402/_0_  = n20856 ;
  assign \g216404/_0_  = ~n20863 ;
  assign \g216405/_0_  = ~n20879 ;
  assign \g216406/_0_  = ~n20895 ;
  assign \g216407/_0_  = ~n20910 ;
  assign \g216408/_0_  = ~n20925 ;
  assign \g216409/_0_  = ~n20942 ;
  assign \g216410/_0_  = ~n20958 ;
  assign \g216411/_0_  = ~n20968 ;
  assign \g216412/_0_  = ~n20986 ;
  assign \g216413/_0_  = ~n20997 ;
  assign \g216414/_0_  = ~n21013 ;
  assign \g216415/_0_  = ~n21042 ;
  assign \g216416/_0_  = ~n21059 ;
  assign \g216417/_0_  = ~n21075 ;
  assign \g216418/_0_  = ~n21085 ;
  assign \g216419/_0_  = ~n21096 ;
  assign \g216420/_0_  = ~n21106 ;
  assign \g216421/_0_  = ~n21117 ;
  assign \g216422/_0_  = ~n21127 ;
  assign \g216423/_0_  = ~n21129 ;
  assign \g216424/_0_  = ~n21131 ;
  assign \g216425/_0_  = ~n21645 ;
  assign \g216426/_0_  = ~n21647 ;
  assign \g216427/_0_  = ~n21649 ;
  assign \g216428/_0_  = ~n21651 ;
  assign \g216429/_0_  = ~n21656 ;
  assign \g216430/_0_  = ~n21658 ;
  assign \g216431/_0_  = ~n21660 ;
  assign \g216432/_0_  = ~n22174 ;
  assign \g216433/_0_  = ~n22176 ;
  assign \g216434/_0_  = ~n22690 ;
  assign \g216435/_0_  = ~n23204 ;
  assign \g216436/_0_  = ~n23206 ;
  assign \g216437/_0_  = ~n23720 ;
  assign \g216438/_0_  = ~n23722 ;
  assign \g216439/_3_  = ~n23760 ;
  assign \g216447/_3_  = ~n23775 ;
  assign \g216448/_3_  = ~n24332 ;
  assign \g216452/_0_  = ~n24353 ;
  assign \g216453/_0_  = ~n24385 ;
  assign \g216454/_0_  = ~n24389 ;
  assign \g216455/_0_  = ~n24904 ;
  assign \g216456/_0_  = ~n24906 ;
  assign \g216457/_0_  = ~n24909 ;
  assign \g216458/_3_  = ~n24924 ;
  assign \g216459/_3_  = ~n24939 ;
  assign \g216461/_3_  = ~n24954 ;
  assign \g216462/_3_  = ~n24969 ;
  assign \g216463/_3_  = ~n24984 ;
  assign \g216464/_3_  = ~n24999 ;
  assign \g216465/_3_  = ~n25014 ;
  assign \g216466/_0_  = ~n25016 ;
  assign \g216467/_3_  = ~n25031 ;
  assign \g216468/_3_  = ~n25046 ;
  assign \g216469/_3_  = ~n25615 ;
  assign \g216470/_3_  = ~n26171 ;
  assign \g216471/_3_  = ~n26725 ;
  assign \g216473/_3_  = ~n27267 ;
  assign \g216474/_3_  = ~n27809 ;
  assign \g216475/_3_  = ~n28349 ;
  assign \g216476/_3_  = ~n28364 ;
  assign \g216477/_3_  = ~n28904 ;
  assign \g216478/_0_  = ~n28912 ;
  assign \g216479/_3_  = ~n29478 ;
  assign \g216480/_3_  = ~n29529 ;
  assign \g216481/_3_  = ~n29589 ;
  assign \g216492/_0_  = ~n29594 ;
  assign \g216494/_0_  = ~n29621 ;
  assign \g216495/_3_  = ~n29642 ;
  assign \g216496/_3_  = ~n30194 ;
  assign \g216498/_3_  = ~n30211 ;
  assign \g216499/_3_  = ~n30228 ;
  assign \g216500/_3_  = ~n30245 ;
  assign \g216513/_3_  = ~n30256 ;
  assign \g216514/_3_  = ~n30261 ;
  assign \g216515/_3_  = ~n30268 ;
  assign \g216516/_3_  = ~n30275 ;
  assign \g216517/_3_  = ~n30282 ;
  assign \g216518/_3_  = ~n30287 ;
  assign \g216519/_3_  = ~n30294 ;
  assign \g216520/_3_  = ~n30302 ;
  assign \g216521/_3_  = ~n30310 ;
  assign \g216522/_3_  = ~n30317 ;
  assign \g216523/_3_  = ~n30322 ;
  assign \g216524/_3_  = ~n30331 ;
  assign \g216525/_3_  = ~n30340 ;
  assign \g216526/_3_  = ~n30349 ;
  assign \g216527/_3_  = ~n30355 ;
  assign \g216528/_3_  = ~n30363 ;
  assign \g216529/_3_  = ~n30368 ;
  assign \g216530/_3_  = ~n30375 ;
  assign \g216531/_3_  = ~n30382 ;
  assign \g216532/_3_  = ~n30391 ;
  assign \g216533/_3_  = ~n30398 ;
  assign \g216534/_3_  = ~n30406 ;
  assign \g216535/_3_  = ~n30413 ;
  assign \g216536/_3_  = ~n30418 ;
  assign \g216537/_3_  = ~n30428 ;
  assign \g216538/_3_  = ~n30435 ;
  assign \g216555/_3_  = ~n30973 ;
  assign \g216556/_3_  = ~n31511 ;
  assign \g216557/_3_  = ~n31538 ;
  assign \g216560/_3_  = ~n31546 ;
  assign \g216561/_3_  = ~n31553 ;
  assign \g216562/_3_  = ~n31559 ;
  assign \g216563/_3_  = ~n31566 ;
  assign \g216564/_3_  = ~n31573 ;
  assign \g216565/_3_  = ~n31578 ;
  assign \g216566/_3_  = ~n31585 ;
  assign \g216567/_3_  = ~n31592 ;
  assign \g216568/_3_  = ~n31598 ;
  assign \g216569/_3_  = ~n31605 ;
  assign \g216570/_3_  = ~n31610 ;
  assign \g216571/_3_  = ~n31617 ;
  assign \g216575/_3_  = ~n31624 ;
  assign \g216576/_3_  = ~n31629 ;
  assign \g216577/_3_  = ~n31636 ;
  assign \g216578/_3_  = ~n31644 ;
  assign \g216579/_3_  = ~n31649 ;
  assign \g216580/_3_  = ~n31656 ;
  assign \g216581/_3_  = ~n31662 ;
  assign \g216582/_3_  = ~n31667 ;
  assign \g216583/_3_  = ~n31673 ;
  assign \g216586/_3_  = ~n32191 ;
  assign \g216587/_3_  = ~n32197 ;
  assign \g216588/_3_  = ~n32204 ;
  assign \g216589/_3_  = ~n32211 ;
  assign \g216590/_3_  = ~n32218 ;
  assign \g216591/_3_  = ~n32223 ;
  assign \g216592/_3_  = ~n32229 ;
  assign \g216593/_3_  = ~n32235 ;
  assign \g216594/_3_  = ~n32240 ;
  assign \g216595/_3_  = ~n32246 ;
  assign \g216600/_3_  = n32267 ;
  assign \g216683/_0_  = n32281 ;
  assign \g216689/_0_  = n32285 ;
  assign \g216693/_0_  = n32297 ;
  assign \g216694/_0_  = n32308 ;
  assign \g216727/_0_  = n32316 ;
  assign \g216728/_0_  = ~n32321 ;
  assign \g216729/_0_  = n32325 ;
  assign \g216732/_0_  = ~n32330 ;
  assign \g216733/_0_  = n32336 ;
  assign \g216734/_0_  = n32343 ;
  assign \g216735/_0_  = n32349 ;
  assign \g216736/_0_  = n32353 ;
  assign \g216737/_0_  = n32356 ;
  assign \g216738/_0_  = ~n32363 ;
  assign \g216739/_0_  = n32369 ;
  assign \g216740/_0_  = n32375 ;
  assign \g216741/_0_  = ~n32380 ;
  assign \g216742/_0_  = n32385 ;
  assign \g216743/_0_  = n32390 ;
  assign \g216744/_0_  = n32398 ;
  assign \g216745/_0_  = ~n32403 ;
  assign \g216746/_0_  = ~n32410 ;
  assign \g216748/_0_  = ~n32433 ;
  assign \g216751/_0_  = ~n32443 ;
  assign \g216754/_0_  = n32455 ;
  assign \g216762/_0_  = n32458 ;
  assign \g216934/_2_  = ~n32460 ;
  assign \g216952/_0_  = ~n32481 ;
  assign \g216955/_0_  = ~n32483 ;
  assign \g216969/_0_  = ~n32492 ;
  assign \g216979/_0_  = n32496 ;
  assign \g216984/_0_  = n32500 ;
  assign \g216996/_0_  = n32504 ;
  assign \g217002/_0_  = n32512 ;
  assign \g217014/_0_  = n32550 ;
  assign \g217015/_0_  = n32566 ;
  assign \g217016/_0_  = n32582 ;
  assign \g217017/_0_  = n32598 ;
  assign \g217018/_0_  = n32614 ;
  assign \g217019/_0_  = ~n32627 ;
  assign \g217023/_0_  = n32631 ;
  assign \g217116/_0_  = n32815 ;
  assign \g217146/_3_  = n32859 ;
  assign \g217149/_0_  = ~n32861 ;
  assign \g217151/_0_  = ~n32867 ;
  assign \g217160/_0_  = ~n32874 ;
  assign \g217167/_0_  = ~n32879 ;
  assign \g217168/_0_  = ~n32886 ;
  assign \g217169/_0_  = ~n32893 ;
  assign \g217170/_0_  = ~n32898 ;
  assign \g217171/_0_  = ~n32903 ;
  assign \g217172/_0_  = ~n32908 ;
  assign \g217173/_0_  = ~n32913 ;
  assign \g217174/_0_  = ~n32918 ;
  assign \g217175/_0_  = ~n32923 ;
  assign \g217176/_0_  = ~n32927 ;
  assign \g217177/_0_  = ~n32931 ;
  assign \g217178/_0_  = ~n32935 ;
  assign \g217179/_0_  = ~n32939 ;
  assign \g217180/_0_  = ~n32943 ;
  assign \g217181/_0_  = ~n32947 ;
  assign \g217182/_0_  = ~n32951 ;
  assign \g217183/_0_  = ~n32955 ;
  assign \g217187/_0_  = ~n32961 ;
  assign \g217188/_0_  = ~n32965 ;
  assign \g217189/_0_  = ~n32970 ;
  assign \g217193/_0_  = ~n32974 ;
  assign \g217194/_0_  = ~n32976 ;
  assign \g217195/_0_  = n33016 ;
  assign \g217196/_0_  = ~n33026 ;
  assign \g217202/_0_  = ~n33029 ;
  assign \g217205/_0_  = ~n33035 ;
  assign \g217206/_0_  = ~n33040 ;
  assign \g217207/_0_  = ~n33045 ;
  assign \g217208/_0_  = ~n33050 ;
  assign \g217209/_0_  = ~n33055 ;
  assign \g217210/_0_  = ~n33060 ;
  assign \g217211/_0_  = ~n33065 ;
  assign \g217212/_0_  = ~n33070 ;
  assign \g217213/_0_  = ~n33075 ;
  assign \g217214/_0_  = ~n33080 ;
  assign \g217215/_0_  = ~n33085 ;
  assign \g217216/_0_  = ~n33090 ;
  assign \g217217/_0_  = ~n33095 ;
  assign \g217218/_0_  = ~n33100 ;
  assign \g217219/_0_  = ~n33105 ;
  assign \g217220/_0_  = ~n33110 ;
  assign \g217223/_0_  = n33119 ;
  assign \g217231/_0_  = ~n33125 ;
  assign \g217237/_0_  = n33139 ;
  assign \g217238/_0_  = ~n33152 ;
  assign \g217242/_0_  = ~n33156 ;
  assign \g217243/_0_  = ~n33163 ;
  assign \g217250/_3_  = ~n33221 ;
  assign \g217251/_3_  = ~n33255 ;
  assign \g217252/_3_  = ~n33287 ;
  assign \g217253/_3_  = ~n33321 ;
  assign \g217254/_3_  = ~n33353 ;
  assign \g217255/_3_  = ~n33387 ;
  assign \g217256/_3_  = ~n33419 ;
  assign \g217257/_3_  = ~n33453 ;
  assign \g217258/_3_  = ~n33485 ;
  assign \g217259/_3_  = ~n33517 ;
  assign \g217260/_3_  = ~n33549 ;
  assign \g217261/_3_  = ~n33583 ;
  assign \g217262/_3_  = ~n33617 ;
  assign \g217263/_3_  = ~n33649 ;
  assign \g217264/_3_  = ~n33681 ;
  assign \g217265/_3_  = ~n33713 ;
  assign \g217266/_3_  = ~n33745 ;
  assign \g217267/_3_  = ~n33777 ;
  assign \g217268/_3_  = ~n33809 ;
  assign \g217269/_3_  = ~n33843 ;
  assign \g217270/_3_  = ~n33877 ;
  assign \g217271/_3_  = ~n33911 ;
  assign \g217272/_3_  = ~n33943 ;
  assign \g217273/_3_  = ~n33975 ;
  assign \g217274/_3_  = ~n34009 ;
  assign \g217275/_3_  = ~n34041 ;
  assign \g217276/_3_  = ~n34075 ;
  assign \g217277/_3_  = ~n34109 ;
  assign \g217278/_3_  = ~n34141 ;
  assign \g217279/_3_  = ~n34175 ;
  assign \g217280/_3_  = ~n34207 ;
  assign \g217281/_3_  = ~n34241 ;
  assign \g217282/_3_  = ~n34299 ;
  assign \g217283/_3_  = ~n34331 ;
  assign \g217284/_3_  = ~n34363 ;
  assign \g217285/_3_  = ~n34395 ;
  assign \g217286/_3_  = ~n34427 ;
  assign \g217287/_3_  = ~n34459 ;
  assign \g217288/_3_  = ~n34491 ;
  assign \g217289/_3_  = ~n34523 ;
  assign \g217290/_3_  = ~n34555 ;
  assign \g217291/_3_  = ~n34587 ;
  assign \g217292/_3_  = ~n34619 ;
  assign \g217293/_3_  = ~n34651 ;
  assign \g217294/_3_  = ~n34683 ;
  assign \g217295/_3_  = ~n34715 ;
  assign \g217296/_3_  = ~n34747 ;
  assign \g217297/_3_  = ~n34779 ;
  assign \g217298/_3_  = ~n34811 ;
  assign \g217299/_3_  = ~n34843 ;
  assign \g217300/_3_  = ~n34875 ;
  assign \g217301/_3_  = ~n34907 ;
  assign \g217302/_3_  = ~n34939 ;
  assign \g217303/_3_  = ~n34971 ;
  assign \g217304/_3_  = ~n35003 ;
  assign \g217305/_3_  = ~n35035 ;
  assign \g217306/_3_  = ~n35067 ;
  assign \g217307/_3_  = ~n35099 ;
  assign \g217308/_3_  = ~n35131 ;
  assign \g217309/_3_  = ~n35163 ;
  assign \g217310/_3_  = ~n35195 ;
  assign \g217311/_3_  = ~n35227 ;
  assign \g217312/_3_  = ~n35259 ;
  assign \g217313/_3_  = ~n35291 ;
  assign \g217318/_0_  = ~n35297 ;
  assign \g217662/_0_  = n35322 ;
  assign \g217663/_0_  = n35326 ;
  assign \g217682/_0_  = ~n35342 ;
  assign \g217697/_0_  = ~n35358 ;
  assign \g217698/_0_  = ~n35381 ;
  assign \g217699/_0_  = ~n35389 ;
  assign \g217700/_0_  = n35393 ;
  assign \g217701/_0_  = ~n35396 ;
  assign \g217705/_0_  = ~n35406 ;
  assign \g217711/_0_  = ~n35413 ;
  assign \g217747/_0_  = n35419 ;
  assign \g217753/_00_  = ~n35424 ;
  assign \g217775/_0_  = ~n35443 ;
  assign \g217781/_0_  = ~n35460 ;
  assign \g217784/_0_  = n35463 ;
  assign \g217785/_0_  = ~n35468 ;
  assign \g217786/_0_  = ~n35475 ;
  assign \g217787/_0_  = ~n35481 ;
  assign \g217788/_0_  = ~n35486 ;
  assign \g217790/_0_  = ~n35491 ;
  assign \g217815/_0_  = ~n35503 ;
  assign \g217817/_0_  = ~n35507 ;
  assign \g218145/_0_  = n35509 ;
  assign \g218148/_0_  = n35514 ;
  assign \g218150/_0_  = n35543 ;
  assign \g218167/_0_  = ~n35555 ;
  assign \g218168/_0_  = ~n35560 ;
  assign \g218234/_0_  = ~n35561 ;
  assign \g218235/_0_  = ~n35562 ;
  assign \g218236/_0_  = ~n35567 ;
  assign \g218238/_0_  = n35573 ;
  assign \g218242/_0_  = ~n35577 ;
  assign \g218332/_0_  = n35586 ;
  assign \g218335/_0_  = ~n35596 ;
  assign \g218336/_0_  = ~n35606 ;
  assign \g218337/_0_  = n35617 ;
  assign \g218338/_0_  = n35622 ;
  assign \g218339/_0_  = n35627 ;
  assign \g218340/_0_  = n35632 ;
  assign \g218341/_0_  = n35637 ;
  assign \g218342/_0_  = n35642 ;
  assign \g218343/_0_  = n35653 ;
  assign \g218344/_0_  = n35658 ;
  assign \g218345/_0_  = n35661 ;
  assign \g218346/_0_  = n35664 ;
  assign \g218347/_0_  = n35667 ;
  assign \g218348/_0_  = n35670 ;
  assign \g218349/_0_  = n35673 ;
  assign \g218350/_0_  = n35676 ;
  assign \g218351/_0_  = n35683 ;
  assign \g218352/_0_  = n35686 ;
  assign \g218353/_0_  = n35689 ;
  assign \g218354/_0_  = n35692 ;
  assign \g218355/_0_  = n35695 ;
  assign \g218356/_0_  = n35698 ;
  assign \g218357/_0_  = n35701 ;
  assign \g218358/_0_  = n35704 ;
  assign \g218359/_0_  = n35707 ;
  assign \g218360/_0_  = n35710 ;
  assign \g218398/_3_  = ~n35714 ;
  assign \g218430/_0_  = ~n35721 ;
  assign \g218440/_0_  = ~n35729 ;
  assign \g218452/u3_syn_4  = n35736 ;
  assign \g218495/u3_syn_4  = n35740 ;
  assign \g218517/u3_syn_4  = n35742 ;
  assign \g218554/u3_syn_4  = n35748 ;
  assign \g218575/u3_syn_4  = n35750 ;
  assign \g218600/u3_syn_4  = n35752 ;
  assign \g218621/u3_syn_4  = n35753 ;
  assign \g218638/u3_syn_4  = n35754 ;
  assign \g218659/u3_syn_4  = n35759 ;
  assign \g218673/u3_syn_4  = n35765 ;
  assign \g218707/u3_syn_4  = n35769 ;
  assign \g218735/_3_  = ~n35773 ;
  assign \g219186/_0_  = n35785 ;
  assign \g219187/_0_  = n35792 ;
  assign \g219188/_0_  = n35798 ;
  assign \g219189/_0_  = n35804 ;
  assign \g219190/_0_  = n35816 ;
  assign \g219196/_0_  = n35823 ;
  assign \g219198/_0_  = n35831 ;
  assign \g219199/_0_  = n35841 ;
  assign \g219200/_0_  = n35848 ;
  assign \g219308/_0_  = ~n35855 ;
  assign \g219314/_0_  = ~n35860 ;
  assign \g219326/_0_  = n35864 ;
  assign \g219328/_0_  = n35867 ;
  assign \g219348/_0_  = ~n35881 ;
  assign \g219351/_0_  = ~n35883 ;
  assign \g219363/_0_  = n35887 ;
  assign \g219364/_0_  = ~n35894 ;
  assign \g219365/_0_  = ~n35898 ;
  assign \g219366/_0_  = ~n35902 ;
  assign \g219367/_0_  = ~n35906 ;
  assign \g219368/_0_  = ~n35910 ;
  assign \g219369/_0_  = ~n35914 ;
  assign \g219376/_0_  = n35919 ;
  assign \g219381/_0_  = ~n35922 ;
  assign \g219382/_0_  = ~n35930 ;
  assign \g219384/_0_  = ~n35936 ;
  assign \g219385/_0_  = ~n35946 ;
  assign \g219391/_0_  = n35952 ;
  assign \g219394/_0_  = ~n35961 ;
  assign \g219395/_0_  = ~n35965 ;
  assign \g219396/_0_  = ~n35969 ;
  assign \g219397/_0_  = ~n35973 ;
  assign \g219398/_0_  = ~n35977 ;
  assign \g219399/_0_  = ~n35984 ;
  assign \g219400/_0_  = ~n35987 ;
  assign \g219401/_0_  = ~n35990 ;
  assign \g219402/_0_  = ~n35994 ;
  assign \g219403/_0_  = ~n35998 ;
  assign \g219404/_0_  = ~n36001 ;
  assign \g219405/_0_  = ~n36005 ;
  assign \g219406/_0_  = ~n36009 ;
  assign \g219407/_0_  = ~n36012 ;
  assign \g219408/_0_  = ~n36016 ;
  assign \g219409/_0_  = ~n36022 ;
  assign \g219410/_0_  = ~n36026 ;
  assign \g219411/_0_  = ~n36030 ;
  assign \g219412/_0_  = ~n36034 ;
  assign \g219413/_0_  = ~n36038 ;
  assign \g219414/_0_  = ~n36042 ;
  assign \g219415/_0_  = ~n36046 ;
  assign \g219416/_0_  = ~n36050 ;
  assign \g219417/_0_  = ~n36054 ;
  assign \g219418/_0_  = ~n36058 ;
  assign \g219419/_0_  = ~n36062 ;
  assign \g219420/_0_  = ~n36066 ;
  assign \g219421/_0_  = ~n36069 ;
  assign \g219422/_0_  = ~n36072 ;
  assign \g219423/_0_  = ~n36076 ;
  assign \g219424/_0_  = ~n36080 ;
  assign \g219425/_0_  = ~n36084 ;
  assign \g219426/_0_  = ~n36087 ;
  assign \g219427/_0_  = ~n36091 ;
  assign \g219428/_0_  = ~n36095 ;
  assign \g219429/_0_  = ~n36099 ;
  assign \g219430/_0_  = ~n36102 ;
  assign \g219431/_0_  = ~n36109 ;
  assign \g219432/_0_  = ~n36113 ;
  assign \g219433/_0_  = ~n36117 ;
  assign \g219434/_0_  = ~n36121 ;
  assign \g219435/_0_  = ~n36125 ;
  assign \g219436/_0_  = ~n36129 ;
  assign \g219437/_0_  = ~n36133 ;
  assign \g219438/_0_  = ~n36137 ;
  assign \g219439/_0_  = ~n36141 ;
  assign \g219440/_0_  = ~n36145 ;
  assign \g219441/_0_  = ~n36149 ;
  assign \g219442/_0_  = ~n36153 ;
  assign \g219443/_0_  = ~n36157 ;
  assign \g219444/_0_  = ~n36161 ;
  assign \g219445/_0_  = ~n36165 ;
  assign \g219446/_0_  = ~n36169 ;
  assign \g219447/_0_  = ~n36173 ;
  assign \g219449/_0_  = ~n36179 ;
  assign \g219450/_0_  = ~n36183 ;
  assign \g219451/_0_  = ~n36187 ;
  assign \g219452/_0_  = ~n36191 ;
  assign \g219453/_0_  = ~n36195 ;
  assign \g219454/_0_  = ~n36199 ;
  assign \g219455/_0_  = ~n36203 ;
  assign \g219456/_0_  = ~n36207 ;
  assign \g219457/_0_  = ~n36211 ;
  assign \g219458/_0_  = ~n36215 ;
  assign \g219464/u3_syn_7  = ~n36219 ;
  assign \g219496/u3_syn_4  = n36220 ;
  assign \g219512/u3_syn_4  = n35742 ;
  assign \g219526/u3_syn_4  = n36223 ;
  assign \g219549/u3_syn_4  = n36225 ;
  assign \g219571/u3_syn_4  = n35748 ;
  assign \g219588/u3_syn_4  = n35753 ;
  assign \g219603/u3_syn_4  = n35765 ;
  assign \g219621/u3_syn_4  = n36227 ;
  assign \g219636/_3_  = ~n36232 ;
  assign \g219652/u3_syn_4  = n36236 ;
  assign \g219676/_3_  = n36240 ;
  assign \g219686/_0_  = n36247 ;
  assign \g219689/_0_  = n36249 ;
  assign \g219694/_3_  = n36250 ;
  assign \g220062/_0_  = ~n36251 ;
  assign \g220068/_0_  = ~n36252 ;
  assign \g220069/_0_  = ~n36254 ;
  assign \g220072/_0_  = ~n36262 ;
  assign \g220084/_0_  = n36264 ;
  assign \g220149/_0_  = n36276 ;
  assign \g220162/_0_  = n36284 ;
  assign \g220317/_0_  = n36289 ;
  assign \g220360/_2_  = ~n12169 ;
  assign \g220368/_2_  = ~n36292 ;
  assign \g220369/_0_  = ~n36317 ;
  assign \g220370/_0_  = ~n36327 ;
  assign \g220371/_0_  = ~n36334 ;
  assign \g220372/_0_  = ~n36344 ;
  assign \g220376/_0_  = ~n36357 ;
  assign \g220390/_0_  = ~n36398 ;
  assign \g220395/_0_  = ~n36405 ;
  assign \g220499/_0_  = ~n36430 ;
  assign \g220500/_0_  = ~n36440 ;
  assign \g220501/_0_  = ~n36450 ;
  assign \g220502/_0_  = ~n36460 ;
  assign \g220503/_0_  = ~n36470 ;
  assign \g220504/_0_  = ~n36480 ;
  assign \g220505/_0_  = ~n36490 ;
  assign \g220506/_0_  = ~n36500 ;
  assign \g220507/_0_  = ~n36510 ;
  assign \g220508/_0_  = ~n36520 ;
  assign \g220509/_0_  = ~n36530 ;
  assign \g220510/_0_  = ~n36540 ;
  assign \g220511/_0_  = ~n36550 ;
  assign \g220512/_0_  = ~n36560 ;
  assign \g220513/_0_  = ~n36570 ;
  assign \g220514/_0_  = ~n36580 ;
  assign \g220515/_0_  = ~n36590 ;
  assign \g220516/_0_  = ~n36600 ;
  assign \g220517/_0_  = ~n36610 ;
  assign \g220518/_0_  = ~n36620 ;
  assign \g220519/_0_  = ~n36630 ;
  assign \g220520/_0_  = ~n36640 ;
  assign \g220521/_0_  = ~n36650 ;
  assign \g220522/_0_  = ~n36660 ;
  assign \g220523/_0_  = ~n36670 ;
  assign \g220524/_0_  = ~n36680 ;
  assign \g220525/_0_  = ~n36690 ;
  assign \g220526/_0_  = ~n36700 ;
  assign \g220527/_0_  = ~n36710 ;
  assign \g220528/_0_  = ~n36720 ;
  assign \g220529/_0_  = ~n36730 ;
  assign \g220530/_0_  = ~n36740 ;
  assign \g220531/_0_  = ~n36750 ;
  assign \g220532/_0_  = ~n36760 ;
  assign \g220533/_0_  = ~n36770 ;
  assign \g220534/_0_  = ~n36776 ;
  assign \g220535/_0_  = ~n36784 ;
  assign \g220557/_0_  = ~n36794 ;
  assign \g220558/_0_  = ~n36798 ;
  assign \g220559/_0_  = ~n36802 ;
  assign \g220560/_0_  = ~n36806 ;
  assign \g220561/_0_  = ~n36810 ;
  assign \g220562/_0_  = ~n36814 ;
  assign \g220563/_0_  = ~n36818 ;
  assign \g220564/_0_  = ~n36822 ;
  assign \g220565/_0_  = ~n36826 ;
  assign \g220566/_0_  = ~n36830 ;
  assign \g220567/_0_  = ~n36834 ;
  assign \g220568/_0_  = ~n36838 ;
  assign \g220569/_0_  = ~n36842 ;
  assign \g220570/_0_  = ~n36846 ;
  assign \g220571/_0_  = ~n36856 ;
  assign \g220572/_0_  = ~n36861 ;
  assign \g220573/_0_  = ~n36866 ;
  assign \g220574/_0_  = ~n36871 ;
  assign \g220575/_0_  = ~n36876 ;
  assign \g220576/_0_  = ~n36881 ;
  assign \g220577/_0_  = ~n36886 ;
  assign \g220578/_0_  = ~n36891 ;
  assign \g220579/_0_  = ~n36896 ;
  assign \g220580/_0_  = ~n36901 ;
  assign \g220581/_0_  = ~n36906 ;
  assign \g220582/_0_  = ~n36911 ;
  assign \g220583/_0_  = ~n36916 ;
  assign \g220584/_0_  = ~n36921 ;
  assign \g220585/_0_  = ~n36926 ;
  assign \g220586/_0_  = ~n36931 ;
  assign \g220587/_0_  = ~n36937 ;
  assign \g220588/_0_  = ~n36941 ;
  assign \g220589/_0_  = ~n36945 ;
  assign \g220590/_0_  = ~n36949 ;
  assign \g220591/_0_  = ~n36953 ;
  assign \g220592/_0_  = ~n36957 ;
  assign \g220593/_0_  = ~n36961 ;
  assign \g220594/_0_  = ~n36965 ;
  assign \g220595/_0_  = ~n36969 ;
  assign \g220596/_0_  = ~n36973 ;
  assign \g220597/_0_  = ~n36977 ;
  assign \g220598/_0_  = ~n36981 ;
  assign \g220599/_0_  = ~n36985 ;
  assign \g220600/_0_  = ~n36989 ;
  assign \g220601/_0_  = ~n36993 ;
  assign \g220602/_0_  = ~n36997 ;
  assign \g220603/_0_  = ~n37001 ;
  assign \g220604/_0_  = ~n37008 ;
  assign \g220605/_0_  = ~n37013 ;
  assign \g220606/_0_  = ~n37017 ;
  assign \g220607/_0_  = ~n37021 ;
  assign \g220608/_0_  = ~n37025 ;
  assign \g220609/_0_  = ~n37030 ;
  assign \g220610/_0_  = ~n37034 ;
  assign \g220611/_0_  = ~n37038 ;
  assign \g220612/_0_  = ~n37043 ;
  assign \g220613/_0_  = ~n37047 ;
  assign \g220614/_0_  = ~n37051 ;
  assign \g220615/_0_  = ~n37056 ;
  assign \g220616/_0_  = ~n37060 ;
  assign \g220617/_0_  = ~n37065 ;
  assign \g220618/_0_  = ~n37070 ;
  assign \g220619/_0_  = ~n37075 ;
  assign \g220620/_0_  = ~n37083 ;
  assign \g220621/_0_  = ~n37088 ;
  assign \g220622/_0_  = ~n37093 ;
  assign \g220623/_0_  = ~n37098 ;
  assign \g220624/_0_  = ~n37103 ;
  assign \g220625/_0_  = ~n37108 ;
  assign \g220626/_0_  = ~n37113 ;
  assign \g220627/_0_  = ~n37118 ;
  assign \g220628/_0_  = ~n37123 ;
  assign \g220629/_0_  = ~n37128 ;
  assign \g220630/_0_  = ~n37133 ;
  assign \g220631/_0_  = ~n37138 ;
  assign \g220632/_0_  = ~n37143 ;
  assign \g220633/_0_  = ~n37148 ;
  assign \g220634/_0_  = ~n37153 ;
  assign \g220635/_0_  = ~n37158 ;
  assign \g220636/_0_  = ~n37163 ;
  assign \g220637/_0_  = ~n37168 ;
  assign \g220638/_0_  = ~n37173 ;
  assign \g220639/_0_  = ~n37178 ;
  assign \g220640/_0_  = ~n37183 ;
  assign \g220641/_0_  = ~n37188 ;
  assign \g220642/_0_  = ~n37193 ;
  assign \g220643/_0_  = ~n37202 ;
  assign \g220644/_0_  = ~n37205 ;
  assign \g220645/_0_  = ~n37208 ;
  assign \g220646/_0_  = ~n37211 ;
  assign \g220647/_0_  = ~n37214 ;
  assign \g220648/_0_  = ~n37217 ;
  assign \g220649/_0_  = ~n37220 ;
  assign \g220650/_0_  = ~n37223 ;
  assign \g220651/_0_  = ~n37226 ;
  assign \g220652/_0_  = ~n37229 ;
  assign \g220653/_0_  = ~n37232 ;
  assign \g220654/_0_  = ~n37235 ;
  assign \g220655/_0_  = ~n37238 ;
  assign \g220656/_0_  = ~n37241 ;
  assign \g220657/_0_  = ~n37244 ;
  assign \g220658/_0_  = ~n37247 ;
  assign \g220659/_0_  = ~n37250 ;
  assign \g220660/_0_  = ~n37253 ;
  assign \g220661/_0_  = ~n37256 ;
  assign \g220662/_0_  = ~n37259 ;
  assign \g220663/_0_  = ~n37262 ;
  assign \g220664/_0_  = ~n37265 ;
  assign \g220665/_0_  = ~n37268 ;
  assign \g220666/_0_  = ~n37271 ;
  assign \g220674/_0_  = ~n37275 ;
  assign \g220679/u3_syn_7  = n37278 ;
  assign \g220711/u3_syn_4  = n37279 ;
  assign \g220726/u3_syn_4  = n37281 ;
  assign \g220739/u3_syn_4  = n37283 ;
  assign \g220751/u3_syn_4  = n37285 ;
  assign \g220759/u3_syn_4  = n37288 ;
  assign \g220773/u3_syn_4  = n37289 ;
  assign \g220782/u3_syn_4  = n37291 ;
  assign \g220805/u3_syn_4  = n37293 ;
  assign \g220828/u3_syn_4  = n37296 ;
  assign \g220921/_0_  = n35570 ;
  assign \g220930/u3_syn_4  = n37299 ;
  assign \g220949/_3_  = ~n37305 ;
  assign \g220994/_3_  = n37306 ;
  assign \g221207/_0_  = ~n37339 ;
  assign \g221213/_0_  = ~n11551 ;
  assign \g221223/_0_  = ~n37347 ;
  assign \g221224/_0_  = ~n37355 ;
  assign \g221225/_0_  = n37364 ;
  assign \g221226/_0_  = n37372 ;
  assign \g221231/_0_  = ~n37380 ;
  assign \g221232/_0_  = n37386 ;
  assign \g221234/_0_  = ~n37391 ;
  assign \g221235/_0_  = ~n37396 ;
  assign \g221246/_2_  = n11553 ;
  assign \g221249/_2_  = n11556 ;
  assign \g221265/_0_  = ~n37399 ;
  assign \g221287/_0_  = n37402 ;
  assign \g221325/_0_  = n37407 ;
  assign \g221326/_0_  = n37415 ;
  assign \g221447/_0_  = n37420 ;
  assign \g221449/_0_  = n37423 ;
  assign \g221452/_0_  = n37424 ;
  assign \g221469/_0_  = ~n37425 ;
  assign \g221473/_0_  = n37437 ;
  assign \g221503/_0_  = ~n37440 ;
  assign \g221510/_0_  = n37452 ;
  assign \g221512/_0_  = ~n37462 ;
  assign \g221516/_0_  = ~n37470 ;
  assign \g221517/_0_  = ~n37478 ;
  assign \g221524/_0_  = ~n37485 ;
  assign \g221530/_0_  = ~n37495 ;
  assign \g221592/_0_  = n37498 ;
  assign \g221593/_0_  = n37501 ;
  assign \g221634/u3_syn_4  = n36790 ;
  assign \g221669/u3_syn_4  = n36851 ;
  assign \g221789/u3_syn_4  = n36933 ;
  assign \g221813/u3_syn_4  = n37003 ;
  assign \g221829/u3_syn_4  = n37078 ;
  assign \g221861/u3_syn_4  = n37199 ;
  assign \g221876/_0_  = ~n37504 ;
  assign \g221935/_0_  = n37511 ;
  assign \g221944/_3_  = ~n11524 ;
  assign \g230200/_0_  = n37514 ;
  assign \g230201/_0_  = n37516 ;
  assign \g230205/_0_  = ~n37521 ;
  assign \g230295/_0_  = n37526 ;
  assign \g230297/_0_  = n37532 ;
  assign \g230298/_0_  = n37538 ;
  assign \g230300/_0_  = n37544 ;
  assign \g230302/_0_  = n37557 ;
  assign \g230303/_0_  = ~n37567 ;
  assign \g230343/_0_  = ~n37572 ;
  assign \g230368/_0_  = ~n37574 ;
  assign \g230511/_0_  = n37578 ;
  assign \g230531/_0_  = n37580 ;
  assign \g230635/_2_  = n37581 ;
  assign \g230661/_0_  = n37585 ;
  assign \g230715/_1__syn_2  = n37586 ;
  assign \g230731/_0_  = ~n37621 ;
  assign \g230766/_0_  = n37623 ;
  assign \g230784/_0_  = n37630 ;
  assign \g230785/_0_  = n37635 ;
  assign \g230786/_0_  = n37640 ;
  assign \g230787/_0_  = n37645 ;
  assign \g230797/_0_  = n37648 ;
  assign \g230798/_0_  = ~n37650 ;
  assign \g230803/_0_  = ~n37652 ;
  assign \g230804/_00_  = ~n37657 ;
  assign \g230805/_00_  = ~n37662 ;
  assign \g230806/_00_  = ~n37667 ;
  assign \g230807/_00_  = ~n37672 ;
  assign \g230808/_00_  = ~n37677 ;
  assign \g230809/_00_  = ~n37682 ;
  assign \g230815/_0_  = n37690 ;
  assign \g230816/_2_  = n37692 ;
  assign \g230817/_2_  = n37697 ;
  assign \g230829/_0_  = n37711 ;
  assign \g230834/_0_  = ~n37720 ;
  assign \g230835/_0_  = ~n37729 ;
  assign \g230836/_0_  = ~n37735 ;
  assign \g230837/_0_  = ~n37744 ;
  assign \g230844/_0_  = n37749 ;
  assign \g230863/_3_  = ~n37756 ;
  assign \g230864/_3_  = ~n37761 ;
  assign \g230870/_0_  = ~n37771 ;
  assign \g230988/_3_  = ~n37776 ;
  assign \g231010/_3_  = ~n37781 ;
  assign \g231016/_3_  = ~n37786 ;
  assign \g231042/_3_  = ~n37791 ;
  assign \g231471/_0_  = ~n37798 ;
  assign \g231472/_0_  = n37805 ;
  assign \g231476/_3_  = n37806 ;
  assign \g231480/_3_  = n37807 ;
  assign \g231484/_3_  = n37809 ;
  assign \g231504/_0_  = ~n37813 ;
  assign \g231532/_0_  = n32513 ;
  assign \g231542/_0_  = n37816 ;
  assign \g231560/_1_  = n37821 ;
  assign \g231578/_1_  = n37823 ;
  assign \g231580/_0_  = n37827 ;
  assign \g231590/_1__syn_2  = n35338 ;
  assign \g231615/_0_  = n37831 ;
  assign \g231623/_1_  = n37832 ;
  assign \g231634/_2_  = n37833 ;
  assign \g231635/_0_  = n37836 ;
  assign \g231638/_2_  = n37838 ;
  assign \g231640/_0_  = n37841 ;
  assign \g231653/_2_  = n37843 ;
  assign \g231787/_0_  = n37845 ;
  assign \g231931/_0_  = ~n37850 ;
  assign \g231939/_3_  = n37853 ;
  assign \g231940/_0_  = n37857 ;
  assign \g231951/_0_  = n37863 ;
  assign \g231955/_0_  = ~n37864 ;
  assign \g231956/_0_  = ~n37870 ;
  assign \g231959/_2_  = n37873 ;
  assign \g231960/_0_  = ~n37874 ;
  assign \g231964/_0_  = ~n37883 ;
  assign \g231965/_0_  = n37889 ;
  assign \g231975/_0_  = n37895 ;
  assign \g231986/_1_  = n37897 ;
  assign \g231987/_1_  = n37898 ;
  assign \g231989/_1_  = n37900 ;
  assign \g231990/_1_  = n37901 ;
  assign \g231991/_0_  = ~n37934 ;
  assign \g231992/_0_  = ~n37966 ;
  assign \g231995/_0_  = n37973 ;
  assign \g231998/_0_  = n37979 ;
  assign \g231999/_0_  = n37986 ;
  assign \g232002/_3_  = n38004 ;
  assign \g232035/u3_syn_4  = n38016 ;
  assign \g232038/u3_syn_4  = n38024 ;
  assign \g232046/u3_syn_4  = n38029 ;
  assign \g232054/u3_syn_4  = n38034 ;
  assign \g232062/u3_syn_4  = n38037 ;
  assign \g232070/u3_syn_4  = n38039 ;
  assign \g232078/u3_syn_4  = n38048 ;
  assign \g232079/u3_syn_4  = n38052 ;
  assign \g232087/u3_syn_4  = n38055 ;
  assign \g232096/u3_syn_4  = n38057 ;
  assign \g232104/u3_syn_4  = n38060 ;
  assign \g232112/u3_syn_4  = n38062 ;
  assign \g232120/u3_syn_4  = n38069 ;
  assign \g232128/u3_syn_4  = n38073 ;
  assign \g232136/u3_syn_4  = n38077 ;
  assign \g232144/u3_syn_4  = n38081 ;
  assign \g232152/u3_syn_4  = n38084 ;
  assign \g232161/u3_syn_4  = n38087 ;
  assign \g232169/u3_syn_4  = n38089 ;
  assign \g232177/u3_syn_4  = n38092 ;
  assign \g232185/u3_syn_4  = n38093 ;
  assign \g232186/u3_syn_4  = n38097 ;
  assign \g232194/u3_syn_4  = n38100 ;
  assign \g232202/u3_syn_4  = n38102 ;
  assign \g232210/u3_syn_4  = n38105 ;
  assign \g232218/u3_syn_4  = n38108 ;
  assign \g232226/u3_syn_4  = n38110 ;
  assign \g232234/u3_syn_4  = n38113 ;
  assign \g232242/u3_syn_4  = n38115 ;
  assign \g232251/u3_syn_4  = n38118 ;
  assign \g232259/u3_syn_4  = n38120 ;
  assign \g232267/u3_syn_4  = n38123 ;
  assign \g232275/u3_syn_4  = n38125 ;
  assign \g232283/u3_syn_4  = n38127 ;
  assign \g232291/u3_syn_4  = n38129 ;
  assign \g232299/u3_syn_4  = n38131 ;
  assign \g232307/u3_syn_4  = n38133 ;
  assign \g232315/u3_syn_4  = n38135 ;
  assign \g232324/u3_syn_4  = n38137 ;
  assign \g232332/u3_syn_4  = n38139 ;
  assign \g232341/u3_syn_4  = n38141 ;
  assign \g232349/u3_syn_4  = n38143 ;
  assign \g232357/u3_syn_4  = n38145 ;
  assign \g232366/u3_syn_4  = n38147 ;
  assign \g232374/u3_syn_4  = n38149 ;
  assign \g232382/u3_syn_4  = n38151 ;
  assign \g232390/u3_syn_4  = n38153 ;
  assign \g232398/u3_syn_4  = n38155 ;
  assign \g232406/u3_syn_4  = n38157 ;
  assign \g232414/u3_syn_4  = n38159 ;
  assign \g232422/u3_syn_4  = n38161 ;
  assign \g232427/u3_syn_4  = n38162 ;
  assign \g232431/u3_syn_4  = n38164 ;
  assign \g232439/u3_syn_4  = n38166 ;
  assign \g232444/u3_syn_4  = n38167 ;
  assign \g232452/u3_syn_4  = n38169 ;
  assign \g232461/u3_syn_4  = n38170 ;
  assign \g232471/u3_syn_4  = n38172 ;
  assign \g232479/u3_syn_4  = n38174 ;
  assign \g232487/u3_syn_4  = n38175 ;
  assign \g232495/u3_syn_4  = n38176 ;
  assign \g232503/u3_syn_4  = n38178 ;
  assign \g232506/u3_syn_4  = n38179 ;
  assign \g232514/u3_syn_4  = n38181 ;
  assign \g232527/u3_syn_4  = n38182 ;
  assign \g232530/u3_syn_4  = n38185 ;
  assign \g232536/u3_syn_4  = n38186 ;
  assign \g232544/u3_syn_4  = n38189 ;
  assign \g232551/u3_syn_4  = n38190 ;
  assign \g232557/u3_syn_4  = n38192 ;
  assign \g232568/u3_syn_4  = n38194 ;
  assign \g232576/u3_syn_4  = n38196 ;
  assign \g232585/u3_syn_4  = n38197 ;
  assign \g232593/u3_syn_4  = n38198 ;
  assign \g232597/u3_syn_4  = n38200 ;
  assign \g232609/u3_syn_4  = n38202 ;
  assign \g232617/u3_syn_4  = n38204 ;
  assign \g232625/u3_syn_4  = n38206 ;
  assign \g232633/u3_syn_4  = n38208 ;
  assign \g232641/u3_syn_4  = n38210 ;
  assign \g232649/u3_syn_4  = n38212 ;
  assign \g232657/u3_syn_4  = n38214 ;
  assign \g232665/u3_syn_4  = n38216 ;
  assign \g232673/u3_syn_4  = n38218 ;
  assign \g232681/u3_syn_4  = n38220 ;
  assign \g232689/u3_syn_4  = n38221 ;
  assign \g232697/u3_syn_4  = n38222 ;
  assign \g232705/u3_syn_4  = n38224 ;
  assign \g232713/u3_syn_4  = n38225 ;
  assign \g232717/u3_syn_4  = n38227 ;
  assign \g232729/u3_syn_4  = n38229 ;
  assign \g232737/u3_syn_4  = n38230 ;
  assign \g232745/u3_syn_4  = n38232 ;
  assign \g232749/u3_syn_4  = n38233 ;
  assign \g232761/u3_syn_4  = n38234 ;
  assign \g232768/u3_syn_4  = n38236 ;
  assign \g232777/u3_syn_4  = n38238 ;
  assign \g232785/u3_syn_4  = n38240 ;
  assign \g232793/u3_syn_4  = n38242 ;
  assign \g232801/u3_syn_4  = n38244 ;
  assign \g232809/u3_syn_4  = n38246 ;
  assign \g232815/u3_syn_4  = n38247 ;
  assign \g232823/u3_syn_4  = n38249 ;
  assign \g232833/u3_syn_4  = n38250 ;
  assign \g232841/u3_syn_4  = n38252 ;
  assign \g232846/u3_syn_4  = n38253 ;
  assign \g232851/u3_syn_4  = n38255 ;
  assign \g232865/u3_syn_4  = n38256 ;
  assign \g232873/u3_syn_4  = n38257 ;
  assign \g232881/u3_syn_4  = n38258 ;
  assign \g232882/u3_syn_4  = n38262 ;
  assign \g232895/u3_syn_4  = n38263 ;
  assign \g232904/u3_syn_4  = n38264 ;
  assign \g232913/u3_syn_4  = n38265 ;
  assign \g232921/u3_syn_4  = n38266 ;
  assign \g232928/u3_syn_4  = n38267 ;
  assign \g232934/u3_syn_4  = n38268 ;
  assign \g232945/u3_syn_4  = n38269 ;
  assign \g232953/u3_syn_4  = n38270 ;
  assign \g232954/u3_syn_4  = n38271 ;
  assign \g232969/u3_syn_4  = n38272 ;
  assign \g232977/u3_syn_4  = n38273 ;
  assign \g232981/u3_syn_4  = n38274 ;
  assign \g232993/u3_syn_4  = n38275 ;
  assign \g232995/u3_syn_4  = n38276 ;
  assign \g233009/u3_syn_4  = n38277 ;
  assign \g233017/u3_syn_4  = n38278 ;
  assign \g233025/u3_syn_4  = n38279 ;
  assign \g233033/u3_syn_4  = n38280 ;
  assign \g233041/u3_syn_4  = n38281 ;
  assign \g233047/u3_syn_4  = n38282 ;
  assign \g233057/u3_syn_4  = n38283 ;
  assign \g233065/u3_syn_4  = n38284 ;
  assign \g233073/u3_syn_4  = n38285 ;
  assign \g233081/u3_syn_4  = n38286 ;
  assign \g233087/u3_syn_4  = n38287 ;
  assign \g233097/u3_syn_4  = n38288 ;
  assign \g233105/u3_syn_4  = n38289 ;
  assign \g233113/u3_syn_4  = n38290 ;
  assign \g233121/u3_syn_4  = n38291 ;
  assign \g233128/u3_syn_4  = n38292 ;
  assign \g233134/u3_syn_4  = n38293 ;
  assign \g233144/u3_syn_4  = n38294 ;
  assign \g233153/u3_syn_4  = n38295 ;
  assign \g233161/u3_syn_4  = n38296 ;
  assign \g233169/u3_syn_4  = n38297 ;
  assign \g233177/u3_syn_4  = n38298 ;
  assign \g233185/u3_syn_4  = n38299 ;
  assign \g233193/u3_syn_4  = n38300 ;
  assign \g233201/u3_syn_4  = n38301 ;
  assign \g233209/u3_syn_4  = n38302 ;
  assign \g233217/u3_syn_4  = n38303 ;
  assign \g233219/u3_syn_4  = n38304 ;
  assign \g233229/u3_syn_4  = n38305 ;
  assign \g233241/u3_syn_4  = n38306 ;
  assign \g233249/u3_syn_4  = n38307 ;
  assign \g233257/u3_syn_4  = n38308 ;
  assign \g233265/u3_syn_4  = n38309 ;
  assign \g233273/u3_syn_4  = n38310 ;
  assign \g233281/u3_syn_4  = n38311 ;
  assign \g233289/u3_syn_4  = n38312 ;
  assign \g233297/u3_syn_4  = n38313 ;
  assign \g233305/u3_syn_4  = n38314 ;
  assign \g233313/u3_syn_4  = n38315 ;
  assign \g233321/u3_syn_4  = n38316 ;
  assign \g233329/u3_syn_4  = n38317 ;
  assign \g233337/u3_syn_4  = n38318 ;
  assign \g233345/u3_syn_4  = n38319 ;
  assign \g233353/u3_syn_4  = n38320 ;
  assign \g233361/u3_syn_4  = n38321 ;
  assign \g233369/u3_syn_4  = n38322 ;
  assign \g233377/u3_syn_4  = n38323 ;
  assign \g233382/u3_syn_4  = n38324 ;
  assign \g233392/u3_syn_4  = n38325 ;
  assign \g233394/u3_syn_4  = n38326 ;
  assign \g233409/u3_syn_4  = n38327 ;
  assign \g233417/u3_syn_4  = n38328 ;
  assign \g233425/u3_syn_4  = n38329 ;
  assign \g233433/u3_syn_4  = n38330 ;
  assign \g233441/u3_syn_4  = n38331 ;
  assign \g233449/u3_syn_4  = n38332 ;
  assign \g233453/u3_syn_4  = n38333 ;
  assign \g233465/u3_syn_4  = n38334 ;
  assign \g233473/u3_syn_4  = n38335 ;
  assign \g233481/u3_syn_4  = n38336 ;
  assign \g233489/u3_syn_4  = n38337 ;
  assign \g233497/u3_syn_4  = n38338 ;
  assign \g233505/u3_syn_4  = n38339 ;
  assign \g233513/u3_syn_4  = n38340 ;
  assign \g233516/u3_syn_4  = n38341 ;
  assign \g233529/u3_syn_4  = n38342 ;
  assign \g233531/u3_syn_4  = n38343 ;
  assign \g233546/u3_syn_4  = n38344 ;
  assign \g233554/u3_syn_4  = n38345 ;
  assign \g233562/u3_syn_4  = n38346 ;
  assign \g233570/u3_syn_4  = n38347 ;
  assign \g233578/u3_syn_4  = n38348 ;
  assign \g233586/u3_syn_4  = n38349 ;
  assign \g233594/u3_syn_4  = n38350 ;
  assign \g233602/u3_syn_4  = n38351 ;
  assign \g233603/u3_syn_4  = n38352 ;
  assign \g233618/u3_syn_4  = n38353 ;
  assign \g233626/u3_syn_4  = n38354 ;
  assign \g233634/u3_syn_4  = n38355 ;
  assign \g233642/u3_syn_4  = n38356 ;
  assign \g233650/u3_syn_4  = n38357 ;
  assign \g233658/u3_syn_4  = n38358 ;
  assign \g233666/u3_syn_4  = n38359 ;
  assign \g233674/u3_syn_4  = n38360 ;
  assign \g233682/u3_syn_4  = n38361 ;
  assign \g233690/u3_syn_4  = n38362 ;
  assign \g233698/u3_syn_4  = n38363 ;
  assign \g233706/u3_syn_4  = n38364 ;
  assign \g233714/u3_syn_4  = n38365 ;
  assign \g233722/u3_syn_4  = n38366 ;
  assign \g233730/u3_syn_4  = n38367 ;
  assign \g233738/u3_syn_4  = n38368 ;
  assign \g233746/u3_syn_4  = n38369 ;
  assign \g233754/u3_syn_4  = n38370 ;
  assign \g233762/u3_syn_4  = n38371 ;
  assign \g233770/u3_syn_4  = n38372 ;
  assign \g233778/u3_syn_4  = n38373 ;
  assign \g233783/u3_syn_4  = n38374 ;
  assign \g233794/u3_syn_4  = n38375 ;
  assign \g233802/u3_syn_4  = n38376 ;
  assign \g233806/u3_syn_4  = n38377 ;
  assign \g233818/u3_syn_4  = n38378 ;
  assign \g233826/u3_syn_4  = n38379 ;
  assign \g233828/u3_syn_4  = n38380 ;
  assign \g233838/u3_syn_4  = n38381 ;
  assign \g233850/u3_syn_4  = n38382 ;
  assign \g233858/u3_syn_4  = n38383 ;
  assign \g233860/u3_syn_4  = n38384 ;
  assign \g233870/u3_syn_4  = n38385 ;
  assign \g233881/u3_syn_4  = n38386 ;
  assign \g233890/u3_syn_4  = n38387 ;
  assign \g233899/u3_syn_4  = n38388 ;
  assign \g233908/u3_syn_4  = n38389 ;
  assign \g233917/u3_syn_4  = n38390 ;
  assign \g233919/u3_syn_4  = n38391 ;
  assign \g233927/u3_syn_4  = n38392 ;
  assign \g233935/u3_syn_4  = n38393 ;
  assign \g233943/u3_syn_4  = n38394 ;
  assign \g233945/u3_syn_4  = n38395 ;
  assign \g233953/u3_syn_4  = n38396 ;
  assign \g233961/u3_syn_4  = n38397 ;
  assign \g233969/u3_syn_4  = n38398 ;
  assign \g233977/u3_syn_4  = n38399 ;
  assign \g233985/u3_syn_4  = n38400 ;
  assign \g233993/u3_syn_4  = n38401 ;
  assign \g234001/u3_syn_4  = n38402 ;
  assign \g234008/u3_syn_4  = n38403 ;
  assign \g234009/u3_syn_4  = n38404 ;
  assign \g234024/u3_syn_4  = n38405 ;
  assign \g234032/u3_syn_4  = n38406 ;
  assign \g234038/u3_syn_4  = n38407 ;
  assign \g234056/u3_syn_4  = n38408 ;
  assign \g234063/u3_syn_4  = n38409 ;
  assign \g234071/u3_syn_4  = n38410 ;
  assign \g234079/u3_syn_4  = n38411 ;
  assign \g234098/u3_syn_4  = n38412 ;
  assign \g234106/u3_syn_4  = n38413 ;
  assign \g234114/u3_syn_4  = n38414 ;
  assign \g234122/u3_syn_4  = n38415 ;
  assign \g234130/u3_syn_4  = n38416 ;
  assign \g234138/u3_syn_4  = n38417 ;
  assign \g234145/u3_syn_4  = n38418 ;
  assign \g234156/u3_syn_4  = n38419 ;
  assign \g234162/u3_syn_4  = n38420 ;
  assign \g234171/u3_syn_4  = n38421 ;
  assign \g234183/u3_syn_4  = n38422 ;
  assign \g234248/u3_syn_4  = n38423 ;
  assign \g234265/u3_syn_4  = n38424 ;
  assign \g234273/u3_syn_4  = n38425 ;
  assign \g234281/u3_syn_4  = n38426 ;
  assign \g234289/u3_syn_4  = n38427 ;
  assign \g234297/u3_syn_4  = n38428 ;
  assign \g234306/u3_syn_4  = n38429 ;
  assign \g234314/u3_syn_4  = n38430 ;
  assign \g234322/u3_syn_4  = n38431 ;
  assign \g234331/u3_syn_4  = n38432 ;
  assign \g234339/u3_syn_4  = n38433 ;
  assign \g234347/u3_syn_4  = n38434 ;
  assign \g234355/u3_syn_4  = n38435 ;
  assign \g234363/u3_syn_4  = n38436 ;
  assign \g234371/u3_syn_4  = n38437 ;
  assign \g234379/u3_syn_4  = n38438 ;
  assign \g234387/u3_syn_4  = n38439 ;
  assign \g234395/u3_syn_4  = n38440 ;
  assign \g234403/u3_syn_4  = n38441 ;
  assign \g234411/u3_syn_4  = n38442 ;
  assign \g234419/u3_syn_4  = n38443 ;
  assign \g234427/u3_syn_4  = n38444 ;
  assign \g234435/u3_syn_4  = n38445 ;
  assign \g234443/u3_syn_4  = n38446 ;
  assign \g234451/u3_syn_4  = n38447 ;
  assign \g234459/u3_syn_4  = n38448 ;
  assign \g234467/u3_syn_4  = n38449 ;
  assign \g234475/u3_syn_4  = n38450 ;
  assign \g234483/u3_syn_4  = n38451 ;
  assign \g234491/u3_syn_4  = n38452 ;
  assign \g234499/u3_syn_4  = n38453 ;
  assign \g234507/u3_syn_4  = n38454 ;
  assign \g234515/u3_syn_4  = n38455 ;
  assign \g234523/u3_syn_4  = n38456 ;
  assign \g234531/u3_syn_4  = n38457 ;
  assign \g234539/u3_syn_4  = n38458 ;
  assign \g234547/u3_syn_4  = n38459 ;
  assign \g234555/u3_syn_4  = n38460 ;
  assign \g234563/u3_syn_4  = n38461 ;
  assign \g234571/u3_syn_4  = n38462 ;
  assign \g234579/u3_syn_4  = n38463 ;
  assign \g234587/u3_syn_4  = n38464 ;
  assign \g234595/u3_syn_4  = n38465 ;
  assign \g234604/u3_syn_4  = n38466 ;
  assign \g234612/u3_syn_4  = n38467 ;
  assign \g234620/u3_syn_4  = n38468 ;
  assign \g234628/u3_syn_4  = n38469 ;
  assign \g234636/u3_syn_4  = n38470 ;
  assign \g234644/u3_syn_4  = n38471 ;
  assign \g234652/u3_syn_4  = n38472 ;
  assign \g234660/u3_syn_4  = n38473 ;
  assign \g234668/u3_syn_4  = n38474 ;
  assign \g234676/u3_syn_4  = n38475 ;
  assign \g234684/u3_syn_4  = n38476 ;
  assign \g234692/u3_syn_4  = n38477 ;
  assign \g234700/u3_syn_4  = n38478 ;
  assign \g234708/u3_syn_4  = n38479 ;
  assign \g234716/u3_syn_4  = n38480 ;
  assign \g234725/u3_syn_4  = n38481 ;
  assign \g234733/u3_syn_4  = n38482 ;
  assign \g234741/u3_syn_4  = n38483 ;
  assign \g234749/u3_syn_4  = n38484 ;
  assign \g234757/u3_syn_4  = n38485 ;
  assign \g234765/u3_syn_4  = n38486 ;
  assign \g234773/u3_syn_4  = n38487 ;
  assign \g234781/u3_syn_4  = n38488 ;
  assign \g234789/u3_syn_4  = n38489 ;
  assign \g234798/u3_syn_4  = n38490 ;
  assign \g234806/u3_syn_4  = n38491 ;
  assign \g234814/u3_syn_4  = n38492 ;
  assign \g234822/u3_syn_4  = n38493 ;
  assign \g234830/u3_syn_4  = n38494 ;
  assign \g234838/u3_syn_4  = n38495 ;
  assign \g235911/u3_syn_4  = n38497 ;
  assign \g235912/u3_syn_4  = n38499 ;
  assign \g235920/u3_syn_4  = n38501 ;
  assign \g235928/u3_syn_4  = n38503 ;
  assign \g235936/u3_syn_4  = n38505 ;
  assign \g235944/u3_syn_4  = n38507 ;
  assign \g235952/u3_syn_4  = n38509 ;
  assign \g235960/u3_syn_4  = n38511 ;
  assign \g235968/u3_syn_4  = n38513 ;
  assign \g235976/u3_syn_4  = n38515 ;
  assign \g235984/u3_syn_4  = n38517 ;
  assign \g235992/u3_syn_4  = n38519 ;
  assign \g236000/u3_syn_4  = n38520 ;
  assign \g236008/u3_syn_4  = n38522 ;
  assign \g236016/u3_syn_4  = n38524 ;
  assign \g236021/u3_syn_4  = n38526 ;
  assign \g236025/u3_syn_4  = n38528 ;
  assign \g236033/u3_syn_4  = n38530 ;
  assign \g236041/u3_syn_4  = n38532 ;
  assign \g236049/u3_syn_4  = n38534 ;
  assign \g236057/u3_syn_4  = n38536 ;
  assign \g236065/u3_syn_4  = n38538 ;
  assign \g236073/u3_syn_4  = n38540 ;
  assign \g236081/u3_syn_4  = n38542 ;
  assign \g236089/u3_syn_4  = n38544 ;
  assign \g236097/u3_syn_4  = n38546 ;
  assign \g236105/u3_syn_4  = n38548 ;
  assign \g236113/u3_syn_4  = n38550 ;
  assign \g236121/u3_syn_4  = n38552 ;
  assign \g236129/u3_syn_4  = n38554 ;
  assign \g236137/u3_syn_4  = n38556 ;
  assign \g236145/u3_syn_4  = n38558 ;
  assign \g236153/u3_syn_4  = n38560 ;
  assign \g236161/u3_syn_4  = n38562 ;
  assign \g236169/u3_syn_4  = n38564 ;
  assign \g236177/u3_syn_4  = n38566 ;
  assign \g236185/u3_syn_4  = n38568 ;
  assign \g236193/u3_syn_4  = n38570 ;
  assign \g236196/u3_syn_4  = n38571 ;
  assign \g236198/u3_syn_4  = n38572 ;
  assign \g236203/u3_syn_4  = n38574 ;
  assign \g236211/u3_syn_4  = n38576 ;
  assign \g236219/u3_syn_4  = n38577 ;
  assign \g236220/u3_syn_4  = n38579 ;
  assign \g236229/u3_syn_4  = n38581 ;
  assign \g236232/u3_syn_4  = n38582 ;
  assign \g236238/u3_syn_4  = n38584 ;
  assign \g236246/u3_syn_4  = n38586 ;
  assign \g236255/u3_syn_4  = n38588 ;
  assign \g236263/u3_syn_4  = n38590 ;
  assign \g236271/u3_syn_4  = n38592 ;
  assign \g236275/u3_syn_4  = n38593 ;
  assign \g236280/u3_syn_4  = n38595 ;
  assign \g236288/u3_syn_4  = n38597 ;
  assign \g236296/u3_syn_4  = n38599 ;
  assign \g236304/u3_syn_4  = n38600 ;
  assign \g236305/u3_syn_4  = n38601 ;
  assign \g236306/u3_syn_4  = n38603 ;
  assign \g236315/u3_syn_4  = n38605 ;
  assign \g236323/u3_syn_4  = n38607 ;
  assign \g236331/u3_syn_4  = n38609 ;
  assign \g236334/u3_syn_4  = n38610 ;
  assign \g236340/u3_syn_4  = n38612 ;
  assign \g236348/u3_syn_4  = n38614 ;
  assign \g236357/u3_syn_4  = n38615 ;
  assign \g236359/u3_syn_4  = n38617 ;
  assign \g236367/u3_syn_4  = n38619 ;
  assign \g236374/u3_syn_4  = n38620 ;
  assign \g236376/u3_syn_4  = n38622 ;
  assign \g236377/u3_syn_4  = n38624 ;
  assign \g236385/u3_syn_4  = n38626 ;
  assign \g236393/u3_syn_4  = n38628 ;
  assign \g236402/u3_syn_4  = n38630 ;
  assign \g236410/u3_syn_4  = n38632 ;
  assign \g236419/u3_syn_4  = n38634 ;
  assign \g236427/u3_syn_4  = n38636 ;
  assign \g236433/u3_syn_4  = n38637 ;
  assign \g236436/u3_syn_4  = n38639 ;
  assign \g236444/u3_syn_4  = n38641 ;
  assign \g236452/u3_syn_4  = n38643 ;
  assign \g236460/u3_syn_4  = n38645 ;
  assign \g236468/u3_syn_4  = n38647 ;
  assign \g236476/u3_syn_4  = n38649 ;
  assign \g236484/u3_syn_4  = n38651 ;
  assign \g236492/u3_syn_4  = n38653 ;
  assign \g236500/u3_syn_4  = n38655 ;
  assign \g236508/u3_syn_4  = n38657 ;
  assign \g236516/u3_syn_4  = n38659 ;
  assign \g236518/u3_syn_4  = n38660 ;
  assign \g236525/u3_syn_4  = n38662 ;
  assign \g236533/u3_syn_4  = n38664 ;
  assign \g236542/u3_syn_4  = n38666 ;
  assign \g236550/u3_syn_4  = n38668 ;
  assign \g236559/u3_syn_4  = n38670 ;
  assign \g236567/u3_syn_4  = n38672 ;
  assign \g236575/u3_syn_4  = n38674 ;
  assign \g236583/u3_syn_4  = n38676 ;
  assign \g236591/u3_syn_4  = n38678 ;
  assign \g236599/u3_syn_4  = n38680 ;
  assign \g236607/u3_syn_4  = n38682 ;
  assign \g236608/u3_syn_4  = n38684 ;
  assign \g236616/u3_syn_4  = n38686 ;
  assign \g236624/u3_syn_4  = n38688 ;
  assign \g236632/u3_syn_4  = n38690 ;
  assign \g236640/u3_syn_4  = n38692 ;
  assign \g236647/u3_syn_4  = n38693 ;
  assign \g236649/u3_syn_4  = n38695 ;
  assign \g236659/u3_syn_4  = n38697 ;
  assign \g236671/u3_syn_4  = n38699 ;
  assign \g236677/u3_syn_4  = n38700 ;
  assign \g236688/u3_syn_4  = n38702 ;
  assign \g236696/u3_syn_4  = n38704 ;
  assign \g236705/u3_syn_4  = n38706 ;
  assign \g236712/u3_syn_4  = n38707 ;
  assign \g236718/u3_syn_4  = n38709 ;
  assign \g236729/u3_syn_4  = n38710 ;
  assign \g236732/u3_syn_4  = n38712 ;
  assign \g236745/u3_syn_4  = n38714 ;
  assign \g236753/u3_syn_4  = n38716 ;
  assign \g236761/u3_syn_4  = n38718 ;
  assign \g236769/u3_syn_4  = n38720 ;
  assign \g236777/u3_syn_4  = n38722 ;
  assign \g236779/u3_syn_4  = n38723 ;
  assign \g236788/u3_syn_4  = n38725 ;
  assign \g236800/u3_syn_4  = n38727 ;
  assign \g236802/u3_syn_4  = n38729 ;
  assign \g236805/u3_syn_4  = n38730 ;
  assign \g236813/u3_syn_4  = n38732 ;
  assign \g236825/u3_syn_4  = n38734 ;
  assign \g236829/u3_syn_4  = n38735 ;
  assign \g236837/u3_syn_4  = n38737 ;
  assign \g236849/u3_syn_4  = n38739 ;
  assign \g236854/u3_syn_4  = n38740 ;
  assign \g236860/u3_syn_4  = n38742 ;
  assign \g236872/u3_syn_4  = n38744 ;
  assign \g236878/u3_syn_4  = n38745 ;
  assign \g236884/u3_syn_4  = n38747 ;
  assign \g236896/u3_syn_4  = n38749 ;
  assign \g236903/u3_syn_4  = n38750 ;
  assign \g236908/u3_syn_4  = n38752 ;
  assign \g236920/u3_syn_4  = n38754 ;
  assign \g236930/u3_syn_4  = n38756 ;
  assign \g236939/u3_syn_4  = n38758 ;
  assign \g236947/u3_syn_4  = n38760 ;
  assign \g236949/u3_syn_4  = n38761 ;
  assign \g236956/u3_syn_4  = n38763 ;
  assign \g236962/u3_syn_4  = n38764 ;
  assign \g236965/u3_syn_4  = n38766 ;
  assign \g236980/u3_syn_4  = n38768 ;
  assign \g236988/u3_syn_4  = n38769 ;
  assign \g236989/u3_syn_4  = n38771 ;
  assign \g237004/u3_syn_4  = n38773 ;
  assign \g237005/u3_syn_4  = n38774 ;
  assign \g237020/u3_syn_4  = n38775 ;
  assign \g237021/u3_syn_4  = n38777 ;
  assign \g237033/u3_syn_4  = n38779 ;
  assign \g237044/u3_syn_4  = n38780 ;
  assign \g237045/u3_syn_4  = n38782 ;
  assign \g237056/u3_syn_4  = n38784 ;
  assign \g237068/u3_syn_4  = n38786 ;
  assign \g237076/u3_syn_4  = n38788 ;
  assign \g237084/u3_syn_4  = n38790 ;
  assign \g237092/u3_syn_4  = n38791 ;
  assign \g237095/u3_syn_4  = n38793 ;
  assign \g237107/u3_syn_4  = n38795 ;
  assign \g237110/u3_syn_4  = n38796 ;
  assign \g237119/u3_syn_4  = n38798 ;
  assign \g237131/u3_syn_4  = n38800 ;
  assign \g237135/u3_syn_4  = n38801 ;
  assign \g237148/u3_syn_4  = n38802 ;
  assign \g237152/u3_syn_4  = n38803 ;
  assign \g237165/u3_syn_4  = n38804 ;
  assign \g237168/u3_syn_4  = n38806 ;
  assign \g237180/u3_syn_4  = n38808 ;
  assign \g237185/u3_syn_4  = n38809 ;
  assign \g237192/u3_syn_4  = n38811 ;
  assign \g237204/u3_syn_4  = n38813 ;
  assign \g237209/u3_syn_4  = n38814 ;
  assign \g237215/u3_syn_4  = n38816 ;
  assign \g237229/u3_syn_4  = n38817 ;
  assign \g237231/u3_syn_4  = n38819 ;
  assign \g237245/u3_syn_4  = n38820 ;
  assign \g237251/u3_syn_4  = n38822 ;
  assign \g237260/u3_syn_4  = n38823 ;
  assign \g237262/u3_syn_4  = n38825 ;
  assign \g237277/u3_syn_4  = n38826 ;
  assign \g237281/u3_syn_4  = n38828 ;
  assign \g237293/u3_syn_4  = n38829 ;
  assign \g237294/u3_syn_4  = n38831 ;
  assign \g237310/u3_syn_4  = n38832 ;
  assign \g237311/u3_syn_4  = n38834 ;
  assign \g237323/u3_syn_4  = n38836 ;
  assign \g237334/u3_syn_4  = n38838 ;
  assign \g237342/u3_syn_4  = n38839 ;
  assign \g237350/u3_syn_4  = n38841 ;
  assign \g237353/u3_syn_4  = n38842 ;
  assign \g237359/u3_syn_4  = n38844 ;
  assign \g237367/u3_syn_4  = n38846 ;
  assign \g237368/u3_syn_4  = n38847 ;
  assign \g237378/u3_syn_4  = n38849 ;
  assign \g237391/u3_syn_4  = n38851 ;
  assign \g237392/u3_syn_4  = n38852 ;
  assign \g237403/u3_syn_4  = n38854 ;
  assign \g237415/u3_syn_4  = n38856 ;
  assign \g237417/u3_syn_4  = n38857 ;
  assign \g237431/u3_syn_4  = n38859 ;
  assign \g237439/u3_syn_4  = n38861 ;
  assign \g237440/u3_syn_4  = n38862 ;
  assign \g237454/u3_syn_4  = n38864 ;
  assign \g237457/u3_syn_4  = n38865 ;
  assign \g237472/u3_syn_4  = n38867 ;
  assign \g237480/u3_syn_4  = n38868 ;
  assign \g237488/u3_syn_4  = n38870 ;
  assign \g237496/u3_syn_4  = n38871 ;
  assign \g237499/u3_syn_4  = n38872 ;
  assign \g237512/u3_syn_4  = n38873 ;
  assign \g237515/u3_syn_4  = n38875 ;
  assign \g237525/u3_syn_4  = n38877 ;
  assign \g237529/u3_syn_4  = n38878 ;
  assign \g237535/u3_syn_4  = n38880 ;
  assign \g237541/u3_syn_4  = n38881 ;
  assign \g237553/u3_syn_4  = n38883 ;
  assign \g237561/u3_syn_4  = n38884 ;
  assign \g237569/u3_syn_4  = n38886 ;
  assign \g237575/u3_syn_4  = n38887 ;
  assign \g237578/u3_syn_4  = n38888 ;
  assign \g237581/u3_syn_4  = n38889 ;
  assign \g237591/u3_syn_4  = n38891 ;
  assign \g237602/u3_syn_4  = n38893 ;
  assign \g237610/u3_syn_4  = n38895 ;
  assign \g237617/u3_syn_4  = n38896 ;
  assign \g237623/u3_syn_4  = n38897 ;
  assign \g237633/u3_syn_4  = n38898 ;
  assign \g237635/u3_syn_4  = n38899 ;
  assign \g237648/u3_syn_4  = n38900 ;
  assign \g237658/u3_syn_4  = n38901 ;
  assign \g237659/u3_syn_4  = n38902 ;
  assign \g237660/u3_syn_4  = n38903 ;
  assign \g237668/u3_syn_4  = n38904 ;
  assign \g237675/u3_syn_4  = n38905 ;
  assign \g237684/u3_syn_4  = n38906 ;
  assign \g237692/u3_syn_4  = n38907 ;
  assign \g237693/u3_syn_4  = n38908 ;
  assign \g237705/u3_syn_4  = n38909 ;
  assign \g237716/u3_syn_4  = n38910 ;
  assign \g237717/u3_syn_4  = n38911 ;
  assign \g237729/u3_syn_4  = n38912 ;
  assign \g237740/u3_syn_4  = n38913 ;
  assign \g237741/u3_syn_4  = n38914 ;
  assign \g237756/u3_syn_4  = n38915 ;
  assign \g237764/u3_syn_4  = n38916 ;
  assign \g237768/u3_syn_4  = n38917 ;
  assign \g237780/u3_syn_4  = n38918 ;
  assign \g237782/u3_syn_4  = n38919 ;
  assign \g237792/u3_syn_4  = n38920 ;
  assign \g237804/u3_syn_4  = n38921 ;
  assign \g237812/u3_syn_4  = n38922 ;
  assign \g237820/u3_syn_4  = n38923 ;
  assign \g237828/u3_syn_4  = n38924 ;
  assign \g237836/u3_syn_4  = n38925 ;
  assign \g237844/u3_syn_4  = n38926 ;
  assign \g237852/u3_syn_4  = n38927 ;
  assign \g237860/u3_syn_4  = n38928 ;
  assign \g237868/u3_syn_4  = n38929 ;
  assign \g237876/u3_syn_4  = n38930 ;
  assign \g237884/u3_syn_4  = n38931 ;
  assign \g237888/u3_syn_4  = n38932 ;
  assign \g237895/u3_syn_4  = n38933 ;
  assign \g237907/u3_syn_4  = n38934 ;
  assign \g237916/u3_syn_4  = n38935 ;
  assign \g237924/u3_syn_4  = n38936 ;
  assign \g237931/u3_syn_4  = n38937 ;
  assign \g237940/u3_syn_4  = n38938 ;
  assign \g237949/u3_syn_4  = n38939 ;
  assign \g237950/u3_syn_4  = n38940 ;
  assign \g237955/u3_syn_4  = n38941 ;
  assign \g237961/u3_syn_4  = n38942 ;
  assign \g237965/u3_syn_4  = n38943 ;
  assign \g237975/u3_syn_4  = n38944 ;
  assign \g237983/u3_syn_4  = n38945 ;
  assign \g237989/u3_syn_4  = n38946 ;
  assign \g237999/u3_syn_4  = n38947 ;
  assign \g238007/u3_syn_4  = n38948 ;
  assign \g238015/u3_syn_4  = n38949 ;
  assign \g238017/u3_syn_4  = n38950 ;
  assign \g238033/u3_syn_4  = n38951 ;
  assign \g238035/u3_syn_4  = n38952 ;
  assign \g238049/u3_syn_4  = n38953 ;
  assign \g238057/u3_syn_4  = n38954 ;
  assign \g238065/u3_syn_4  = n38955 ;
  assign \g238072/u3_syn_4  = n38956 ;
  assign \g238081/u3_syn_4  = n38957 ;
  assign \g238082/u3_syn_4  = n38958 ;
  assign \g238097/u3_syn_4  = n38959 ;
  assign \g238105/u3_syn_4  = n38960 ;
  assign \g238113/u3_syn_4  = n38961 ;
  assign \g238114/u3_syn_4  = n38962 ;
  assign \g238129/u3_syn_4  = n38963 ;
  assign \g238137/u3_syn_4  = n38964 ;
  assign \g238145/u3_syn_4  = n38965 ;
  assign \g238153/u3_syn_4  = n38966 ;
  assign \g238161/u3_syn_4  = n38967 ;
  assign \g238163/u3_syn_4  = n38968 ;
  assign \g238177/u3_syn_4  = n38969 ;
  assign \g238179/u3_syn_4  = n38970 ;
  assign \g238194/u3_syn_4  = n38971 ;
  assign \g238197/u3_syn_4  = n38972 ;
  assign \g238209/u3_syn_4  = n38973 ;
  assign \g238213/u3_syn_4  = n38974 ;
  assign \g238225/u3_syn_4  = n38975 ;
  assign \g238229/u3_syn_4  = n38976 ;
  assign \g238237/u3_syn_4  = n38977 ;
  assign \g238250/u3_syn_4  = n38978 ;
  assign \g238257/u3_syn_4  = n38979 ;
  assign \g238263/u3_syn_4  = n38980 ;
  assign \g238269/u3_syn_4  = n38981 ;
  assign \g238282/u3_syn_4  = n38982 ;
  assign \g238285/u3_syn_4  = n38983 ;
  assign \g238298/u3_syn_4  = n38984 ;
  assign \g238301/u3_syn_4  = n38985 ;
  assign \g238314/u3_syn_4  = n38986 ;
  assign \g238316/u3_syn_4  = n38987 ;
  assign \g238329/u3_syn_4  = n38988 ;
  assign \g238338/u3_syn_4  = n38989 ;
  assign \g238346/u3_syn_4  = n38990 ;
  assign \g238351/u3_syn_4  = n38991 ;
  assign \g238356/u3_syn_4  = n38992 ;
  assign \g238368/u3_syn_4  = n38993 ;
  assign \g238378/u3_syn_4  = n38994 ;
  assign \g238386/u3_syn_4  = n38995 ;
  assign \g238394/u3_syn_4  = n38996 ;
  assign \g238402/u3_syn_4  = n38997 ;
  assign \g238409/u3_syn_4  = n38998 ;
  assign \g238412/u3_syn_4  = n38999 ;
  assign \g238427/u3_syn_4  = n39000 ;
  assign \g238429/u3_syn_4  = n39001 ;
  assign \g238443/u3_syn_4  = n39002 ;
  assign \g238448/u3_syn_4  = n39003 ;
  assign \g238457/u3_syn_4  = n39004 ;
  assign \g238460/u3_syn_4  = n39005 ;
  assign \g238472/u3_syn_4  = n39006 ;
  assign \g238484/u3_syn_4  = n39007 ;
  assign \g238492/u3_syn_4  = n39008 ;
  assign \g238500/u3_syn_4  = n39009 ;
  assign \g238505/u3_syn_4  = n39010 ;
  assign \g238516/u3_syn_4  = n39011 ;
  assign \g238524/u3_syn_4  = n39012 ;
  assign \g238532/u3_syn_4  = n39013 ;
  assign \g238534/u3_syn_4  = n39014 ;
  assign \g238544/u3_syn_4  = n39015 ;
  assign \g238549/u3_syn_4  = n39016 ;
  assign \g238550/u3_syn_4  = n39017 ;
  assign \g238565/u3_syn_4  = n39018 ;
  assign \g238566/u3_syn_4  = n39019 ;
  assign \g238582/u3_syn_4  = n39020 ;
  assign \g238583/u3_syn_4  = n39021 ;
  assign \g238594/u3_syn_4  = n39022 ;
  assign \g238606/u3_syn_4  = n39023 ;
  assign \g238614/u3_syn_4  = n39024 ;
  assign \g238615/u3_syn_4  = n39025 ;
  assign \g238619/u3_syn_4  = n39026 ;
  assign \g238631/u3_syn_4  = n39027 ;
  assign \g238639/u3_syn_4  = n39028 ;
  assign \g238647/u3_syn_4  = n39029 ;
  assign \g238649/u3_syn_4  = n39030 ;
  assign \g238659/u3_syn_4  = n39031 ;
  assign \g238670/u3_syn_4  = n39032 ;
  assign \g238671/u3_syn_4  = n39033 ;
  assign \g238680/u3_syn_4  = n39034 ;
  assign \g238688/u3_syn_4  = n39035 ;
  assign \g238691/u3_syn_4  = n39036 ;
  assign \g238696/u3_syn_4  = n39037 ;
  assign \g238705/u3_syn_4  = n39038 ;
  assign \g238708/u3_syn_4  = n39039 ;
  assign \g238721/u3_syn_4  = n39040 ;
  assign \g238724/u3_syn_4  = n39041 ;
  assign \g238736/u3_syn_4  = n39042 ;
  assign \g238745/u3_syn_4  = n39043 ;
  assign \g238753/u3_syn_4  = n39044 ;
  assign \g238757/u3_syn_4  = n39045 ;
  assign \g238764/u3_syn_4  = n39046 ;
  assign \g238776/u3_syn_4  = n39047 ;
  assign \g238781/u3_syn_4  = n39048 ;
  assign \g238787/u3_syn_4  = n39049 ;
  assign \g238799/u3_syn_4  = n39050 ;
  assign \g238807/u3_syn_4  = n39051 ;
  assign \g238811/u3_syn_4  = n39052 ;
  assign \g238824/u3_syn_4  = n39053 ;
  assign \g238830/u3_syn_4  = n39054 ;
  assign \g238841/u3_syn_4  = n39055 ;
  assign \g238843/u3_syn_4  = n39056 ;
  assign \g238855/u3_syn_4  = n39057 ;
  assign \g238859/u3_syn_4  = n39058 ;
  assign \g238863/u3_syn_4  = n39059 ;
  assign \g238868/u3_syn_4  = n39060 ;
  assign \g238880/u3_syn_4  = n39061 ;
  assign \g238888/u3_syn_4  = n39062 ;
  assign \g238892/u3_syn_4  = n39063 ;
  assign \g238903/u3_syn_4  = n39064 ;
  assign \g238911/u3_syn_4  = n39065 ;
  assign \g238915/u3_syn_4  = n39066 ;
  assign \g238927/u3_syn_4  = n39067 ;
  assign \g238937/u3_syn_4  = n39068 ;
  assign \g238945/u3_syn_4  = n39069 ;
  assign \g238953/u3_syn_4  = n39070 ;
  assign \g238961/u3_syn_4  = n39071 ;
  assign \g238970/u3_syn_4  = n39072 ;
  assign \g238971/u3_syn_4  = n39073 ;
  assign \g238983/u3_syn_4  = n39074 ;
  assign \g238994/u3_syn_4  = n39075 ;
  assign \g239002/u3_syn_4  = n39076 ;
  assign \g239009/u3_syn_4  = n39077 ;
  assign \g239015/u3_syn_4  = n39078 ;
  assign \g239025/u3_syn_4  = n39079 ;
  assign \g239030/u3_syn_4  = n39080 ;
  assign \g239041/u3_syn_4  = n39081 ;
  assign \g239048/u3_syn_4  = n39082 ;
  assign \g239053/u3_syn_4  = n39083 ;
  assign \g239065/u3_syn_4  = n39084 ;
  assign \g239073/u3_syn_4  = n39085 ;
  assign \g239081/u3_syn_4  = n39086 ;
  assign \g239082/u3_syn_4  = n39087 ;
  assign \g239093/u3_syn_4  = n39088 ;
  assign \g239105/u3_syn_4  = n39089 ;
  assign \g239108/u3_syn_4  = n39090 ;
  assign \g239117/u3_syn_4  = n39091 ;
  assign \g239129/u3_syn_4  = n39092 ;
  assign \g239137/u3_syn_4  = n39093 ;
  assign \g239139/u3_syn_4  = n39094 ;
  assign \g239148/u3_syn_4  = n39095 ;
  assign \g239160/u3_syn_4  = n39096 ;
  assign \g239162/u3_syn_4  = n39097 ;
  assign \g239172/u3_syn_4  = n39098 ;
  assign \g239184/u3_syn_4  = n39099 ;
  assign \g239187/u3_syn_4  = n39100 ;
  assign \g239189/u3_syn_4  = n39101 ;
  assign \g239201/u3_syn_4  = n39102 ;
  assign \g239208/u3_syn_4  = n39103 ;
  assign \g239217/u3_syn_4  = n39104 ;
  assign \g239219/u3_syn_4  = n39105 ;
  assign \g239226/u3_syn_4  = n39106 ;
  assign \g239234/u3_syn_4  = n39107 ;
  assign \g239242/u3_syn_4  = n39108 ;
  assign \g239246/u3_syn_4  = n39109 ;
  assign \g239257/u3_syn_4  = n39110 ;
  assign \g239258/u3_syn_4  = n39111 ;
  assign \g239263/u3_syn_4  = n39112 ;
  assign \g239275/u3_syn_4  = n39113 ;
  assign \g239277/u3_syn_4  = n39114 ;
  assign \g239291/u3_syn_4  = n39115 ;
  assign \g239296/u3_syn_4  = n39116 ;
  assign \g239308/u3_syn_4  = n39117 ;
  assign \g239311/u3_syn_4  = n39118 ;
  assign \g239322/u3_syn_4  = n39119 ;
  assign \g239329/u3_syn_4  = n39120 ;
  assign \g239338/u3_syn_4  = n39121 ;
  assign \g239339/u3_syn_4  = n39122 ;
  assign \g239346/u3_syn_4  = n39123 ;
  assign \g239351/u3_syn_4  = n39124 ;
  assign \g239363/u3_syn_4  = n39125 ;
  assign \g239370/u3_syn_4  = n39126 ;
  assign \g239375/u3_syn_4  = n39127 ;
  assign \g239387/u3_syn_4  = n39128 ;
  assign \g239395/u3_syn_4  = n39129 ;
  assign \g239418/u3_syn_4  = n39130 ;
  assign \g239439/u3_syn_4  = n39131 ;
  assign \g239442/u3_syn_4  = n39132 ;
  assign \g239454/u3_syn_4  = n39133 ;
  assign \g239464/u3_syn_4  = n39134 ;
  assign \g239470/u3_syn_4  = n39135 ;
  assign \g239481/u3_syn_4  = n39136 ;
  assign \g239487/u3_syn_4  = n39137 ;
  assign \g239497/u3_syn_4  = n39138 ;
  assign \g239520/u3_syn_4  = n39139 ;
  assign \g239532/u3_syn_4  = n39140 ;
  assign \g239543/u3_syn_4  = n39141 ;
  assign \g239551/u3_syn_4  = n39142 ;
  assign \g239552/u3_syn_4  = n39143 ;
  assign \g239567/u3_syn_4  = n39144 ;
  assign \g239575/u3_syn_4  = n39145 ;
  assign \g239579/u3_syn_4  = n39146 ;
  assign \g239592/u3_syn_4  = n39147 ;
  assign \g239594/u3_syn_4  = n39148 ;
  assign \g239608/u3_syn_4  = n39149 ;
  assign \g239626/u3_syn_4  = n39150 ;
  assign \g239634/u3_syn_4  = n39151 ;
  assign \g239646/u3_syn_4  = n39152 ;
  assign \g239649/u3_syn_4  = n39153 ;
  assign \g239657/u3_syn_4  = n39154 ;
  assign \g239670/u3_syn_4  = n39155 ;
  assign \g239673/u3_syn_4  = n39156 ;
  assign \g239686/u3_syn_4  = n39157 ;
  assign \g239694/u3_syn_4  = n39158 ;
  assign \g239695/u3_syn_4  = n39159 ;
  assign \g239701/u3_syn_4  = n39160 ;
  assign \g239705/u3_syn_4  = n39161 ;
  assign \g239709/u3_syn_4  = n39162 ;
  assign \g239715/u3_syn_4  = n39163 ;
  assign \g239717/u3_syn_4  = n39164 ;
  assign \g239726/u3_syn_4  = n39165 ;
  assign \g239734/u3_syn_4  = n39166 ;
  assign \g239735/u3_syn_4  = n39167 ;
  assign \g239743/u3_syn_4  = n39168 ;
  assign \g239760/u3_syn_4  = n39169 ;
  assign \g239768/u3_syn_4  = n39170 ;
  assign \g239776/u3_syn_4  = n39171 ;
  assign \g239784/u3_syn_4  = n39172 ;
  assign \g239793/u3_syn_4  = n39173 ;
  assign \g239801/u3_syn_4  = n39174 ;
  assign \g239817/u3_syn_4  = n39175 ;
  assign \g239818/u3_syn_4  = n39176 ;
  assign \g239848/u3_syn_4  = n39177 ;
  assign \g239856/u3_syn_4  = n39178 ;
  assign \g239872/u3_syn_4  = n39179 ;
  assign \g239880/u3_syn_4  = n39180 ;
  assign \g239888/u3_syn_4  = n39181 ;
  assign \g239896/u3_syn_4  = n39182 ;
  assign \g239904/u3_syn_4  = n39183 ;
  assign \g239912/u3_syn_4  = n39184 ;
  assign \g239920/u3_syn_4  = n39185 ;
  assign \g239928/u3_syn_4  = n39186 ;
  assign \g239936/u3_syn_4  = n39187 ;
  assign \g239951/u3_syn_4  = n39188 ;
  assign \g239963/u3_syn_4  = n39189 ;
  assign \g239979/u3_syn_4  = n39190 ;
  assign \g239986/u3_syn_4  = n39191 ;
  assign \g239999/u3_syn_4  = n39192 ;
  assign \g240000/u3_syn_4  = n39193 ;
  assign \g240008/u3_syn_4  = n39194 ;
  assign \g240012/u3_syn_4  = n39195 ;
  assign \g240018/u3_syn_4  = n39196 ;
  assign \g240026/u3_syn_4  = n39197 ;
  assign \g240034/u3_syn_4  = n39198 ;
  assign \g240042/u3_syn_4  = n39199 ;
  assign \g240050/u3_syn_4  = n39200 ;
  assign \g240074/u3_syn_4  = n39201 ;
  assign \g240091/u3_syn_4  = n39202 ;
  assign \g240122/u3_syn_4  = n39203 ;
  assign \g240147/u3_syn_4  = n39204 ;
  assign \g240209/u3_syn_4  = n39205 ;
  assign \g240219/u3_syn_4  = n39206 ;
  assign \g240259/u3_syn_4  = n39207 ;
  assign \g240334/u3_syn_4  = n39208 ;
  assign \g240406/u3_syn_4  = n39209 ;
  assign \g240416/u3_syn_4  = n39210 ;
  assign \g240424/u3_syn_4  = n39211 ;
  assign \g240432/u3_syn_4  = n39212 ;
  assign \g240440/u3_syn_4  = n39213 ;
  assign \g240448/u3_syn_4  = n39214 ;
  assign \g240456/u3_syn_4  = n39215 ;
  assign \g240464/u3_syn_4  = n39216 ;
  assign \g240472/u3_syn_4  = n39217 ;
  assign \g240480/u3_syn_4  = n39218 ;
  assign \g240488/u3_syn_4  = n39219 ;
  assign \g240496/u3_syn_4  = n39220 ;
  assign \g240504/u3_syn_4  = n39221 ;
  assign \g240512/u3_syn_4  = n39222 ;
  assign \g240520/u3_syn_4  = n39223 ;
  assign \g240530/u3_syn_4  = n39224 ;
  assign \g240538/u3_syn_4  = n39225 ;
  assign \g240547/u3_syn_4  = n39226 ;
  assign \g240555/u3_syn_4  = n39227 ;
  assign \g240563/u3_syn_4  = n39228 ;
  assign \g240571/u3_syn_4  = n39229 ;
  assign \g240579/u3_syn_4  = n39230 ;
  assign \g240587/u3_syn_4  = n39231 ;
  assign \g240595/u3_syn_4  = n39232 ;
  assign \g240603/u3_syn_4  = n39233 ;
  assign \g240611/u3_syn_4  = n39234 ;
  assign \g240619/u3_syn_4  = n39235 ;
  assign \g240627/u3_syn_4  = n39236 ;
  assign \g240635/u3_syn_4  = n39237 ;
  assign \g240643/u3_syn_4  = n39238 ;
  assign \g240651/u3_syn_4  = n39239 ;
  assign \g240659/u3_syn_4  = n39240 ;
  assign \g240667/u3_syn_4  = n39241 ;
  assign \g240675/u3_syn_4  = n39242 ;
  assign \g240683/u3_syn_4  = n39243 ;
  assign \g240691/u3_syn_4  = n39244 ;
  assign \g240699/u3_syn_4  = n39245 ;
  assign \g240707/u3_syn_4  = n39246 ;
  assign \g240715/u3_syn_4  = n39247 ;
  assign \g240723/u3_syn_4  = n39248 ;
  assign \g240731/u3_syn_4  = n39249 ;
  assign \g240739/u3_syn_4  = n39250 ;
  assign \g240747/u3_syn_4  = n39251 ;
  assign \g240755/u3_syn_4  = n39252 ;
  assign \g240763/u3_syn_4  = n39253 ;
  assign \g240771/u3_syn_4  = n39254 ;
  assign \g240779/u3_syn_4  = n39255 ;
  assign \g240787/u3_syn_4  = n39256 ;
  assign \g240795/u3_syn_4  = n39257 ;
  assign \g240803/u3_syn_4  = n39258 ;
  assign \g240811/u3_syn_4  = n39259 ;
  assign \g240819/u3_syn_4  = n39260 ;
  assign \g240827/u3_syn_4  = n39261 ;
  assign \g240835/u3_syn_4  = n39262 ;
  assign \g240843/u3_syn_4  = n39263 ;
  assign \g240851/u3_syn_4  = n39264 ;
  assign \g240859/u3_syn_4  = n39265 ;
  assign \g240867/u3_syn_4  = n39266 ;
  assign \g240875/u3_syn_4  = n39267 ;
  assign \g240883/u3_syn_4  = n39268 ;
  assign \g240891/u3_syn_4  = n39269 ;
  assign \g240899/u3_syn_4  = n39270 ;
  assign \g240907/u3_syn_4  = n39271 ;
  assign \g240915/u3_syn_4  = n39272 ;
  assign \g240923/u3_syn_4  = n39273 ;
  assign \g240931/u3_syn_4  = n39274 ;
  assign \g240939/u3_syn_4  = n39275 ;
  assign \g240947/u3_syn_4  = n39276 ;
  assign \g240955/u3_syn_4  = n39277 ;
  assign \g240963/u3_syn_4  = n39278 ;
  assign \g240971/u3_syn_4  = n39279 ;
  assign \g240979/u3_syn_4  = n39280 ;
  assign \g240987/u3_syn_4  = n39281 ;
  assign \g240995/u3_syn_4  = n39282 ;
  assign \g241003/u3_syn_4  = n39283 ;
  assign \g241011/u3_syn_4  = n39284 ;
  assign \g241019/u3_syn_4  = n39285 ;
  assign \g241027/u3_syn_4  = n39286 ;
  assign \g241036/u3_syn_4  = n39287 ;
  assign \g241044/u3_syn_4  = n39288 ;
  assign \g241052/u3_syn_4  = n39289 ;
  assign \g241060/u3_syn_4  = n39290 ;
  assign \g241068/u3_syn_4  = n39291 ;
  assign \g241076/u3_syn_4  = n39292 ;
  assign \g241084/u3_syn_4  = n39293 ;
  assign \g241092/u3_syn_4  = n39294 ;
  assign \g241100/u3_syn_4  = n39295 ;
  assign \g241108/u3_syn_4  = n39296 ;
  assign \g241116/u3_syn_4  = n39297 ;
  assign \g241124/u3_syn_4  = n39298 ;
  assign \g241132/u3_syn_4  = n39299 ;
  assign \g241140/u3_syn_4  = n39300 ;
  assign \g241148/u3_syn_4  = n39301 ;
  assign \g241156/u3_syn_4  = n39302 ;
  assign \g241164/u3_syn_4  = n39303 ;
  assign \g241172/u3_syn_4  = n39304 ;
  assign \g241180/u3_syn_4  = n39305 ;
  assign \g241188/u3_syn_4  = n39306 ;
  assign \g241196/u3_syn_4  = n39307 ;
  assign \g241205/u3_syn_4  = n39308 ;
  assign \g241213/u3_syn_4  = n39309 ;
  assign \g241221/u3_syn_4  = n39310 ;
  assign \g241229/u3_syn_4  = n39311 ;
  assign \g241237/u3_syn_4  = n39312 ;
  assign \g241245/u3_syn_4  = n39313 ;
  assign \g241253/u3_syn_4  = n39314 ;
  assign \g241261/u3_syn_4  = n39315 ;
  assign \g241269/u3_syn_4  = n39316 ;
  assign \g241277/u3_syn_4  = n39317 ;
  assign \g241285/u3_syn_4  = n39318 ;
  assign \g241293/u3_syn_4  = n39319 ;
  assign \g241301/u3_syn_4  = n39320 ;
  assign \g241309/u3_syn_4  = n39321 ;
  assign \g241317/u3_syn_4  = n39322 ;
  assign \g241325/u3_syn_4  = n39323 ;
  assign \g241333/u3_syn_4  = n39324 ;
  assign \g241341/u3_syn_4  = n39325 ;
  assign \g241349/u3_syn_4  = n39326 ;
  assign \g241358/u3_syn_4  = n39327 ;
  assign \g241366/u3_syn_4  = n39328 ;
  assign \g241374/u3_syn_4  = n39329 ;
  assign \g241382/u3_syn_4  = n39330 ;
  assign \g241390/u3_syn_4  = n39331 ;
  assign \g241398/u3_syn_4  = n39332 ;
  assign \g241406/u3_syn_4  = n39333 ;
  assign \g241415/u3_syn_4  = n39334 ;
  assign \g241424/u3_syn_4  = n39335 ;
  assign \g241433/u3_syn_4  = n39336 ;
  assign \g241441/u3_syn_4  = n39337 ;
  assign \g241449/u3_syn_4  = n39338 ;
  assign \g241459/u3_syn_4  = n39339 ;
  assign \g241470/u3_syn_4  = n39340 ;
  assign \g241480/u3_syn_4  = n39341 ;
  assign \g241489/u3_syn_4  = n39342 ;
  assign \g241497/u3_syn_4  = n39343 ;
  assign \g241505/u3_syn_4  = n39344 ;
  assign \g241513/u3_syn_4  = n39345 ;
  assign \g241545/_3_  = n39346 ;
  assign \g241580/_00_  = ~n39351 ;
  assign \g241737/_0_  = n39353 ;
  assign \g241752/_0_  = n39355 ;
  assign \g241755/_0_  = n39356 ;
  assign \g241767/_2__syn_2  = ~n39358 ;
  assign \g241781/_1__syn_2  = n39359 ;
  assign \g241782/_0_  = n39360 ;
  assign \g241803/_1__syn_2  = n39361 ;
  assign \g241805/_0_  = n39362 ;
  assign \g241812/_1__syn_2  = n39363 ;
  assign \g241814/_1__syn_2  = n39364 ;
  assign \g241816/_1__syn_2  = n39365 ;
  assign \g241819/_1__syn_2  = n39366 ;
  assign \g241822/_1__syn_2  = n39367 ;
  assign \g241823/_0_  = n39368 ;
  assign \g241833/_1__syn_2  = n39369 ;
  assign \g241843/_1__syn_2  = n39371 ;
  assign \g241844/_1__syn_2  = n39372 ;
  assign \g241848/_1__syn_2  = n39374 ;
  assign \g241855/_1__syn_2  = n39375 ;
  assign \g241868/_1__syn_2  = n39376 ;
  assign \g242013/_1__syn_2  = n39377 ;
  assign \g242015/_1__syn_2  = n39379 ;
  assign \g242017/_1__syn_2  = n39380 ;
  assign \g242021/_1__syn_2  = n39381 ;
  assign \g242039/_1__syn_2  = n39382 ;
  assign \g242081/_0_  = ~n39388 ;
  assign \g242086/_0_  = n39389 ;
  assign \g242101/_3_  = n11977 ;
  assign \g242116/_0_  = n39396 ;
  assign \g242135/_2_  = n33021 ;
  assign \g242147/_0_  = ~n39402 ;
  assign \g242158/_0_  = ~n39407 ;
  assign \g242196/_0_  = ~n39413 ;
  assign \g242202/_0_  = ~n39444 ;
  assign \g242203/_0_  = ~n39475 ;
  assign \g242204/_0_  = ~n39506 ;
  assign \g242212/_0_  = n39509 ;
  assign \g242226/_01_  = n39537 ;
  assign \g242281/_0_  = n39538 ;
  assign \g242407/_0_  = ~n39544 ;
  assign \g242410/_0_  = ~n39549 ;
  assign \g242426/_0_  = n39561 ;
  assign \g242438/_2_  = n39563 ;
  assign \g242466/_0_  = n39566 ;
  assign \g242530/_0_  = n39574 ;
  assign \g242532/_0_  = ~n39577 ;
  assign \g243397/_0_  = ~n39585 ;
  assign \g245925/_0_  = ~n39591 ;
  assign \g245932/_0_  = n39597 ;
  assign \g245933/_0_  = ~n39604 ;
  assign \g245986/_3_  = n39613 ;
  assign \g250157/_3_  = n39614 ;
  assign \g250202/_0_  = ~n39620 ;
  assign \g250246/_1_  = n39621 ;
  assign \g250248/_0_  = n39627 ;
  assign \g250250/_0_  = n39628 ;
  assign \g250305/_0_  = n39631 ;
  assign \g250323/_0_  = n39635 ;
  assign \g250373/_0_  = n39639 ;
  assign \g250377/_0_  = n39640 ;
  assign \g250412/_0_  = n39647 ;
  assign \g250413/_0_  = ~n39650 ;
  assign \g250418/_0_  = ~n39654 ;
  assign \g250419/_0_  = ~n39658 ;
  assign \g250421/_0_  = n39661 ;
  assign \g250433/_0_  = ~n39669 ;
  assign \g250448/_3_  = ~n39673 ;
  assign \g250567/_3_  = n11760 ;
  assign \g258965/_0_  = n39676 ;
  assign \g259006/_0_  = ~n39681 ;
  assign \g259471/_0_  = ~n39686 ;
  assign \g259473/_2_  = n39687 ;
  assign \g260557/_0_  = n39688 ;
  assign \g261035/_0_  = n39689 ;
  assign \g261095/_3_  = ~n39695 ;
  assign \g261207/_2__syn_2  = n39697 ;
  assign \g261754/_0_  = n39698 ;
  assign \g262017/_0_  = ~n39703 ;
  assign \g262045/_0_  = n39708 ;
  assign \g262046/_0_  = n39711 ;
  assign \g262100/_3_  = ~n39714 ;
  assign \g263539/_1_  = n15780 ;
  assign \g263574/_0_  = n14046 ;
  assign \g263858/_0_  = ~n11203 ;
  assign \g264104/_1_  = n39609 ;
  assign \g264107/_1_  = n38000 ;
  assign \g264117/_0_  = n39716 ;
  assign \g264282/_0_  = n39576 ;
  assign \g264511/_0_  = ~n39718 ;
  assign \g264541/_0_  = n39722 ;
  assign \g264562/_0_  = n39725 ;
  assign \g264618/_0_  = n39727 ;
  assign \g264660/_0_  = ~n39729 ;
  assign \g264681/_3_  = ~n39732 ;
  assign \g264727/_0_  = ~n39734 ;
  assign \g265013/_0_  = n39736 ;
  assign \g265084/_0_  = ~n39738 ;
  assign \g265378/_0_  = n39740 ;
  assign \g265413/_0_  = ~n39742 ;
  assign \g265446/_0_  = n39744 ;
  assign \g265486/_0_  = ~n39747 ;
  assign \g265524/_3_  = ~n10671 ;
  assign \g265528/_3_  = ~n11356 ;
  assign \g265548/_3_  = ~n10657 ;
  assign \g265579/_0_  = n11754 ;
  assign \g265768/_0_  = n39638 ;
  assign \g265801/_0_  = n12725 ;
  assign \g265819/_1_  = n35444 ;
  assign \g265853/_0_  = n39739 ;
  assign \g265933/_0_  = ~n39748 ;
  assign \g266022/_0_  = n39749 ;
  assign \g266183/_1_  = n36399 ;
  assign \g281909/_0_  = ~n39783 ;
  assign \g281965/_1_  = n39784 ;
  assign \g282284/_1_  = n39785 ;
  assign \g282639/_1_  = n39786 ;
  assign \g283047/_0_  = ~n39792 ;
  assign \g283157/_1_  = n39793 ;
  assign \g283184/_0_  = ~n39822 ;
  assign \g283334/_3_  = ~n39827 ;
  assign int_o_pad = ~n39840 ;
  assign \m_wb_adr_o[0]_pad  = 1'b0 ;
  assign \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2  = ~\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  ;
  assign \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3  = ~n39844 ;
  assign \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3  = ~n39848 ;
  assign \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3  = ~n39852 ;
  assign \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3  = ~n39856 ;
  assign \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3  = ~n39860 ;
  assign \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3  = ~n39864 ;
  assign \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3  = ~n39868 ;
endmodule
