module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G1_pad , \G22_reg/NET0131 , \G23_reg/NET0131 , \G24_reg/NET0131 , \G25_reg/NET0131 , \G26_reg/NET0131 , \G27_reg/NET0131 , \G28_reg/NET0131 , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \G31_reg/NET0131 , \G32_reg/NET0131 , \G33_reg/NET0131 , \G34_reg/NET0131 , \G35_reg/NET0131 , \G36_reg/NET0131 , \G37_reg/NET0131 , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G43_reg/NET0131 , \G44_reg/NET0131 , \G45_reg/NET0131 , \G46_reg/NET0131 , \G47_reg/NET0131 , \G48_reg/NET0131 , \G49_reg/NET0131 , \G4_pad , \G50_reg/NET0131 , \G51_reg/NET0131 , \G52_reg/NET0131 , \G53_reg/NET0131 , \G55_reg/NET0131 , \G56_reg/NET0131 , \G57_reg/NET0131 , \G58_reg/NET0131 , \G59_reg/NET0131 , \G5_pad , \G60_reg/NET0131 , \G61_reg/NET0131 , \G62_reg/NET0131 , \G63_reg/NET0131 , \G64_reg/NET0131 , \G65_reg/NET0131 , \G66_reg/NET0131 , \G67_reg/NET0131 , \G68_reg/NET0131 , \G69_reg/NET0131 , \G6_pad , \G70_reg/NET0131 , \G71_reg/NET0131 , \G72_reg/NET0131 , \G73_reg/NET0131 , \G74_reg/NET0131 , \G75_reg/NET0131 , \G76_reg/NET0131 , \G77_reg/NET0131 , \G78_reg/NET0131 , \G79_reg/NET0131 , \G7_pad , \G80_reg/NET0131 , \G81_reg/NET0131 , \G82_reg/NET0131 , \G83_reg/NET0131 , \G84_reg/NET0131 , \G85_reg/NET0131 , \G86_reg/NET0131 , \G87_reg/NET0131 , \G88_reg/NET0131 , \G89_reg/NET0131 , \G8_pad , \G90_reg/NET0131 , \G91_reg/NET0131 , \G92_reg/NET0131 , \G94_reg/NET0131 , \G9_pad , \G701BF_pad , \G702_pad , \G727_pad , \_al_n0 , \_al_n1 , \g2503/_0_ , \g2514/_0_ , \g2516/_0_ , \g2542/_0_ , \g2549/_0_ , \g2553/_0_ , \g2554/_0_ , \g2570/_0_ , \g2574/_0_ , \g2576/_0_ , \g2583/_0_ , \g2588/_0_ , \g2602/_0_ , \g2603/_0_ , \g2604/_0_ , \g2605/_0_ , \g2611/_0_ , \g2614/_0_ , \g2615/_0_ , \g2644/_0_ , \g2657/_0_ , \g2663/_0_ , \g2664/_0_ , \g2666/_0_ , \g2672/_0_ , \g2678/_0_ , \g2681/_0_ , \g2696/_00_ , \g2698/_0_ , \g2699/_0_ , \g2700/_00_ , \g2717/_0_ , \g2719/_0_ , \g2723/_0_ , \g2726/_3_ , \g2735/_0_ , \g2737/_0_ , \g2740/_0_ , \g2785/_0_ , \g2786/_0_ , \g2787/_1__syn_2 , \g2790/_1__syn_2 , \g2798/_2_ , \g2801/_0_ , \g2841/_0_ , \g2844/_0_ , \g2845/_0_ , \g2846/_0_ , \g2860/_0_ , \g2861/_0_ , \g2862/_0_ , \g2864/_0_ , \g2882/_3_ , \g2883/_3_ , \g2887/_3_ , \g2906/_0_ , \g2911/_0_ , \g3282/_0_ , \g3406/_0_ , \g3409/_0_ , \g3506/_0_ , \g3685/_3_ , \g3694/_0_ , \g3743/_0_ , \g3753/_0_ , \g3785/_0_ , \g3835/_0_ , \g3946/_2_ , \g3976/_0_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G1_pad  ;
	input \G22_reg/NET0131  ;
	input \G23_reg/NET0131  ;
	input \G24_reg/NET0131  ;
	input \G25_reg/NET0131  ;
	input \G26_reg/NET0131  ;
	input \G27_reg/NET0131  ;
	input \G28_reg/NET0131  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	input \G31_reg/NET0131  ;
	input \G32_reg/NET0131  ;
	input \G33_reg/NET0131  ;
	input \G34_reg/NET0131  ;
	input \G35_reg/NET0131  ;
	input \G36_reg/NET0131  ;
	input \G37_reg/NET0131  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G43_reg/NET0131  ;
	input \G44_reg/NET0131  ;
	input \G45_reg/NET0131  ;
	input \G46_reg/NET0131  ;
	input \G47_reg/NET0131  ;
	input \G48_reg/NET0131  ;
	input \G49_reg/NET0131  ;
	input \G4_pad  ;
	input \G50_reg/NET0131  ;
	input \G51_reg/NET0131  ;
	input \G52_reg/NET0131  ;
	input \G53_reg/NET0131  ;
	input \G55_reg/NET0131  ;
	input \G56_reg/NET0131  ;
	input \G57_reg/NET0131  ;
	input \G58_reg/NET0131  ;
	input \G59_reg/NET0131  ;
	input \G5_pad  ;
	input \G60_reg/NET0131  ;
	input \G61_reg/NET0131  ;
	input \G62_reg/NET0131  ;
	input \G63_reg/NET0131  ;
	input \G64_reg/NET0131  ;
	input \G65_reg/NET0131  ;
	input \G66_reg/NET0131  ;
	input \G67_reg/NET0131  ;
	input \G68_reg/NET0131  ;
	input \G69_reg/NET0131  ;
	input \G6_pad  ;
	input \G70_reg/NET0131  ;
	input \G71_reg/NET0131  ;
	input \G72_reg/NET0131  ;
	input \G73_reg/NET0131  ;
	input \G74_reg/NET0131  ;
	input \G75_reg/NET0131  ;
	input \G76_reg/NET0131  ;
	input \G77_reg/NET0131  ;
	input \G78_reg/NET0131  ;
	input \G79_reg/NET0131  ;
	input \G7_pad  ;
	input \G80_reg/NET0131  ;
	input \G81_reg/NET0131  ;
	input \G82_reg/NET0131  ;
	input \G83_reg/NET0131  ;
	input \G84_reg/NET0131  ;
	input \G85_reg/NET0131  ;
	input \G86_reg/NET0131  ;
	input \G87_reg/NET0131  ;
	input \G88_reg/NET0131  ;
	input \G89_reg/NET0131  ;
	input \G8_pad  ;
	input \G90_reg/NET0131  ;
	input \G91_reg/NET0131  ;
	input \G92_reg/NET0131  ;
	input \G94_reg/NET0131  ;
	input \G9_pad  ;
	output \G701BF_pad  ;
	output \G702_pad  ;
	output \G727_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g2503/_0_  ;
	output \g2514/_0_  ;
	output \g2516/_0_  ;
	output \g2542/_0_  ;
	output \g2549/_0_  ;
	output \g2553/_0_  ;
	output \g2554/_0_  ;
	output \g2570/_0_  ;
	output \g2574/_0_  ;
	output \g2576/_0_  ;
	output \g2583/_0_  ;
	output \g2588/_0_  ;
	output \g2602/_0_  ;
	output \g2603/_0_  ;
	output \g2604/_0_  ;
	output \g2605/_0_  ;
	output \g2611/_0_  ;
	output \g2614/_0_  ;
	output \g2615/_0_  ;
	output \g2644/_0_  ;
	output \g2657/_0_  ;
	output \g2663/_0_  ;
	output \g2664/_0_  ;
	output \g2666/_0_  ;
	output \g2672/_0_  ;
	output \g2678/_0_  ;
	output \g2681/_0_  ;
	output \g2696/_00_  ;
	output \g2698/_0_  ;
	output \g2699/_0_  ;
	output \g2700/_00_  ;
	output \g2717/_0_  ;
	output \g2719/_0_  ;
	output \g2723/_0_  ;
	output \g2726/_3_  ;
	output \g2735/_0_  ;
	output \g2737/_0_  ;
	output \g2740/_0_  ;
	output \g2785/_0_  ;
	output \g2786/_0_  ;
	output \g2787/_1__syn_2  ;
	output \g2790/_1__syn_2  ;
	output \g2798/_2_  ;
	output \g2801/_0_  ;
	output \g2841/_0_  ;
	output \g2844/_0_  ;
	output \g2845/_0_  ;
	output \g2846/_0_  ;
	output \g2860/_0_  ;
	output \g2861/_0_  ;
	output \g2862/_0_  ;
	output \g2864/_0_  ;
	output \g2882/_3_  ;
	output \g2883/_3_  ;
	output \g2887/_3_  ;
	output \g2906/_0_  ;
	output \g2911/_0_  ;
	output \g3282/_0_  ;
	output \g3406/_0_  ;
	output \g3409/_0_  ;
	output \g3506/_0_  ;
	output \g3685/_3_  ;
	output \g3694/_0_  ;
	output \g3743/_0_  ;
	output \g3753/_0_  ;
	output \g3785/_0_  ;
	output \g3835/_0_  ;
	output \g3946/_2_  ;
	output \g3976/_0_  ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\G4_pad ,
		\G90_reg/NET0131 ,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\G64_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\G8_pad ,
		\G90_reg/NET0131 ,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w90_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\G84_reg/NET0131 ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\G85_reg/NET0131 ,
		_w92_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\G78_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w95_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w89_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\G46_reg/NET0131 ,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\G3_pad ,
		\G90_reg/NET0131 ,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\G77_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w95_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w100_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\G45_reg/NET0131 ,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\G2_pad ,
		\G90_reg/NET0131 ,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\G76_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w95_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w105_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\G44_reg/NET0131 ,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\G45_reg/NET0131 ,
		_w103_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w109_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\G0_pad ,
		\G90_reg/NET0131 ,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\G74_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w95_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w112_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\G42_reg/NET0131 ,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\G1_pad ,
		\G90_reg/NET0131 ,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\G75_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w95_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w117_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\G43_reg/NET0131 ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w116_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\G44_reg/NET0131 ,
		_w108_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\G43_reg/NET0131 ,
		_w120_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		_w122_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		_w111_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w104_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\G46_reg/NET0131 ,
		_w98_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w99_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\G24_reg/NET0131 ,
		\G25_reg/NET0131 ,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\G26_reg/NET0131 ,
		\G27_reg/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\G28_reg/NET0131 ,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w131_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\G94_reg/NET0131 ,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\G32_reg/NET0131 ,
		\G33_reg/NET0131 ,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\G29_reg/NET0131 ,
		\G30_reg/NET0131 ,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\G31_reg/NET0131 ,
		\G34_reg/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w138_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w139_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w136_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\G92_reg/NET0131 ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\G75_reg/NET0131 ,
		\G80_reg/NET0131 ,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\G75_reg/NET0131 ,
		\G80_reg/NET0131 ,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\G79_reg/NET0131 ,
		\G80_reg/NET0131 ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\G81_reg/NET0131 ,
		\G82_reg/NET0131 ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		\G78_reg/NET0131 ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\G78_reg/NET0131 ,
		_w150_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\G77_reg/NET0131 ,
		\G82_reg/NET0131 ,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\G77_reg/NET0131 ,
		\G82_reg/NET0131 ,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\G74_reg/NET0131 ,
		\G79_reg/NET0131 ,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		\G74_reg/NET0131 ,
		\G79_reg/NET0131 ,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\G76_reg/NET0131 ,
		\G81_reg/NET0131 ,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\G76_reg/NET0131 ,
		\G81_reg/NET0131 ,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w158_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w154_,
		_w155_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w156_,
		_w157_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w161_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w147_,
		_w160_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w153_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\G16_pad ,
		\G66_reg/NET0131 ,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\G83_reg/NET0131 ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w166_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\G90_reg/NET0131 ,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w144_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\G58_reg/NET0131 ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\G91_reg/NET0131 ,
		_w144_,
		_w173_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\G36_reg/NET0131 ,
		\G37_reg/NET0131 ,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\G38_reg/NET0131 ,
		_w170_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w174_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\G41_reg/NET0131 ,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		\G91_reg/NET0131 ,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\G58_reg/NET0131 ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w176_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w173_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w172_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\G59_reg/NET0131 ,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\G91_reg/NET0131 ,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\G53_reg/NET0131 ,
		\G61_reg/NET0131 ,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\G62_reg/NET0131 ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w185_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\G89_reg/NET0131 ,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w144_,
		_w178_,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\G88_reg/NET0131 ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\G92_reg/NET0131 ,
		_w136_,
		_w192_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		_w142_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\G87_reg/NET0131 ,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\G90_reg/NET0131 ,
		_w137_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w191_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w189_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\G68_reg/NET0131 ,
		\G72_reg/NET0131 ,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\G71_reg/NET0131 ,
		\G72_reg/NET0131 ,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		\G73_reg/NET0131 ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		\G70_reg/NET0131 ,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\G70_reg/NET0131 ,
		_w201_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\G67_reg/NET0131 ,
		\G71_reg/NET0131 ,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\G69_reg/NET0131 ,
		\G73_reg/NET0131 ,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		\G69_reg/NET0131 ,
		\G73_reg/NET0131 ,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\G67_reg/NET0131 ,
		\G71_reg/NET0131 ,
		_w207_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\G68_reg/NET0131 ,
		\G72_reg/NET0131 ,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w199_,
		_w204_,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w205_,
		_w206_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w207_,
		_w208_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w209_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w202_,
		_w203_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w213_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\G14_pad ,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		\G90_reg/NET0131 ,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w185_,
		_w186_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\G62_reg/NET0131 ,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\G14_pad ,
		_w188_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w219_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\G51_reg/NET0131 ,
		_w185_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		\G53_reg/NET0131 ,
		_w185_,
		_w223_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		\G14_pad ,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		\G51_reg/NET0131 ,
		_w185_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w222_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w224_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		\G52_reg/NET0131 ,
		_w222_,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\G52_reg/NET0131 ,
		_w222_,
		_w229_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		_w224_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w228_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\G90_reg/NET0131 ,
		\G9_pad ,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\G90_reg/NET0131 ,
		_w216_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\G91_reg/NET0131 ,
		_w190_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		_w174_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\G38_reg/NET0131 ,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h2)
	) name149 (
		_w170_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		_w139_,
		_w192_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\G31_reg/NET0131 ,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\G34_reg/NET0131 ,
		_w138_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		\G92_reg/NET0131 ,
		_w170_,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w242_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w166_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		_w238_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		\G74_reg/NET0131 ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\G74_reg/NET0131 ,
		_w246_,
		_w248_
	);
	LUT2 #(
		.INIT('h2)
	) name160 (
		_w234_,
		_w247_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w248_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\G14_pad ,
		_w183_,
		_w251_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		_w176_,
		_w235_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w171_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		\G57_reg/NET0131 ,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\G58_reg/NET0131 ,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\G58_reg/NET0131 ,
		_w254_,
		_w256_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		_w251_,
		_w255_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		\G57_reg/NET0131 ,
		_w253_,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		_w251_,
		_w254_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		_w259_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\G59_reg/NET0131 ,
		_w183_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name174 (
		\G14_pad ,
		_w184_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w262_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\G38_reg/NET0131 ,
		_w236_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w237_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		\G14_pad ,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\G36_reg/NET0131 ,
		_w235_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\G37_reg/NET0131 ,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\G14_pad ,
		_w236_,
		_w270_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		\G36_reg/NET0131 ,
		_w235_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w268_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\G14_pad ,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\G39_reg/NET0131 ,
		_w144_,
		_w275_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		\G40_reg/NET0131 ,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\G41_reg/NET0131 ,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\G14_pad ,
		_w190_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\G40_reg/NET0131 ,
		_w275_,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w276_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\G14_pad ,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		\G39_reg/NET0131 ,
		_w144_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\G56_reg/NET0131 ,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		\G91_reg/NET0131 ,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\G12_pad ,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		\G47_reg/NET0131 ,
		_w285_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		\G14_pad ,
		_w286_,
		_w288_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\G48_reg/NET0131 ,
		_w285_,
		_w290_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		\G49_reg/NET0131 ,
		_w285_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\G14_pad ,
		_w290_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w291_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		\G47_reg/NET0131 ,
		_w285_,
		_w294_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		\G48_reg/NET0131 ,
		_w285_,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		\G14_pad ,
		_w294_,
		_w296_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\G49_reg/NET0131 ,
		_w285_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		\G50_reg/NET0131 ,
		_w285_,
		_w299_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\G14_pad ,
		_w298_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\G55_reg/NET0131 ,
		_w283_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\G56_reg/NET0131 ,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		\G14_pad ,
		_w284_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		_w303_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		\G55_reg/NET0131 ,
		_w283_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w302_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w304_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\G39_reg/NET0131 ,
		_w144_,
		_w309_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\G14_pad ,
		_w283_,
		_w310_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w309_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\G32_reg/NET0131 ,
		_w240_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\G33_reg/NET0131 ,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		\G34_reg/NET0131 ,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		_w193_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		\G14_pad ,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\G33_reg/NET0131 ,
		_w312_,
		_w317_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\G14_pad ,
		_w313_,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		\G29_reg/NET0131 ,
		_w192_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		\G30_reg/NET0131 ,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		\G14_pad ,
		_w239_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		_w321_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		\G32_reg/NET0131 ,
		_w240_,
		_w324_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\G14_pad ,
		_w312_,
		_w325_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\G29_reg/NET0131 ,
		_w192_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w320_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\G14_pad ,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\G31_reg/NET0131 ,
		_w239_,
		_w330_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\G14_pad ,
		_w240_,
		_w331_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w131_,
		_w134_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\G28_reg/NET0131 ,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\G14_pad ,
		_w136_,
		_w335_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w334_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\G24_reg/NET0131 ,
		_w131_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\G25_reg/NET0131 ,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		\G26_reg/NET0131 ,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\G27_reg/NET0131 ,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w333_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		\G14_pad ,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		\G25_reg/NET0131 ,
		_w337_,
		_w343_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		\G14_pad ,
		_w338_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		\G26_reg/NET0131 ,
		_w338_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name258 (
		\G14_pad ,
		_w339_,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\G24_reg/NET0131 ,
		_w131_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w337_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		\G14_pad ,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		\G6_pad ,
		\G90_reg/NET0131 ,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w170_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		\G59_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\G62_reg/NET0131 ,
		\G91_reg/NET0131 ,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		\G90_reg/NET0131 ,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\G35_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w357_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w353_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		\G5_pad ,
		\G90_reg/NET0131 ,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		\G83_reg/NET0131 ,
		\G90_reg/NET0131 ,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w166_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w361_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		\G42_reg/NET0131 ,
		_w115_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w99_,
		_w104_,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w129_,
		_w365_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w366_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w111_,
		_w122_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w125_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w368_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w364_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		\G35_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		\G34_reg/NET0131 ,
		\G92_reg/NET0131 ,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w373_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		_w170_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w175_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w372_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w131_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w353_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		\G14_pad ,
		_w360_,
		_w381_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		_w380_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		\G7_pad ,
		\G90_reg/NET0131 ,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w233_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		\G15_pad ,
		\G23_reg/NET0131 ,
		_w385_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\G15_pad ,
		\G22_reg/NET0131 ,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w385_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		\G47_reg/NET0131 ,
		\G48_reg/NET0131 ,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		\G49_reg/NET0131 ,
		\G50_reg/NET0131 ,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w388_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w387_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		\G42_reg/NET0131 ,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		\G43_reg/NET0131 ,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		\G44_reg/NET0131 ,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\G45_reg/NET0131 ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		\G46_reg/NET0131 ,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		\G46_reg/NET0131 ,
		_w395_,
		_w397_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		_w384_,
		_w396_,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w397_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		\G63_reg/NET0131 ,
		_w377_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		\G14_pad ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		\G45_reg/NET0131 ,
		_w394_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w395_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		_w384_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		\G14_pad ,
		\G83_reg/NET0131 ,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w95_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w377_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		\G44_reg/NET0131 ,
		_w393_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w394_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w384_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		\G42_reg/NET0131 ,
		_w391_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w392_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w384_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		\G43_reg/NET0131 ,
		_w392_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w393_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w384_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		\G64_reg/NET0131 ,
		_w215_,
		_w417_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		\G63_reg/NET0131 ,
		_w215_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		\G14_pad ,
		_w417_,
		_w419_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		_w418_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		\G66_reg/NET0131 ,
		_w215_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		\G65_reg/NET0131 ,
		_w215_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		\G14_pad ,
		_w421_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		\G14_pad ,
		_w233_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\G91_reg/NET0131 ,
		_w215_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		\G14_pad ,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		\G65_reg/NET0131 ,
		_w215_,
		_w428_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		\G14_pad ,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\G13_pad ,
		\G14_pad ,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		\G10_pad ,
		\G90_reg/NET0131 ,
		_w431_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\G86_reg/NET0131 ,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		_w430_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		_w386_,
		_w390_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		\G15_pad ,
		\G47_reg/NET0131 ,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\G48_reg/NET0131 ,
		\G49_reg/NET0131 ,
		_w436_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		\G50_reg/NET0131 ,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w435_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		\G22_reg/NET0131 ,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w434_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		\G10_pad ,
		\G91_reg/NET0131 ,
		_w441_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\G13_pad ,
		\G86_reg/NET0131 ,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		\G10_pad ,
		\G92_reg/NET0131 ,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w441_,
		_w442_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w443_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		_w430_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		\G10_pad ,
		\G91_reg/NET0131 ,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\G10_pad ,
		\G90_reg/NET0131 ,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w442_,
		_w447_,
		_w449_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w448_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		_w430_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		\G11_pad ,
		\G87_reg/NET0131 ,
		_w452_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\G11_pad ,
		\G94_reg/NET0131 ,
		_w453_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		\G14_pad ,
		_w452_,
		_w454_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w453_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		\G11_pad ,
		\G88_reg/NET0131 ,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		\G11_pad ,
		\G87_reg/NET0131 ,
		_w457_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		\G14_pad ,
		_w456_,
		_w458_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w457_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		\G11_pad ,
		\G89_reg/NET0131 ,
		_w460_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		\G11_pad ,
		\G88_reg/NET0131 ,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\G14_pad ,
		_w460_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w461_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		\G11_pad ,
		\G94_reg/NET0131 ,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		\G11_pad ,
		\G89_reg/NET0131 ,
		_w465_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		\G14_pad ,
		_w464_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		\G4_pad ,
		\G63_reg/NET0131 ,
		_w468_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		\G1_pad ,
		\G63_reg/NET0131 ,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w468_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name382 (
		\G3_pad ,
		\G63_reg/NET0131 ,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\G0_pad ,
		\G63_reg/NET0131 ,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		\G5_pad ,
		\G63_reg/NET0131 ,
		_w474_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		\G2_pad ,
		\G63_reg/NET0131 ,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w474_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\G14_pad ,
		\G35_reg/NET0131 ,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		\G74_reg/NET0131 ,
		\G75_reg/NET0131 ,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		_w245_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		_w238_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\G76_reg/NET0131 ,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		\G77_reg/NET0131 ,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		\G78_reg/NET0131 ,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		\G78_reg/NET0131 ,
		_w482_,
		_w484_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w234_,
		_w483_,
		_w485_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w484_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		\G75_reg/NET0131 ,
		_w247_,
		_w487_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		_w234_,
		_w480_,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name400 (
		_w487_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w166_,
		_w377_,
		_w490_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		\G83_reg/NET0131 ,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w246_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		_w234_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		\G77_reg/NET0131 ,
		_w481_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		_w234_,
		_w482_,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		\G91_reg/NET0131 ,
		_w187_,
		_w497_
	);
	LUT2 #(
		.INIT('h2)
	) name409 (
		_w184_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		\G90_reg/NET0131 ,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		\G67_reg/NET0131 ,
		\G68_reg/NET0131 ,
		_w500_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w499_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\G67_reg/NET0131 ,
		_w499_,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		\G68_reg/NET0131 ,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		_w216_,
		_w501_,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w503_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\G60_reg/NET0131 ,
		_w223_,
		_w506_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\G14_pad ,
		_w218_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		\G60_reg/NET0131 ,
		_w223_,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w506_,
		_w507_,
		_w509_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w508_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\G53_reg/NET0131 ,
		_w230_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		\G14_pad ,
		\G53_reg/NET0131 ,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		_w229_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w511_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		\G61_reg/NET0131 ,
		_w506_,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		_w507_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		\G76_reg/NET0131 ,
		_w480_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		_w234_,
		_w481_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		_w517_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		\G67_reg/NET0131 ,
		_w499_,
		_w520_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		_w216_,
		_w502_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name433 (
		_w520_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\G69_reg/NET0131 ,
		_w501_,
		_w523_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		\G69_reg/NET0131 ,
		_w501_,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		_w216_,
		_w523_,
		_w525_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w524_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		\G70_reg/NET0131 ,
		_w524_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\G70_reg/NET0131 ,
		_w524_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name440 (
		_w216_,
		_w527_,
		_w529_
	);
	LUT2 #(
		.INIT('h4)
	) name441 (
		_w528_,
		_w529_,
		_w530_
	);
	assign \G701BF_pad  = \G15_pad ;
	assign \G702_pad  = _w198_ ;
	assign \G727_pad  = _w217_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g2503/_0_  = _w221_ ;
	assign \g2514/_0_  = _w227_ ;
	assign \g2516/_0_  = _w231_ ;
	assign \g2542/_0_  = _w250_ ;
	assign \g2549/_0_  = _w258_ ;
	assign \g2553/_0_  = _w261_ ;
	assign \g2554/_0_  = _w264_ ;
	assign \g2570/_0_  = _w267_ ;
	assign \g2574/_0_  = _w271_ ;
	assign \g2576/_0_  = _w274_ ;
	assign \g2583/_0_  = _w279_ ;
	assign \g2588/_0_  = _w282_ ;
	assign \g2602/_0_  = _w289_ ;
	assign \g2603/_0_  = _w293_ ;
	assign \g2604/_0_  = _w297_ ;
	assign \g2605/_0_  = _w301_ ;
	assign \g2611/_0_  = _w305_ ;
	assign \g2614/_0_  = _w308_ ;
	assign \g2615/_0_  = _w311_ ;
	assign \g2644/_0_  = _w316_ ;
	assign \g2657/_0_  = _w319_ ;
	assign \g2663/_0_  = _w323_ ;
	assign \g2664/_0_  = _w326_ ;
	assign \g2666/_0_  = _w329_ ;
	assign \g2672/_0_  = _w332_ ;
	assign \g2678/_0_  = _w336_ ;
	assign \g2681/_0_  = _w342_ ;
	assign \g2696/_00_  = _w345_ ;
	assign \g2698/_0_  = _w348_ ;
	assign \g2699/_0_  = _w351_ ;
	assign \g2700/_00_  = _w382_ ;
	assign \g2717/_0_  = _w399_ ;
	assign \g2719/_0_  = _w401_ ;
	assign \g2723/_0_  = _w404_ ;
	assign \g2726/_3_  = _w407_ ;
	assign \g2735/_0_  = _w410_ ;
	assign \g2737/_0_  = _w413_ ;
	assign \g2740/_0_  = _w416_ ;
	assign \g2785/_0_  = _w420_ ;
	assign \g2786/_0_  = _w424_ ;
	assign \g2787/_1__syn_2  = _w425_ ;
	assign \g2790/_1__syn_2  = _w427_ ;
	assign \g2798/_2_  = _w387_ ;
	assign \g2801/_0_  = _w429_ ;
	assign \g2841/_0_  = _w433_ ;
	assign \g2844/_0_  = _w440_ ;
	assign \g2845/_0_  = _w446_ ;
	assign \g2846/_0_  = _w451_ ;
	assign \g2860/_0_  = _w455_ ;
	assign \g2861/_0_  = _w459_ ;
	assign \g2862/_0_  = _w463_ ;
	assign \g2864/_0_  = _w467_ ;
	assign \g2882/_3_  = _w470_ ;
	assign \g2883/_3_  = _w473_ ;
	assign \g2887/_3_  = _w476_ ;
	assign \g2906/_0_  = _w477_ ;
	assign \g2911/_0_  = _w430_ ;
	assign \g3282/_0_  = _w486_ ;
	assign \g3406/_0_  = _w489_ ;
	assign \g3409/_0_  = _w493_ ;
	assign \g3506/_0_  = _w496_ ;
	assign \g3685/_3_  = _w505_ ;
	assign \g3694/_0_  = _w510_ ;
	assign \g3743/_0_  = _w514_ ;
	assign \g3753/_0_  = _w516_ ;
	assign \g3785/_0_  = _w519_ ;
	assign \g3835/_0_  = _w522_ ;
	assign \g3946/_2_  = _w526_ ;
	assign \g3976/_0_  = _w530_ ;
endmodule;