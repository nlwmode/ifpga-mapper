module top( \P1_B_reg/NET0131  , \P1_IR_reg[0]/NET0131  , \P1_IR_reg[10]/NET0131  , \P1_IR_reg[11]/NET0131  , \P1_IR_reg[12]/NET0131  , \P1_IR_reg[13]/NET0131  , \P1_IR_reg[14]/NET0131  , \P1_IR_reg[15]/NET0131  , \P1_IR_reg[16]/NET0131  , \P1_IR_reg[17]/NET0131  , \P1_IR_reg[18]/NET0131  , \P1_IR_reg[19]/NET0131  , \P1_IR_reg[1]/NET0131  , \P1_IR_reg[20]/NET0131  , \P1_IR_reg[21]/NET0131  , \P1_IR_reg[22]/NET0131  , \P1_IR_reg[23]/NET0131  , \P1_IR_reg[24]/NET0131  , \P1_IR_reg[25]/NET0131  , \P1_IR_reg[26]/NET0131  , \P1_IR_reg[27]/NET0131  , \P1_IR_reg[28]/NET0131  , \P1_IR_reg[29]/NET0131  , \P1_IR_reg[2]/NET0131  , \P1_IR_reg[30]/NET0131  , \P1_IR_reg[31]/NET0131  , \P1_IR_reg[3]/NET0131  , \P1_IR_reg[4]/NET0131  , \P1_IR_reg[5]/NET0131  , \P1_IR_reg[6]/NET0131  , \P1_IR_reg[7]/NET0131  , \P1_IR_reg[8]/NET0131  , \P1_IR_reg[9]/NET0131  , \P1_addr_reg[0]/NET0131  , \P1_addr_reg[10]/NET0131  , \P1_addr_reg[11]/NET0131  , \P1_addr_reg[12]/NET0131  , \P1_addr_reg[13]/NET0131  , \P1_addr_reg[14]/NET0131  , \P1_addr_reg[15]/NET0131  , \P1_addr_reg[16]/NET0131  , \P1_addr_reg[17]/NET0131  , \P1_addr_reg[18]/NET0131  , \P1_addr_reg[19]/NET0131  , \P1_addr_reg[1]/NET0131  , \P1_addr_reg[2]/NET0131  , \P1_addr_reg[3]/NET0131  , \P1_addr_reg[4]/NET0131  , \P1_addr_reg[5]/NET0131  , \P1_addr_reg[6]/NET0131  , \P1_addr_reg[7]/NET0131  , \P1_addr_reg[8]/NET0131  , \P1_addr_reg[9]/NET0131  , \P1_d_reg[0]/NET0131  , \P1_d_reg[1]/NET0131  , \P1_datao_reg[0]/NET0131  , \P1_datao_reg[10]/NET0131  , \P1_datao_reg[11]/NET0131  , \P1_datao_reg[12]/NET0131  , \P1_datao_reg[13]/NET0131  , \P1_datao_reg[14]/NET0131  , \P1_datao_reg[15]/NET0131  , \P1_datao_reg[16]/NET0131  , \P1_datao_reg[17]/NET0131  , \P1_datao_reg[18]/NET0131  , \P1_datao_reg[19]/NET0131  , \P1_datao_reg[1]/NET0131  , \P1_datao_reg[20]/NET0131  , \P1_datao_reg[21]/NET0131  , \P1_datao_reg[22]/NET0131  , \P1_datao_reg[23]/NET0131  , \P1_datao_reg[24]/NET0131  , \P1_datao_reg[25]/NET0131  , \P1_datao_reg[26]/NET0131  , \P1_datao_reg[27]/NET0131  , \P1_datao_reg[28]/NET0131  , \P1_datao_reg[29]/NET0131  , \P1_datao_reg[2]/NET0131  , \P1_datao_reg[30]/NET0131  , \P1_datao_reg[31]/NET0131  , \P1_datao_reg[3]/NET0131  , \P1_datao_reg[4]/NET0131  , \P1_datao_reg[5]/NET0131  , \P1_datao_reg[6]/NET0131  , \P1_datao_reg[7]/NET0131  , \P1_datao_reg[8]/NET0131  , \P1_datao_reg[9]/NET0131  , \P1_rd_reg/NET0131  , \P1_reg0_reg[0]/NET0131  , \P1_reg0_reg[10]/NET0131  , \P1_reg0_reg[11]/NET0131  , \P1_reg0_reg[12]/NET0131  , \P1_reg0_reg[13]/NET0131  , \P1_reg0_reg[14]/NET0131  , \P1_reg0_reg[15]/NET0131  , \P1_reg0_reg[16]/NET0131  , \P1_reg0_reg[17]/NET0131  , \P1_reg0_reg[18]/NET0131  , \P1_reg0_reg[19]/NET0131  , \P1_reg0_reg[1]/NET0131  , \P1_reg0_reg[20]/NET0131  , \P1_reg0_reg[21]/NET0131  , \P1_reg0_reg[22]/NET0131  , \P1_reg0_reg[23]/NET0131  , \P1_reg0_reg[24]/NET0131  , \P1_reg0_reg[25]/NET0131  , \P1_reg0_reg[26]/NET0131  , \P1_reg0_reg[27]/NET0131  , \P1_reg0_reg[28]/NET0131  , \P1_reg0_reg[29]/NET0131  , \P1_reg0_reg[2]/NET0131  , \P1_reg0_reg[30]/NET0131  , \P1_reg0_reg[31]/NET0131  , \P1_reg0_reg[3]/NET0131  , \P1_reg0_reg[4]/NET0131  , \P1_reg0_reg[5]/NET0131  , \P1_reg0_reg[6]/NET0131  , \P1_reg0_reg[7]/NET0131  , \P1_reg0_reg[8]/NET0131  , \P1_reg0_reg[9]/NET0131  , \P1_reg1_reg[0]/NET0131  , \P1_reg1_reg[10]/NET0131  , \P1_reg1_reg[11]/NET0131  , \P1_reg1_reg[12]/NET0131  , \P1_reg1_reg[13]/NET0131  , \P1_reg1_reg[14]/NET0131  , \P1_reg1_reg[15]/NET0131  , \P1_reg1_reg[16]/NET0131  , \P1_reg1_reg[17]/NET0131  , \P1_reg1_reg[18]/NET0131  , \P1_reg1_reg[19]/NET0131  , \P1_reg1_reg[1]/NET0131  , \P1_reg1_reg[20]/NET0131  , \P1_reg1_reg[21]/NET0131  , \P1_reg1_reg[22]/NET0131  , \P1_reg1_reg[23]/NET0131  , \P1_reg1_reg[24]/NET0131  , \P1_reg1_reg[25]/NET0131  , \P1_reg1_reg[26]/NET0131  , \P1_reg1_reg[27]/NET0131  , \P1_reg1_reg[28]/NET0131  , \P1_reg1_reg[29]/NET0131  , \P1_reg1_reg[2]/NET0131  , \P1_reg1_reg[30]/NET0131  , \P1_reg1_reg[31]/NET0131  , \P1_reg1_reg[3]/NET0131  , \P1_reg1_reg[4]/NET0131  , \P1_reg1_reg[5]/NET0131  , \P1_reg1_reg[6]/NET0131  , \P1_reg1_reg[7]/NET0131  , \P1_reg1_reg[8]/NET0131  , \P1_reg1_reg[9]/NET0131  , \P1_reg2_reg[0]/NET0131  , \P1_reg2_reg[10]/NET0131  , \P1_reg2_reg[11]/NET0131  , \P1_reg2_reg[12]/NET0131  , \P1_reg2_reg[13]/NET0131  , \P1_reg2_reg[14]/NET0131  , \P1_reg2_reg[15]/NET0131  , \P1_reg2_reg[16]/NET0131  , \P1_reg2_reg[17]/NET0131  , \P1_reg2_reg[18]/NET0131  , \P1_reg2_reg[19]/NET0131  , \P1_reg2_reg[1]/NET0131  , \P1_reg2_reg[20]/NET0131  , \P1_reg2_reg[21]/NET0131  , \P1_reg2_reg[22]/NET0131  , \P1_reg2_reg[23]/NET0131  , \P1_reg2_reg[24]/NET0131  , \P1_reg2_reg[25]/NET0131  , \P1_reg2_reg[26]/NET0131  , \P1_reg2_reg[27]/NET0131  , \P1_reg2_reg[28]/NET0131  , \P1_reg2_reg[29]/NET0131  , \P1_reg2_reg[2]/NET0131  , \P1_reg2_reg[30]/NET0131  , \P1_reg2_reg[31]/NET0131  , \P1_reg2_reg[3]/NET0131  , \P1_reg2_reg[4]/NET0131  , \P1_reg2_reg[5]/NET0131  , \P1_reg2_reg[6]/NET0131  , \P1_reg2_reg[7]/NET0131  , \P1_reg2_reg[8]/NET0131  , \P1_reg2_reg[9]/NET0131  , \P1_reg3_reg[0]/NET0131  , \P1_reg3_reg[10]/NET0131  , \P1_reg3_reg[11]/NET0131  , \P1_reg3_reg[12]/NET0131  , \P1_reg3_reg[13]/NET0131  , \P1_reg3_reg[14]/NET0131  , \P1_reg3_reg[15]/NET0131  , \P1_reg3_reg[16]/NET0131  , \P1_reg3_reg[17]/NET0131  , \P1_reg3_reg[18]/NET0131  , \P1_reg3_reg[19]/NET0131  , \P1_reg3_reg[1]/NET0131  , \P1_reg3_reg[20]/NET0131  , \P1_reg3_reg[21]/NET0131  , \P1_reg3_reg[22]/NET0131  , \P1_reg3_reg[23]/NET0131  , \P1_reg3_reg[24]/NET0131  , \P1_reg3_reg[25]/NET0131  , \P1_reg3_reg[26]/NET0131  , \P1_reg3_reg[27]/NET0131  , \P1_reg3_reg[28]/NET0131  , \P1_reg3_reg[2]/NET0131  , \P1_reg3_reg[3]/NET0131  , \P1_reg3_reg[4]/NET0131  , \P1_reg3_reg[5]/NET0131  , \P1_reg3_reg[6]/NET0131  , \P1_reg3_reg[7]/NET0131  , \P1_reg3_reg[8]/NET0131  , \P1_reg3_reg[9]/NET0131  , \P1_state_reg[0]/NET0131  , \P1_wr_reg/NET0131  , \P2_B_reg/NET0131  , \P2_IR_reg[0]/NET0131  , \P2_IR_reg[10]/NET0131  , \P2_IR_reg[11]/NET0131  , \P2_IR_reg[12]/NET0131  , \P2_IR_reg[13]/NET0131  , \P2_IR_reg[14]/NET0131  , \P2_IR_reg[15]/NET0131  , \P2_IR_reg[16]/NET0131  , \P2_IR_reg[17]/NET0131  , \P2_IR_reg[18]/NET0131  , \P2_IR_reg[19]/NET0131  , \P2_IR_reg[1]/NET0131  , \P2_IR_reg[20]/NET0131  , \P2_IR_reg[21]/NET0131  , \P2_IR_reg[22]/NET0131  , \P2_IR_reg[23]/NET0131  , \P2_IR_reg[24]/NET0131  , \P2_IR_reg[25]/NET0131  , \P2_IR_reg[26]/NET0131  , \P2_IR_reg[27]/NET0131  , \P2_IR_reg[28]/NET0131  , \P2_IR_reg[29]/NET0131  , \P2_IR_reg[2]/NET0131  , \P2_IR_reg[30]/NET0131  , \P2_IR_reg[31]/NET0131  , \P2_IR_reg[3]/NET0131  , \P2_IR_reg[4]/NET0131  , \P2_IR_reg[5]/NET0131  , \P2_IR_reg[6]/NET0131  , \P2_IR_reg[7]/NET0131  , \P2_IR_reg[8]/NET0131  , \P2_IR_reg[9]/NET0131  , \P2_addr_reg[0]/NET0131  , \P2_addr_reg[10]/NET0131  , \P2_addr_reg[11]/NET0131  , \P2_addr_reg[12]/NET0131  , \P2_addr_reg[13]/NET0131  , \P2_addr_reg[14]/NET0131  , \P2_addr_reg[15]/NET0131  , \P2_addr_reg[16]/NET0131  , \P2_addr_reg[17]/NET0131  , \P2_addr_reg[18]/NET0131  , \P2_addr_reg[19]/NET0131  , \P2_addr_reg[1]/NET0131  , \P2_addr_reg[2]/NET0131  , \P2_addr_reg[3]/NET0131  , \P2_addr_reg[4]/NET0131  , \P2_addr_reg[5]/NET0131  , \P2_addr_reg[6]/NET0131  , \P2_addr_reg[7]/NET0131  , \P2_addr_reg[8]/NET0131  , \P2_addr_reg[9]/NET0131  , \P2_d_reg[0]/NET0131  , \P2_d_reg[1]/NET0131  , \P2_datao_reg[0]/NET0131  , \P2_datao_reg[10]/NET0131  , \P2_datao_reg[11]/NET0131  , \P2_datao_reg[12]/NET0131  , \P2_datao_reg[13]/NET0131  , \P2_datao_reg[14]/NET0131  , \P2_datao_reg[15]/NET0131  , \P2_datao_reg[16]/NET0131  , \P2_datao_reg[17]/NET0131  , \P2_datao_reg[18]/NET0131  , \P2_datao_reg[19]/NET0131  , \P2_datao_reg[1]/NET0131  , \P2_datao_reg[20]/NET0131  , \P2_datao_reg[21]/NET0131  , \P2_datao_reg[22]/NET0131  , \P2_datao_reg[23]/NET0131  , \P2_datao_reg[24]/NET0131  , \P2_datao_reg[25]/NET0131  , \P2_datao_reg[26]/NET0131  , \P2_datao_reg[27]/NET0131  , \P2_datao_reg[28]/NET0131  , \P2_datao_reg[29]/NET0131  , \P2_datao_reg[2]/NET0131  , \P2_datao_reg[30]/NET0131  , \P2_datao_reg[31]/NET0131  , \P2_datao_reg[3]/NET0131  , \P2_datao_reg[4]/NET0131  , \P2_datao_reg[5]/NET0131  , \P2_datao_reg[6]/NET0131  , \P2_datao_reg[7]/NET0131  , \P2_datao_reg[8]/NET0131  , \P2_datao_reg[9]/NET0131  , \P2_rd_reg/NET0131  , \P2_reg0_reg[0]/NET0131  , \P2_reg0_reg[10]/NET0131  , \P2_reg0_reg[11]/NET0131  , \P2_reg0_reg[12]/NET0131  , \P2_reg0_reg[13]/NET0131  , \P2_reg0_reg[14]/NET0131  , \P2_reg0_reg[15]/NET0131  , \P2_reg0_reg[16]/NET0131  , \P2_reg0_reg[17]/NET0131  , \P2_reg0_reg[18]/NET0131  , \P2_reg0_reg[19]/NET0131  , \P2_reg0_reg[1]/NET0131  , \P2_reg0_reg[20]/NET0131  , \P2_reg0_reg[21]/NET0131  , \P2_reg0_reg[22]/NET0131  , \P2_reg0_reg[23]/NET0131  , \P2_reg0_reg[24]/NET0131  , \P2_reg0_reg[25]/NET0131  , \P2_reg0_reg[26]/NET0131  , \P2_reg0_reg[27]/NET0131  , \P2_reg0_reg[28]/NET0131  , \P2_reg0_reg[29]/NET0131  , \P2_reg0_reg[2]/NET0131  , \P2_reg0_reg[30]/NET0131  , \P2_reg0_reg[31]/NET0131  , \P2_reg0_reg[3]/NET0131  , \P2_reg0_reg[4]/NET0131  , \P2_reg0_reg[5]/NET0131  , \P2_reg0_reg[6]/NET0131  , \P2_reg0_reg[7]/NET0131  , \P2_reg0_reg[8]/NET0131  , \P2_reg0_reg[9]/NET0131  , \P2_reg1_reg[0]/NET0131  , \P2_reg1_reg[10]/NET0131  , \P2_reg1_reg[11]/NET0131  , \P2_reg1_reg[12]/NET0131  , \P2_reg1_reg[13]/NET0131  , \P2_reg1_reg[14]/NET0131  , \P2_reg1_reg[15]/NET0131  , \P2_reg1_reg[16]/NET0131  , \P2_reg1_reg[17]/NET0131  , \P2_reg1_reg[18]/NET0131  , \P2_reg1_reg[19]/NET0131  , \P2_reg1_reg[1]/NET0131  , \P2_reg1_reg[20]/NET0131  , \P2_reg1_reg[21]/NET0131  , \P2_reg1_reg[22]/NET0131  , \P2_reg1_reg[23]/NET0131  , \P2_reg1_reg[24]/NET0131  , \P2_reg1_reg[25]/NET0131  , \P2_reg1_reg[26]/NET0131  , \P2_reg1_reg[27]/NET0131  , \P2_reg1_reg[28]/NET0131  , \P2_reg1_reg[29]/NET0131  , \P2_reg1_reg[2]/NET0131  , \P2_reg1_reg[30]/NET0131  , \P2_reg1_reg[31]/NET0131  , \P2_reg1_reg[3]/NET0131  , \P2_reg1_reg[4]/NET0131  , \P2_reg1_reg[5]/NET0131  , \P2_reg1_reg[6]/NET0131  , \P2_reg1_reg[7]/NET0131  , \P2_reg1_reg[8]/NET0131  , \P2_reg1_reg[9]/NET0131  , \P2_reg2_reg[0]/NET0131  , \P2_reg2_reg[10]/NET0131  , \P2_reg2_reg[11]/NET0131  , \P2_reg2_reg[12]/NET0131  , \P2_reg2_reg[13]/NET0131  , \P2_reg2_reg[14]/NET0131  , \P2_reg2_reg[15]/NET0131  , \P2_reg2_reg[16]/NET0131  , \P2_reg2_reg[17]/NET0131  , \P2_reg2_reg[18]/NET0131  , \P2_reg2_reg[19]/NET0131  , \P2_reg2_reg[1]/NET0131  , \P2_reg2_reg[20]/NET0131  , \P2_reg2_reg[21]/NET0131  , \P2_reg2_reg[22]/NET0131  , \P2_reg2_reg[23]/NET0131  , \P2_reg2_reg[24]/NET0131  , \P2_reg2_reg[25]/NET0131  , \P2_reg2_reg[26]/NET0131  , \P2_reg2_reg[27]/NET0131  , \P2_reg2_reg[28]/NET0131  , \P2_reg2_reg[29]/NET0131  , \P2_reg2_reg[2]/NET0131  , \P2_reg2_reg[30]/NET0131  , \P2_reg2_reg[31]/NET0131  , \P2_reg2_reg[3]/NET0131  , \P2_reg2_reg[4]/NET0131  , \P2_reg2_reg[5]/NET0131  , \P2_reg2_reg[6]/NET0131  , \P2_reg2_reg[7]/NET0131  , \P2_reg2_reg[8]/NET0131  , \P2_reg2_reg[9]/NET0131  , \P2_reg3_reg[0]/NET0131  , \P2_reg3_reg[10]/NET0131  , \P2_reg3_reg[11]/NET0131  , \P2_reg3_reg[12]/NET0131  , \P2_reg3_reg[13]/NET0131  , \P2_reg3_reg[14]/NET0131  , \P2_reg3_reg[15]/NET0131  , \P2_reg3_reg[16]/NET0131  , \P2_reg3_reg[17]/NET0131  , \P2_reg3_reg[18]/NET0131  , \P2_reg3_reg[19]/NET0131  , \P2_reg3_reg[1]/NET0131  , \P2_reg3_reg[20]/NET0131  , \P2_reg3_reg[21]/NET0131  , \P2_reg3_reg[22]/NET0131  , \P2_reg3_reg[23]/NET0131  , \P2_reg3_reg[24]/NET0131  , \P2_reg3_reg[25]/NET0131  , \P2_reg3_reg[26]/NET0131  , \P2_reg3_reg[27]/NET0131  , \P2_reg3_reg[28]/NET0131  , \P2_reg3_reg[2]/NET0131  , \P2_reg3_reg[3]/NET0131  , \P2_reg3_reg[4]/NET0131  , \P2_reg3_reg[5]/NET0131  , \P2_reg3_reg[6]/NET0131  , \P2_reg3_reg[7]/NET0131  , \P2_reg3_reg[8]/NET0131  , \P2_reg3_reg[9]/NET0131  , \P2_wr_reg/NET0131  , \si[0]_pad  , \si[10]_pad  , \si[11]_pad  , \si[12]_pad  , \si[13]_pad  , \si[14]_pad  , \si[15]_pad  , \si[16]_pad  , \si[17]_pad  , \si[18]_pad  , \si[19]_pad  , \si[1]_pad  , \si[20]_pad  , \si[21]_pad  , \si[22]_pad  , \si[23]_pad  , \si[24]_pad  , \si[25]_pad  , \si[26]_pad  , \si[27]_pad  , \si[28]_pad  , \si[29]_pad  , \si[2]_pad  , \si[30]_pad  , \si[31]_pad  , \si[3]_pad  , \si[4]_pad  , \si[5]_pad  , \si[6]_pad  , \si[7]_pad  , \si[8]_pad  , \si[9]_pad  , \P1_state_reg[0]/NET0131_syn_2  , \_al_n0  , \_al_n1  , \g70791/_0_  , \g70792/_0_  , \g70793/_0_  , \g70794/_0_  , \g70795/_0_  , \g70796/_0_  , \g70813/_0_  , \g70814/_0_  , \g70848/_0_  , \g70849/_0_  , \g70850/_0_  , \g70851/_0_  , \g70852/_0_  , \g70856/_0_  , \g70857/_0_  , \g70858/_0_  , \g70859/_0_  , \g70860/_0_  , \g70861/_0_  , \g70862/_0_  , \g70896/_0_  , \g70902/_0_  , \g70903/_0_  , \g70904/_0_  , \g70906/_0_  , \g70907/_0_  , \g70908/_0_  , \g70909/_0_  , \g70910/_0_  , \g70911/_0_  , \g70912/_0_  , \g70913/_0_  , \g70914/_0_  , \g70915/_0_  , \g70916/_0_  , \g70917/_0_  , \g70918/_0_  , \g70919/_0_  , \g70920/_0_  , \g70921/_0_  , \g70922/_0_  , \g70923/_0_  , \g70924/_0_  , \g70925/_0_  , \g70926/_0_  , \g70927/_0_  , \g70987/_0_  , \g70988/_0_  , \g70989/_0_  , \g70990/_0_  , \g70991/_0_  , \g71006/_0_  , \g71007/_0_  , \g71009/_0_  , \g71010/_0_  , \g71011/_0_  , \g71012/_0_  , \g71013/_0_  , \g71014/_0_  , \g71015/_0_  , \g71016/_0_  , \g71017/_0_  , \g71018/_0_  , \g71019/_0_  , \g71020/_0_  , \g71021/_0_  , \g71022/_0_  , \g71023/_0_  , \g71090/_0_  , \g71091/_0_  , \g71092/_0_  , \g71093/_0_  , \g71094/_0_  , \g71125/_0_  , \g71130/_0_  , \g71131/_0_  , \g71132/_0_  , \g71133/_0_  , \g71134/_0_  , \g71135/_0_  , \g71136/_0_  , \g71137/_0_  , \g71138/_0_  , \g71139/_0_  , \g71140/_0_  , \g71141/_0_  , \g71142/_0_  , \g71143/_0_  , \g71144/_0_  , \g71145/_0_  , \g71150/_0_  , \g71151/_0_  , \g71152/_0_  , \g71153/_0_  , \g71154/_0_  , \g71155/_0_  , \g71156/_0_  , \g71157/_0_  , \g71158/_0_  , \g71230/_0_  , \g71231/_0_  , \g71232/_0_  , \g71233/_0_  , \g71234/_0_  , \g71235/_0_  , \g71236/_0_  , \g71238/_0_  , \g71239/_0_  , \g71270/_0_  , \g71275/_0_  , \g71276/_0_  , \g71277/_0_  , \g71278/_0_  , \g71279/_0_  , \g71280/_0_  , \g71281/_0_  , \g71282/_0_  , \g71283/_0_  , \g71284/_0_  , \g71285/_0_  , \g71286/_0_  , \g71287/_0_  , \g71288/_0_  , \g71289/_0_  , \g71290/_0_  , \g71291/_0_  , \g71292/_0_  , \g71293/_0_  , \g71294/_0_  , \g71295/_0_  , \g71296/_0_  , \g71297/_0_  , \g71298/_0_  , \g71299/_0_  , \g71300/_0_  , \g71301/_0_  , \g71302/_0_  , \g71303/_0_  , \g71304/_0_  , \g71305/_0_  , \g71306/_0_  , \g71307/_0_  , \g71382/_0_  , \g71384/_0_  , \g71385/_0_  , \g71387/_0_  , \g71388/_0_  , \g71389/_0_  , \g71439/_0_  , \g71440/_0_  , \g71441/_0_  , \g71442/_0_  , \g71443/_0_  , \g71444/_0_  , \g71445/_0_  , \g71446/_0_  , \g71447/_0_  , \g71448/_0_  , \g71449/_0_  , \g71450/_0_  , \g71451/_0_  , \g71452/_0_  , \g71453/_0_  , \g71454/_0_  , \g71455/_0_  , \g71456/_0_  , \g71457/_0_  , \g71458/_0_  , \g71459/_0_  , \g71460/_0_  , \g71461/_0_  , \g71536/_0_  , \g71537/_0_  , \g71538/_0_  , \g71540/_0_  , \g71541/_0_  , \g71542/_0_  , \g71602/_0_  , \g71604/_0_  , \g71610/_0_  , \g71611/_0_  , \g71618/_0_  , \g71619/_0_  , \g71620/_0_  , \g71621/_0_  , \g71622/_0_  , \g71623/_0_  , \g71624/_0_  , \g71625/_0_  , \g71626/_0_  , \g71627/_0_  , \g71629/_0_  , \g71630/_0_  , \g71631/_0_  , \g71632/_0_  , \g71633/_0_  , \g71634/_0_  , \g71635/_0_  , \g71636/_0_  , \g71710/_0_  , \g71711/_0_  , \g71782/_0_  , \g71785/_0_  , \g71786/_0_  , \g71787/_0_  , \g71788/_0_  , \g71789/_0_  , \g71790/_0_  , \g71791/_0_  , \g71792/_0_  , \g71793/_0_  , \g71794/_0_  , \g71795/_0_  , \g71796/_0_  , \g71797/_0_  , \g71798/_0_  , \g71799/_0_  , \g71883/_0_  , \g72000/_0_  , \g72001/_0_  , \g72002/_0_  , \g72003/_0_  , \g72004/_0_  , \g72005/_0_  , \g72236/_0_  , \g72237/_0_  , \g72238/_0_  , \g72239/_0_  , \g72240/_0_  , \g72372/_0_  , \g72376/_0_  , \g72383/_0_  , \g72561/_0_  , \g72562/_0_  , \g72563/_0_  , \g72564/_0_  , \g72970/_0_  , \g72980/_0_  , \g72981/_0_  , \g72982/_0_  , \g72983/_0_  , \g74234/_0_  , \g74260/_0_  , \g75086/_0_  , \g75087/_0_  , \g75088/_0_  , \g75089/_0_  , \g75091/_0_  , \g75092/_0_  , \g80304/_3_  , \g80305/_3_  , \g80306/_3_  , \g80307/_3_  , \g80308/_0_  , \g80309/_0_  , \g80815/_0_  , \g80816/_0_  , \g80817/_0_  , \g80818/_0_  , \g80819/_0_  , \g80820/_0_  , \g80821/_0_  , \g80822/_0_  , \g80823/_0_  , \g80824/_0_  , \g80825/_0_  , \g80826/_3_  , \g80827/_0_  , \g80828/_0_  , \g80829/_0_  , \g80830/_0_  , \g80831/_0_  , \g80832/_0_  , \g80833/_0_  , \g80834/_0_  , \g80835/_0_  , \g80836/_0_  , \g80837/_0_  , \g80838/_3_  , \g80839/_0_  , \g80840/_3_  , \g80841/_0_  , \g80859/_3_  , \g80860/_3_  , \g80861/_3_  , \g80862/_3_  , \g80863/_3_  , \g80864/_3_  , \g80865/_3_  , \g80866/_3_  , \g80867/_3_  , \g80868/_3_  , \g80869/_3_  , \g80870/_3_  , \g80871/_3_  , \g80872/_3_  , \g80873/_3_  , \g80874/_3_  , \g80875/_3_  , \g80876/_3_  , \g80877/_3_  , \g80878/_3_  , \g80879/_0_  , \g80880/_3_  , \g80881/_3_  , \g80882/_3_  , \g80883/_3_  , \g80884/_3_  , \g80885/_3_  , \g80886/_3_  , \g80888/_0_  , \g81262/_0_  , \g81278/_0_  , \g81884/_0_  , \g81893/_0_  , \g81896/_0_  , \g81897/_0_  , \g81898/_0_  , \g81899/_0_  , \g81900/_0_  , \g81901/_0_  , \g81902/_0_  , \g81903/_0_  , \g81904/_0_  , \g81905/_0_  , \g81906/_0_  , \g81907/_0_  , \g81908/_0_  , \g81909/_0_  , \g81910/_0_  , \g81911/_0_  , \g81923/_0_  , \g81924/_0_  , \g81925/_0_  , \g81926/_0_  , \g82414/_0_  , \g82532/_0_  , \g83134/_0_  , \g83135/_0_  , \g83141/_0_  , \g83142/_0_  , \g83145/_0_  , \g83146/_0_  , \g83147/_0_  , \g83148/_0_  , \g83152/_0_  , \g83153/_0_  , \g83154/_0_  , \g83155/_0_  , \g83156/_0_  , \g83157/_0_  , \g83158/_0_  , \g83159/_0_  , \g83164/_0_  , \g83165/_0_  , \g83177/_0_  , \g83178/_0_  , \g83409/_0_  , \g83411/_0_  , \g83807/u3_syn_4  , \g84138/u3_syn_4  , \g85062/_0_  , \g85079/_2_  , \g85113/_0_  , \g85121/_0_  , \g85594/_0_  , \g85663/_0_  , \g85669/_0_  , \g85749/_0_  , \g85784/_0_  , \g85809/_0_  , \g85817/_0_  , \g85828/_0_  , \g85845/_0_  , \g85851/_0_  , \g85858/_0_  , \g85871/_0_  , \g85882_dup/_0_  , \g85891/_0_  , \g85900/_0_  , \g85905/_0_  , \g85917/_0_  , \g85934/_0_  , \g85949/_0_  , \g85971/_0_  , \g85997/_0_  , \g86044/_0_  , \g86053/_0_  , \g86063/_0_  , \g86082/_0_  , \g86088/_0_  , \g86098/_0_  , \g86105/_0_  , \g86179/_0_  , \g86256_dup/_0_  , \g86264/_0_  , \g86273/_0_  , \g86281/_0_  , \g86288/_0_  , \g86297/_0_  , \g86304/_0_  , \g86310/_0_  , \g86320/_0_  , \g86328/_0_  , \g86339/_0_  , \g86353/_0_  , \g86360/_0_  , \g86368/_0_  , \g86373/_0_  , \g86385/_0_  , \g86392/_0_  , \g86399/_0_  , \g86421/_0_  , \g86432/_0_  , \g87592/_1__syn_2  , \g87632/_1_  , \g92847/_0_  , \g92957/_0_  , \g93056/_0_  , \g93289/_0_  , \g93538_dup95061/_0_  , \g93856/_0_  , \g93870/_0_  , \g94004/_0_  , \g94128/_0_  , \g94173/_0_  , \g94187/_0_  , \g94191/_0_  , \g94318/_0_  , \g94505/_0_  , rd_pad , \so[0]_pad  , \so[10]_pad  , \so[11]_pad  , \so[12]_pad  , \so[13]_pad  , \so[14]_pad  , \so[15]_pad  , \so[16]_pad  , \so[17]_pad  , \so[18]_pad  , \so[19]_pad  , \so[1]_pad  , \so[2]_pad  , \so[3]_pad  , \so[4]_pad  , \so[5]_pad  , \so[6]_pad  , \so[7]_pad  , \so[8]_pad  , \so[9]_pad  , wr_pad );
  input \P1_B_reg/NET0131  ;
  input \P1_IR_reg[0]/NET0131  ;
  input \P1_IR_reg[10]/NET0131  ;
  input \P1_IR_reg[11]/NET0131  ;
  input \P1_IR_reg[12]/NET0131  ;
  input \P1_IR_reg[13]/NET0131  ;
  input \P1_IR_reg[14]/NET0131  ;
  input \P1_IR_reg[15]/NET0131  ;
  input \P1_IR_reg[16]/NET0131  ;
  input \P1_IR_reg[17]/NET0131  ;
  input \P1_IR_reg[18]/NET0131  ;
  input \P1_IR_reg[19]/NET0131  ;
  input \P1_IR_reg[1]/NET0131  ;
  input \P1_IR_reg[20]/NET0131  ;
  input \P1_IR_reg[21]/NET0131  ;
  input \P1_IR_reg[22]/NET0131  ;
  input \P1_IR_reg[23]/NET0131  ;
  input \P1_IR_reg[24]/NET0131  ;
  input \P1_IR_reg[25]/NET0131  ;
  input \P1_IR_reg[26]/NET0131  ;
  input \P1_IR_reg[27]/NET0131  ;
  input \P1_IR_reg[28]/NET0131  ;
  input \P1_IR_reg[29]/NET0131  ;
  input \P1_IR_reg[2]/NET0131  ;
  input \P1_IR_reg[30]/NET0131  ;
  input \P1_IR_reg[31]/NET0131  ;
  input \P1_IR_reg[3]/NET0131  ;
  input \P1_IR_reg[4]/NET0131  ;
  input \P1_IR_reg[5]/NET0131  ;
  input \P1_IR_reg[6]/NET0131  ;
  input \P1_IR_reg[7]/NET0131  ;
  input \P1_IR_reg[8]/NET0131  ;
  input \P1_IR_reg[9]/NET0131  ;
  input \P1_addr_reg[0]/NET0131  ;
  input \P1_addr_reg[10]/NET0131  ;
  input \P1_addr_reg[11]/NET0131  ;
  input \P1_addr_reg[12]/NET0131  ;
  input \P1_addr_reg[13]/NET0131  ;
  input \P1_addr_reg[14]/NET0131  ;
  input \P1_addr_reg[15]/NET0131  ;
  input \P1_addr_reg[16]/NET0131  ;
  input \P1_addr_reg[17]/NET0131  ;
  input \P1_addr_reg[18]/NET0131  ;
  input \P1_addr_reg[19]/NET0131  ;
  input \P1_addr_reg[1]/NET0131  ;
  input \P1_addr_reg[2]/NET0131  ;
  input \P1_addr_reg[3]/NET0131  ;
  input \P1_addr_reg[4]/NET0131  ;
  input \P1_addr_reg[5]/NET0131  ;
  input \P1_addr_reg[6]/NET0131  ;
  input \P1_addr_reg[7]/NET0131  ;
  input \P1_addr_reg[8]/NET0131  ;
  input \P1_addr_reg[9]/NET0131  ;
  input \P1_d_reg[0]/NET0131  ;
  input \P1_d_reg[1]/NET0131  ;
  input \P1_datao_reg[0]/NET0131  ;
  input \P1_datao_reg[10]/NET0131  ;
  input \P1_datao_reg[11]/NET0131  ;
  input \P1_datao_reg[12]/NET0131  ;
  input \P1_datao_reg[13]/NET0131  ;
  input \P1_datao_reg[14]/NET0131  ;
  input \P1_datao_reg[15]/NET0131  ;
  input \P1_datao_reg[16]/NET0131  ;
  input \P1_datao_reg[17]/NET0131  ;
  input \P1_datao_reg[18]/NET0131  ;
  input \P1_datao_reg[19]/NET0131  ;
  input \P1_datao_reg[1]/NET0131  ;
  input \P1_datao_reg[20]/NET0131  ;
  input \P1_datao_reg[21]/NET0131  ;
  input \P1_datao_reg[22]/NET0131  ;
  input \P1_datao_reg[23]/NET0131  ;
  input \P1_datao_reg[24]/NET0131  ;
  input \P1_datao_reg[25]/NET0131  ;
  input \P1_datao_reg[26]/NET0131  ;
  input \P1_datao_reg[27]/NET0131  ;
  input \P1_datao_reg[28]/NET0131  ;
  input \P1_datao_reg[29]/NET0131  ;
  input \P1_datao_reg[2]/NET0131  ;
  input \P1_datao_reg[30]/NET0131  ;
  input \P1_datao_reg[31]/NET0131  ;
  input \P1_datao_reg[3]/NET0131  ;
  input \P1_datao_reg[4]/NET0131  ;
  input \P1_datao_reg[5]/NET0131  ;
  input \P1_datao_reg[6]/NET0131  ;
  input \P1_datao_reg[7]/NET0131  ;
  input \P1_datao_reg[8]/NET0131  ;
  input \P1_datao_reg[9]/NET0131  ;
  input \P1_rd_reg/NET0131  ;
  input \P1_reg0_reg[0]/NET0131  ;
  input \P1_reg0_reg[10]/NET0131  ;
  input \P1_reg0_reg[11]/NET0131  ;
  input \P1_reg0_reg[12]/NET0131  ;
  input \P1_reg0_reg[13]/NET0131  ;
  input \P1_reg0_reg[14]/NET0131  ;
  input \P1_reg0_reg[15]/NET0131  ;
  input \P1_reg0_reg[16]/NET0131  ;
  input \P1_reg0_reg[17]/NET0131  ;
  input \P1_reg0_reg[18]/NET0131  ;
  input \P1_reg0_reg[19]/NET0131  ;
  input \P1_reg0_reg[1]/NET0131  ;
  input \P1_reg0_reg[20]/NET0131  ;
  input \P1_reg0_reg[21]/NET0131  ;
  input \P1_reg0_reg[22]/NET0131  ;
  input \P1_reg0_reg[23]/NET0131  ;
  input \P1_reg0_reg[24]/NET0131  ;
  input \P1_reg0_reg[25]/NET0131  ;
  input \P1_reg0_reg[26]/NET0131  ;
  input \P1_reg0_reg[27]/NET0131  ;
  input \P1_reg0_reg[28]/NET0131  ;
  input \P1_reg0_reg[29]/NET0131  ;
  input \P1_reg0_reg[2]/NET0131  ;
  input \P1_reg0_reg[30]/NET0131  ;
  input \P1_reg0_reg[31]/NET0131  ;
  input \P1_reg0_reg[3]/NET0131  ;
  input \P1_reg0_reg[4]/NET0131  ;
  input \P1_reg0_reg[5]/NET0131  ;
  input \P1_reg0_reg[6]/NET0131  ;
  input \P1_reg0_reg[7]/NET0131  ;
  input \P1_reg0_reg[8]/NET0131  ;
  input \P1_reg0_reg[9]/NET0131  ;
  input \P1_reg1_reg[0]/NET0131  ;
  input \P1_reg1_reg[10]/NET0131  ;
  input \P1_reg1_reg[11]/NET0131  ;
  input \P1_reg1_reg[12]/NET0131  ;
  input \P1_reg1_reg[13]/NET0131  ;
  input \P1_reg1_reg[14]/NET0131  ;
  input \P1_reg1_reg[15]/NET0131  ;
  input \P1_reg1_reg[16]/NET0131  ;
  input \P1_reg1_reg[17]/NET0131  ;
  input \P1_reg1_reg[18]/NET0131  ;
  input \P1_reg1_reg[19]/NET0131  ;
  input \P1_reg1_reg[1]/NET0131  ;
  input \P1_reg1_reg[20]/NET0131  ;
  input \P1_reg1_reg[21]/NET0131  ;
  input \P1_reg1_reg[22]/NET0131  ;
  input \P1_reg1_reg[23]/NET0131  ;
  input \P1_reg1_reg[24]/NET0131  ;
  input \P1_reg1_reg[25]/NET0131  ;
  input \P1_reg1_reg[26]/NET0131  ;
  input \P1_reg1_reg[27]/NET0131  ;
  input \P1_reg1_reg[28]/NET0131  ;
  input \P1_reg1_reg[29]/NET0131  ;
  input \P1_reg1_reg[2]/NET0131  ;
  input \P1_reg1_reg[30]/NET0131  ;
  input \P1_reg1_reg[31]/NET0131  ;
  input \P1_reg1_reg[3]/NET0131  ;
  input \P1_reg1_reg[4]/NET0131  ;
  input \P1_reg1_reg[5]/NET0131  ;
  input \P1_reg1_reg[6]/NET0131  ;
  input \P1_reg1_reg[7]/NET0131  ;
  input \P1_reg1_reg[8]/NET0131  ;
  input \P1_reg1_reg[9]/NET0131  ;
  input \P1_reg2_reg[0]/NET0131  ;
  input \P1_reg2_reg[10]/NET0131  ;
  input \P1_reg2_reg[11]/NET0131  ;
  input \P1_reg2_reg[12]/NET0131  ;
  input \P1_reg2_reg[13]/NET0131  ;
  input \P1_reg2_reg[14]/NET0131  ;
  input \P1_reg2_reg[15]/NET0131  ;
  input \P1_reg2_reg[16]/NET0131  ;
  input \P1_reg2_reg[17]/NET0131  ;
  input \P1_reg2_reg[18]/NET0131  ;
  input \P1_reg2_reg[19]/NET0131  ;
  input \P1_reg2_reg[1]/NET0131  ;
  input \P1_reg2_reg[20]/NET0131  ;
  input \P1_reg2_reg[21]/NET0131  ;
  input \P1_reg2_reg[22]/NET0131  ;
  input \P1_reg2_reg[23]/NET0131  ;
  input \P1_reg2_reg[24]/NET0131  ;
  input \P1_reg2_reg[25]/NET0131  ;
  input \P1_reg2_reg[26]/NET0131  ;
  input \P1_reg2_reg[27]/NET0131  ;
  input \P1_reg2_reg[28]/NET0131  ;
  input \P1_reg2_reg[29]/NET0131  ;
  input \P1_reg2_reg[2]/NET0131  ;
  input \P1_reg2_reg[30]/NET0131  ;
  input \P1_reg2_reg[31]/NET0131  ;
  input \P1_reg2_reg[3]/NET0131  ;
  input \P1_reg2_reg[4]/NET0131  ;
  input \P1_reg2_reg[5]/NET0131  ;
  input \P1_reg2_reg[6]/NET0131  ;
  input \P1_reg2_reg[7]/NET0131  ;
  input \P1_reg2_reg[8]/NET0131  ;
  input \P1_reg2_reg[9]/NET0131  ;
  input \P1_reg3_reg[0]/NET0131  ;
  input \P1_reg3_reg[10]/NET0131  ;
  input \P1_reg3_reg[11]/NET0131  ;
  input \P1_reg3_reg[12]/NET0131  ;
  input \P1_reg3_reg[13]/NET0131  ;
  input \P1_reg3_reg[14]/NET0131  ;
  input \P1_reg3_reg[15]/NET0131  ;
  input \P1_reg3_reg[16]/NET0131  ;
  input \P1_reg3_reg[17]/NET0131  ;
  input \P1_reg3_reg[18]/NET0131  ;
  input \P1_reg3_reg[19]/NET0131  ;
  input \P1_reg3_reg[1]/NET0131  ;
  input \P1_reg3_reg[20]/NET0131  ;
  input \P1_reg3_reg[21]/NET0131  ;
  input \P1_reg3_reg[22]/NET0131  ;
  input \P1_reg3_reg[23]/NET0131  ;
  input \P1_reg3_reg[24]/NET0131  ;
  input \P1_reg3_reg[25]/NET0131  ;
  input \P1_reg3_reg[26]/NET0131  ;
  input \P1_reg3_reg[27]/NET0131  ;
  input \P1_reg3_reg[28]/NET0131  ;
  input \P1_reg3_reg[2]/NET0131  ;
  input \P1_reg3_reg[3]/NET0131  ;
  input \P1_reg3_reg[4]/NET0131  ;
  input \P1_reg3_reg[5]/NET0131  ;
  input \P1_reg3_reg[6]/NET0131  ;
  input \P1_reg3_reg[7]/NET0131  ;
  input \P1_reg3_reg[8]/NET0131  ;
  input \P1_reg3_reg[9]/NET0131  ;
  input \P1_state_reg[0]/NET0131  ;
  input \P1_wr_reg/NET0131  ;
  input \P2_B_reg/NET0131  ;
  input \P2_IR_reg[0]/NET0131  ;
  input \P2_IR_reg[10]/NET0131  ;
  input \P2_IR_reg[11]/NET0131  ;
  input \P2_IR_reg[12]/NET0131  ;
  input \P2_IR_reg[13]/NET0131  ;
  input \P2_IR_reg[14]/NET0131  ;
  input \P2_IR_reg[15]/NET0131  ;
  input \P2_IR_reg[16]/NET0131  ;
  input \P2_IR_reg[17]/NET0131  ;
  input \P2_IR_reg[18]/NET0131  ;
  input \P2_IR_reg[19]/NET0131  ;
  input \P2_IR_reg[1]/NET0131  ;
  input \P2_IR_reg[20]/NET0131  ;
  input \P2_IR_reg[21]/NET0131  ;
  input \P2_IR_reg[22]/NET0131  ;
  input \P2_IR_reg[23]/NET0131  ;
  input \P2_IR_reg[24]/NET0131  ;
  input \P2_IR_reg[25]/NET0131  ;
  input \P2_IR_reg[26]/NET0131  ;
  input \P2_IR_reg[27]/NET0131  ;
  input \P2_IR_reg[28]/NET0131  ;
  input \P2_IR_reg[29]/NET0131  ;
  input \P2_IR_reg[2]/NET0131  ;
  input \P2_IR_reg[30]/NET0131  ;
  input \P2_IR_reg[31]/NET0131  ;
  input \P2_IR_reg[3]/NET0131  ;
  input \P2_IR_reg[4]/NET0131  ;
  input \P2_IR_reg[5]/NET0131  ;
  input \P2_IR_reg[6]/NET0131  ;
  input \P2_IR_reg[7]/NET0131  ;
  input \P2_IR_reg[8]/NET0131  ;
  input \P2_IR_reg[9]/NET0131  ;
  input \P2_addr_reg[0]/NET0131  ;
  input \P2_addr_reg[10]/NET0131  ;
  input \P2_addr_reg[11]/NET0131  ;
  input \P2_addr_reg[12]/NET0131  ;
  input \P2_addr_reg[13]/NET0131  ;
  input \P2_addr_reg[14]/NET0131  ;
  input \P2_addr_reg[15]/NET0131  ;
  input \P2_addr_reg[16]/NET0131  ;
  input \P2_addr_reg[17]/NET0131  ;
  input \P2_addr_reg[18]/NET0131  ;
  input \P2_addr_reg[19]/NET0131  ;
  input \P2_addr_reg[1]/NET0131  ;
  input \P2_addr_reg[2]/NET0131  ;
  input \P2_addr_reg[3]/NET0131  ;
  input \P2_addr_reg[4]/NET0131  ;
  input \P2_addr_reg[5]/NET0131  ;
  input \P2_addr_reg[6]/NET0131  ;
  input \P2_addr_reg[7]/NET0131  ;
  input \P2_addr_reg[8]/NET0131  ;
  input \P2_addr_reg[9]/NET0131  ;
  input \P2_d_reg[0]/NET0131  ;
  input \P2_d_reg[1]/NET0131  ;
  input \P2_datao_reg[0]/NET0131  ;
  input \P2_datao_reg[10]/NET0131  ;
  input \P2_datao_reg[11]/NET0131  ;
  input \P2_datao_reg[12]/NET0131  ;
  input \P2_datao_reg[13]/NET0131  ;
  input \P2_datao_reg[14]/NET0131  ;
  input \P2_datao_reg[15]/NET0131  ;
  input \P2_datao_reg[16]/NET0131  ;
  input \P2_datao_reg[17]/NET0131  ;
  input \P2_datao_reg[18]/NET0131  ;
  input \P2_datao_reg[19]/NET0131  ;
  input \P2_datao_reg[1]/NET0131  ;
  input \P2_datao_reg[20]/NET0131  ;
  input \P2_datao_reg[21]/NET0131  ;
  input \P2_datao_reg[22]/NET0131  ;
  input \P2_datao_reg[23]/NET0131  ;
  input \P2_datao_reg[24]/NET0131  ;
  input \P2_datao_reg[25]/NET0131  ;
  input \P2_datao_reg[26]/NET0131  ;
  input \P2_datao_reg[27]/NET0131  ;
  input \P2_datao_reg[28]/NET0131  ;
  input \P2_datao_reg[29]/NET0131  ;
  input \P2_datao_reg[2]/NET0131  ;
  input \P2_datao_reg[30]/NET0131  ;
  input \P2_datao_reg[31]/NET0131  ;
  input \P2_datao_reg[3]/NET0131  ;
  input \P2_datao_reg[4]/NET0131  ;
  input \P2_datao_reg[5]/NET0131  ;
  input \P2_datao_reg[6]/NET0131  ;
  input \P2_datao_reg[7]/NET0131  ;
  input \P2_datao_reg[8]/NET0131  ;
  input \P2_datao_reg[9]/NET0131  ;
  input \P2_rd_reg/NET0131  ;
  input \P2_reg0_reg[0]/NET0131  ;
  input \P2_reg0_reg[10]/NET0131  ;
  input \P2_reg0_reg[11]/NET0131  ;
  input \P2_reg0_reg[12]/NET0131  ;
  input \P2_reg0_reg[13]/NET0131  ;
  input \P2_reg0_reg[14]/NET0131  ;
  input \P2_reg0_reg[15]/NET0131  ;
  input \P2_reg0_reg[16]/NET0131  ;
  input \P2_reg0_reg[17]/NET0131  ;
  input \P2_reg0_reg[18]/NET0131  ;
  input \P2_reg0_reg[19]/NET0131  ;
  input \P2_reg0_reg[1]/NET0131  ;
  input \P2_reg0_reg[20]/NET0131  ;
  input \P2_reg0_reg[21]/NET0131  ;
  input \P2_reg0_reg[22]/NET0131  ;
  input \P2_reg0_reg[23]/NET0131  ;
  input \P2_reg0_reg[24]/NET0131  ;
  input \P2_reg0_reg[25]/NET0131  ;
  input \P2_reg0_reg[26]/NET0131  ;
  input \P2_reg0_reg[27]/NET0131  ;
  input \P2_reg0_reg[28]/NET0131  ;
  input \P2_reg0_reg[29]/NET0131  ;
  input \P2_reg0_reg[2]/NET0131  ;
  input \P2_reg0_reg[30]/NET0131  ;
  input \P2_reg0_reg[31]/NET0131  ;
  input \P2_reg0_reg[3]/NET0131  ;
  input \P2_reg0_reg[4]/NET0131  ;
  input \P2_reg0_reg[5]/NET0131  ;
  input \P2_reg0_reg[6]/NET0131  ;
  input \P2_reg0_reg[7]/NET0131  ;
  input \P2_reg0_reg[8]/NET0131  ;
  input \P2_reg0_reg[9]/NET0131  ;
  input \P2_reg1_reg[0]/NET0131  ;
  input \P2_reg1_reg[10]/NET0131  ;
  input \P2_reg1_reg[11]/NET0131  ;
  input \P2_reg1_reg[12]/NET0131  ;
  input \P2_reg1_reg[13]/NET0131  ;
  input \P2_reg1_reg[14]/NET0131  ;
  input \P2_reg1_reg[15]/NET0131  ;
  input \P2_reg1_reg[16]/NET0131  ;
  input \P2_reg1_reg[17]/NET0131  ;
  input \P2_reg1_reg[18]/NET0131  ;
  input \P2_reg1_reg[19]/NET0131  ;
  input \P2_reg1_reg[1]/NET0131  ;
  input \P2_reg1_reg[20]/NET0131  ;
  input \P2_reg1_reg[21]/NET0131  ;
  input \P2_reg1_reg[22]/NET0131  ;
  input \P2_reg1_reg[23]/NET0131  ;
  input \P2_reg1_reg[24]/NET0131  ;
  input \P2_reg1_reg[25]/NET0131  ;
  input \P2_reg1_reg[26]/NET0131  ;
  input \P2_reg1_reg[27]/NET0131  ;
  input \P2_reg1_reg[28]/NET0131  ;
  input \P2_reg1_reg[29]/NET0131  ;
  input \P2_reg1_reg[2]/NET0131  ;
  input \P2_reg1_reg[30]/NET0131  ;
  input \P2_reg1_reg[31]/NET0131  ;
  input \P2_reg1_reg[3]/NET0131  ;
  input \P2_reg1_reg[4]/NET0131  ;
  input \P2_reg1_reg[5]/NET0131  ;
  input \P2_reg1_reg[6]/NET0131  ;
  input \P2_reg1_reg[7]/NET0131  ;
  input \P2_reg1_reg[8]/NET0131  ;
  input \P2_reg1_reg[9]/NET0131  ;
  input \P2_reg2_reg[0]/NET0131  ;
  input \P2_reg2_reg[10]/NET0131  ;
  input \P2_reg2_reg[11]/NET0131  ;
  input \P2_reg2_reg[12]/NET0131  ;
  input \P2_reg2_reg[13]/NET0131  ;
  input \P2_reg2_reg[14]/NET0131  ;
  input \P2_reg2_reg[15]/NET0131  ;
  input \P2_reg2_reg[16]/NET0131  ;
  input \P2_reg2_reg[17]/NET0131  ;
  input \P2_reg2_reg[18]/NET0131  ;
  input \P2_reg2_reg[19]/NET0131  ;
  input \P2_reg2_reg[1]/NET0131  ;
  input \P2_reg2_reg[20]/NET0131  ;
  input \P2_reg2_reg[21]/NET0131  ;
  input \P2_reg2_reg[22]/NET0131  ;
  input \P2_reg2_reg[23]/NET0131  ;
  input \P2_reg2_reg[24]/NET0131  ;
  input \P2_reg2_reg[25]/NET0131  ;
  input \P2_reg2_reg[26]/NET0131  ;
  input \P2_reg2_reg[27]/NET0131  ;
  input \P2_reg2_reg[28]/NET0131  ;
  input \P2_reg2_reg[29]/NET0131  ;
  input \P2_reg2_reg[2]/NET0131  ;
  input \P2_reg2_reg[30]/NET0131  ;
  input \P2_reg2_reg[31]/NET0131  ;
  input \P2_reg2_reg[3]/NET0131  ;
  input \P2_reg2_reg[4]/NET0131  ;
  input \P2_reg2_reg[5]/NET0131  ;
  input \P2_reg2_reg[6]/NET0131  ;
  input \P2_reg2_reg[7]/NET0131  ;
  input \P2_reg2_reg[8]/NET0131  ;
  input \P2_reg2_reg[9]/NET0131  ;
  input \P2_reg3_reg[0]/NET0131  ;
  input \P2_reg3_reg[10]/NET0131  ;
  input \P2_reg3_reg[11]/NET0131  ;
  input \P2_reg3_reg[12]/NET0131  ;
  input \P2_reg3_reg[13]/NET0131  ;
  input \P2_reg3_reg[14]/NET0131  ;
  input \P2_reg3_reg[15]/NET0131  ;
  input \P2_reg3_reg[16]/NET0131  ;
  input \P2_reg3_reg[17]/NET0131  ;
  input \P2_reg3_reg[18]/NET0131  ;
  input \P2_reg3_reg[19]/NET0131  ;
  input \P2_reg3_reg[1]/NET0131  ;
  input \P2_reg3_reg[20]/NET0131  ;
  input \P2_reg3_reg[21]/NET0131  ;
  input \P2_reg3_reg[22]/NET0131  ;
  input \P2_reg3_reg[23]/NET0131  ;
  input \P2_reg3_reg[24]/NET0131  ;
  input \P2_reg3_reg[25]/NET0131  ;
  input \P2_reg3_reg[26]/NET0131  ;
  input \P2_reg3_reg[27]/NET0131  ;
  input \P2_reg3_reg[28]/NET0131  ;
  input \P2_reg3_reg[2]/NET0131  ;
  input \P2_reg3_reg[3]/NET0131  ;
  input \P2_reg3_reg[4]/NET0131  ;
  input \P2_reg3_reg[5]/NET0131  ;
  input \P2_reg3_reg[6]/NET0131  ;
  input \P2_reg3_reg[7]/NET0131  ;
  input \P2_reg3_reg[8]/NET0131  ;
  input \P2_reg3_reg[9]/NET0131  ;
  input \P2_wr_reg/NET0131  ;
  input \si[0]_pad  ;
  input \si[10]_pad  ;
  input \si[11]_pad  ;
  input \si[12]_pad  ;
  input \si[13]_pad  ;
  input \si[14]_pad  ;
  input \si[15]_pad  ;
  input \si[16]_pad  ;
  input \si[17]_pad  ;
  input \si[18]_pad  ;
  input \si[19]_pad  ;
  input \si[1]_pad  ;
  input \si[20]_pad  ;
  input \si[21]_pad  ;
  input \si[22]_pad  ;
  input \si[23]_pad  ;
  input \si[24]_pad  ;
  input \si[25]_pad  ;
  input \si[26]_pad  ;
  input \si[27]_pad  ;
  input \si[28]_pad  ;
  input \si[29]_pad  ;
  input \si[2]_pad  ;
  input \si[30]_pad  ;
  input \si[31]_pad  ;
  input \si[3]_pad  ;
  input \si[4]_pad  ;
  input \si[5]_pad  ;
  input \si[6]_pad  ;
  input \si[7]_pad  ;
  input \si[8]_pad  ;
  input \si[9]_pad  ;
  output \P1_state_reg[0]/NET0131_syn_2  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g70791/_0_  ;
  output \g70792/_0_  ;
  output \g70793/_0_  ;
  output \g70794/_0_  ;
  output \g70795/_0_  ;
  output \g70796/_0_  ;
  output \g70813/_0_  ;
  output \g70814/_0_  ;
  output \g70848/_0_  ;
  output \g70849/_0_  ;
  output \g70850/_0_  ;
  output \g70851/_0_  ;
  output \g70852/_0_  ;
  output \g70856/_0_  ;
  output \g70857/_0_  ;
  output \g70858/_0_  ;
  output \g70859/_0_  ;
  output \g70860/_0_  ;
  output \g70861/_0_  ;
  output \g70862/_0_  ;
  output \g70896/_0_  ;
  output \g70902/_0_  ;
  output \g70903/_0_  ;
  output \g70904/_0_  ;
  output \g70906/_0_  ;
  output \g70907/_0_  ;
  output \g70908/_0_  ;
  output \g70909/_0_  ;
  output \g70910/_0_  ;
  output \g70911/_0_  ;
  output \g70912/_0_  ;
  output \g70913/_0_  ;
  output \g70914/_0_  ;
  output \g70915/_0_  ;
  output \g70916/_0_  ;
  output \g70917/_0_  ;
  output \g70918/_0_  ;
  output \g70919/_0_  ;
  output \g70920/_0_  ;
  output \g70921/_0_  ;
  output \g70922/_0_  ;
  output \g70923/_0_  ;
  output \g70924/_0_  ;
  output \g70925/_0_  ;
  output \g70926/_0_  ;
  output \g70927/_0_  ;
  output \g70987/_0_  ;
  output \g70988/_0_  ;
  output \g70989/_0_  ;
  output \g70990/_0_  ;
  output \g70991/_0_  ;
  output \g71006/_0_  ;
  output \g71007/_0_  ;
  output \g71009/_0_  ;
  output \g71010/_0_  ;
  output \g71011/_0_  ;
  output \g71012/_0_  ;
  output \g71013/_0_  ;
  output \g71014/_0_  ;
  output \g71015/_0_  ;
  output \g71016/_0_  ;
  output \g71017/_0_  ;
  output \g71018/_0_  ;
  output \g71019/_0_  ;
  output \g71020/_0_  ;
  output \g71021/_0_  ;
  output \g71022/_0_  ;
  output \g71023/_0_  ;
  output \g71090/_0_  ;
  output \g71091/_0_  ;
  output \g71092/_0_  ;
  output \g71093/_0_  ;
  output \g71094/_0_  ;
  output \g71125/_0_  ;
  output \g71130/_0_  ;
  output \g71131/_0_  ;
  output \g71132/_0_  ;
  output \g71133/_0_  ;
  output \g71134/_0_  ;
  output \g71135/_0_  ;
  output \g71136/_0_  ;
  output \g71137/_0_  ;
  output \g71138/_0_  ;
  output \g71139/_0_  ;
  output \g71140/_0_  ;
  output \g71141/_0_  ;
  output \g71142/_0_  ;
  output \g71143/_0_  ;
  output \g71144/_0_  ;
  output \g71145/_0_  ;
  output \g71150/_0_  ;
  output \g71151/_0_  ;
  output \g71152/_0_  ;
  output \g71153/_0_  ;
  output \g71154/_0_  ;
  output \g71155/_0_  ;
  output \g71156/_0_  ;
  output \g71157/_0_  ;
  output \g71158/_0_  ;
  output \g71230/_0_  ;
  output \g71231/_0_  ;
  output \g71232/_0_  ;
  output \g71233/_0_  ;
  output \g71234/_0_  ;
  output \g71235/_0_  ;
  output \g71236/_0_  ;
  output \g71238/_0_  ;
  output \g71239/_0_  ;
  output \g71270/_0_  ;
  output \g71275/_0_  ;
  output \g71276/_0_  ;
  output \g71277/_0_  ;
  output \g71278/_0_  ;
  output \g71279/_0_  ;
  output \g71280/_0_  ;
  output \g71281/_0_  ;
  output \g71282/_0_  ;
  output \g71283/_0_  ;
  output \g71284/_0_  ;
  output \g71285/_0_  ;
  output \g71286/_0_  ;
  output \g71287/_0_  ;
  output \g71288/_0_  ;
  output \g71289/_0_  ;
  output \g71290/_0_  ;
  output \g71291/_0_  ;
  output \g71292/_0_  ;
  output \g71293/_0_  ;
  output \g71294/_0_  ;
  output \g71295/_0_  ;
  output \g71296/_0_  ;
  output \g71297/_0_  ;
  output \g71298/_0_  ;
  output \g71299/_0_  ;
  output \g71300/_0_  ;
  output \g71301/_0_  ;
  output \g71302/_0_  ;
  output \g71303/_0_  ;
  output \g71304/_0_  ;
  output \g71305/_0_  ;
  output \g71306/_0_  ;
  output \g71307/_0_  ;
  output \g71382/_0_  ;
  output \g71384/_0_  ;
  output \g71385/_0_  ;
  output \g71387/_0_  ;
  output \g71388/_0_  ;
  output \g71389/_0_  ;
  output \g71439/_0_  ;
  output \g71440/_0_  ;
  output \g71441/_0_  ;
  output \g71442/_0_  ;
  output \g71443/_0_  ;
  output \g71444/_0_  ;
  output \g71445/_0_  ;
  output \g71446/_0_  ;
  output \g71447/_0_  ;
  output \g71448/_0_  ;
  output \g71449/_0_  ;
  output \g71450/_0_  ;
  output \g71451/_0_  ;
  output \g71452/_0_  ;
  output \g71453/_0_  ;
  output \g71454/_0_  ;
  output \g71455/_0_  ;
  output \g71456/_0_  ;
  output \g71457/_0_  ;
  output \g71458/_0_  ;
  output \g71459/_0_  ;
  output \g71460/_0_  ;
  output \g71461/_0_  ;
  output \g71536/_0_  ;
  output \g71537/_0_  ;
  output \g71538/_0_  ;
  output \g71540/_0_  ;
  output \g71541/_0_  ;
  output \g71542/_0_  ;
  output \g71602/_0_  ;
  output \g71604/_0_  ;
  output \g71610/_0_  ;
  output \g71611/_0_  ;
  output \g71618/_0_  ;
  output \g71619/_0_  ;
  output \g71620/_0_  ;
  output \g71621/_0_  ;
  output \g71622/_0_  ;
  output \g71623/_0_  ;
  output \g71624/_0_  ;
  output \g71625/_0_  ;
  output \g71626/_0_  ;
  output \g71627/_0_  ;
  output \g71629/_0_  ;
  output \g71630/_0_  ;
  output \g71631/_0_  ;
  output \g71632/_0_  ;
  output \g71633/_0_  ;
  output \g71634/_0_  ;
  output \g71635/_0_  ;
  output \g71636/_0_  ;
  output \g71710/_0_  ;
  output \g71711/_0_  ;
  output \g71782/_0_  ;
  output \g71785/_0_  ;
  output \g71786/_0_  ;
  output \g71787/_0_  ;
  output \g71788/_0_  ;
  output \g71789/_0_  ;
  output \g71790/_0_  ;
  output \g71791/_0_  ;
  output \g71792/_0_  ;
  output \g71793/_0_  ;
  output \g71794/_0_  ;
  output \g71795/_0_  ;
  output \g71796/_0_  ;
  output \g71797/_0_  ;
  output \g71798/_0_  ;
  output \g71799/_0_  ;
  output \g71883/_0_  ;
  output \g72000/_0_  ;
  output \g72001/_0_  ;
  output \g72002/_0_  ;
  output \g72003/_0_  ;
  output \g72004/_0_  ;
  output \g72005/_0_  ;
  output \g72236/_0_  ;
  output \g72237/_0_  ;
  output \g72238/_0_  ;
  output \g72239/_0_  ;
  output \g72240/_0_  ;
  output \g72372/_0_  ;
  output \g72376/_0_  ;
  output \g72383/_0_  ;
  output \g72561/_0_  ;
  output \g72562/_0_  ;
  output \g72563/_0_  ;
  output \g72564/_0_  ;
  output \g72970/_0_  ;
  output \g72980/_0_  ;
  output \g72981/_0_  ;
  output \g72982/_0_  ;
  output \g72983/_0_  ;
  output \g74234/_0_  ;
  output \g74260/_0_  ;
  output \g75086/_0_  ;
  output \g75087/_0_  ;
  output \g75088/_0_  ;
  output \g75089/_0_  ;
  output \g75091/_0_  ;
  output \g75092/_0_  ;
  output \g80304/_3_  ;
  output \g80305/_3_  ;
  output \g80306/_3_  ;
  output \g80307/_3_  ;
  output \g80308/_0_  ;
  output \g80309/_0_  ;
  output \g80815/_0_  ;
  output \g80816/_0_  ;
  output \g80817/_0_  ;
  output \g80818/_0_  ;
  output \g80819/_0_  ;
  output \g80820/_0_  ;
  output \g80821/_0_  ;
  output \g80822/_0_  ;
  output \g80823/_0_  ;
  output \g80824/_0_  ;
  output \g80825/_0_  ;
  output \g80826/_3_  ;
  output \g80827/_0_  ;
  output \g80828/_0_  ;
  output \g80829/_0_  ;
  output \g80830/_0_  ;
  output \g80831/_0_  ;
  output \g80832/_0_  ;
  output \g80833/_0_  ;
  output \g80834/_0_  ;
  output \g80835/_0_  ;
  output \g80836/_0_  ;
  output \g80837/_0_  ;
  output \g80838/_3_  ;
  output \g80839/_0_  ;
  output \g80840/_3_  ;
  output \g80841/_0_  ;
  output \g80859/_3_  ;
  output \g80860/_3_  ;
  output \g80861/_3_  ;
  output \g80862/_3_  ;
  output \g80863/_3_  ;
  output \g80864/_3_  ;
  output \g80865/_3_  ;
  output \g80866/_3_  ;
  output \g80867/_3_  ;
  output \g80868/_3_  ;
  output \g80869/_3_  ;
  output \g80870/_3_  ;
  output \g80871/_3_  ;
  output \g80872/_3_  ;
  output \g80873/_3_  ;
  output \g80874/_3_  ;
  output \g80875/_3_  ;
  output \g80876/_3_  ;
  output \g80877/_3_  ;
  output \g80878/_3_  ;
  output \g80879/_0_  ;
  output \g80880/_3_  ;
  output \g80881/_3_  ;
  output \g80882/_3_  ;
  output \g80883/_3_  ;
  output \g80884/_3_  ;
  output \g80885/_3_  ;
  output \g80886/_3_  ;
  output \g80888/_0_  ;
  output \g81262/_0_  ;
  output \g81278/_0_  ;
  output \g81884/_0_  ;
  output \g81893/_0_  ;
  output \g81896/_0_  ;
  output \g81897/_0_  ;
  output \g81898/_0_  ;
  output \g81899/_0_  ;
  output \g81900/_0_  ;
  output \g81901/_0_  ;
  output \g81902/_0_  ;
  output \g81903/_0_  ;
  output \g81904/_0_  ;
  output \g81905/_0_  ;
  output \g81906/_0_  ;
  output \g81907/_0_  ;
  output \g81908/_0_  ;
  output \g81909/_0_  ;
  output \g81910/_0_  ;
  output \g81911/_0_  ;
  output \g81923/_0_  ;
  output \g81924/_0_  ;
  output \g81925/_0_  ;
  output \g81926/_0_  ;
  output \g82414/_0_  ;
  output \g82532/_0_  ;
  output \g83134/_0_  ;
  output \g83135/_0_  ;
  output \g83141/_0_  ;
  output \g83142/_0_  ;
  output \g83145/_0_  ;
  output \g83146/_0_  ;
  output \g83147/_0_  ;
  output \g83148/_0_  ;
  output \g83152/_0_  ;
  output \g83153/_0_  ;
  output \g83154/_0_  ;
  output \g83155/_0_  ;
  output \g83156/_0_  ;
  output \g83157/_0_  ;
  output \g83158/_0_  ;
  output \g83159/_0_  ;
  output \g83164/_0_  ;
  output \g83165/_0_  ;
  output \g83177/_0_  ;
  output \g83178/_0_  ;
  output \g83409/_0_  ;
  output \g83411/_0_  ;
  output \g83807/u3_syn_4  ;
  output \g84138/u3_syn_4  ;
  output \g85062/_0_  ;
  output \g85079/_2_  ;
  output \g85113/_0_  ;
  output \g85121/_0_  ;
  output \g85594/_0_  ;
  output \g85663/_0_  ;
  output \g85669/_0_  ;
  output \g85749/_0_  ;
  output \g85784/_0_  ;
  output \g85809/_0_  ;
  output \g85817/_0_  ;
  output \g85828/_0_  ;
  output \g85845/_0_  ;
  output \g85851/_0_  ;
  output \g85858/_0_  ;
  output \g85871/_0_  ;
  output \g85882_dup/_0_  ;
  output \g85891/_0_  ;
  output \g85900/_0_  ;
  output \g85905/_0_  ;
  output \g85917/_0_  ;
  output \g85934/_0_  ;
  output \g85949/_0_  ;
  output \g85971/_0_  ;
  output \g85997/_0_  ;
  output \g86044/_0_  ;
  output \g86053/_0_  ;
  output \g86063/_0_  ;
  output \g86082/_0_  ;
  output \g86088/_0_  ;
  output \g86098/_0_  ;
  output \g86105/_0_  ;
  output \g86179/_0_  ;
  output \g86256_dup/_0_  ;
  output \g86264/_0_  ;
  output \g86273/_0_  ;
  output \g86281/_0_  ;
  output \g86288/_0_  ;
  output \g86297/_0_  ;
  output \g86304/_0_  ;
  output \g86310/_0_  ;
  output \g86320/_0_  ;
  output \g86328/_0_  ;
  output \g86339/_0_  ;
  output \g86353/_0_  ;
  output \g86360/_0_  ;
  output \g86368/_0_  ;
  output \g86373/_0_  ;
  output \g86385/_0_  ;
  output \g86392/_0_  ;
  output \g86399/_0_  ;
  output \g86421/_0_  ;
  output \g86432/_0_  ;
  output \g87592/_1__syn_2  ;
  output \g87632/_1_  ;
  output \g92847/_0_  ;
  output \g92957/_0_  ;
  output \g93056/_0_  ;
  output \g93289/_0_  ;
  output \g93538_dup95061/_0_  ;
  output \g93856/_0_  ;
  output \g93870/_0_  ;
  output \g94004/_0_  ;
  output \g94128/_0_  ;
  output \g94173/_0_  ;
  output \g94187/_0_  ;
  output \g94191/_0_  ;
  output \g94318/_0_  ;
  output \g94505/_0_  ;
  output rd_pad ;
  output \so[0]_pad  ;
  output \so[10]_pad  ;
  output \so[11]_pad  ;
  output \so[12]_pad  ;
  output \so[13]_pad  ;
  output \so[14]_pad  ;
  output \so[15]_pad  ;
  output \so[16]_pad  ;
  output \so[17]_pad  ;
  output \so[18]_pad  ;
  output \so[19]_pad  ;
  output \so[1]_pad  ;
  output \so[2]_pad  ;
  output \so[3]_pad  ;
  output \so[4]_pad  ;
  output \so[5]_pad  ;
  output \so[6]_pad  ;
  output \so[7]_pad  ;
  output \so[8]_pad  ;
  output \so[9]_pad  ;
  output wr_pad ;
  wire n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 ;
  assign n462 = ~\P1_IR_reg[8]/NET0131  & ~\P1_IR_reg[9]/NET0131  ;
  assign n463 = ~\P1_IR_reg[10]/NET0131  & n462 ;
  assign n464 = ~\P1_IR_reg[0]/NET0131  & ~\P1_IR_reg[1]/NET0131  ;
  assign n465 = ~\P1_IR_reg[2]/NET0131  & n464 ;
  assign n466 = ~\P1_IR_reg[3]/NET0131  & n465 ;
  assign n467 = ~\P1_IR_reg[4]/NET0131  & n466 ;
  assign n468 = ~\P1_IR_reg[5]/NET0131  & ~\P1_IR_reg[6]/NET0131  ;
  assign n469 = ~\P1_IR_reg[7]/NET0131  & n468 ;
  assign n470 = n467 & n469 ;
  assign n471 = n463 & n470 ;
  assign n472 = ~\P1_IR_reg[11]/NET0131  & ~\P1_IR_reg[12]/NET0131  ;
  assign n487 = ~\P1_IR_reg[13]/NET0131  & n472 ;
  assign n508 = ~\P1_IR_reg[14]/NET0131  & n487 ;
  assign n507 = ~\P1_IR_reg[16]/NET0131  & ~\P1_IR_reg[17]/NET0131  ;
  assign n509 = ~\P1_IR_reg[15]/NET0131  & ~\P1_IR_reg[18]/NET0131  ;
  assign n510 = n507 & n509 ;
  assign n511 = n508 & n510 ;
  assign n512 = n471 & n511 ;
  assign n500 = ~\P1_IR_reg[20]/NET0131  & ~\P1_IR_reg[21]/NET0131  ;
  assign n519 = ~\P1_IR_reg[19]/NET0131  & ~\P1_IR_reg[22]/NET0131  ;
  assign n520 = n500 & n519 ;
  assign n521 = n512 & n520 ;
  assign n517 = ~\P1_IR_reg[24]/NET0131  & ~\P1_IR_reg[25]/NET0131  ;
  assign n518 = ~\P1_IR_reg[26]/NET0131  & n517 ;
  assign n522 = ~\P1_IR_reg[23]/NET0131  & n518 ;
  assign n523 = n521 & n522 ;
  assign n524 = \P1_IR_reg[31]/NET0131  & ~n523 ;
  assign n525 = \P1_IR_reg[27]/NET0131  & ~n524 ;
  assign n526 = ~\P1_IR_reg[27]/NET0131  & n524 ;
  assign n527 = ~n525 & ~n526 ;
  assign n474 = ~\P1_IR_reg[14]/NET0131  & ~\P1_IR_reg[15]/NET0131  ;
  assign n488 = n463 & n487 ;
  assign n489 = n470 & n488 ;
  assign n490 = n474 & n489 ;
  assign n491 = \P1_IR_reg[31]/NET0131  & ~n490 ;
  assign n479 = ~\P1_IR_reg[17]/NET0131  & ~\P1_IR_reg[18]/NET0131  ;
  assign n492 = ~\P1_IR_reg[16]/NET0131  & ~\P1_IR_reg[19]/NET0131  ;
  assign n493 = n479 & n492 ;
  assign n501 = n493 & n500 ;
  assign n528 = ~\P1_IR_reg[22]/NET0131  & ~\P1_IR_reg[23]/NET0131  ;
  assign n529 = n501 & n528 ;
  assign n530 = ~\P1_IR_reg[27]/NET0131  & n518 ;
  assign n531 = n529 & n530 ;
  assign n532 = \P1_IR_reg[31]/NET0131  & ~n531 ;
  assign n533 = ~n491 & ~n532 ;
  assign n534 = \P1_IR_reg[28]/NET0131  & ~n533 ;
  assign n535 = ~\P1_IR_reg[28]/NET0131  & n533 ;
  assign n536 = ~n534 & ~n535 ;
  assign n537 = n527 & ~n536 ;
  assign n570 = ~\P2_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n571 = ~\P2_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n572 = \P2_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n573 = \P2_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n574 = ~n572 & ~n573 ;
  assign n575 = ~n571 & ~n574 ;
  assign n576 = ~n570 & n575 ;
  assign n577 = \P2_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = ~\P2_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n580 = ~\P2_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n581 = ~n579 & ~n580 ;
  assign n582 = ~\P2_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n583 = ~\P2_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n584 = ~n582 & ~n583 ;
  assign n585 = n581 & n584 ;
  assign n586 = ~n578 & n585 ;
  assign n587 = \P2_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n588 = \P2_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n589 = ~n587 & ~n588 ;
  assign n590 = ~n579 & ~n589 ;
  assign n591 = \P2_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n592 = \P2_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = n581 & ~n582 ;
  assign n595 = ~n593 & n594 ;
  assign n596 = ~n590 & ~n595 ;
  assign n597 = ~n586 & n596 ;
  assign n557 = ~\P2_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n562 = ~\P2_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n563 = ~n557 & ~n562 ;
  assign n564 = ~\P2_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n598 = ~\P2_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n599 = ~n564 & ~n598 ;
  assign n600 = n563 & n599 ;
  assign n601 = ~n597 & n600 ;
  assign n558 = \P2_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n559 = \P2_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n560 = ~n558 & ~n559 ;
  assign n561 = ~n557 & ~n560 ;
  assign n565 = n563 & ~n564 ;
  assign n566 = \P2_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n567 = \P2_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n568 = ~n566 & ~n567 ;
  assign n569 = n565 & ~n568 ;
  assign n602 = ~n561 & ~n569 ;
  assign n603 = ~n601 & n602 ;
  assign n549 = ~\P2_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n544 = ~\P2_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n550 = ~\P2_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n551 = ~n544 & ~n550 ;
  assign n552 = ~n549 & n551 ;
  assign n604 = ~\P2_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n605 = n552 & ~n604 ;
  assign n606 = ~n603 & n605 ;
  assign n545 = \P2_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n546 = \P2_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = ~n544 & ~n547 ;
  assign n553 = \P2_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n554 = \P2_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n555 = ~n553 & ~n554 ;
  assign n556 = n552 & ~n555 ;
  assign n607 = ~n548 & ~n556 ;
  assign n608 = ~n606 & n607 ;
  assign n609 = ~\P2_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n610 = ~\P2_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n611 = ~n609 & ~n610 ;
  assign n612 = ~\P2_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n613 = ~\P2_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n614 = ~n612 & ~n613 ;
  assign n615 = n611 & n614 ;
  assign n616 = ~n608 & n615 ;
  assign n849 = ~\P2_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n867 = ~\P2_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n890 = ~n849 & ~n867 ;
  assign n628 = ~\P2_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n850 = ~\P2_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n891 = ~n628 & ~n850 ;
  assign n892 = n890 & n891 ;
  assign n893 = n616 & n892 ;
  assign n856 = \P2_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n868 = \P2_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n894 = ~n856 & ~n868 ;
  assign n895 = ~n867 & ~n894 ;
  assign n629 = \P2_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n857 = \P2_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n896 = ~n629 & ~n857 ;
  assign n897 = ~n850 & ~n896 ;
  assign n898 = n890 & n897 ;
  assign n899 = ~n895 & ~n898 ;
  assign n617 = \P2_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n618 = \P2_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n619 = ~n617 & ~n618 ;
  assign n620 = ~n609 & ~n619 ;
  assign n621 = \P2_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n622 = \P2_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = ~n612 & ~n623 ;
  assign n625 = n611 & n624 ;
  assign n626 = ~n620 & ~n625 ;
  assign n900 = ~n626 & n892 ;
  assign n901 = n899 & ~n900 ;
  assign n902 = ~n893 & n901 ;
  assign n903 = ~\P2_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n1434 = ~\P2_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n1437 = ~\P2_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n1442 = ~\P2_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n1443 = ~n1437 & ~n1442 ;
  assign n1486 = ~n1434 & n1443 ;
  assign n1490 = ~n903 & n1486 ;
  assign n1650 = ~\P2_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n1586 = ~\P2_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n1481 = ~\P2_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n1589 = ~\P2_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n1597 = ~n1481 & ~n1589 ;
  assign n1651 = ~n1586 & n1597 ;
  assign n1652 = ~n1650 & n1651 ;
  assign n1653 = n1490 & n1652 ;
  assign n1654 = ~n902 & n1653 ;
  assign n1435 = \P2_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n1438 = \P2_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n1484 = ~n1435 & ~n1438 ;
  assign n1485 = ~n1434 & ~n1484 ;
  assign n904 = \P2_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n1439 = \P2_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n1487 = ~n904 & ~n1439 ;
  assign n1488 = n1486 & ~n1487 ;
  assign n1489 = ~n1485 & ~n1488 ;
  assign n1659 = ~n1489 & n1652 ;
  assign n1587 = \P2_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n1482 = \P2_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n1590 = \P2_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n1591 = ~n1482 & ~n1590 ;
  assign n1655 = ~n1586 & ~n1589 ;
  assign n1656 = ~n1591 & n1655 ;
  assign n1657 = ~n1587 & ~n1656 ;
  assign n1658 = ~n1650 & ~n1657 ;
  assign n1660 = \P2_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n1661 = ~n1658 & ~n1660 ;
  assign n1662 = ~n1659 & n1661 ;
  assign n1663 = ~n1654 & n1662 ;
  assign n1665 = ~\si[31]_pad  & n1663 ;
  assign n538 = ~\P1_addr_reg[19]/NET0131  & ~\P2_addr_reg[19]/NET0131  ;
  assign n539 = ~\P1_rd_reg/NET0131  & n538 ;
  assign n540 = \P1_addr_reg[19]/NET0131  & \P2_addr_reg[19]/NET0131  ;
  assign n541 = ~\P2_rd_reg/NET0131  & n540 ;
  assign n542 = ~n539 & ~n541 ;
  assign n1664 = \si[31]_pad  & ~n1663 ;
  assign n1666 = ~n542 & ~n1664 ;
  assign n1667 = ~n1665 & n1666 ;
  assign n1668 = \P2_datao_reg[31]/NET0131  & n1667 ;
  assign n1669 = ~\P2_datao_reg[31]/NET0131  & ~n1667 ;
  assign n1670 = ~n1668 & ~n1669 ;
  assign n1671 = ~n537 & n1670 ;
  assign n639 = n474 & n517 ;
  assign n640 = n529 & n639 ;
  assign n641 = n489 & n640 ;
  assign n642 = \P1_IR_reg[31]/NET0131  & ~n641 ;
  assign n643 = ~\P1_IR_reg[27]/NET0131  & ~\P1_IR_reg[28]/NET0131  ;
  assign n644 = ~\P1_IR_reg[26]/NET0131  & n643 ;
  assign n645 = ~\P1_IR_reg[29]/NET0131  & n644 ;
  assign n646 = \P1_IR_reg[31]/NET0131  & ~n645 ;
  assign n647 = ~n642 & ~n646 ;
  assign n648 = \P1_IR_reg[30]/NET0131  & ~n647 ;
  assign n649 = ~\P1_IR_reg[30]/NET0131  & n647 ;
  assign n650 = ~n648 & ~n649 ;
  assign n473 = n471 & n472 ;
  assign n651 = \P1_IR_reg[31]/NET0131  & ~n473 ;
  assign n480 = ~\P1_IR_reg[19]/NET0131  & ~\P1_IR_reg[20]/NET0131  ;
  assign n481 = n479 & n480 ;
  assign n475 = ~\P1_IR_reg[13]/NET0131  & ~\P1_IR_reg[16]/NET0131  ;
  assign n476 = n474 & n475 ;
  assign n652 = ~\P1_IR_reg[21]/NET0131  & ~\P1_IR_reg[24]/NET0131  ;
  assign n653 = n528 & n652 ;
  assign n654 = n476 & n653 ;
  assign n655 = n481 & n654 ;
  assign n656 = ~\P1_IR_reg[25]/NET0131  & n644 ;
  assign n657 = n655 & n656 ;
  assign n658 = \P1_IR_reg[31]/NET0131  & ~n657 ;
  assign n659 = ~n651 & ~n658 ;
  assign n660 = \P1_IR_reg[29]/NET0131  & ~n659 ;
  assign n661 = ~\P1_IR_reg[29]/NET0131  & n659 ;
  assign n662 = ~n660 & ~n661 ;
  assign n669 = n650 & n662 ;
  assign n670 = \P1_reg3_reg[3]/NET0131  & \P1_reg3_reg[4]/NET0131  ;
  assign n671 = \P1_reg3_reg[5]/NET0131  & n670 ;
  assign n672 = \P1_reg3_reg[6]/NET0131  & n671 ;
  assign n673 = \P1_reg3_reg[7]/NET0131  & n672 ;
  assign n674 = \P1_reg3_reg[8]/NET0131  & n673 ;
  assign n675 = \P1_reg3_reg[9]/NET0131  & n674 ;
  assign n676 = \P1_reg3_reg[10]/NET0131  & n675 ;
  assign n677 = \P1_reg3_reg[11]/NET0131  & n676 ;
  assign n678 = \P1_reg3_reg[12]/NET0131  & n677 ;
  assign n679 = \P1_reg3_reg[13]/NET0131  & \P1_reg3_reg[14]/NET0131  ;
  assign n680 = n678 & n679 ;
  assign n681 = \P1_reg3_reg[15]/NET0131  & \P1_reg3_reg[16]/NET0131  ;
  assign n682 = \P1_reg3_reg[17]/NET0131  & n681 ;
  assign n683 = n680 & n682 ;
  assign n684 = \P1_reg3_reg[18]/NET0131  & \P1_reg3_reg[19]/NET0131  ;
  assign n685 = n683 & n684 ;
  assign n879 = \P1_reg3_reg[20]/NET0131  & \P1_reg3_reg[21]/NET0131  ;
  assign n1467 = \P1_reg3_reg[22]/NET0131  & \P1_reg3_reg[23]/NET0131  ;
  assign n1468 = \P1_reg3_reg[24]/NET0131  & n1467 ;
  assign n1469 = n879 & n1468 ;
  assign n1470 = n685 & n1469 ;
  assign n1609 = \P1_reg3_reg[25]/NET0131  & \P1_reg3_reg[26]/NET0131  ;
  assign n1610 = \P1_reg3_reg[27]/NET0131  & \P1_reg3_reg[28]/NET0131  ;
  assign n1611 = n1609 & n1610 ;
  assign n1612 = n1470 & n1611 ;
  assign n1613 = n669 & n1612 ;
  assign n665 = ~n650 & ~n662 ;
  assign n1674 = \P1_reg0_reg[31]/NET0131  & n665 ;
  assign n667 = n650 & ~n662 ;
  assign n1672 = \P1_reg2_reg[31]/NET0131  & n667 ;
  assign n663 = ~n650 & n662 ;
  assign n1673 = \P1_reg1_reg[31]/NET0131  & n663 ;
  assign n1675 = ~n1672 & ~n1673 ;
  assign n1676 = ~n1674 & n1675 ;
  assign n1677 = ~n1613 & n1676 ;
  assign n1722 = n1671 & n1677 ;
  assign n1678 = ~n1671 & ~n1677 ;
  assign n1679 = \P2_datao_reg[30]/NET0131  & n542 ;
  assign n1680 = ~n1650 & ~n1660 ;
  assign n708 = ~n577 & ~n592 ;
  assign n709 = ~n576 & n708 ;
  assign n710 = n584 & ~n709 ;
  assign n711 = ~n588 & ~n591 ;
  assign n712 = ~n710 & n711 ;
  assign n705 = ~n562 & n599 ;
  assign n713 = n581 & n705 ;
  assign n714 = ~n712 & n713 ;
  assign n703 = ~n559 & ~n566 ;
  assign n704 = ~n562 & ~n703 ;
  assign n706 = ~n567 & ~n587 ;
  assign n707 = n705 & ~n706 ;
  assign n715 = ~n704 & ~n707 ;
  assign n716 = ~n714 & n715 ;
  assign n717 = ~n549 & ~n604 ;
  assign n718 = ~n550 & n717 ;
  assign n719 = ~n557 & n718 ;
  assign n720 = ~n716 & n719 ;
  assign n721 = ~n546 & ~n553 ;
  assign n722 = ~n550 & ~n721 ;
  assign n723 = ~n554 & ~n558 ;
  assign n724 = n718 & ~n723 ;
  assign n725 = ~n722 & ~n724 ;
  assign n726 = ~n720 & n725 ;
  assign n698 = ~n610 & ~n612 ;
  assign n727 = ~n544 & ~n613 ;
  assign n728 = n698 & n727 ;
  assign n851 = ~n849 & ~n850 ;
  assign n852 = ~n609 & ~n628 ;
  assign n853 = n851 & n852 ;
  assign n854 = n728 & n853 ;
  assign n855 = ~n726 & n854 ;
  assign n858 = ~n856 & ~n857 ;
  assign n859 = ~n849 & ~n858 ;
  assign n860 = ~n617 & ~n629 ;
  assign n861 = ~n628 & ~n860 ;
  assign n862 = n851 & n861 ;
  assign n863 = ~n859 & ~n862 ;
  assign n696 = ~n618 & ~n621 ;
  assign n697 = ~n610 & ~n696 ;
  assign n699 = ~n545 & ~n622 ;
  assign n700 = ~n613 & ~n699 ;
  assign n701 = n698 & n700 ;
  assign n702 = ~n697 & ~n701 ;
  assign n864 = ~n702 & n853 ;
  assign n865 = n863 & ~n864 ;
  assign n866 = ~n855 & n865 ;
  assign n1448 = ~n867 & ~n903 ;
  assign n1449 = n1443 & n1448 ;
  assign n1682 = ~n1434 & n1651 ;
  assign n1685 = n1449 & n1682 ;
  assign n1686 = ~n866 & n1685 ;
  assign n1440 = ~n1438 & ~n1439 ;
  assign n1441 = ~n1437 & ~n1440 ;
  assign n1444 = ~n868 & ~n904 ;
  assign n1445 = ~n903 & ~n1444 ;
  assign n1446 = n1443 & n1445 ;
  assign n1447 = ~n1441 & ~n1446 ;
  assign n1683 = ~n1447 & n1682 ;
  assign n1625 = ~n1435 & ~n1482 ;
  assign n1684 = ~n1625 & n1651 ;
  assign n1681 = ~n1586 & n1590 ;
  assign n1687 = ~n1587 & ~n1681 ;
  assign n1688 = ~n1684 & n1687 ;
  assign n1689 = ~n1683 & n1688 ;
  assign n1690 = ~n1686 & n1689 ;
  assign n1692 = ~n1680 & n1690 ;
  assign n1691 = n1680 & ~n1690 ;
  assign n1693 = ~n542 & ~n1691 ;
  assign n1694 = ~n1692 & n1693 ;
  assign n1695 = ~n1679 & ~n1694 ;
  assign n1696 = ~n537 & ~n1695 ;
  assign n1699 = \P1_reg2_reg[30]/NET0131  & n667 ;
  assign n1697 = \P1_reg0_reg[30]/NET0131  & n665 ;
  assign n1698 = \P1_reg1_reg[30]/NET0131  & n663 ;
  assign n1700 = ~n1697 & ~n1698 ;
  assign n1701 = ~n1699 & n1700 ;
  assign n1702 = ~n1613 & n1701 ;
  assign n1723 = n1696 & n1702 ;
  assign n1724 = ~n1678 & ~n1723 ;
  assign n1585 = \P2_datao_reg[29]/NET0131  & n542 ;
  assign n1588 = ~n1586 & ~n1587 ;
  assign n1515 = n895 & ~n903 ;
  assign n1516 = n1487 & ~n1515 ;
  assign n1592 = n1486 & ~n1516 ;
  assign n1593 = ~n1485 & ~n1592 ;
  assign n1594 = ~n1481 & ~n1593 ;
  assign n1595 = n1591 & ~n1594 ;
  assign n1596 = ~n1589 & ~n1595 ;
  assign n759 = ~n554 & ~n561 ;
  assign n760 = n717 & ~n759 ;
  assign n761 = ~n553 & ~n760 ;
  assign n762 = ~n591 & ~n710 ;
  assign n763 = n581 & n599 ;
  assign n764 = ~n762 & n763 ;
  assign n765 = ~n567 & ~n590 ;
  assign n766 = n599 & ~n765 ;
  assign n767 = ~n566 & ~n766 ;
  assign n768 = ~n764 & n767 ;
  assign n769 = n563 & n717 ;
  assign n770 = ~n768 & n769 ;
  assign n771 = n761 & ~n770 ;
  assign n772 = n551 & n614 ;
  assign n925 = n611 & n891 ;
  assign n926 = n772 & n925 ;
  assign n927 = ~n771 & n926 ;
  assign n928 = n620 & n891 ;
  assign n929 = ~n897 & ~n928 ;
  assign n757 = n548 & n614 ;
  assign n758 = ~n624 & ~n757 ;
  assign n930 = ~n758 & n925 ;
  assign n931 = n929 & ~n930 ;
  assign n932 = ~n927 & n931 ;
  assign n1598 = n890 & n1597 ;
  assign n1599 = n1490 & n1598 ;
  assign n1600 = ~n932 & n1599 ;
  assign n1601 = ~n1596 & ~n1600 ;
  assign n1603 = ~n1588 & n1601 ;
  assign n1602 = n1588 & ~n1601 ;
  assign n1604 = ~n542 & ~n1602 ;
  assign n1605 = ~n1603 & n1604 ;
  assign n1606 = ~n1585 & ~n1605 ;
  assign n1607 = ~n537 & ~n1606 ;
  assign n1615 = \P1_reg2_reg[29]/NET0131  & n667 ;
  assign n1608 = \P1_reg0_reg[29]/NET0131  & n665 ;
  assign n1614 = \P1_reg1_reg[29]/NET0131  & n663 ;
  assign n1616 = ~n1608 & ~n1614 ;
  assign n1617 = ~n1615 & n1616 ;
  assign n1618 = ~n1613 & n1617 ;
  assign n1619 = n1607 & n1618 ;
  assign n1620 = \P2_datao_reg[28]/NET0131  & n542 ;
  assign n1621 = ~n1589 & ~n1590 ;
  assign n953 = n697 & n852 ;
  assign n954 = ~n861 & ~n953 ;
  assign n800 = n552 & ~n613 ;
  assign n802 = n581 & n710 ;
  assign n801 = n581 & ~n711 ;
  assign n803 = n706 & ~n801 ;
  assign n804 = ~n802 & n803 ;
  assign n805 = ~n598 & ~n804 ;
  assign n806 = n565 & ~n604 ;
  assign n807 = n805 & n806 ;
  assign n808 = n800 & n807 ;
  assign n810 = ~n558 & ~n704 ;
  assign n811 = ~n557 & ~n604 ;
  assign n812 = ~n810 & n811 ;
  assign n813 = ~n554 & ~n812 ;
  assign n814 = n800 & ~n813 ;
  assign n809 = n722 & n727 ;
  assign n815 = ~n700 & ~n809 ;
  assign n816 = ~n814 & n815 ;
  assign n817 = ~n808 & n816 ;
  assign n955 = n698 & n852 ;
  assign n956 = ~n817 & n955 ;
  assign n957 = n954 & ~n956 ;
  assign n1548 = n851 & n1448 ;
  assign n1622 = ~n1481 & n1486 ;
  assign n1623 = n1548 & n1622 ;
  assign n1624 = ~n957 & n1623 ;
  assign n1546 = n859 & n1448 ;
  assign n1547 = ~n1445 & ~n1546 ;
  assign n1626 = n1486 & ~n1547 ;
  assign n1627 = ~n1434 & n1441 ;
  assign n1628 = n1625 & ~n1627 ;
  assign n1629 = ~n1626 & n1628 ;
  assign n1630 = ~n1481 & ~n1629 ;
  assign n1631 = ~n1624 & ~n1630 ;
  assign n1633 = ~n1621 & n1631 ;
  assign n1632 = n1621 & ~n1631 ;
  assign n1634 = ~n542 & ~n1632 ;
  assign n1635 = ~n1633 & n1634 ;
  assign n1636 = ~n1620 & ~n1635 ;
  assign n1637 = ~n537 & ~n1636 ;
  assign n1471 = \P1_reg3_reg[25]/NET0131  & n1470 ;
  assign n1472 = \P1_reg3_reg[26]/NET0131  & n1471 ;
  assign n1504 = \P1_reg3_reg[27]/NET0131  & n1472 ;
  assign n1641 = ~\P1_reg3_reg[28]/NET0131  & ~n1504 ;
  assign n1642 = ~n1612 & ~n1641 ;
  assign n1643 = n669 & n1642 ;
  assign n1640 = \P1_reg2_reg[28]/NET0131  & n667 ;
  assign n1638 = \P1_reg1_reg[28]/NET0131  & n663 ;
  assign n1639 = \P1_reg0_reg[28]/NET0131  & n665 ;
  assign n1644 = ~n1638 & ~n1639 ;
  assign n1645 = ~n1640 & n1644 ;
  assign n1646 = ~n1643 & n1645 ;
  assign n1710 = ~n1637 & ~n1646 ;
  assign n1711 = ~n1619 & n1710 ;
  assign n1707 = ~n1696 & ~n1702 ;
  assign n1712 = ~n1607 & ~n1618 ;
  assign n1725 = ~n1707 & ~n1712 ;
  assign n1726 = ~n1711 & n1725 ;
  assign n1727 = n1724 & ~n1726 ;
  assign n1728 = ~n1722 & ~n1727 ;
  assign n543 = \P2_datao_reg[19]/NET0131  & n542 ;
  assign n627 = ~n616 & n626 ;
  assign n630 = ~n628 & ~n629 ;
  assign n632 = ~n627 & n630 ;
  assign n631 = n627 & ~n630 ;
  assign n633 = ~n542 & ~n631 ;
  assign n634 = ~n632 & n633 ;
  assign n635 = ~n543 & ~n634 ;
  assign n636 = ~n537 & ~n635 ;
  assign n513 = \P1_IR_reg[31]/NET0131  & ~n512 ;
  assign n514 = ~\P1_IR_reg[19]/NET0131  & n513 ;
  assign n515 = \P1_IR_reg[19]/NET0131  & ~n513 ;
  assign n516 = ~n514 & ~n515 ;
  assign n637 = ~n516 & n537 ;
  assign n638 = ~n636 & ~n637 ;
  assign n686 = \P1_reg3_reg[18]/NET0131  & n683 ;
  assign n687 = ~\P1_reg3_reg[19]/NET0131  & ~n686 ;
  assign n688 = ~n685 & ~n687 ;
  assign n689 = n669 & n688 ;
  assign n668 = \P1_reg2_reg[19]/NET0131  & n667 ;
  assign n664 = \P1_reg1_reg[19]/NET0131  & n663 ;
  assign n666 = \P1_reg0_reg[19]/NET0131  & n665 ;
  assign n690 = ~n664 & ~n666 ;
  assign n691 = ~n668 & n690 ;
  assign n692 = ~n689 & n691 ;
  assign n693 = ~n638 & n692 ;
  assign n694 = \P2_datao_reg[18]/NET0131  & n542 ;
  assign n695 = ~n609 & ~n617 ;
  assign n729 = ~n726 & n728 ;
  assign n730 = n702 & ~n729 ;
  assign n732 = ~n695 & n730 ;
  assign n731 = n695 & ~n730 ;
  assign n733 = ~n542 & ~n731 ;
  assign n734 = ~n732 & n733 ;
  assign n735 = ~n694 & ~n734 ;
  assign n736 = ~n537 & ~n735 ;
  assign n737 = \P1_IR_reg[31]/NET0131  & ~n507 ;
  assign n738 = ~n491 & ~n737 ;
  assign n739 = \P1_IR_reg[18]/NET0131  & ~n738 ;
  assign n740 = ~\P1_IR_reg[18]/NET0131  & n738 ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = n537 & n741 ;
  assign n743 = ~n736 & ~n742 ;
  assign n747 = ~\P1_reg3_reg[18]/NET0131  & ~n683 ;
  assign n748 = ~n686 & ~n747 ;
  assign n749 = n669 & n748 ;
  assign n746 = \P1_reg1_reg[18]/NET0131  & n663 ;
  assign n744 = \P1_reg0_reg[18]/NET0131  & n665 ;
  assign n745 = \P1_reg2_reg[18]/NET0131  & n667 ;
  assign n750 = ~n744 & ~n745 ;
  assign n751 = ~n746 & n750 ;
  assign n752 = ~n749 & n751 ;
  assign n753 = ~n743 & n752 ;
  assign n754 = ~n693 & ~n753 ;
  assign n755 = \P2_datao_reg[17]/NET0131  & n542 ;
  assign n756 = ~n610 & ~n618 ;
  assign n773 = ~n771 & n772 ;
  assign n774 = n758 & ~n773 ;
  assign n776 = ~n756 & n774 ;
  assign n775 = n756 & ~n774 ;
  assign n777 = ~n542 & ~n775 ;
  assign n778 = ~n776 & n777 ;
  assign n779 = ~n755 & ~n778 ;
  assign n780 = ~n537 & ~n779 ;
  assign n477 = n473 & n476 ;
  assign n478 = \P1_IR_reg[31]/NET0131  & ~n477 ;
  assign n781 = ~\P1_IR_reg[17]/NET0131  & ~n478 ;
  assign n782 = \P1_IR_reg[17]/NET0131  & n478 ;
  assign n783 = ~n781 & ~n782 ;
  assign n784 = n537 & n783 ;
  assign n785 = ~n780 & ~n784 ;
  assign n789 = \P1_reg3_reg[15]/NET0131  & n680 ;
  assign n790 = \P1_reg3_reg[16]/NET0131  & n789 ;
  assign n791 = ~\P1_reg3_reg[17]/NET0131  & ~n790 ;
  assign n792 = ~n683 & ~n791 ;
  assign n793 = n669 & n792 ;
  assign n788 = \P1_reg1_reg[17]/NET0131  & n663 ;
  assign n786 = \P1_reg2_reg[17]/NET0131  & n667 ;
  assign n787 = \P1_reg0_reg[17]/NET0131  & n665 ;
  assign n794 = ~n786 & ~n787 ;
  assign n795 = ~n788 & n794 ;
  assign n796 = ~n793 & n795 ;
  assign n797 = ~n785 & n796 ;
  assign n798 = n785 & ~n796 ;
  assign n799 = \P2_datao_reg[16]/NET0131  & n542 ;
  assign n818 = ~n612 & ~n621 ;
  assign n820 = n817 & ~n818 ;
  assign n819 = ~n817 & n818 ;
  assign n821 = ~n542 & ~n819 ;
  assign n822 = ~n820 & n821 ;
  assign n823 = ~n799 & ~n822 ;
  assign n824 = ~n537 & ~n823 ;
  assign n825 = ~\P1_IR_reg[16]/NET0131  & ~n491 ;
  assign n826 = \P1_IR_reg[16]/NET0131  & n491 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = n537 & n827 ;
  assign n829 = ~n824 & ~n828 ;
  assign n833 = ~\P1_reg3_reg[16]/NET0131  & ~n789 ;
  assign n834 = ~n790 & ~n833 ;
  assign n835 = n669 & n834 ;
  assign n832 = \P1_reg2_reg[16]/NET0131  & n667 ;
  assign n830 = \P1_reg1_reg[16]/NET0131  & n663 ;
  assign n831 = \P1_reg0_reg[16]/NET0131  & n665 ;
  assign n836 = ~n830 & ~n831 ;
  assign n837 = ~n832 & n836 ;
  assign n838 = ~n835 & n837 ;
  assign n839 = n829 & ~n838 ;
  assign n840 = ~n798 & ~n839 ;
  assign n841 = ~n797 & ~n840 ;
  assign n842 = n754 & n841 ;
  assign n843 = n743 & ~n752 ;
  assign n844 = n638 & ~n692 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = ~n693 & ~n845 ;
  assign n847 = ~n842 & ~n846 ;
  assign n848 = \P2_datao_reg[22]/NET0131  & n542 ;
  assign n869 = ~n867 & ~n868 ;
  assign n871 = n866 & ~n869 ;
  assign n870 = ~n866 & n869 ;
  assign n872 = ~n542 & ~n870 ;
  assign n873 = ~n871 & n872 ;
  assign n874 = ~n848 & ~n873 ;
  assign n875 = ~n537 & ~n874 ;
  assign n880 = n685 & n879 ;
  assign n881 = ~\P1_reg3_reg[22]/NET0131  & ~n880 ;
  assign n882 = \P1_reg3_reg[22]/NET0131  & n880 ;
  assign n883 = ~n881 & ~n882 ;
  assign n884 = n669 & n883 ;
  assign n878 = \P1_reg0_reg[22]/NET0131  & n665 ;
  assign n876 = \P1_reg1_reg[22]/NET0131  & n663 ;
  assign n877 = \P1_reg2_reg[22]/NET0131  & n667 ;
  assign n885 = ~n876 & ~n877 ;
  assign n886 = ~n878 & n885 ;
  assign n887 = ~n884 & n886 ;
  assign n888 = n875 & n887 ;
  assign n889 = \P2_datao_reg[23]/NET0131  & n542 ;
  assign n905 = ~n903 & ~n904 ;
  assign n907 = n902 & ~n905 ;
  assign n906 = ~n902 & n905 ;
  assign n908 = ~n542 & ~n906 ;
  assign n909 = ~n907 & n908 ;
  assign n910 = ~n889 & ~n909 ;
  assign n911 = ~n537 & ~n910 ;
  assign n915 = ~\P1_reg3_reg[23]/NET0131  & ~n882 ;
  assign n916 = \P1_reg3_reg[23]/NET0131  & n882 ;
  assign n917 = ~n915 & ~n916 ;
  assign n918 = n669 & n917 ;
  assign n914 = \P1_reg2_reg[23]/NET0131  & n667 ;
  assign n912 = \P1_reg1_reg[23]/NET0131  & n663 ;
  assign n913 = \P1_reg0_reg[23]/NET0131  & n665 ;
  assign n919 = ~n912 & ~n913 ;
  assign n920 = ~n914 & n919 ;
  assign n921 = ~n918 & n920 ;
  assign n922 = n911 & n921 ;
  assign n923 = ~n888 & ~n922 ;
  assign n924 = \P2_datao_reg[21]/NET0131  & n542 ;
  assign n933 = ~n849 & ~n856 ;
  assign n935 = n932 & ~n933 ;
  assign n934 = ~n932 & n933 ;
  assign n936 = ~n542 & ~n934 ;
  assign n937 = ~n935 & n936 ;
  assign n938 = ~n924 & ~n937 ;
  assign n939 = ~n537 & ~n938 ;
  assign n943 = \P1_reg3_reg[20]/NET0131  & n685 ;
  assign n944 = ~\P1_reg3_reg[21]/NET0131  & ~n943 ;
  assign n945 = ~n880 & ~n944 ;
  assign n946 = n669 & n945 ;
  assign n942 = \P1_reg2_reg[21]/NET0131  & n667 ;
  assign n940 = \P1_reg1_reg[21]/NET0131  & n663 ;
  assign n941 = \P1_reg0_reg[21]/NET0131  & n665 ;
  assign n947 = ~n940 & ~n941 ;
  assign n948 = ~n942 & n947 ;
  assign n949 = ~n946 & n948 ;
  assign n950 = n939 & n949 ;
  assign n951 = ~n939 & ~n949 ;
  assign n952 = \P2_datao_reg[20]/NET0131  & n542 ;
  assign n958 = ~n850 & ~n857 ;
  assign n960 = n957 & ~n958 ;
  assign n959 = ~n957 & n958 ;
  assign n961 = ~n542 & ~n959 ;
  assign n962 = ~n960 & n961 ;
  assign n963 = ~n952 & ~n962 ;
  assign n964 = ~n537 & ~n963 ;
  assign n968 = ~\P1_reg3_reg[20]/NET0131  & ~n685 ;
  assign n969 = ~n943 & ~n968 ;
  assign n970 = n669 & n969 ;
  assign n967 = \P1_reg0_reg[20]/NET0131  & n665 ;
  assign n965 = \P1_reg2_reg[20]/NET0131  & n667 ;
  assign n966 = \P1_reg1_reg[20]/NET0131  & n663 ;
  assign n971 = ~n965 & ~n966 ;
  assign n972 = ~n967 & n971 ;
  assign n973 = ~n970 & n972 ;
  assign n974 = ~n964 & ~n973 ;
  assign n975 = ~n951 & ~n974 ;
  assign n976 = ~n950 & ~n975 ;
  assign n977 = n923 & n976 ;
  assign n978 = ~n911 & ~n921 ;
  assign n979 = ~n875 & ~n887 ;
  assign n980 = ~n978 & ~n979 ;
  assign n981 = ~n922 & ~n980 ;
  assign n982 = ~n977 & ~n981 ;
  assign n983 = n847 & n982 ;
  assign n984 = n964 & n973 ;
  assign n985 = ~n950 & ~n984 ;
  assign n986 = ~n951 & ~n979 ;
  assign n987 = ~n985 & n986 ;
  assign n988 = n923 & ~n987 ;
  assign n989 = ~n978 & ~n988 ;
  assign n990 = ~n983 & ~n989 ;
  assign n991 = \P1_reg1_reg[15]/NET0131  & n663 ;
  assign n992 = \P1_reg2_reg[15]/NET0131  & n667 ;
  assign n997 = ~n991 & ~n992 ;
  assign n993 = ~\P1_reg3_reg[15]/NET0131  & ~n680 ;
  assign n994 = ~n789 & ~n993 ;
  assign n995 = n669 & n994 ;
  assign n996 = \P1_reg0_reg[15]/NET0131  & n665 ;
  assign n998 = ~n995 & ~n996 ;
  assign n999 = n997 & n998 ;
  assign n1000 = \P2_datao_reg[15]/NET0131  & n542 ;
  assign n1001 = ~n613 & ~n622 ;
  assign n1003 = n608 & ~n1001 ;
  assign n1002 = ~n608 & n1001 ;
  assign n1004 = ~n542 & ~n1002 ;
  assign n1005 = ~n1003 & n1004 ;
  assign n1006 = ~n1000 & ~n1005 ;
  assign n1007 = ~n537 & ~n1006 ;
  assign n1008 = \P1_IR_reg[31]/NET0131  & ~n471 ;
  assign n1009 = \P1_IR_reg[31]/NET0131  & ~n508 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = \P1_IR_reg[15]/NET0131  & ~n1010 ;
  assign n1012 = ~\P1_IR_reg[15]/NET0131  & n1010 ;
  assign n1013 = ~n1011 & ~n1012 ;
  assign n1014 = n537 & n1013 ;
  assign n1015 = ~n1007 & ~n1014 ;
  assign n1016 = n999 & ~n1015 ;
  assign n1017 = \P1_reg2_reg[14]/NET0131  & n667 ;
  assign n1018 = \P1_reg0_reg[14]/NET0131  & n665 ;
  assign n1024 = ~n1017 & ~n1018 ;
  assign n1019 = \P1_reg3_reg[13]/NET0131  & n678 ;
  assign n1020 = ~\P1_reg3_reg[14]/NET0131  & ~n1019 ;
  assign n1021 = ~n680 & ~n1020 ;
  assign n1022 = n669 & n1021 ;
  assign n1023 = \P1_reg1_reg[14]/NET0131  & n663 ;
  assign n1025 = ~n1022 & ~n1023 ;
  assign n1026 = n1024 & n1025 ;
  assign n1027 = \P2_datao_reg[14]/NET0131  & n542 ;
  assign n1028 = ~n544 & ~n545 ;
  assign n1030 = n726 & ~n1028 ;
  assign n1029 = ~n726 & n1028 ;
  assign n1031 = ~n542 & ~n1029 ;
  assign n1032 = ~n1030 & n1031 ;
  assign n1033 = ~n1027 & ~n1032 ;
  assign n1034 = ~n537 & ~n1033 ;
  assign n1035 = \P1_IR_reg[31]/NET0131  & ~n489 ;
  assign n1036 = \P1_IR_reg[14]/NET0131  & ~n1035 ;
  assign n1037 = ~\P1_IR_reg[14]/NET0131  & n1035 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = n537 & ~n1038 ;
  assign n1040 = ~n1034 & ~n1039 ;
  assign n1041 = n1026 & ~n1040 ;
  assign n1042 = ~n1016 & ~n1041 ;
  assign n1043 = \P1_reg0_reg[13]/NET0131  & n665 ;
  assign n1044 = ~\P1_reg3_reg[13]/NET0131  & ~n678 ;
  assign n1045 = ~n1019 & ~n1044 ;
  assign n1046 = n669 & n1045 ;
  assign n1049 = ~n1043 & ~n1046 ;
  assign n1047 = \P1_reg2_reg[13]/NET0131  & n667 ;
  assign n1048 = \P1_reg1_reg[13]/NET0131  & n663 ;
  assign n1050 = ~n1047 & ~n1048 ;
  assign n1051 = n1049 & n1050 ;
  assign n1052 = \P2_datao_reg[13]/NET0131  & n542 ;
  assign n1053 = ~n546 & ~n550 ;
  assign n1055 = n771 & ~n1053 ;
  assign n1054 = ~n771 & n1053 ;
  assign n1056 = ~n542 & ~n1054 ;
  assign n1057 = ~n1055 & n1056 ;
  assign n1058 = ~n1052 & ~n1057 ;
  assign n1059 = ~n537 & ~n1058 ;
  assign n1060 = ~\P1_IR_reg[13]/NET0131  & ~n651 ;
  assign n1061 = \P1_IR_reg[13]/NET0131  & n651 ;
  assign n1062 = ~n1060 & ~n1061 ;
  assign n1063 = n537 & n1062 ;
  assign n1064 = ~n1059 & ~n1063 ;
  assign n1065 = n1051 & ~n1064 ;
  assign n1066 = ~n1051 & n1064 ;
  assign n1067 = ~\P1_reg3_reg[12]/NET0131  & ~n677 ;
  assign n1068 = ~n678 & ~n1067 ;
  assign n1069 = n669 & n1068 ;
  assign n1070 = \P1_reg1_reg[12]/NET0131  & n663 ;
  assign n1073 = ~n1069 & ~n1070 ;
  assign n1071 = \P1_reg2_reg[12]/NET0131  & n667 ;
  assign n1072 = \P1_reg0_reg[12]/NET0131  & n665 ;
  assign n1074 = ~n1071 & ~n1072 ;
  assign n1075 = n1073 & n1074 ;
  assign n1076 = \P2_datao_reg[12]/NET0131  & n542 ;
  assign n1077 = ~n549 & ~n553 ;
  assign n1078 = ~n807 & n813 ;
  assign n1080 = ~n1077 & n1078 ;
  assign n1079 = n1077 & ~n1078 ;
  assign n1081 = ~n542 & ~n1079 ;
  assign n1082 = ~n1080 & n1081 ;
  assign n1083 = ~n1076 & ~n1082 ;
  assign n1084 = ~n537 & ~n1083 ;
  assign n1085 = n462 & n470 ;
  assign n1086 = \P1_IR_reg[31]/NET0131  & ~n1085 ;
  assign n1087 = ~\P1_IR_reg[10]/NET0131  & ~\P1_IR_reg[11]/NET0131  ;
  assign n1088 = \P1_IR_reg[31]/NET0131  & ~n1087 ;
  assign n1089 = ~n1086 & ~n1088 ;
  assign n1090 = \P1_IR_reg[12]/NET0131  & ~n1089 ;
  assign n1091 = ~\P1_IR_reg[12]/NET0131  & n1089 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1093 = n537 & n1092 ;
  assign n1094 = ~n1084 & ~n1093 ;
  assign n1095 = ~n1075 & n1094 ;
  assign n1096 = ~n1066 & ~n1095 ;
  assign n1097 = ~n1065 & ~n1096 ;
  assign n1098 = n1042 & n1097 ;
  assign n1099 = ~n1026 & n1040 ;
  assign n1100 = ~n999 & n1015 ;
  assign n1101 = ~n1099 & ~n1100 ;
  assign n1102 = ~n1016 & ~n1101 ;
  assign n1103 = ~n1098 & ~n1102 ;
  assign n1104 = n1075 & ~n1094 ;
  assign n1105 = ~n1065 & ~n1104 ;
  assign n1106 = n1042 & n1105 ;
  assign n1107 = \P1_reg0_reg[11]/NET0131  & n665 ;
  assign n1108 = \P1_reg1_reg[11]/NET0131  & n663 ;
  assign n1113 = ~n1107 & ~n1108 ;
  assign n1109 = \P1_reg2_reg[11]/NET0131  & n667 ;
  assign n1110 = ~\P1_reg3_reg[11]/NET0131  & ~n676 ;
  assign n1111 = ~n677 & ~n1110 ;
  assign n1112 = n669 & n1111 ;
  assign n1114 = ~n1109 & ~n1112 ;
  assign n1115 = n1113 & n1114 ;
  assign n1116 = \P2_datao_reg[11]/NET0131  & n542 ;
  assign n1117 = ~n554 & ~n604 ;
  assign n1119 = n603 & ~n1117 ;
  assign n1118 = ~n603 & n1117 ;
  assign n1120 = ~n542 & ~n1118 ;
  assign n1121 = ~n1119 & n1120 ;
  assign n1122 = ~n1116 & ~n1121 ;
  assign n1123 = ~n537 & ~n1122 ;
  assign n1124 = ~\P1_IR_reg[11]/NET0131  & ~n1008 ;
  assign n1125 = \P1_IR_reg[11]/NET0131  & n1008 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = n537 & n1126 ;
  assign n1128 = ~n1123 & ~n1127 ;
  assign n1129 = n1115 & ~n1128 ;
  assign n1130 = \P1_reg0_reg[10]/NET0131  & n665 ;
  assign n1131 = ~\P1_reg3_reg[10]/NET0131  & ~n675 ;
  assign n1132 = ~n676 & ~n1131 ;
  assign n1133 = n669 & n1132 ;
  assign n1136 = ~n1130 & ~n1133 ;
  assign n1134 = \P1_reg1_reg[10]/NET0131  & n663 ;
  assign n1135 = \P1_reg2_reg[10]/NET0131  & n667 ;
  assign n1137 = ~n1134 & ~n1135 ;
  assign n1138 = n1136 & n1137 ;
  assign n1139 = \P2_datao_reg[10]/NET0131  & n542 ;
  assign n1140 = ~n557 & ~n558 ;
  assign n1142 = n716 & ~n1140 ;
  assign n1141 = ~n716 & n1140 ;
  assign n1143 = ~n542 & ~n1141 ;
  assign n1144 = ~n1142 & n1143 ;
  assign n1145 = ~n1139 & ~n1144 ;
  assign n1146 = ~n537 & ~n1145 ;
  assign n1147 = \P1_IR_reg[10]/NET0131  & ~n1086 ;
  assign n1148 = ~\P1_IR_reg[10]/NET0131  & n1086 ;
  assign n1149 = ~n1147 & ~n1148 ;
  assign n1150 = n537 & ~n1149 ;
  assign n1151 = ~n1146 & ~n1150 ;
  assign n1152 = n1138 & ~n1151 ;
  assign n1153 = ~n1129 & ~n1152 ;
  assign n1154 = \P1_reg2_reg[9]/NET0131  & n667 ;
  assign n1155 = \P1_reg1_reg[9]/NET0131  & n663 ;
  assign n1160 = ~n1154 & ~n1155 ;
  assign n1156 = \P1_reg0_reg[9]/NET0131  & n665 ;
  assign n1157 = ~\P1_reg3_reg[9]/NET0131  & ~n674 ;
  assign n1158 = ~n675 & ~n1157 ;
  assign n1159 = n669 & n1158 ;
  assign n1161 = ~n1156 & ~n1159 ;
  assign n1162 = n1160 & n1161 ;
  assign n1163 = \P2_datao_reg[9]/NET0131  & n542 ;
  assign n1164 = ~n559 & ~n562 ;
  assign n1166 = n768 & ~n1164 ;
  assign n1165 = ~n768 & n1164 ;
  assign n1167 = ~n542 & ~n1165 ;
  assign n1168 = ~n1166 & n1167 ;
  assign n1169 = ~n1163 & ~n1168 ;
  assign n1170 = ~n537 & ~n1169 ;
  assign n1171 = \P1_IR_reg[31]/NET0131  & ~n470 ;
  assign n1172 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[8]/NET0131  ;
  assign n1173 = ~n1171 & ~n1172 ;
  assign n1174 = \P1_IR_reg[9]/NET0131  & ~n1173 ;
  assign n1175 = ~\P1_IR_reg[9]/NET0131  & n1173 ;
  assign n1176 = ~n1174 & ~n1175 ;
  assign n1177 = n537 & n1176 ;
  assign n1178 = ~n1170 & ~n1177 ;
  assign n1179 = n1162 & ~n1178 ;
  assign n1180 = ~n1162 & n1178 ;
  assign n1181 = ~\P1_reg3_reg[8]/NET0131  & ~n673 ;
  assign n1182 = ~n674 & ~n1181 ;
  assign n1183 = n669 & n1182 ;
  assign n1184 = \P1_reg2_reg[8]/NET0131  & n667 ;
  assign n1187 = ~n1183 & ~n1184 ;
  assign n1185 = \P1_reg1_reg[8]/NET0131  & n663 ;
  assign n1186 = \P1_reg0_reg[8]/NET0131  & n665 ;
  assign n1188 = ~n1185 & ~n1186 ;
  assign n1189 = n1187 & n1188 ;
  assign n1190 = \P2_datao_reg[8]/NET0131  & n542 ;
  assign n1191 = ~n564 & ~n566 ;
  assign n1193 = n805 & n1191 ;
  assign n1192 = ~n805 & ~n1191 ;
  assign n1194 = ~n542 & ~n1192 ;
  assign n1195 = ~n1193 & n1194 ;
  assign n1196 = ~n1190 & ~n1195 ;
  assign n1197 = ~n537 & ~n1196 ;
  assign n1198 = \P1_IR_reg[8]/NET0131  & ~n1171 ;
  assign n1199 = ~\P1_IR_reg[8]/NET0131  & n1171 ;
  assign n1200 = ~n1198 & ~n1199 ;
  assign n1201 = n537 & ~n1200 ;
  assign n1202 = ~n1197 & ~n1201 ;
  assign n1203 = ~n1189 & n1202 ;
  assign n1204 = ~n1180 & ~n1203 ;
  assign n1205 = ~n1179 & ~n1204 ;
  assign n1206 = n1153 & n1205 ;
  assign n1207 = ~n1138 & n1151 ;
  assign n1208 = ~n1115 & n1128 ;
  assign n1209 = ~n1207 & ~n1208 ;
  assign n1210 = ~n1129 & ~n1209 ;
  assign n1211 = ~n1206 & ~n1210 ;
  assign n1212 = n1106 & ~n1211 ;
  assign n1213 = n1103 & ~n1212 ;
  assign n1214 = \P1_reg0_reg[6]/NET0131  & n665 ;
  assign n1215 = \P1_reg2_reg[6]/NET0131  & n667 ;
  assign n1220 = ~n1214 & ~n1215 ;
  assign n1216 = \P1_reg1_reg[6]/NET0131  & n663 ;
  assign n1217 = ~\P1_reg3_reg[6]/NET0131  & ~n671 ;
  assign n1218 = ~n672 & ~n1217 ;
  assign n1219 = n669 & n1218 ;
  assign n1221 = ~n1216 & ~n1219 ;
  assign n1222 = n1220 & n1221 ;
  assign n1223 = \P2_datao_reg[6]/NET0131  & n542 ;
  assign n1224 = ~n579 & ~n587 ;
  assign n1225 = ~n580 & ~n712 ;
  assign n1227 = n1224 & n1225 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1228 = ~n542 & ~n1226 ;
  assign n1229 = ~n1227 & n1228 ;
  assign n1230 = ~n1223 & ~n1229 ;
  assign n1231 = ~n537 & ~n1230 ;
  assign n1232 = ~\P1_IR_reg[5]/NET0131  & n467 ;
  assign n1233 = \P1_IR_reg[31]/NET0131  & ~n1232 ;
  assign n1234 = ~\P1_IR_reg[6]/NET0131  & ~n1233 ;
  assign n1235 = \P1_IR_reg[6]/NET0131  & n1233 ;
  assign n1236 = ~n1234 & ~n1235 ;
  assign n1237 = n537 & n1236 ;
  assign n1238 = ~n1231 & ~n1237 ;
  assign n1239 = n1222 & ~n1238 ;
  assign n1240 = \P1_reg0_reg[7]/NET0131  & n665 ;
  assign n1241 = \P1_reg2_reg[7]/NET0131  & n667 ;
  assign n1246 = ~n1240 & ~n1241 ;
  assign n1242 = ~\P1_reg3_reg[7]/NET0131  & ~n672 ;
  assign n1243 = ~n673 & ~n1242 ;
  assign n1244 = n669 & n1243 ;
  assign n1245 = \P1_reg1_reg[7]/NET0131  & n663 ;
  assign n1247 = ~n1244 & ~n1245 ;
  assign n1248 = n1246 & n1247 ;
  assign n1249 = \P2_datao_reg[7]/NET0131  & n542 ;
  assign n1250 = ~n567 & ~n598 ;
  assign n1252 = n597 & ~n1250 ;
  assign n1251 = ~n597 & n1250 ;
  assign n1253 = ~n542 & ~n1251 ;
  assign n1254 = ~n1252 & n1253 ;
  assign n1255 = ~n1249 & ~n1254 ;
  assign n1256 = ~n537 & ~n1255 ;
  assign n1257 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[6]/NET0131  ;
  assign n1258 = ~n1233 & ~n1257 ;
  assign n1259 = \P1_IR_reg[7]/NET0131  & ~n1258 ;
  assign n1260 = ~\P1_IR_reg[7]/NET0131  & n1258 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1262 = n537 & n1261 ;
  assign n1263 = ~n1256 & ~n1262 ;
  assign n1264 = n1248 & ~n1263 ;
  assign n1265 = ~n1239 & ~n1264 ;
  assign n1266 = \P1_reg0_reg[5]/NET0131  & n665 ;
  assign n1267 = \P1_reg2_reg[5]/NET0131  & n667 ;
  assign n1272 = ~n1266 & ~n1267 ;
  assign n1268 = \P1_reg1_reg[5]/NET0131  & n663 ;
  assign n1269 = ~\P1_reg3_reg[5]/NET0131  & ~n670 ;
  assign n1270 = ~n671 & ~n1269 ;
  assign n1271 = n669 & n1270 ;
  assign n1273 = ~n1268 & ~n1271 ;
  assign n1274 = n1272 & n1273 ;
  assign n1275 = \P2_datao_reg[5]/NET0131  & n542 ;
  assign n1276 = ~n580 & ~n588 ;
  assign n1278 = n762 & ~n1276 ;
  assign n1277 = ~n762 & n1276 ;
  assign n1279 = ~n542 & ~n1277 ;
  assign n1280 = ~n1278 & n1279 ;
  assign n1281 = ~n1275 & ~n1280 ;
  assign n1282 = ~n537 & ~n1281 ;
  assign n1283 = \P1_IR_reg[31]/NET0131  & ~n467 ;
  assign n1284 = \P1_IR_reg[5]/NET0131  & ~n1283 ;
  assign n1285 = ~\P1_IR_reg[5]/NET0131  & n1283 ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = n537 & ~n1286 ;
  assign n1288 = ~n1282 & ~n1287 ;
  assign n1289 = n1274 & ~n1288 ;
  assign n1290 = ~\P1_reg3_reg[3]/NET0131  & ~\P1_reg3_reg[4]/NET0131  ;
  assign n1291 = ~n670 & ~n1290 ;
  assign n1292 = n669 & n1291 ;
  assign n1293 = \P1_reg1_reg[4]/NET0131  & n663 ;
  assign n1296 = ~n1292 & ~n1293 ;
  assign n1294 = \P1_reg2_reg[4]/NET0131  & n667 ;
  assign n1295 = \P1_reg0_reg[4]/NET0131  & n665 ;
  assign n1297 = ~n1294 & ~n1295 ;
  assign n1298 = n1296 & n1297 ;
  assign n1299 = \P1_IR_reg[31]/NET0131  & ~n466 ;
  assign n1300 = \P1_IR_reg[4]/NET0131  & n1299 ;
  assign n1301 = ~\P1_IR_reg[4]/NET0131  & ~n1299 ;
  assign n1302 = ~n1300 & ~n1301 ;
  assign n1303 = n537 & n1302 ;
  assign n1304 = ~\P2_datao_reg[4]/NET0131  & n542 ;
  assign n1305 = ~n583 & ~n709 ;
  assign n1306 = ~n582 & ~n591 ;
  assign n1308 = ~n1305 & n1306 ;
  assign n1307 = n1305 & ~n1306 ;
  assign n1309 = ~n542 & ~n1307 ;
  assign n1310 = ~n1308 & n1309 ;
  assign n1311 = ~n1304 & ~n1310 ;
  assign n1312 = ~n537 & n1311 ;
  assign n1313 = ~n1303 & ~n1312 ;
  assign n1314 = n1298 & ~n1313 ;
  assign n1315 = ~n1289 & ~n1314 ;
  assign n1316 = \P1_reg0_reg[3]/NET0131  & n665 ;
  assign n1317 = ~\P1_reg3_reg[3]/NET0131  & n669 ;
  assign n1320 = ~n1316 & ~n1317 ;
  assign n1318 = \P1_reg1_reg[3]/NET0131  & n663 ;
  assign n1319 = \P1_reg2_reg[3]/NET0131  & n667 ;
  assign n1321 = ~n1318 & ~n1319 ;
  assign n1322 = n1320 & n1321 ;
  assign n1323 = \P2_datao_reg[3]/NET0131  & n542 ;
  assign n1324 = ~n583 & ~n592 ;
  assign n1326 = n578 & ~n1324 ;
  assign n1325 = ~n578 & n1324 ;
  assign n1327 = ~n542 & ~n1325 ;
  assign n1328 = ~n1326 & n1327 ;
  assign n1329 = ~n1323 & ~n1328 ;
  assign n1330 = ~n537 & ~n1329 ;
  assign n1331 = \P1_IR_reg[31]/NET0131  & ~n465 ;
  assign n1332 = \P1_IR_reg[3]/NET0131  & n1331 ;
  assign n1333 = ~\P1_IR_reg[3]/NET0131  & ~n1331 ;
  assign n1334 = ~n1332 & ~n1333 ;
  assign n1335 = n537 & n1334 ;
  assign n1336 = ~n1330 & ~n1335 ;
  assign n1337 = n1322 & ~n1336 ;
  assign n1338 = \P1_reg0_reg[2]/NET0131  & n665 ;
  assign n1339 = \P1_reg1_reg[2]/NET0131  & n663 ;
  assign n1342 = ~n1338 & ~n1339 ;
  assign n1340 = \P1_reg2_reg[2]/NET0131  & n667 ;
  assign n1341 = \P1_reg3_reg[2]/NET0131  & n669 ;
  assign n1343 = ~n1340 & ~n1341 ;
  assign n1344 = n1342 & n1343 ;
  assign n1345 = \P2_datao_reg[2]/NET0131  & n542 ;
  assign n1346 = ~n570 & ~n577 ;
  assign n1348 = n575 & n1346 ;
  assign n1347 = ~n575 & ~n1346 ;
  assign n1349 = ~n542 & ~n1347 ;
  assign n1350 = ~n1348 & n1349 ;
  assign n1351 = ~n1345 & ~n1350 ;
  assign n1352 = ~n537 & ~n1351 ;
  assign n1353 = \P1_IR_reg[31]/NET0131  & ~n464 ;
  assign n1354 = ~\P1_IR_reg[2]/NET0131  & ~n1353 ;
  assign n1355 = \P1_IR_reg[2]/NET0131  & n1353 ;
  assign n1356 = ~n1354 & ~n1355 ;
  assign n1357 = n537 & n1356 ;
  assign n1358 = ~n1352 & ~n1357 ;
  assign n1359 = n1344 & ~n1358 ;
  assign n1360 = ~n1337 & ~n1359 ;
  assign n1361 = \P1_reg3_reg[1]/NET0131  & n669 ;
  assign n1362 = \P1_reg2_reg[1]/NET0131  & n667 ;
  assign n1365 = ~n1361 & ~n1362 ;
  assign n1363 = \P1_reg1_reg[1]/NET0131  & n663 ;
  assign n1364 = \P1_reg0_reg[1]/NET0131  & n665 ;
  assign n1366 = ~n1363 & ~n1364 ;
  assign n1367 = n1365 & n1366 ;
  assign n1368 = \P1_IR_reg[1]/NET0131  & ~\P1_IR_reg[31]/NET0131  ;
  assign n1369 = \P1_IR_reg[0]/NET0131  & \P1_IR_reg[1]/NET0131  ;
  assign n1370 = n1353 & ~n1369 ;
  assign n1371 = ~n1368 & ~n1370 ;
  assign n1372 = n537 & ~n1371 ;
  assign n1373 = ~\P2_datao_reg[1]/NET0131  & n542 ;
  assign n1374 = ~n571 & ~n572 ;
  assign n1376 = ~n573 & n1374 ;
  assign n1375 = n573 & ~n1374 ;
  assign n1377 = ~n542 & ~n1375 ;
  assign n1378 = ~n1376 & n1377 ;
  assign n1379 = ~n1373 & ~n1378 ;
  assign n1380 = ~n537 & n1379 ;
  assign n1381 = ~n1372 & ~n1380 ;
  assign n1382 = ~n1367 & n1381 ;
  assign n1383 = n1367 & ~n1381 ;
  assign n1384 = \P1_reg1_reg[0]/NET0131  & n663 ;
  assign n1385 = \P1_reg0_reg[0]/NET0131  & n665 ;
  assign n1388 = ~n1384 & ~n1385 ;
  assign n1386 = \P1_reg3_reg[0]/NET0131  & n669 ;
  assign n1387 = \P1_reg2_reg[0]/NET0131  & n667 ;
  assign n1389 = ~n1386 & ~n1387 ;
  assign n1390 = n1388 & n1389 ;
  assign n1391 = \si[0]_pad  & ~n542 ;
  assign n1392 = ~\P2_datao_reg[0]/NET0131  & ~n1391 ;
  assign n1393 = ~n542 & n573 ;
  assign n1394 = ~n1392 & ~n1393 ;
  assign n1395 = ~n537 & n1394 ;
  assign n1396 = \P1_IR_reg[0]/NET0131  & n537 ;
  assign n1397 = ~n1395 & ~n1396 ;
  assign n1398 = n1390 & ~n1397 ;
  assign n1399 = ~n1383 & ~n1398 ;
  assign n1400 = ~n1382 & ~n1399 ;
  assign n1401 = n1360 & ~n1400 ;
  assign n1402 = ~n1322 & n1336 ;
  assign n1403 = ~n1344 & n1358 ;
  assign n1404 = ~n1337 & n1403 ;
  assign n1405 = ~n1402 & ~n1404 ;
  assign n1406 = ~n1401 & n1405 ;
  assign n1407 = n1315 & ~n1406 ;
  assign n1408 = n1265 & n1407 ;
  assign n1409 = ~n1274 & n1288 ;
  assign n1410 = ~n1298 & n1313 ;
  assign n1411 = ~n1289 & n1410 ;
  assign n1412 = ~n1409 & ~n1411 ;
  assign n1413 = n1265 & ~n1412 ;
  assign n1414 = ~n1248 & n1263 ;
  assign n1415 = ~n1222 & n1238 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = ~n1264 & ~n1416 ;
  assign n1418 = ~n1413 & ~n1417 ;
  assign n1419 = ~n1408 & n1418 ;
  assign n1420 = n1189 & ~n1202 ;
  assign n1421 = ~n1179 & ~n1420 ;
  assign n1422 = n1153 & n1421 ;
  assign n1423 = ~n1419 & n1422 ;
  assign n1424 = n1106 & n1423 ;
  assign n1425 = n1213 & ~n1424 ;
  assign n1426 = n923 & n985 ;
  assign n1427 = ~n829 & n838 ;
  assign n1428 = ~n797 & ~n1427 ;
  assign n1429 = n754 & n1428 ;
  assign n1430 = n1426 & n1429 ;
  assign n1431 = ~n1425 & n1430 ;
  assign n1432 = ~n990 & ~n1431 ;
  assign n1433 = \P2_datao_reg[26]/NET0131  & n542 ;
  assign n1436 = ~n1434 & ~n1435 ;
  assign n1450 = n720 & n854 ;
  assign n1451 = ~n725 & n728 ;
  assign n1452 = n702 & ~n1451 ;
  assign n1453 = n853 & ~n1452 ;
  assign n1454 = n863 & ~n1453 ;
  assign n1455 = ~n1450 & n1454 ;
  assign n1456 = n1449 & ~n1455 ;
  assign n1457 = n1447 & ~n1456 ;
  assign n1459 = ~n1436 & n1457 ;
  assign n1458 = n1436 & ~n1457 ;
  assign n1460 = ~n542 & ~n1458 ;
  assign n1461 = ~n1459 & n1460 ;
  assign n1462 = ~n1433 & ~n1461 ;
  assign n1463 = ~n537 & ~n1462 ;
  assign n1473 = ~\P1_reg3_reg[26]/NET0131  & ~n1471 ;
  assign n1474 = ~n1472 & ~n1473 ;
  assign n1475 = n669 & n1474 ;
  assign n1466 = \P1_reg1_reg[26]/NET0131  & n663 ;
  assign n1464 = \P1_reg0_reg[26]/NET0131  & n665 ;
  assign n1465 = \P1_reg2_reg[26]/NET0131  & n667 ;
  assign n1476 = ~n1464 & ~n1465 ;
  assign n1477 = ~n1466 & n1476 ;
  assign n1478 = ~n1475 & n1477 ;
  assign n1479 = n1463 & n1478 ;
  assign n1480 = \P2_datao_reg[27]/NET0131  & n542 ;
  assign n1483 = ~n1481 & ~n1482 ;
  assign n1491 = ~n627 & n892 ;
  assign n1492 = n899 & ~n1491 ;
  assign n1493 = n1490 & ~n1492 ;
  assign n1494 = n1489 & ~n1493 ;
  assign n1496 = ~n1483 & n1494 ;
  assign n1495 = n1483 & ~n1494 ;
  assign n1497 = ~n542 & ~n1495 ;
  assign n1498 = ~n1496 & n1497 ;
  assign n1499 = ~n1480 & ~n1498 ;
  assign n1500 = ~n537 & ~n1499 ;
  assign n1505 = ~\P1_reg3_reg[27]/NET0131  & ~n1472 ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = n669 & n1506 ;
  assign n1503 = \P1_reg2_reg[27]/NET0131  & n667 ;
  assign n1501 = \P1_reg0_reg[27]/NET0131  & n665 ;
  assign n1502 = \P1_reg1_reg[27]/NET0131  & n663 ;
  assign n1508 = ~n1501 & ~n1502 ;
  assign n1509 = ~n1503 & n1508 ;
  assign n1510 = ~n1507 & n1509 ;
  assign n1511 = n1500 & n1510 ;
  assign n1512 = ~n1479 & ~n1511 ;
  assign n1513 = \P2_datao_reg[25]/NET0131  & n542 ;
  assign n1514 = ~n1437 & ~n1438 ;
  assign n1517 = ~n1442 & ~n1516 ;
  assign n1521 = n770 & n926 ;
  assign n1518 = ~n761 & n772 ;
  assign n1519 = n758 & ~n1518 ;
  assign n1520 = n925 & ~n1519 ;
  assign n1522 = n929 & ~n1520 ;
  assign n1523 = ~n1521 & n1522 ;
  assign n1524 = ~n903 & ~n1442 ;
  assign n1525 = n890 & n1524 ;
  assign n1526 = ~n1523 & n1525 ;
  assign n1527 = ~n1517 & ~n1526 ;
  assign n1529 = ~n1514 & n1527 ;
  assign n1528 = n1514 & ~n1527 ;
  assign n1530 = ~n542 & ~n1528 ;
  assign n1531 = ~n1529 & n1530 ;
  assign n1532 = ~n1513 & ~n1531 ;
  assign n1533 = ~n537 & ~n1532 ;
  assign n1537 = ~\P1_reg3_reg[25]/NET0131  & ~n1470 ;
  assign n1538 = ~n1471 & ~n1537 ;
  assign n1539 = n669 & n1538 ;
  assign n1536 = \P1_reg2_reg[25]/NET0131  & n667 ;
  assign n1534 = \P1_reg1_reg[25]/NET0131  & n663 ;
  assign n1535 = \P1_reg0_reg[25]/NET0131  & n665 ;
  assign n1540 = ~n1534 & ~n1535 ;
  assign n1541 = ~n1536 & n1540 ;
  assign n1542 = ~n1539 & n1541 ;
  assign n1543 = n1533 & n1542 ;
  assign n1544 = \P2_datao_reg[24]/NET0131  & n542 ;
  assign n1545 = ~n1439 & ~n1442 ;
  assign n1552 = n955 & n1548 ;
  assign n1553 = n808 & n1552 ;
  assign n1549 = ~n816 & n955 ;
  assign n1550 = n954 & ~n1549 ;
  assign n1551 = n1548 & ~n1550 ;
  assign n1554 = n1547 & ~n1551 ;
  assign n1555 = ~n1553 & n1554 ;
  assign n1557 = ~n1545 & n1555 ;
  assign n1556 = n1545 & ~n1555 ;
  assign n1558 = ~n542 & ~n1556 ;
  assign n1559 = ~n1557 & n1558 ;
  assign n1560 = ~n1544 & ~n1559 ;
  assign n1561 = ~n537 & ~n1560 ;
  assign n1562 = ~\P1_reg3_reg[24]/NET0131  & ~n916 ;
  assign n1563 = ~n1470 & ~n1562 ;
  assign n1564 = n669 & n1563 ;
  assign n1567 = \P1_reg0_reg[24]/NET0131  & n665 ;
  assign n1565 = \P1_reg2_reg[24]/NET0131  & n667 ;
  assign n1566 = \P1_reg1_reg[24]/NET0131  & n663 ;
  assign n1568 = ~n1565 & ~n1566 ;
  assign n1569 = ~n1567 & n1568 ;
  assign n1570 = ~n1564 & n1569 ;
  assign n1571 = n1561 & n1570 ;
  assign n1572 = ~n1543 & ~n1571 ;
  assign n1573 = n1512 & n1572 ;
  assign n1574 = ~n1432 & n1573 ;
  assign n1575 = ~n1500 & ~n1510 ;
  assign n1576 = ~n1463 & ~n1478 ;
  assign n1577 = ~n1533 & ~n1542 ;
  assign n1578 = ~n1561 & ~n1570 ;
  assign n1579 = ~n1543 & n1578 ;
  assign n1580 = ~n1577 & ~n1579 ;
  assign n1581 = ~n1576 & n1580 ;
  assign n1582 = n1512 & ~n1581 ;
  assign n1583 = ~n1575 & ~n1582 ;
  assign n1584 = ~n1574 & n1583 ;
  assign n1647 = n1637 & n1646 ;
  assign n1648 = ~n1619 & ~n1647 ;
  assign n1649 = ~n1584 & n1648 ;
  assign n1729 = n1649 & n1724 ;
  assign n1730 = n1728 & ~n1729 ;
  assign n1918 = ~\P1_B_reg/NET0131  & n1730 ;
  assign n482 = \P1_IR_reg[31]/NET0131  & ~n481 ;
  assign n483 = ~n478 & ~n482 ;
  assign n484 = \P1_IR_reg[21]/NET0131  & ~n483 ;
  assign n485 = ~\P1_IR_reg[21]/NET0131  & n483 ;
  assign n486 = ~n484 & ~n485 ;
  assign n502 = \P1_IR_reg[31]/NET0131  & ~n501 ;
  assign n503 = ~n491 & ~n502 ;
  assign n504 = \P1_IR_reg[22]/NET0131  & ~n503 ;
  assign n505 = ~\P1_IR_reg[22]/NET0131  & n503 ;
  assign n506 = ~n504 & ~n505 ;
  assign n494 = \P1_IR_reg[31]/NET0131  & ~n493 ;
  assign n495 = ~n491 & ~n494 ;
  assign n496 = \P1_IR_reg[20]/NET0131  & ~n495 ;
  assign n497 = ~\P1_IR_reg[20]/NET0131  & n495 ;
  assign n498 = ~n496 & ~n497 ;
  assign n1734 = ~n498 & ~n516 ;
  assign n1901 = n506 & n1734 ;
  assign n1919 = ~n486 & n1901 ;
  assign n1920 = ~n1918 & n1919 ;
  assign n1703 = ~n1677 & ~n1702 ;
  assign n1704 = n1696 & ~n1703 ;
  assign n1705 = ~n1678 & ~n1704 ;
  assign n1706 = n1649 & n1705 ;
  assign n1708 = ~n1677 & ~n1707 ;
  assign n1709 = n1671 & ~n1708 ;
  assign n1713 = ~n1711 & ~n1712 ;
  assign n1714 = n1705 & ~n1713 ;
  assign n1715 = ~n1709 & ~n1714 ;
  assign n1716 = ~n1706 & n1715 ;
  assign n1910 = ~\P1_B_reg/NET0131  & n1716 ;
  assign n499 = n486 & n498 ;
  assign n1911 = n506 & ~n516 ;
  assign n1912 = n499 & n1911 ;
  assign n1913 = ~n1910 & n1912 ;
  assign n1914 = ~\P1_B_reg/NET0131  & ~n1716 ;
  assign n1915 = n506 & n516 ;
  assign n1916 = n499 & n1915 ;
  assign n1917 = ~n1914 & n1916 ;
  assign n1926 = ~n1913 & ~n1917 ;
  assign n1927 = ~n1920 & n1926 ;
  assign n1718 = ~n516 & n1716 ;
  assign n1717 = n516 & ~n1716 ;
  assign n1719 = n499 & ~n506 ;
  assign n1720 = ~n1717 & n1719 ;
  assign n1721 = ~n1718 & n1720 ;
  assign n1735 = ~n486 & ~n506 ;
  assign n1736 = n1734 & n1735 ;
  assign n1737 = ~n1730 & n1736 ;
  assign n1731 = ~n498 & n516 ;
  assign n1732 = ~n486 & n1731 ;
  assign n1733 = n1730 & n1732 ;
  assign n1842 = ~n1648 & n1725 ;
  assign n1843 = n1724 & ~n1842 ;
  assign n1844 = ~n1722 & ~n1843 ;
  assign n1845 = ~n1576 & ~n1577 ;
  assign n1846 = ~n1572 & n1845 ;
  assign n1847 = n1512 & ~n1846 ;
  assign n1848 = ~n1575 & ~n1847 ;
  assign n1849 = ~n1844 & ~n1848 ;
  assign n1850 = n1728 & ~n1849 ;
  assign n1851 = ~n798 & ~n843 ;
  assign n1852 = ~n1428 & n1851 ;
  assign n1853 = n754 & ~n1852 ;
  assign n1854 = ~n844 & ~n1853 ;
  assign n1855 = ~n989 & ~n1854 ;
  assign n1856 = n982 & ~n1855 ;
  assign n1857 = ~n1066 & ~n1099 ;
  assign n1858 = ~n1105 & n1857 ;
  assign n1859 = n1042 & ~n1858 ;
  assign n1860 = ~n1100 & ~n1859 ;
  assign n1861 = ~n1180 & ~n1207 ;
  assign n1862 = ~n1421 & n1861 ;
  assign n1863 = n1153 & ~n1862 ;
  assign n1864 = ~n1208 & ~n1863 ;
  assign n1865 = ~n1860 & ~n1864 ;
  assign n1866 = n1103 & ~n1865 ;
  assign n1738 = ~n1390 & n1397 ;
  assign n1869 = ~n1383 & n1738 ;
  assign n1870 = ~n1382 & ~n1403 ;
  assign n1871 = ~n1869 & n1870 ;
  assign n1872 = n1360 & ~n1871 ;
  assign n1867 = ~n1409 & ~n1415 ;
  assign n1873 = ~n1402 & ~n1410 ;
  assign n1874 = n1867 & n1873 ;
  assign n1875 = ~n1872 & n1874 ;
  assign n1868 = ~n1315 & n1867 ;
  assign n1876 = n1265 & ~n1868 ;
  assign n1877 = ~n1875 & n1876 ;
  assign n1878 = n1204 & ~n1414 ;
  assign n1879 = n1209 & n1878 ;
  assign n1880 = n1096 & n1879 ;
  assign n1881 = n1101 & n1880 ;
  assign n1882 = ~n1877 & n1881 ;
  assign n1883 = ~n1866 & ~n1882 ;
  assign n1884 = n840 & n845 ;
  assign n1885 = n975 & n980 ;
  assign n1886 = n1884 & n1885 ;
  assign n1887 = ~n1883 & n1886 ;
  assign n1888 = ~n1856 & ~n1887 ;
  assign n1889 = ~n1578 & n1845 ;
  assign n1890 = ~n1710 & n1889 ;
  assign n1891 = n1725 & n1890 ;
  assign n1892 = ~n1575 & ~n1722 ;
  assign n1893 = n1891 & n1892 ;
  assign n1894 = ~n1888 & n1893 ;
  assign n1895 = ~n1850 & ~n1894 ;
  assign n1905 = n516 & n1895 ;
  assign n1904 = ~n516 & ~n1895 ;
  assign n1906 = ~n498 & ~n506 ;
  assign n1907 = n486 & n1906 ;
  assign n1908 = ~n1904 & n1907 ;
  assign n1909 = ~n1905 & n1908 ;
  assign n1791 = ~n1637 & n1646 ;
  assign n1792 = n1637 & ~n1646 ;
  assign n1793 = ~n1791 & ~n1792 ;
  assign n1829 = ~n1678 & ~n1722 ;
  assign n1830 = ~n1793 & n1829 ;
  assign n1788 = n1500 & ~n1510 ;
  assign n1789 = ~n1500 & n1510 ;
  assign n1790 = ~n1788 & ~n1789 ;
  assign n1766 = ~n1065 & ~n1066 ;
  assign n1760 = ~n1075 & ~n1094 ;
  assign n1761 = n1075 & n1094 ;
  assign n1762 = ~n1760 & ~n1761 ;
  assign n1763 = n999 & n1015 ;
  assign n1764 = ~n999 & ~n1015 ;
  assign n1765 = ~n1763 & ~n1764 ;
  assign n1812 = ~n1762 & ~n1765 ;
  assign n1813 = n1766 & n1812 ;
  assign n1747 = n1162 & n1178 ;
  assign n1748 = ~n1162 & ~n1178 ;
  assign n1749 = ~n1747 & ~n1748 ;
  assign n1750 = ~n1129 & ~n1208 ;
  assign n1803 = ~n1749 & n1750 ;
  assign n1751 = ~n1298 & ~n1313 ;
  assign n1752 = n1298 & n1313 ;
  assign n1753 = ~n1751 & ~n1752 ;
  assign n1754 = ~n1152 & ~n1207 ;
  assign n1804 = ~n1753 & n1754 ;
  assign n1808 = n1803 & n1804 ;
  assign n1739 = ~n1398 & ~n1738 ;
  assign n1740 = ~n1239 & ~n1415 ;
  assign n1801 = n1739 & n1740 ;
  assign n1741 = n1248 & n1263 ;
  assign n1742 = ~n1248 & ~n1263 ;
  assign n1743 = ~n1741 & ~n1742 ;
  assign n1744 = n1322 & n1336 ;
  assign n1745 = ~n1322 & ~n1336 ;
  assign n1746 = ~n1744 & ~n1745 ;
  assign n1802 = ~n1743 & ~n1746 ;
  assign n1809 = n1801 & n1802 ;
  assign n1810 = n1808 & n1809 ;
  assign n1756 = ~n1041 & ~n1099 ;
  assign n1755 = ~n1382 & ~n1383 ;
  assign n1757 = ~n1203 & ~n1420 ;
  assign n1805 = n1755 & n1757 ;
  assign n1758 = ~n1289 & ~n1409 ;
  assign n1759 = ~n1359 & ~n1403 ;
  assign n1806 = n1758 & n1759 ;
  assign n1807 = n1805 & n1806 ;
  assign n1811 = n1756 & n1807 ;
  assign n1814 = n1810 & n1811 ;
  assign n1817 = n1813 & n1814 ;
  assign n1818 = ~n1707 & ~n1723 ;
  assign n1825 = n1817 & n1818 ;
  assign n1780 = ~n1619 & ~n1712 ;
  assign n1787 = ~n839 & ~n1427 ;
  assign n1777 = ~n875 & n887 ;
  assign n1778 = n875 & ~n887 ;
  assign n1779 = ~n1777 & ~n1778 ;
  assign n1784 = ~n939 & n949 ;
  assign n1785 = n939 & ~n949 ;
  assign n1786 = ~n1784 & ~n1785 ;
  assign n1815 = ~n1779 & ~n1786 ;
  assign n1816 = n1787 & n1815 ;
  assign n1826 = n1780 & n1816 ;
  assign n1827 = n1825 & n1826 ;
  assign n1781 = ~n1561 & n1570 ;
  assign n1782 = n1561 & ~n1570 ;
  assign n1783 = ~n1781 & ~n1782 ;
  assign n1794 = ~n911 & n921 ;
  assign n1795 = n911 & ~n921 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1821 = ~n1783 & ~n1796 ;
  assign n1797 = ~n743 & ~n752 ;
  assign n1798 = n743 & n752 ;
  assign n1799 = ~n1797 & ~n1798 ;
  assign n1800 = ~n693 & ~n844 ;
  assign n1822 = ~n1799 & n1800 ;
  assign n1823 = n1821 & n1822 ;
  assign n1767 = ~n1533 & n1542 ;
  assign n1768 = n1533 & ~n1542 ;
  assign n1769 = ~n1767 & ~n1768 ;
  assign n1770 = ~n1463 & n1478 ;
  assign n1771 = n1463 & ~n1478 ;
  assign n1772 = ~n1770 & ~n1771 ;
  assign n1819 = ~n1769 & ~n1772 ;
  assign n1773 = ~n797 & ~n798 ;
  assign n1774 = n964 & ~n973 ;
  assign n1775 = ~n964 & n973 ;
  assign n1776 = ~n1774 & ~n1775 ;
  assign n1820 = n1773 & ~n1776 ;
  assign n1824 = n1819 & n1820 ;
  assign n1828 = n1823 & n1824 ;
  assign n1831 = n1827 & n1828 ;
  assign n1832 = ~n1790 & n1831 ;
  assign n1833 = n1830 & n1832 ;
  assign n1834 = ~n516 & ~n1833 ;
  assign n1835 = n516 & n1833 ;
  assign n1836 = ~n1834 & ~n1835 ;
  assign n1837 = n498 & ~n1836 ;
  assign n1838 = \P1_B_reg/NET0131  & n506 ;
  assign n1839 = ~n1734 & n1838 ;
  assign n1840 = ~n1837 & ~n1839 ;
  assign n1841 = ~n486 & ~n1840 ;
  assign n1896 = ~\P1_B_reg/NET0131  & n1895 ;
  assign n1897 = n486 & n506 ;
  assign n1898 = n1731 & n1897 ;
  assign n1899 = ~n1896 & n1898 ;
  assign n1900 = ~\P1_B_reg/NET0131  & ~n1895 ;
  assign n1902 = n486 & n1901 ;
  assign n1903 = ~n1900 & n1902 ;
  assign n1921 = ~n1899 & ~n1903 ;
  assign n1922 = ~n1841 & n1921 ;
  assign n1923 = ~n1909 & n1922 ;
  assign n1924 = ~n1733 & n1923 ;
  assign n1925 = ~n1737 & n1924 ;
  assign n1928 = ~n1721 & n1925 ;
  assign n1929 = n1927 & n1928 ;
  assign n1930 = \P1_IR_reg[31]/NET0131  & ~n521 ;
  assign n1931 = \P1_IR_reg[23]/NET0131  & n1930 ;
  assign n1932 = ~\P1_IR_reg[23]/NET0131  & ~n1930 ;
  assign n1933 = ~n1931 & ~n1932 ;
  assign n1934 = \P1_state_reg[0]/NET0131  & n1933 ;
  assign n1935 = ~n1929 & n1934 ;
  assign n1936 = ~n527 & n536 ;
  assign n1945 = \P1_IR_reg[31]/NET0131  & ~n655 ;
  assign n1946 = ~n651 & ~n1945 ;
  assign n1947 = \P1_IR_reg[25]/NET0131  & ~n1946 ;
  assign n1948 = ~\P1_IR_reg[25]/NET0131  & n1946 ;
  assign n1949 = ~n1947 & ~n1948 ;
  assign n1937 = \P1_IR_reg[26]/NET0131  & ~n642 ;
  assign n1938 = ~\P1_IR_reg[26]/NET0131  & n642 ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = \P1_IR_reg[31]/NET0131  & ~n529 ;
  assign n1941 = ~n491 & ~n1940 ;
  assign n1942 = \P1_IR_reg[24]/NET0131  & ~n1941 ;
  assign n1943 = ~\P1_IR_reg[24]/NET0131  & n1941 ;
  assign n1944 = ~n1942 & ~n1943 ;
  assign n1950 = ~n1939 & n1944 ;
  assign n1951 = n1949 & n1950 ;
  assign n1952 = n1936 & ~n1951 ;
  assign n1953 = n1898 & n1952 ;
  assign n1954 = ~n1933 & ~n1953 ;
  assign n1955 = \P1_state_reg[0]/NET0131  & ~n1954 ;
  assign n1956 = \P1_B_reg/NET0131  & ~n1955 ;
  assign n1957 = ~n1935 & ~n1956 ;
  assign n1958 = ~\P2_IR_reg[17]/NET0131  & ~\P2_IR_reg[18]/NET0131  ;
  assign n1959 = ~\P2_IR_reg[8]/NET0131  & ~\P2_IR_reg[9]/NET0131  ;
  assign n1960 = ~\P2_IR_reg[10]/NET0131  & n1959 ;
  assign n1961 = ~\P2_IR_reg[11]/NET0131  & ~\P2_IR_reg[12]/NET0131  ;
  assign n1962 = n1960 & n1961 ;
  assign n1963 = ~\P2_IR_reg[0]/NET0131  & ~\P2_IR_reg[1]/NET0131  ;
  assign n1964 = ~\P2_IR_reg[2]/NET0131  & n1963 ;
  assign n1965 = ~\P2_IR_reg[3]/NET0131  & n1964 ;
  assign n1966 = ~\P2_IR_reg[5]/NET0131  & ~\P2_IR_reg[6]/NET0131  ;
  assign n1967 = ~\P2_IR_reg[4]/NET0131  & ~\P2_IR_reg[7]/NET0131  ;
  assign n1968 = n1966 & n1967 ;
  assign n1969 = n1965 & n1968 ;
  assign n1970 = n1962 & n1969 ;
  assign n1971 = ~\P2_IR_reg[14]/NET0131  & ~\P2_IR_reg[15]/NET0131  ;
  assign n1972 = ~\P2_IR_reg[13]/NET0131  & n1971 ;
  assign n1973 = ~\P2_IR_reg[16]/NET0131  & n1972 ;
  assign n1974 = n1970 & n1973 ;
  assign n1975 = n1958 & n1974 ;
  assign n1976 = \P2_IR_reg[31]/NET0131  & ~n1975 ;
  assign n1977 = ~\P2_IR_reg[20]/NET0131  & ~\P2_IR_reg[21]/NET0131  ;
  assign n1978 = ~\P2_IR_reg[22]/NET0131  & n1977 ;
  assign n1979 = ~\P2_IR_reg[19]/NET0131  & n1978 ;
  assign n1980 = \P2_IR_reg[31]/NET0131  & ~n1979 ;
  assign n1981 = ~n1976 & ~n1980 ;
  assign n1982 = \P2_IR_reg[23]/NET0131  & ~n1981 ;
  assign n1983 = ~\P2_IR_reg[23]/NET0131  & n1981 ;
  assign n1984 = ~n1982 & ~n1983 ;
  assign n1995 = ~\P2_IR_reg[13]/NET0131  & n1962 ;
  assign n1996 = n1969 & n1995 ;
  assign n1997 = ~\P2_IR_reg[16]/NET0131  & ~\P2_IR_reg[17]/NET0131  ;
  assign n1998 = n1971 & n1997 ;
  assign n1999 = ~\P2_IR_reg[18]/NET0131  & ~\P2_IR_reg[19]/NET0131  ;
  assign n2000 = n1998 & n1999 ;
  assign n2001 = n1996 & n2000 ;
  assign n2002 = \P2_IR_reg[31]/NET0131  & ~n2001 ;
  assign n1985 = ~\P2_IR_reg[23]/NET0131  & n1978 ;
  assign n2003 = \P2_IR_reg[31]/NET0131  & ~n1985 ;
  assign n2004 = ~n2002 & ~n2003 ;
  assign n2005 = \P2_IR_reg[24]/NET0131  & ~n2004 ;
  assign n2006 = ~\P2_IR_reg[24]/NET0131  & n2004 ;
  assign n2007 = ~n2005 & ~n2006 ;
  assign n1986 = ~\P2_IR_reg[24]/NET0131  & n1985 ;
  assign n1987 = ~\P2_IR_reg[19]/NET0131  & n1958 ;
  assign n1988 = n1973 & n1987 ;
  assign n1989 = n1986 & n1988 ;
  assign n1990 = n1970 & n1989 ;
  assign n1991 = \P2_IR_reg[31]/NET0131  & ~n1990 ;
  assign n1992 = \P2_IR_reg[25]/NET0131  & ~n1991 ;
  assign n1993 = ~\P2_IR_reg[25]/NET0131  & n1991 ;
  assign n1994 = ~n1992 & ~n1993 ;
  assign n2008 = ~\P2_IR_reg[25]/NET0131  & n2000 ;
  assign n2009 = n1986 & n2008 ;
  assign n2010 = n1996 & n2009 ;
  assign n2011 = \P2_IR_reg[31]/NET0131  & ~n2010 ;
  assign n2012 = \P2_IR_reg[26]/NET0131  & ~n2011 ;
  assign n2013 = ~\P2_IR_reg[26]/NET0131  & n2011 ;
  assign n2014 = ~n2012 & ~n2013 ;
  assign n2015 = ~n1994 & ~n2014 ;
  assign n2016 = n2007 & n2015 ;
  assign n2017 = ~n1984 & ~n2016 ;
  assign n2018 = n1994 & ~n2014 ;
  assign n2022 = \P2_B_reg/NET0131  & ~n2007 ;
  assign n2023 = n2018 & n2022 ;
  assign n2019 = ~\P2_B_reg/NET0131  & n2007 ;
  assign n2020 = n2018 & n2019 ;
  assign n2021 = n2007 & n2014 ;
  assign n2024 = \P2_d_reg[0]/NET0131  & ~n2014 ;
  assign n2025 = ~n2021 & ~n2024 ;
  assign n2026 = ~n2020 & n2025 ;
  assign n2027 = ~n2023 & n2026 ;
  assign n2028 = \P2_d_reg[1]/NET0131  & ~n2014 ;
  assign n2029 = ~n1994 & n2014 ;
  assign n2030 = ~n2028 & ~n2029 ;
  assign n2031 = ~n2020 & n2030 ;
  assign n2032 = ~n2023 & n2031 ;
  assign n2033 = n2027 & ~n2032 ;
  assign n2034 = \P2_reg2_reg[29]/NET0131  & ~n2033 ;
  assign n2035 = ~\P2_IR_reg[25]/NET0131  & ~\P2_IR_reg[26]/NET0131  ;
  assign n2036 = ~\P2_IR_reg[24]/NET0131  & n2035 ;
  assign n2037 = ~\P2_IR_reg[23]/NET0131  & n2036 ;
  assign n2038 = n1979 & n2037 ;
  assign n2039 = n1975 & n2038 ;
  assign n2040 = \P2_IR_reg[31]/NET0131  & ~n2039 ;
  assign n2041 = \P2_IR_reg[27]/NET0131  & n2040 ;
  assign n2042 = ~\P2_IR_reg[27]/NET0131  & ~n2040 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = ~\P2_IR_reg[27]/NET0131  & n2036 ;
  assign n2045 = n2001 & n2044 ;
  assign n2046 = \P2_IR_reg[31]/NET0131  & ~n2045 ;
  assign n2047 = ~n2003 & ~n2046 ;
  assign n2048 = \P2_IR_reg[28]/NET0131  & ~n2047 ;
  assign n2049 = ~\P2_IR_reg[28]/NET0131  & n2047 ;
  assign n2050 = ~n2048 & ~n2049 ;
  assign n2051 = ~n2043 & ~n2050 ;
  assign n2052 = \P1_datao_reg[29]/NET0131  & ~n542 ;
  assign n2053 = \P1_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n2054 = ~\P1_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n2055 = ~n2053 & ~n2054 ;
  assign n2056 = ~\P1_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n2101 = \P1_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n2102 = ~\P1_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n2103 = ~\P1_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n2104 = ~n2102 & ~n2103 ;
  assign n2105 = \P1_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n2106 = ~\P1_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n2107 = \P1_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n2108 = \P1_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n2109 = ~n2107 & ~n2108 ;
  assign n2110 = ~n2106 & ~n2109 ;
  assign n2111 = ~n2105 & ~n2110 ;
  assign n2112 = n2104 & ~n2111 ;
  assign n2113 = ~n2101 & ~n2112 ;
  assign n2126 = ~\P1_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n2127 = ~\P1_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n2128 = ~\P1_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n2129 = ~\P1_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n2130 = \P1_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n2131 = \P1_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n2132 = ~n2130 & ~n2131 ;
  assign n2133 = ~n2129 & ~n2132 ;
  assign n2134 = ~n2128 & n2133 ;
  assign n2135 = \P1_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n2136 = \P1_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n2137 = ~n2135 & ~n2136 ;
  assign n2138 = ~n2134 & n2137 ;
  assign n2139 = ~n2127 & ~n2138 ;
  assign n2140 = \P1_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n2141 = ~n2139 & ~n2140 ;
  assign n2142 = ~n2126 & ~n2141 ;
  assign n2115 = ~\P1_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n2116 = ~\P1_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n2117 = ~n2115 & ~n2116 ;
  assign n2119 = ~\P1_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n2143 = ~\P1_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n2144 = ~n2119 & ~n2143 ;
  assign n2145 = n2117 & n2144 ;
  assign n2146 = n2142 & n2145 ;
  assign n2114 = \P1_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n2118 = \P1_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n2120 = \P1_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n2121 = \P1_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n2122 = ~n2120 & ~n2121 ;
  assign n2123 = ~n2119 & ~n2122 ;
  assign n2124 = ~n2118 & ~n2123 ;
  assign n2125 = n2117 & ~n2124 ;
  assign n2147 = ~n2114 & ~n2125 ;
  assign n2148 = ~n2146 & n2147 ;
  assign n2149 = ~\P1_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n2150 = ~n2106 & ~n2149 ;
  assign n2151 = n2104 & n2150 ;
  assign n2152 = ~n2148 & n2151 ;
  assign n2153 = n2113 & ~n2152 ;
  assign n2069 = ~\P1_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n2074 = ~\P1_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n2075 = ~n2069 & ~n2074 ;
  assign n2076 = ~\P1_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n2083 = ~\P1_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n2084 = ~n2076 & ~n2083 ;
  assign n2085 = n2075 & n2084 ;
  assign n2086 = ~\P1_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n2091 = ~\P1_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n2092 = ~n2086 & ~n2091 ;
  assign n2093 = ~\P1_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n2154 = ~\P1_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n2155 = ~n2093 & ~n2154 ;
  assign n2156 = n2092 & n2155 ;
  assign n2157 = n2085 & n2156 ;
  assign n2158 = ~n2153 & n2157 ;
  assign n2070 = \P1_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n2071 = \P1_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n2072 = ~n2070 & ~n2071 ;
  assign n2073 = ~n2069 & ~n2072 ;
  assign n2077 = \P1_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n2078 = \P1_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n2079 = ~n2077 & ~n2078 ;
  assign n2080 = ~n2076 & ~n2079 ;
  assign n2081 = n2075 & n2080 ;
  assign n2082 = ~n2073 & ~n2081 ;
  assign n2087 = \P1_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n2088 = \P1_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n2089 = ~n2087 & ~n2088 ;
  assign n2090 = ~n2086 & ~n2089 ;
  assign n2094 = \P1_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n2095 = \P1_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n2096 = ~n2094 & ~n2095 ;
  assign n2097 = ~n2093 & ~n2096 ;
  assign n2098 = n2092 & n2097 ;
  assign n2099 = ~n2090 & ~n2098 ;
  assign n2100 = n2085 & ~n2099 ;
  assign n2159 = n2082 & ~n2100 ;
  assign n2160 = ~n2158 & n2159 ;
  assign n2057 = ~\P1_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n2058 = ~\P1_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n2059 = ~\P1_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n2060 = ~n2058 & ~n2059 ;
  assign n2061 = ~n2057 & n2060 ;
  assign n2062 = ~\P1_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n2063 = ~\P1_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n2064 = ~n2062 & ~n2063 ;
  assign n2065 = ~\P1_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n2066 = ~\P1_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n2067 = ~n2065 & ~n2066 ;
  assign n2068 = n2064 & n2067 ;
  assign n2161 = n2061 & n2068 ;
  assign n2162 = ~n2160 & n2161 ;
  assign n2163 = \P1_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n2164 = \P1_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n2165 = ~n2163 & ~n2164 ;
  assign n2166 = \P1_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n2167 = \P1_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n2168 = ~n2166 & ~n2167 ;
  assign n2169 = ~n2058 & ~n2168 ;
  assign n2170 = \P1_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n2171 = \P1_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n2172 = ~n2170 & ~n2171 ;
  assign n2173 = ~n2062 & ~n2172 ;
  assign n2174 = \P1_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n2175 = \P1_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n2176 = ~n2174 & ~n2175 ;
  assign n2177 = ~n2065 & ~n2176 ;
  assign n2178 = n2064 & n2177 ;
  assign n2179 = ~n2173 & ~n2178 ;
  assign n2180 = n2060 & ~n2179 ;
  assign n2181 = ~n2169 & ~n2180 ;
  assign n2182 = ~n2057 & ~n2181 ;
  assign n2183 = n2165 & ~n2182 ;
  assign n2184 = ~n2162 & n2183 ;
  assign n2185 = ~n2056 & ~n2184 ;
  assign n2187 = n2055 & n2185 ;
  assign n2186 = ~n2055 & ~n2185 ;
  assign n2188 = n542 & ~n2186 ;
  assign n2189 = ~n2187 & n2188 ;
  assign n2190 = ~n2052 & ~n2189 ;
  assign n2191 = ~n2051 & ~n2190 ;
  assign n2192 = ~\P2_IR_reg[27]/NET0131  & ~\P2_IR_reg[28]/NET0131  ;
  assign n2193 = ~\P2_IR_reg[26]/NET0131  & ~\P2_IR_reg[29]/NET0131  ;
  assign n2194 = n2192 & n2193 ;
  assign n2195 = \P2_IR_reg[31]/NET0131  & ~n2194 ;
  assign n2196 = ~n2011 & ~n2195 ;
  assign n2197 = \P2_IR_reg[30]/NET0131  & ~n2196 ;
  assign n2198 = ~\P2_IR_reg[30]/NET0131  & n2196 ;
  assign n2199 = ~n2197 & ~n2198 ;
  assign n2200 = n2035 & n2192 ;
  assign n2201 = \P2_IR_reg[31]/NET0131  & ~n2200 ;
  assign n2202 = ~n1991 & ~n2201 ;
  assign n2203 = \P2_IR_reg[29]/NET0131  & ~n2202 ;
  assign n2204 = ~\P2_IR_reg[29]/NET0131  & n2202 ;
  assign n2205 = ~n2203 & ~n2204 ;
  assign n2212 = n2199 & n2205 ;
  assign n2213 = \P2_reg3_reg[3]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n2214 = \P2_reg3_reg[5]/NET0131  & n2213 ;
  assign n2215 = \P2_reg3_reg[6]/NET0131  & n2214 ;
  assign n2216 = \P2_reg3_reg[7]/NET0131  & n2215 ;
  assign n2217 = \P2_reg3_reg[8]/NET0131  & n2216 ;
  assign n2218 = \P2_reg3_reg[9]/NET0131  & n2217 ;
  assign n2219 = \P2_reg3_reg[10]/NET0131  & n2218 ;
  assign n2220 = \P2_reg3_reg[11]/NET0131  & \P2_reg3_reg[12]/NET0131  ;
  assign n2221 = \P2_reg3_reg[13]/NET0131  & n2220 ;
  assign n2222 = n2219 & n2221 ;
  assign n2223 = \P2_reg3_reg[14]/NET0131  & n2222 ;
  assign n2224 = \P2_reg3_reg[15]/NET0131  & \P2_reg3_reg[16]/NET0131  ;
  assign n2225 = n2223 & n2224 ;
  assign n2226 = \P2_reg3_reg[17]/NET0131  & \P2_reg3_reg[18]/NET0131  ;
  assign n2227 = n2225 & n2226 ;
  assign n2228 = \P2_reg3_reg[20]/NET0131  & \P2_reg3_reg[21]/NET0131  ;
  assign n2229 = \P2_reg3_reg[19]/NET0131  & \P2_reg3_reg[22]/NET0131  ;
  assign n2230 = \P2_reg3_reg[23]/NET0131  & \P2_reg3_reg[24]/NET0131  ;
  assign n2231 = n2229 & n2230 ;
  assign n2232 = n2228 & n2231 ;
  assign n2233 = n2227 & n2232 ;
  assign n2234 = \P2_reg3_reg[25]/NET0131  & \P2_reg3_reg[26]/NET0131  ;
  assign n2235 = \P2_reg3_reg[27]/NET0131  & \P2_reg3_reg[28]/NET0131  ;
  assign n2236 = n2234 & n2235 ;
  assign n2237 = n2233 & n2236 ;
  assign n2238 = n2212 & n2237 ;
  assign n2210 = ~n2199 & ~n2205 ;
  assign n2211 = \P2_reg0_reg[29]/NET0131  & n2210 ;
  assign n2206 = ~n2199 & n2205 ;
  assign n2207 = \P2_reg1_reg[29]/NET0131  & n2206 ;
  assign n2208 = n2199 & ~n2205 ;
  assign n2209 = \P2_reg2_reg[29]/NET0131  & n2208 ;
  assign n2239 = ~n2207 & ~n2209 ;
  assign n2240 = ~n2211 & n2239 ;
  assign n2241 = ~n2238 & n2240 ;
  assign n2242 = n2191 & n2241 ;
  assign n2243 = ~n2191 & ~n2241 ;
  assign n2244 = ~n2242 & ~n2243 ;
  assign n2245 = \P1_datao_reg[28]/NET0131  & ~n542 ;
  assign n2246 = ~n2056 & ~n2163 ;
  assign n2247 = ~n2164 & ~n2167 ;
  assign n2248 = ~n2166 & ~n2170 ;
  assign n2249 = ~n2059 & ~n2248 ;
  assign n2250 = ~n2058 & n2249 ;
  assign n2251 = n2247 & ~n2250 ;
  assign n2252 = ~n2057 & ~n2251 ;
  assign n2253 = ~n2103 & n2155 ;
  assign n2254 = ~n2091 & n2253 ;
  assign n2255 = ~n2126 & ~n2143 ;
  assign n2256 = n2139 & n2255 ;
  assign n2257 = ~n2115 & ~n2119 ;
  assign n2258 = n2256 & n2257 ;
  assign n2259 = ~n2120 & ~n2140 ;
  assign n2260 = ~n2143 & ~n2259 ;
  assign n2261 = ~n2121 & ~n2260 ;
  assign n2262 = n2257 & ~n2261 ;
  assign n2263 = ~n2118 & ~n2262 ;
  assign n2264 = ~n2258 & n2263 ;
  assign n2265 = ~n2116 & ~n2149 ;
  assign n2266 = ~n2102 & ~n2106 ;
  assign n2267 = n2265 & n2266 ;
  assign n2268 = ~n2264 & n2267 ;
  assign n2269 = n2254 & n2268 ;
  assign n2274 = ~n2108 & ~n2114 ;
  assign n2275 = ~n2149 & ~n2274 ;
  assign n2276 = ~n2107 & ~n2275 ;
  assign n2277 = n2266 & ~n2276 ;
  assign n2278 = ~n2105 & ~n2277 ;
  assign n2279 = n2254 & ~n2278 ;
  assign n2270 = ~n2091 & ~n2093 ;
  assign n2271 = ~n2094 & ~n2101 ;
  assign n2272 = ~n2154 & ~n2271 ;
  assign n2273 = n2270 & n2272 ;
  assign n2280 = ~n2087 & ~n2095 ;
  assign n2281 = ~n2091 & ~n2280 ;
  assign n2282 = ~n2273 & ~n2281 ;
  assign n2283 = ~n2279 & n2282 ;
  assign n2284 = ~n2269 & n2283 ;
  assign n2285 = ~n2074 & ~n2076 ;
  assign n2286 = ~n2083 & ~n2086 ;
  assign n2287 = n2285 & n2286 ;
  assign n2288 = ~n2284 & n2287 ;
  assign n2289 = ~n2070 & ~n2077 ;
  assign n2290 = ~n2074 & ~n2289 ;
  assign n2291 = ~n2078 & ~n2088 ;
  assign n2292 = ~n2083 & ~n2291 ;
  assign n2293 = n2285 & n2292 ;
  assign n2294 = ~n2290 & ~n2293 ;
  assign n2295 = ~n2288 & n2294 ;
  assign n2296 = ~n2063 & ~n2065 ;
  assign n2297 = ~n2066 & ~n2069 ;
  assign n2298 = n2296 & n2297 ;
  assign n2299 = ~n2295 & n2298 ;
  assign n2300 = ~n2171 & ~n2174 ;
  assign n2301 = ~n2063 & ~n2300 ;
  assign n2302 = ~n2071 & ~n2175 ;
  assign n2303 = ~n2066 & ~n2302 ;
  assign n2304 = n2296 & n2303 ;
  assign n2305 = ~n2301 & ~n2304 ;
  assign n2306 = ~n2299 & n2305 ;
  assign n2307 = n2061 & ~n2062 ;
  assign n2308 = ~n2306 & n2307 ;
  assign n2309 = ~n2252 & ~n2308 ;
  assign n2311 = ~n2246 & n2309 ;
  assign n2310 = n2246 & ~n2309 ;
  assign n2312 = n542 & ~n2310 ;
  assign n2313 = ~n2311 & n2312 ;
  assign n2314 = ~n2245 & ~n2313 ;
  assign n2315 = ~n2051 & ~n2314 ;
  assign n2319 = \P2_reg3_reg[25]/NET0131  & n2233 ;
  assign n2320 = \P2_reg3_reg[26]/NET0131  & n2319 ;
  assign n2321 = \P2_reg3_reg[27]/NET0131  & n2320 ;
  assign n2322 = ~\P2_reg3_reg[28]/NET0131  & ~n2321 ;
  assign n2323 = \P2_reg3_reg[28]/NET0131  & n2321 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = n2212 & n2324 ;
  assign n2318 = \P2_reg0_reg[28]/NET0131  & n2210 ;
  assign n2316 = \P2_reg2_reg[28]/NET0131  & n2208 ;
  assign n2317 = \P2_reg1_reg[28]/NET0131  & n2206 ;
  assign n2326 = ~n2316 & ~n2317 ;
  assign n2327 = ~n2318 & n2326 ;
  assign n2328 = ~n2325 & n2327 ;
  assign n2329 = ~n2315 & n2328 ;
  assign n2330 = \P1_datao_reg[27]/NET0131  & ~n542 ;
  assign n2331 = ~n2057 & ~n2164 ;
  assign n2332 = n2060 & n2173 ;
  assign n2333 = ~n2169 & ~n2332 ;
  assign n2334 = n2060 & n2064 ;
  assign n2337 = n2067 & n2075 ;
  assign n2338 = n2084 & n2092 ;
  assign n2347 = n2337 & n2338 ;
  assign n2348 = ~n2134 & ~n2136 ;
  assign n2349 = ~n2127 & ~n2348 ;
  assign n2350 = ~n2135 & ~n2140 ;
  assign n2351 = ~n2349 & n2350 ;
  assign n2352 = ~n2119 & n2255 ;
  assign n2353 = ~n2351 & n2352 ;
  assign n2354 = ~n2123 & ~n2353 ;
  assign n2355 = n2117 & ~n2149 ;
  assign n2356 = ~n2106 & n2355 ;
  assign n2357 = ~n2354 & n2356 ;
  assign n2358 = ~n2114 & ~n2118 ;
  assign n2359 = ~n2106 & n2265 ;
  assign n2360 = ~n2358 & n2359 ;
  assign n2361 = ~n2110 & ~n2360 ;
  assign n2362 = ~n2357 & n2361 ;
  assign n2363 = n2104 & ~n2154 ;
  assign n2364 = ~n2093 & n2363 ;
  assign n2365 = ~n2362 & n2364 ;
  assign n2366 = n2347 & n2365 ;
  assign n2335 = n2067 & n2073 ;
  assign n2336 = ~n2177 & ~n2335 ;
  assign n2339 = ~n2101 & ~n2105 ;
  assign n2340 = n2253 & ~n2339 ;
  assign n2341 = ~n2097 & ~n2340 ;
  assign n2342 = n2338 & ~n2341 ;
  assign n2343 = n2084 & n2090 ;
  assign n2344 = ~n2080 & ~n2343 ;
  assign n2345 = ~n2342 & n2344 ;
  assign n2346 = n2337 & ~n2345 ;
  assign n2367 = n2336 & ~n2346 ;
  assign n2368 = ~n2366 & n2367 ;
  assign n2369 = n2334 & ~n2368 ;
  assign n2370 = n2333 & ~n2369 ;
  assign n2372 = ~n2331 & n2370 ;
  assign n2371 = n2331 & ~n2370 ;
  assign n2373 = n542 & ~n2371 ;
  assign n2374 = ~n2372 & n2373 ;
  assign n2375 = ~n2330 & ~n2374 ;
  assign n2376 = ~n2051 & ~n2375 ;
  assign n2380 = ~\P2_reg3_reg[27]/NET0131  & ~n2320 ;
  assign n2381 = ~n2321 & ~n2380 ;
  assign n2382 = n2212 & n2381 ;
  assign n2379 = \P2_reg1_reg[27]/NET0131  & n2206 ;
  assign n2377 = \P2_reg2_reg[27]/NET0131  & n2208 ;
  assign n2378 = \P2_reg0_reg[27]/NET0131  & n2210 ;
  assign n2383 = ~n2377 & ~n2378 ;
  assign n2384 = ~n2379 & n2383 ;
  assign n2385 = ~n2382 & n2384 ;
  assign n2386 = ~n2376 & n2385 ;
  assign n2387 = \P1_datao_reg[26]/NET0131  & ~n542 ;
  assign n2388 = ~n2058 & ~n2167 ;
  assign n2389 = ~n2059 & ~n2062 ;
  assign n2390 = n2301 & n2389 ;
  assign n2391 = ~n2249 & ~n2390 ;
  assign n2392 = n2296 & n2389 ;
  assign n2393 = n2290 & n2297 ;
  assign n2394 = ~n2303 & ~n2393 ;
  assign n2395 = n2270 & n2286 ;
  assign n2396 = ~n2256 & ~n2260 ;
  assign n2397 = n2257 & n2265 ;
  assign n2398 = ~n2396 & n2397 ;
  assign n2399 = ~n2118 & ~n2121 ;
  assign n2400 = n2355 & ~n2399 ;
  assign n2401 = ~n2275 & ~n2400 ;
  assign n2402 = ~n2398 & n2401 ;
  assign n2403 = ~n2106 & n2363 ;
  assign n2404 = ~n2402 & n2403 ;
  assign n2405 = n2395 & n2404 ;
  assign n2406 = ~n2105 & ~n2107 ;
  assign n2407 = n2363 & ~n2406 ;
  assign n2408 = ~n2272 & ~n2407 ;
  assign n2409 = n2395 & ~n2408 ;
  assign n2410 = n2281 & n2286 ;
  assign n2411 = ~n2292 & ~n2410 ;
  assign n2412 = ~n2409 & n2411 ;
  assign n2413 = ~n2405 & n2412 ;
  assign n2414 = n2285 & n2297 ;
  assign n2415 = ~n2413 & n2414 ;
  assign n2416 = n2394 & ~n2415 ;
  assign n2417 = n2392 & ~n2416 ;
  assign n2418 = n2391 & ~n2417 ;
  assign n2420 = ~n2388 & n2418 ;
  assign n2419 = n2388 & ~n2418 ;
  assign n2421 = n542 & ~n2419 ;
  assign n2422 = ~n2420 & n2421 ;
  assign n2423 = ~n2387 & ~n2422 ;
  assign n2424 = ~n2051 & ~n2423 ;
  assign n2428 = ~\P2_reg3_reg[26]/NET0131  & ~n2319 ;
  assign n2429 = ~n2320 & ~n2428 ;
  assign n2430 = n2212 & n2429 ;
  assign n2427 = \P2_reg2_reg[26]/NET0131  & n2208 ;
  assign n2425 = \P2_reg0_reg[26]/NET0131  & n2210 ;
  assign n2426 = \P2_reg1_reg[26]/NET0131  & n2206 ;
  assign n2431 = ~n2425 & ~n2426 ;
  assign n2432 = ~n2427 & n2431 ;
  assign n2433 = ~n2430 & n2432 ;
  assign n2434 = ~n2424 & n2433 ;
  assign n2435 = ~n2386 & ~n2434 ;
  assign n2436 = \P1_datao_reg[25]/NET0131  & ~n542 ;
  assign n2437 = ~n2059 & ~n2166 ;
  assign n2438 = n2152 & n2156 ;
  assign n2439 = n2085 & n2438 ;
  assign n2440 = ~n2113 & n2156 ;
  assign n2441 = n2099 & ~n2440 ;
  assign n2442 = n2085 & ~n2441 ;
  assign n2443 = n2082 & ~n2442 ;
  assign n2444 = ~n2439 & n2443 ;
  assign n2445 = n2068 & ~n2444 ;
  assign n2446 = n2179 & ~n2445 ;
  assign n2448 = ~n2437 & n2446 ;
  assign n2447 = n2437 & ~n2446 ;
  assign n2449 = n542 & ~n2447 ;
  assign n2450 = ~n2448 & n2449 ;
  assign n2451 = ~n2436 & ~n2450 ;
  assign n2452 = ~n2051 & ~n2451 ;
  assign n2456 = ~\P2_reg3_reg[25]/NET0131  & ~n2233 ;
  assign n2457 = ~n2319 & ~n2456 ;
  assign n2458 = n2212 & n2457 ;
  assign n2455 = \P2_reg0_reg[25]/NET0131  & n2210 ;
  assign n2453 = \P2_reg1_reg[25]/NET0131  & n2206 ;
  assign n2454 = \P2_reg2_reg[25]/NET0131  & n2208 ;
  assign n2459 = ~n2453 & ~n2454 ;
  assign n2460 = ~n2455 & n2459 ;
  assign n2461 = ~n2458 & n2460 ;
  assign n2462 = ~n2452 & n2461 ;
  assign n2463 = n2435 & ~n2462 ;
  assign n2464 = \P1_datao_reg[24]/NET0131  & ~n542 ;
  assign n2465 = ~n2062 & ~n2170 ;
  assign n2467 = n2306 & ~n2465 ;
  assign n2466 = ~n2306 & n2465 ;
  assign n2468 = n542 & ~n2466 ;
  assign n2469 = ~n2467 & n2468 ;
  assign n2470 = ~n2464 & ~n2469 ;
  assign n2471 = ~n2051 & ~n2470 ;
  assign n2475 = \P2_reg3_reg[19]/NET0131  & n2227 ;
  assign n2476 = n2228 & n2475 ;
  assign n2477 = \P2_reg3_reg[22]/NET0131  & n2476 ;
  assign n2478 = \P2_reg3_reg[23]/NET0131  & n2477 ;
  assign n2479 = ~\P2_reg3_reg[24]/NET0131  & ~n2478 ;
  assign n2480 = ~n2233 & ~n2479 ;
  assign n2481 = n2212 & n2480 ;
  assign n2474 = \P2_reg1_reg[24]/NET0131  & n2206 ;
  assign n2472 = \P2_reg0_reg[24]/NET0131  & n2210 ;
  assign n2473 = \P2_reg2_reg[24]/NET0131  & n2208 ;
  assign n2482 = ~n2472 & ~n2473 ;
  assign n2483 = ~n2474 & n2482 ;
  assign n2484 = ~n2481 & n2483 ;
  assign n2485 = ~n2471 & n2484 ;
  assign n2486 = \P1_datao_reg[23]/NET0131  & ~n542 ;
  assign n2487 = ~n2063 & ~n2171 ;
  assign n2489 = n2341 & ~n2365 ;
  assign n2490 = n2347 & ~n2489 ;
  assign n2488 = n2337 & ~n2344 ;
  assign n2491 = n2336 & ~n2488 ;
  assign n2492 = ~n2490 & n2491 ;
  assign n2494 = ~n2487 & n2492 ;
  assign n2493 = n2487 & ~n2492 ;
  assign n2495 = n542 & ~n2493 ;
  assign n2496 = ~n2494 & n2495 ;
  assign n2497 = ~n2486 & ~n2496 ;
  assign n2498 = ~n2051 & ~n2497 ;
  assign n2502 = ~\P2_reg3_reg[23]/NET0131  & ~n2477 ;
  assign n2503 = ~n2478 & ~n2502 ;
  assign n2504 = n2212 & n2503 ;
  assign n2501 = \P2_reg2_reg[23]/NET0131  & n2208 ;
  assign n2499 = \P2_reg0_reg[23]/NET0131  & n2210 ;
  assign n2500 = \P2_reg1_reg[23]/NET0131  & n2206 ;
  assign n2505 = ~n2499 & ~n2500 ;
  assign n2506 = ~n2501 & n2505 ;
  assign n2507 = ~n2504 & n2506 ;
  assign n2508 = ~n2498 & n2507 ;
  assign n2509 = ~n2485 & ~n2508 ;
  assign n2510 = \P1_datao_reg[22]/NET0131  & ~n542 ;
  assign n2511 = ~n2065 & ~n2174 ;
  assign n2512 = ~n2404 & n2408 ;
  assign n2513 = n2395 & ~n2512 ;
  assign n2514 = n2411 & ~n2513 ;
  assign n2515 = n2414 & ~n2514 ;
  assign n2516 = n2394 & ~n2515 ;
  assign n2518 = ~n2511 & n2516 ;
  assign n2517 = n2511 & ~n2516 ;
  assign n2519 = n542 & ~n2517 ;
  assign n2520 = ~n2518 & n2519 ;
  assign n2521 = ~n2510 & ~n2520 ;
  assign n2522 = ~n2051 & ~n2521 ;
  assign n2526 = ~\P2_reg3_reg[22]/NET0131  & ~n2476 ;
  assign n2527 = ~n2477 & ~n2526 ;
  assign n2528 = n2212 & n2527 ;
  assign n2525 = \P2_reg1_reg[22]/NET0131  & n2206 ;
  assign n2523 = \P2_reg2_reg[22]/NET0131  & n2208 ;
  assign n2524 = \P2_reg0_reg[22]/NET0131  & n2210 ;
  assign n2529 = ~n2523 & ~n2524 ;
  assign n2530 = ~n2525 & n2529 ;
  assign n2531 = ~n2528 & n2530 ;
  assign n2532 = n2522 & ~n2531 ;
  assign n2533 = ~n2522 & n2531 ;
  assign n2534 = \P1_datao_reg[21]/NET0131  & ~n542 ;
  assign n2535 = ~n2066 & ~n2175 ;
  assign n2537 = n2160 & ~n2535 ;
  assign n2536 = ~n2160 & n2535 ;
  assign n2538 = n542 & ~n2536 ;
  assign n2539 = ~n2537 & n2538 ;
  assign n2540 = ~n2534 & ~n2539 ;
  assign n2541 = ~n2051 & ~n2540 ;
  assign n2545 = \P2_reg3_reg[20]/NET0131  & n2475 ;
  assign n2546 = ~\P2_reg3_reg[21]/NET0131  & ~n2545 ;
  assign n2547 = ~n2476 & ~n2546 ;
  assign n2548 = n2212 & n2547 ;
  assign n2544 = \P2_reg0_reg[21]/NET0131  & n2210 ;
  assign n2542 = \P2_reg2_reg[21]/NET0131  & n2208 ;
  assign n2543 = \P2_reg1_reg[21]/NET0131  & n2206 ;
  assign n2549 = ~n2542 & ~n2543 ;
  assign n2550 = ~n2544 & n2549 ;
  assign n2551 = ~n2548 & n2550 ;
  assign n2552 = n2541 & ~n2551 ;
  assign n2553 = ~n2533 & n2552 ;
  assign n2554 = ~n2532 & ~n2553 ;
  assign n2555 = n2509 & ~n2554 ;
  assign n2556 = n2471 & ~n2484 ;
  assign n2557 = n2498 & ~n2507 ;
  assign n2558 = ~n2485 & n2557 ;
  assign n2559 = ~n2556 & ~n2558 ;
  assign n2560 = ~n2555 & n2559 ;
  assign n2561 = n2463 & ~n2560 ;
  assign n2563 = n2424 & ~n2433 ;
  assign n2564 = n2452 & ~n2461 ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = n2435 & ~n2565 ;
  assign n2562 = n2376 & ~n2385 ;
  assign n2567 = n2315 & ~n2328 ;
  assign n2568 = ~n2562 & ~n2567 ;
  assign n2569 = ~n2566 & n2568 ;
  assign n2570 = ~n2561 & n2569 ;
  assign n2571 = ~n2329 & ~n2570 ;
  assign n2572 = \P1_datao_reg[20]/NET0131  & ~n542 ;
  assign n2573 = ~n2069 & ~n2071 ;
  assign n2575 = n2295 & ~n2573 ;
  assign n2574 = ~n2295 & n2573 ;
  assign n2576 = n542 & ~n2574 ;
  assign n2577 = ~n2575 & n2576 ;
  assign n2578 = ~n2572 & ~n2577 ;
  assign n2579 = ~n2051 & ~n2578 ;
  assign n2583 = ~\P2_reg3_reg[20]/NET0131  & ~n2475 ;
  assign n2584 = ~n2545 & ~n2583 ;
  assign n2585 = n2212 & n2584 ;
  assign n2582 = \P2_reg2_reg[20]/NET0131  & n2208 ;
  assign n2580 = \P2_reg1_reg[20]/NET0131  & n2206 ;
  assign n2581 = \P2_reg0_reg[20]/NET0131  & n2210 ;
  assign n2586 = ~n2580 & ~n2581 ;
  assign n2587 = ~n2582 & n2586 ;
  assign n2588 = ~n2585 & n2587 ;
  assign n2589 = ~n2579 & n2588 ;
  assign n2590 = ~\P2_IR_reg[19]/NET0131  & ~n1976 ;
  assign n2591 = \P2_IR_reg[19]/NET0131  & n1976 ;
  assign n2592 = ~n2590 & ~n2591 ;
  assign n2593 = n2051 & ~n2592 ;
  assign n2594 = \P1_datao_reg[19]/NET0131  & ~n542 ;
  assign n2595 = ~n2070 & ~n2074 ;
  assign n2596 = n2338 & n2365 ;
  assign n2597 = n2345 & ~n2596 ;
  assign n2599 = ~n2595 & n2597 ;
  assign n2598 = n2595 & ~n2597 ;
  assign n2600 = n542 & ~n2598 ;
  assign n2601 = ~n2599 & n2600 ;
  assign n2602 = ~n2594 & ~n2601 ;
  assign n2603 = ~n2051 & n2602 ;
  assign n2604 = ~n2593 & ~n2603 ;
  assign n2608 = ~\P2_reg3_reg[19]/NET0131  & ~n2227 ;
  assign n2609 = ~n2475 & ~n2608 ;
  assign n2610 = n2212 & n2609 ;
  assign n2607 = \P2_reg2_reg[19]/NET0131  & n2208 ;
  assign n2605 = \P2_reg1_reg[19]/NET0131  & n2206 ;
  assign n2606 = \P2_reg0_reg[19]/NET0131  & n2210 ;
  assign n2611 = ~n2605 & ~n2606 ;
  assign n2612 = ~n2607 & n2611 ;
  assign n2613 = ~n2610 & n2612 ;
  assign n2614 = ~n2604 & n2613 ;
  assign n2615 = ~n2589 & ~n2614 ;
  assign n2616 = \P2_IR_reg[31]/NET0131  & ~n1974 ;
  assign n2617 = ~\P2_IR_reg[17]/NET0131  & ~n2616 ;
  assign n2618 = \P2_IR_reg[17]/NET0131  & n2616 ;
  assign n2619 = ~n2617 & ~n2618 ;
  assign n2620 = n2051 & ~n2619 ;
  assign n2621 = \P1_datao_reg[17]/NET0131  & ~n542 ;
  assign n2622 = ~n2078 & ~n2083 ;
  assign n2623 = ~n2438 & n2441 ;
  assign n2625 = ~n2622 & n2623 ;
  assign n2624 = n2622 & ~n2623 ;
  assign n2626 = n542 & ~n2624 ;
  assign n2627 = ~n2625 & n2626 ;
  assign n2628 = ~n2621 & ~n2627 ;
  assign n2629 = ~n2051 & n2628 ;
  assign n2630 = ~n2620 & ~n2629 ;
  assign n2634 = ~\P2_reg3_reg[17]/NET0131  & ~n2225 ;
  assign n2635 = \P2_reg3_reg[17]/NET0131  & n2225 ;
  assign n2636 = ~n2634 & ~n2635 ;
  assign n2637 = n2212 & n2636 ;
  assign n2633 = \P2_reg0_reg[17]/NET0131  & n2210 ;
  assign n2631 = \P2_reg2_reg[17]/NET0131  & n2208 ;
  assign n2632 = \P2_reg1_reg[17]/NET0131  & n2206 ;
  assign n2638 = ~n2631 & ~n2632 ;
  assign n2639 = ~n2633 & n2638 ;
  assign n2640 = ~n2637 & n2639 ;
  assign n2641 = ~n2630 & n2640 ;
  assign n2642 = \P2_IR_reg[31]/NET0131  & ~n1996 ;
  assign n2643 = \P2_IR_reg[31]/NET0131  & ~n1998 ;
  assign n2644 = ~n2642 & ~n2643 ;
  assign n2645 = \P2_IR_reg[18]/NET0131  & ~n2644 ;
  assign n2646 = ~\P2_IR_reg[18]/NET0131  & n2644 ;
  assign n2647 = ~n2645 & ~n2646 ;
  assign n2648 = n2051 & ~n2647 ;
  assign n2649 = \P1_datao_reg[18]/NET0131  & ~n542 ;
  assign n2650 = ~n2076 & ~n2077 ;
  assign n2652 = n2413 & ~n2650 ;
  assign n2651 = ~n2413 & n2650 ;
  assign n2653 = n542 & ~n2651 ;
  assign n2654 = ~n2652 & n2653 ;
  assign n2655 = ~n2649 & ~n2654 ;
  assign n2656 = ~n2051 & n2655 ;
  assign n2657 = ~n2648 & ~n2656 ;
  assign n2661 = ~\P2_reg3_reg[18]/NET0131  & ~n2635 ;
  assign n2662 = ~n2227 & ~n2661 ;
  assign n2663 = n2212 & n2662 ;
  assign n2660 = \P2_reg1_reg[18]/NET0131  & n2206 ;
  assign n2658 = \P2_reg2_reg[18]/NET0131  & n2208 ;
  assign n2659 = \P2_reg0_reg[18]/NET0131  & n2210 ;
  assign n2664 = ~n2658 & ~n2659 ;
  assign n2665 = ~n2660 & n2664 ;
  assign n2666 = ~n2663 & n2665 ;
  assign n2667 = ~n2657 & n2666 ;
  assign n2668 = ~n2641 & ~n2667 ;
  assign n2669 = n2615 & n2668 ;
  assign n2771 = \P2_reg2_reg[2]/NET0131  & n2208 ;
  assign n2772 = \P2_reg3_reg[2]/NET0131  & n2212 ;
  assign n2775 = ~n2771 & ~n2772 ;
  assign n2773 = \P2_reg1_reg[2]/NET0131  & n2206 ;
  assign n2774 = \P2_reg0_reg[2]/NET0131  & n2210 ;
  assign n2776 = ~n2773 & ~n2774 ;
  assign n2777 = n2775 & n2776 ;
  assign n2778 = \P1_datao_reg[2]/NET0131  & ~n542 ;
  assign n2779 = ~n2128 & ~n2136 ;
  assign n2781 = n2133 & n2779 ;
  assign n2780 = ~n2133 & ~n2779 ;
  assign n2782 = n542 & ~n2780 ;
  assign n2783 = ~n2781 & n2782 ;
  assign n2784 = ~n2778 & ~n2783 ;
  assign n2785 = ~n2051 & ~n2784 ;
  assign n2786 = \P2_IR_reg[31]/NET0131  & ~n1963 ;
  assign n2787 = ~\P2_IR_reg[2]/NET0131  & ~n2786 ;
  assign n2788 = \P2_IR_reg[2]/NET0131  & n2786 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2790 = n2051 & n2789 ;
  assign n2791 = ~n2785 & ~n2790 ;
  assign n2792 = ~n2777 & ~n2791 ;
  assign n2793 = n2777 & n2791 ;
  assign n2794 = \P2_reg0_reg[1]/NET0131  & n2210 ;
  assign n2795 = \P2_reg1_reg[1]/NET0131  & n2206 ;
  assign n2798 = ~n2794 & ~n2795 ;
  assign n2796 = \P2_reg2_reg[1]/NET0131  & n2208 ;
  assign n2797 = \P2_reg3_reg[1]/NET0131  & n2212 ;
  assign n2799 = ~n2796 & ~n2797 ;
  assign n2800 = n2798 & n2799 ;
  assign n2801 = ~\P1_datao_reg[1]/NET0131  & ~n542 ;
  assign n2802 = ~n2129 & ~n2130 ;
  assign n2804 = ~n2131 & n2802 ;
  assign n2803 = n2131 & ~n2802 ;
  assign n2805 = n542 & ~n2803 ;
  assign n2806 = ~n2804 & n2805 ;
  assign n2807 = ~n2801 & ~n2806 ;
  assign n2808 = ~n2051 & n2807 ;
  assign n2809 = \P2_IR_reg[1]/NET0131  & ~\P2_IR_reg[31]/NET0131  ;
  assign n2810 = \P2_IR_reg[0]/NET0131  & \P2_IR_reg[1]/NET0131  ;
  assign n2811 = n2786 & ~n2810 ;
  assign n2812 = ~n2809 & ~n2811 ;
  assign n2813 = n2051 & ~n2812 ;
  assign n2814 = ~n2808 & ~n2813 ;
  assign n2815 = n2800 & n2814 ;
  assign n2816 = ~n2800 & ~n2814 ;
  assign n2817 = \P2_reg3_reg[0]/NET0131  & n2212 ;
  assign n2818 = \P2_reg1_reg[0]/NET0131  & n2206 ;
  assign n2821 = ~n2817 & ~n2818 ;
  assign n2819 = \P2_reg2_reg[0]/NET0131  & n2208 ;
  assign n2820 = \P2_reg0_reg[0]/NET0131  & n2210 ;
  assign n2822 = ~n2819 & ~n2820 ;
  assign n2823 = n2821 & n2822 ;
  assign n2824 = \si[0]_pad  & n542 ;
  assign n2825 = ~\P1_datao_reg[0]/NET0131  & ~n2824 ;
  assign n2826 = n542 & n2131 ;
  assign n2827 = ~n2825 & ~n2826 ;
  assign n2828 = ~n2051 & n2827 ;
  assign n2829 = \P2_IR_reg[0]/NET0131  & n2051 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = ~n2823 & ~n2830 ;
  assign n2832 = ~n2816 & ~n2831 ;
  assign n2833 = ~n2815 & ~n2832 ;
  assign n2834 = ~n2793 & n2833 ;
  assign n2835 = ~n2792 & ~n2834 ;
  assign n2836 = ~\P1_datao_reg[4]/NET0131  & ~n542 ;
  assign n2837 = ~n2126 & ~n2140 ;
  assign n2839 = ~n2139 & n2837 ;
  assign n2838 = n2139 & ~n2837 ;
  assign n2840 = n542 & ~n2838 ;
  assign n2841 = ~n2839 & n2840 ;
  assign n2842 = ~n2836 & ~n2841 ;
  assign n2843 = ~n2051 & n2842 ;
  assign n2844 = \P2_IR_reg[31]/NET0131  & ~n1965 ;
  assign n2845 = \P2_IR_reg[4]/NET0131  & ~n2844 ;
  assign n2846 = ~\P2_IR_reg[4]/NET0131  & n2844 ;
  assign n2847 = ~n2845 & ~n2846 ;
  assign n2848 = n2051 & ~n2847 ;
  assign n2849 = ~n2843 & ~n2848 ;
  assign n2850 = \P2_reg2_reg[4]/NET0131  & n2208 ;
  assign n2851 = \P2_reg0_reg[4]/NET0131  & n2210 ;
  assign n2856 = ~n2850 & ~n2851 ;
  assign n2852 = ~\P2_reg3_reg[3]/NET0131  & ~\P2_reg3_reg[4]/NET0131  ;
  assign n2853 = ~n2213 & ~n2852 ;
  assign n2854 = n2212 & n2853 ;
  assign n2855 = \P2_reg1_reg[4]/NET0131  & n2206 ;
  assign n2857 = ~n2854 & ~n2855 ;
  assign n2858 = n2856 & n2857 ;
  assign n2859 = n2849 & n2858 ;
  assign n2860 = \P2_reg2_reg[3]/NET0131  & n2208 ;
  assign n2861 = \P2_reg0_reg[3]/NET0131  & n2210 ;
  assign n2864 = ~n2860 & ~n2861 ;
  assign n2862 = ~\P2_reg3_reg[3]/NET0131  & n2212 ;
  assign n2863 = \P2_reg1_reg[3]/NET0131  & n2206 ;
  assign n2865 = ~n2862 & ~n2863 ;
  assign n2866 = n2864 & n2865 ;
  assign n2867 = \P2_IR_reg[31]/NET0131  & ~n1964 ;
  assign n2868 = \P2_IR_reg[3]/NET0131  & n2867 ;
  assign n2869 = ~\P2_IR_reg[3]/NET0131  & ~n2867 ;
  assign n2870 = ~n2868 & ~n2869 ;
  assign n2871 = n2051 & n2870 ;
  assign n2872 = \P1_datao_reg[3]/NET0131  & ~n542 ;
  assign n2873 = ~n2127 & ~n2135 ;
  assign n2875 = ~n2348 & n2873 ;
  assign n2874 = n2348 & ~n2873 ;
  assign n2876 = n542 & ~n2874 ;
  assign n2877 = ~n2875 & n2876 ;
  assign n2878 = ~n2872 & ~n2877 ;
  assign n2879 = ~n2051 & ~n2878 ;
  assign n2880 = ~n2871 & ~n2879 ;
  assign n2881 = n2866 & n2880 ;
  assign n2882 = ~n2859 & ~n2881 ;
  assign n2883 = ~n2835 & n2882 ;
  assign n2884 = ~n2849 & ~n2858 ;
  assign n2885 = ~n2866 & ~n2880 ;
  assign n2886 = ~n2859 & n2885 ;
  assign n2887 = ~n2884 & ~n2886 ;
  assign n2888 = ~n2883 & n2887 ;
  assign n2670 = \P2_reg0_reg[8]/NET0131  & n2210 ;
  assign n2671 = \P2_reg1_reg[8]/NET0131  & n2206 ;
  assign n2676 = ~n2670 & ~n2671 ;
  assign n2672 = \P2_reg2_reg[8]/NET0131  & n2208 ;
  assign n2673 = ~\P2_reg3_reg[8]/NET0131  & ~n2216 ;
  assign n2674 = ~n2217 & ~n2673 ;
  assign n2675 = n2212 & n2674 ;
  assign n2677 = ~n2672 & ~n2675 ;
  assign n2678 = n2676 & n2677 ;
  assign n2679 = \P2_IR_reg[31]/NET0131  & ~n1969 ;
  assign n2680 = ~\P2_IR_reg[8]/NET0131  & ~n2679 ;
  assign n2681 = \P2_IR_reg[8]/NET0131  & n2679 ;
  assign n2682 = ~n2680 & ~n2681 ;
  assign n2683 = n2051 & ~n2682 ;
  assign n2684 = \P1_datao_reg[8]/NET0131  & ~n542 ;
  assign n2685 = ~n2114 & ~n2116 ;
  assign n2687 = n2264 & ~n2685 ;
  assign n2686 = ~n2264 & n2685 ;
  assign n2688 = n542 & ~n2686 ;
  assign n2689 = ~n2687 & n2688 ;
  assign n2690 = ~n2684 & ~n2689 ;
  assign n2691 = ~n2051 & n2690 ;
  assign n2692 = ~n2683 & ~n2691 ;
  assign n2693 = n2678 & ~n2692 ;
  assign n2694 = \P2_reg2_reg[7]/NET0131  & n2208 ;
  assign n2695 = \P2_reg1_reg[7]/NET0131  & n2206 ;
  assign n2700 = ~n2694 & ~n2695 ;
  assign n2696 = \P2_reg0_reg[7]/NET0131  & n2210 ;
  assign n2697 = ~\P2_reg3_reg[7]/NET0131  & ~n2215 ;
  assign n2698 = ~n2216 & ~n2697 ;
  assign n2699 = n2212 & n2698 ;
  assign n2701 = ~n2696 & ~n2699 ;
  assign n2702 = n2700 & n2701 ;
  assign n2703 = ~\P2_IR_reg[4]/NET0131  & n1965 ;
  assign n2704 = \P2_IR_reg[31]/NET0131  & ~n2703 ;
  assign n2705 = \P2_IR_reg[31]/NET0131  & ~n1966 ;
  assign n2706 = ~n2704 & ~n2705 ;
  assign n2707 = \P2_IR_reg[7]/NET0131  & ~n2706 ;
  assign n2708 = ~\P2_IR_reg[7]/NET0131  & n2706 ;
  assign n2709 = ~n2707 & ~n2708 ;
  assign n2710 = n2051 & ~n2709 ;
  assign n2711 = \P1_datao_reg[7]/NET0131  & ~n542 ;
  assign n2712 = ~n2115 & ~n2118 ;
  assign n2714 = n2354 & ~n2712 ;
  assign n2713 = ~n2354 & n2712 ;
  assign n2715 = n542 & ~n2713 ;
  assign n2716 = ~n2714 & n2715 ;
  assign n2717 = ~n2711 & ~n2716 ;
  assign n2718 = ~n2051 & n2717 ;
  assign n2719 = ~n2710 & ~n2718 ;
  assign n2720 = n2702 & ~n2719 ;
  assign n2721 = ~n2693 & ~n2720 ;
  assign n2722 = \P2_reg1_reg[6]/NET0131  & n2206 ;
  assign n2723 = \P2_reg2_reg[6]/NET0131  & n2208 ;
  assign n2728 = ~n2722 & ~n2723 ;
  assign n2724 = \P2_reg0_reg[6]/NET0131  & n2210 ;
  assign n2725 = ~\P2_reg3_reg[6]/NET0131  & ~n2214 ;
  assign n2726 = ~n2215 & ~n2725 ;
  assign n2727 = n2212 & n2726 ;
  assign n2729 = ~n2724 & ~n2727 ;
  assign n2730 = n2728 & n2729 ;
  assign n2731 = \P2_IR_reg[31]/NET0131  & \P2_IR_reg[5]/NET0131  ;
  assign n2732 = ~n2704 & ~n2731 ;
  assign n2733 = \P2_IR_reg[6]/NET0131  & ~n2732 ;
  assign n2734 = ~\P2_IR_reg[6]/NET0131  & n2732 ;
  assign n2735 = ~n2733 & ~n2734 ;
  assign n2736 = n2051 & ~n2735 ;
  assign n2737 = \P1_datao_reg[6]/NET0131  & ~n542 ;
  assign n2738 = ~n2119 & ~n2121 ;
  assign n2740 = n2396 & ~n2738 ;
  assign n2739 = ~n2396 & n2738 ;
  assign n2741 = n542 & ~n2739 ;
  assign n2742 = ~n2740 & n2741 ;
  assign n2743 = ~n2737 & ~n2742 ;
  assign n2744 = ~n2051 & n2743 ;
  assign n2745 = ~n2736 & ~n2744 ;
  assign n2746 = n2730 & ~n2745 ;
  assign n2747 = \P2_reg1_reg[5]/NET0131  & n2206 ;
  assign n2748 = ~\P2_reg3_reg[5]/NET0131  & ~n2213 ;
  assign n2749 = ~n2214 & ~n2748 ;
  assign n2750 = n2212 & n2749 ;
  assign n2753 = ~n2747 & ~n2750 ;
  assign n2751 = \P2_reg0_reg[5]/NET0131  & n2210 ;
  assign n2752 = \P2_reg2_reg[5]/NET0131  & n2208 ;
  assign n2754 = ~n2751 & ~n2752 ;
  assign n2755 = n2753 & n2754 ;
  assign n2756 = ~\P2_IR_reg[5]/NET0131  & n2704 ;
  assign n2757 = \P2_IR_reg[5]/NET0131  & ~n2704 ;
  assign n2758 = ~n2756 & ~n2757 ;
  assign n2759 = n2051 & n2758 ;
  assign n2760 = \P1_datao_reg[5]/NET0131  & ~n542 ;
  assign n2761 = ~n2120 & ~n2143 ;
  assign n2763 = n2142 & n2761 ;
  assign n2762 = ~n2142 & ~n2761 ;
  assign n2764 = n542 & ~n2762 ;
  assign n2765 = ~n2763 & n2764 ;
  assign n2766 = ~n2760 & ~n2765 ;
  assign n2767 = ~n2051 & n2766 ;
  assign n2768 = ~n2759 & ~n2767 ;
  assign n2769 = n2755 & ~n2768 ;
  assign n2770 = ~n2746 & ~n2769 ;
  assign n2889 = n2721 & n2770 ;
  assign n2890 = ~n2888 & n2889 ;
  assign n2891 = ~n2730 & n2745 ;
  assign n2892 = ~n2755 & n2768 ;
  assign n2893 = ~n2746 & n2892 ;
  assign n2894 = ~n2891 & ~n2893 ;
  assign n2895 = n2721 & ~n2894 ;
  assign n2896 = ~n2678 & n2692 ;
  assign n2897 = ~n2702 & n2719 ;
  assign n2898 = ~n2896 & ~n2897 ;
  assign n2899 = ~n2693 & ~n2898 ;
  assign n2900 = ~n2895 & ~n2899 ;
  assign n2901 = ~n2890 & n2900 ;
  assign n2902 = \P2_reg2_reg[11]/NET0131  & n2208 ;
  assign n2903 = \P2_reg3_reg[11]/NET0131  & n2219 ;
  assign n2904 = ~\P2_reg3_reg[11]/NET0131  & ~n2219 ;
  assign n2905 = ~n2903 & ~n2904 ;
  assign n2906 = n2212 & n2905 ;
  assign n2909 = ~n2902 & ~n2906 ;
  assign n2907 = \P2_reg1_reg[11]/NET0131  & n2206 ;
  assign n2908 = \P2_reg0_reg[11]/NET0131  & n2210 ;
  assign n2910 = ~n2907 & ~n2908 ;
  assign n2911 = n2909 & n2910 ;
  assign n2912 = \P2_IR_reg[31]/NET0131  & ~n1960 ;
  assign n2913 = ~n2679 & ~n2912 ;
  assign n2914 = \P2_IR_reg[11]/NET0131  & ~n2913 ;
  assign n2915 = ~\P2_IR_reg[11]/NET0131  & n2913 ;
  assign n2916 = ~n2914 & ~n2915 ;
  assign n2917 = n2051 & ~n2916 ;
  assign n2918 = \P1_datao_reg[11]/NET0131  & ~n542 ;
  assign n2919 = ~n2102 & ~n2105 ;
  assign n2921 = n2362 & ~n2919 ;
  assign n2920 = ~n2362 & n2919 ;
  assign n2922 = n542 & ~n2920 ;
  assign n2923 = ~n2921 & n2922 ;
  assign n2924 = ~n2918 & ~n2923 ;
  assign n2925 = ~n2051 & n2924 ;
  assign n2926 = ~n2917 & ~n2925 ;
  assign n2927 = n2911 & ~n2926 ;
  assign n2928 = \P2_reg2_reg[12]/NET0131  & n2208 ;
  assign n2929 = \P2_reg3_reg[12]/NET0131  & n2903 ;
  assign n2930 = ~\P2_reg3_reg[12]/NET0131  & ~n2903 ;
  assign n2931 = ~n2929 & ~n2930 ;
  assign n2932 = n2212 & n2931 ;
  assign n2935 = ~n2928 & ~n2932 ;
  assign n2933 = \P2_reg1_reg[12]/NET0131  & n2206 ;
  assign n2934 = \P2_reg0_reg[12]/NET0131  & n2210 ;
  assign n2936 = ~n2933 & ~n2934 ;
  assign n2937 = n2935 & n2936 ;
  assign n2938 = ~\P2_IR_reg[11]/NET0131  & n1969 ;
  assign n2939 = \P2_IR_reg[31]/NET0131  & ~n2938 ;
  assign n2940 = ~n2912 & ~n2939 ;
  assign n2941 = \P2_IR_reg[12]/NET0131  & ~n2940 ;
  assign n2942 = ~\P2_IR_reg[12]/NET0131  & n2940 ;
  assign n2943 = ~n2941 & ~n2942 ;
  assign n2944 = n2051 & ~n2943 ;
  assign n2945 = \P1_datao_reg[12]/NET0131  & ~n542 ;
  assign n2946 = ~n2101 & ~n2103 ;
  assign n2947 = ~n2268 & n2278 ;
  assign n2949 = ~n2946 & n2947 ;
  assign n2948 = n2946 & ~n2947 ;
  assign n2950 = n542 & ~n2948 ;
  assign n2951 = ~n2949 & n2950 ;
  assign n2952 = ~n2945 & ~n2951 ;
  assign n2953 = ~n2051 & n2952 ;
  assign n2954 = ~n2944 & ~n2953 ;
  assign n2955 = n2937 & ~n2954 ;
  assign n2956 = ~n2927 & ~n2955 ;
  assign n2957 = \P2_reg1_reg[10]/NET0131  & n2206 ;
  assign n2958 = \P2_reg0_reg[10]/NET0131  & n2210 ;
  assign n2963 = ~n2957 & ~n2958 ;
  assign n2959 = \P2_reg2_reg[10]/NET0131  & n2208 ;
  assign n2960 = ~\P2_reg3_reg[10]/NET0131  & ~n2218 ;
  assign n2961 = ~n2219 & ~n2960 ;
  assign n2962 = n2212 & n2961 ;
  assign n2964 = ~n2959 & ~n2962 ;
  assign n2965 = n2963 & n2964 ;
  assign n2966 = \P2_IR_reg[31]/NET0131  & ~n1959 ;
  assign n2967 = ~n2679 & ~n2966 ;
  assign n2968 = \P2_IR_reg[10]/NET0131  & ~n2967 ;
  assign n2969 = ~\P2_IR_reg[10]/NET0131  & n2967 ;
  assign n2970 = ~n2968 & ~n2969 ;
  assign n2971 = n2051 & ~n2970 ;
  assign n2972 = \P1_datao_reg[10]/NET0131  & ~n542 ;
  assign n2973 = ~n2106 & ~n2107 ;
  assign n2975 = n2402 & ~n2973 ;
  assign n2974 = ~n2402 & n2973 ;
  assign n2976 = n542 & ~n2974 ;
  assign n2977 = ~n2975 & n2976 ;
  assign n2978 = ~n2972 & ~n2977 ;
  assign n2979 = ~n2051 & n2978 ;
  assign n2980 = ~n2971 & ~n2979 ;
  assign n2981 = n2965 & ~n2980 ;
  assign n2982 = \P2_reg1_reg[9]/NET0131  & n2206 ;
  assign n2983 = ~\P2_reg3_reg[9]/NET0131  & ~n2217 ;
  assign n2984 = ~n2218 & ~n2983 ;
  assign n2985 = n2212 & n2984 ;
  assign n2988 = ~n2982 & ~n2985 ;
  assign n2986 = \P2_reg0_reg[9]/NET0131  & n2210 ;
  assign n2987 = \P2_reg2_reg[9]/NET0131  & n2208 ;
  assign n2989 = ~n2986 & ~n2987 ;
  assign n2990 = n2988 & n2989 ;
  assign n2991 = \P2_IR_reg[31]/NET0131  & \P2_IR_reg[8]/NET0131  ;
  assign n2992 = ~n2679 & ~n2991 ;
  assign n2993 = \P2_IR_reg[9]/NET0131  & ~n2992 ;
  assign n2994 = ~\P2_IR_reg[9]/NET0131  & n2992 ;
  assign n2995 = ~n2993 & ~n2994 ;
  assign n2996 = n2051 & ~n2995 ;
  assign n2997 = \P1_datao_reg[9]/NET0131  & ~n542 ;
  assign n2998 = ~n2108 & ~n2149 ;
  assign n3000 = n2148 & ~n2998 ;
  assign n2999 = ~n2148 & n2998 ;
  assign n3001 = n542 & ~n2999 ;
  assign n3002 = ~n3000 & n3001 ;
  assign n3003 = ~n2997 & ~n3002 ;
  assign n3004 = ~n2051 & n3003 ;
  assign n3005 = ~n2996 & ~n3004 ;
  assign n3006 = n2990 & ~n3005 ;
  assign n3007 = ~n2981 & ~n3006 ;
  assign n3008 = n2956 & n3007 ;
  assign n3009 = ~n2901 & n3008 ;
  assign n3010 = ~n2965 & n2980 ;
  assign n3011 = ~n2990 & n3005 ;
  assign n3012 = ~n2981 & n3011 ;
  assign n3013 = ~n3010 & ~n3012 ;
  assign n3014 = n2956 & ~n3013 ;
  assign n3015 = ~n2937 & n2954 ;
  assign n3016 = ~n2911 & n2926 ;
  assign n3017 = ~n3015 & ~n3016 ;
  assign n3018 = ~n2955 & ~n3017 ;
  assign n3019 = ~n3014 & ~n3018 ;
  assign n3020 = ~n3009 & n3019 ;
  assign n3021 = \P2_IR_reg[31]/NET0131  & ~n1970 ;
  assign n3022 = \P2_IR_reg[31]/NET0131  & ~n1972 ;
  assign n3023 = ~n3021 & ~n3022 ;
  assign n3024 = \P2_IR_reg[16]/NET0131  & ~n3023 ;
  assign n3025 = ~\P2_IR_reg[16]/NET0131  & n3023 ;
  assign n3026 = ~n3024 & ~n3025 ;
  assign n3027 = n2051 & ~n3026 ;
  assign n3028 = \P1_datao_reg[16]/NET0131  & ~n542 ;
  assign n3029 = ~n2086 & ~n2088 ;
  assign n3031 = n2284 & ~n3029 ;
  assign n3030 = ~n2284 & n3029 ;
  assign n3032 = n542 & ~n3030 ;
  assign n3033 = ~n3031 & n3032 ;
  assign n3034 = ~n3028 & ~n3033 ;
  assign n3035 = ~n2051 & n3034 ;
  assign n3036 = ~n3027 & ~n3035 ;
  assign n3040 = \P2_reg3_reg[15]/NET0131  & n2223 ;
  assign n3041 = ~\P2_reg3_reg[16]/NET0131  & ~n3040 ;
  assign n3042 = ~n2225 & ~n3041 ;
  assign n3043 = n2212 & n3042 ;
  assign n3039 = \P2_reg1_reg[16]/NET0131  & n2206 ;
  assign n3037 = \P2_reg2_reg[16]/NET0131  & n2208 ;
  assign n3038 = \P2_reg0_reg[16]/NET0131  & n2210 ;
  assign n3044 = ~n3037 & ~n3038 ;
  assign n3045 = ~n3039 & n3044 ;
  assign n3046 = ~n3043 & n3045 ;
  assign n3047 = ~n3036 & n3046 ;
  assign n3048 = \P2_reg0_reg[15]/NET0131  & n2210 ;
  assign n3049 = \P2_reg1_reg[15]/NET0131  & n2206 ;
  assign n3054 = ~n3048 & ~n3049 ;
  assign n3050 = ~\P2_reg3_reg[15]/NET0131  & ~n2223 ;
  assign n3051 = ~n3040 & ~n3050 ;
  assign n3052 = n2212 & n3051 ;
  assign n3053 = \P2_reg2_reg[15]/NET0131  & n2208 ;
  assign n3055 = ~n3052 & ~n3053 ;
  assign n3056 = n3054 & n3055 ;
  assign n3057 = \P2_IR_reg[14]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n3058 = ~n2642 & ~n3057 ;
  assign n3059 = \P2_IR_reg[15]/NET0131  & ~n3058 ;
  assign n3060 = ~\P2_IR_reg[15]/NET0131  & n3058 ;
  assign n3061 = ~n3059 & ~n3060 ;
  assign n3062 = n2051 & ~n3061 ;
  assign n3063 = \P1_datao_reg[15]/NET0131  & ~n542 ;
  assign n3064 = ~n2087 & ~n2091 ;
  assign n3066 = n2489 & ~n3064 ;
  assign n3065 = ~n2489 & n3064 ;
  assign n3067 = n542 & ~n3065 ;
  assign n3068 = ~n3066 & n3067 ;
  assign n3069 = ~n3063 & ~n3068 ;
  assign n3070 = ~n2051 & n3069 ;
  assign n3071 = ~n3062 & ~n3070 ;
  assign n3072 = n3056 & ~n3071 ;
  assign n3073 = ~n3047 & ~n3072 ;
  assign n3074 = \P2_reg2_reg[14]/NET0131  & n2208 ;
  assign n3075 = \P2_reg0_reg[14]/NET0131  & n2210 ;
  assign n3080 = ~n3074 & ~n3075 ;
  assign n3076 = ~\P2_reg3_reg[14]/NET0131  & ~n2222 ;
  assign n3077 = ~n2223 & ~n3076 ;
  assign n3078 = n2212 & n3077 ;
  assign n3079 = \P2_reg1_reg[14]/NET0131  & n2206 ;
  assign n3081 = ~n3078 & ~n3079 ;
  assign n3082 = n3080 & n3081 ;
  assign n3083 = ~\P2_IR_reg[14]/NET0131  & ~n2642 ;
  assign n3084 = ~n1996 & n3057 ;
  assign n3085 = ~n3083 & ~n3084 ;
  assign n3086 = n2051 & ~n3085 ;
  assign n3087 = \P1_datao_reg[14]/NET0131  & ~n542 ;
  assign n3088 = ~n2093 & ~n2095 ;
  assign n3090 = n2512 & ~n3088 ;
  assign n3089 = ~n2512 & n3088 ;
  assign n3091 = n542 & ~n3089 ;
  assign n3092 = ~n3090 & n3091 ;
  assign n3093 = ~n3087 & ~n3092 ;
  assign n3094 = ~n2051 & n3093 ;
  assign n3095 = ~n3086 & ~n3094 ;
  assign n3096 = n3082 & ~n3095 ;
  assign n3097 = \P2_reg0_reg[13]/NET0131  & n2210 ;
  assign n3098 = ~\P2_reg3_reg[13]/NET0131  & ~n2929 ;
  assign n3099 = ~n2222 & ~n3098 ;
  assign n3100 = n2212 & n3099 ;
  assign n3103 = ~n3097 & ~n3100 ;
  assign n3101 = \P2_reg1_reg[13]/NET0131  & n2206 ;
  assign n3102 = \P2_reg2_reg[13]/NET0131  & n2208 ;
  assign n3104 = ~n3101 & ~n3102 ;
  assign n3105 = n3103 & n3104 ;
  assign n3106 = \P2_IR_reg[13]/NET0131  & ~n3021 ;
  assign n3107 = ~\P2_IR_reg[13]/NET0131  & n3021 ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3109 = n2051 & n3108 ;
  assign n3110 = \P1_datao_reg[13]/NET0131  & ~n542 ;
  assign n3111 = ~n2094 & ~n2154 ;
  assign n3113 = n2153 & ~n3111 ;
  assign n3112 = ~n2153 & n3111 ;
  assign n3114 = n542 & ~n3112 ;
  assign n3115 = ~n3113 & n3114 ;
  assign n3116 = ~n3110 & ~n3115 ;
  assign n3117 = ~n2051 & n3116 ;
  assign n3118 = ~n3109 & ~n3117 ;
  assign n3119 = n3105 & ~n3118 ;
  assign n3120 = ~n3096 & ~n3119 ;
  assign n3121 = n3073 & n3120 ;
  assign n3122 = ~n3020 & n3121 ;
  assign n3123 = n2669 & n3122 ;
  assign n3124 = ~n3082 & n3095 ;
  assign n3125 = ~n3105 & n3118 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = ~n3096 & ~n3126 ;
  assign n3128 = n3073 & n3127 ;
  assign n3129 = n3036 & ~n3046 ;
  assign n3130 = ~n3056 & n3071 ;
  assign n3131 = ~n3047 & n3130 ;
  assign n3132 = ~n3129 & ~n3131 ;
  assign n3133 = ~n3128 & n3132 ;
  assign n3134 = n2669 & ~n3133 ;
  assign n3135 = n2657 & ~n2666 ;
  assign n3136 = n2630 & ~n2640 ;
  assign n3137 = ~n3135 & ~n3136 ;
  assign n3138 = ~n2667 & ~n3137 ;
  assign n3139 = n2615 & n3138 ;
  assign n3140 = n2579 & ~n2588 ;
  assign n3141 = n2604 & ~n2613 ;
  assign n3142 = ~n2589 & n3141 ;
  assign n3143 = ~n3140 & ~n3142 ;
  assign n3144 = ~n3139 & n3143 ;
  assign n3145 = ~n3134 & n3144 ;
  assign n3146 = ~n3123 & n3145 ;
  assign n3147 = ~n2541 & n2551 ;
  assign n3148 = ~n2533 & ~n3147 ;
  assign n3149 = n2509 & n3148 ;
  assign n3150 = ~n2329 & n3149 ;
  assign n3151 = n2463 & n3150 ;
  assign n3152 = ~n3146 & n3151 ;
  assign n3153 = ~n2571 & ~n3152 ;
  assign n3154 = n2244 & ~n3153 ;
  assign n3155 = ~n2244 & n3153 ;
  assign n3156 = ~n3154 & ~n3155 ;
  assign n3157 = n2033 & ~n3156 ;
  assign n3158 = ~n2034 & ~n3157 ;
  assign n3159 = ~\P2_IR_reg[20]/NET0131  & ~n2002 ;
  assign n3160 = \P2_IR_reg[20]/NET0131  & n2002 ;
  assign n3161 = ~n3159 & ~n3160 ;
  assign n3162 = ~\P2_IR_reg[20]/NET0131  & n1987 ;
  assign n3163 = \P2_IR_reg[31]/NET0131  & ~n3162 ;
  assign n3164 = ~n2616 & ~n3163 ;
  assign n3165 = \P2_IR_reg[21]/NET0131  & ~n3164 ;
  assign n3166 = ~\P2_IR_reg[21]/NET0131  & n3164 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = n3161 & n3167 ;
  assign n3169 = \P2_IR_reg[31]/NET0131  & ~n1977 ;
  assign n3170 = ~n2002 & ~n3169 ;
  assign n3171 = \P2_IR_reg[22]/NET0131  & ~n3170 ;
  assign n3172 = ~\P2_IR_reg[22]/NET0131  & n3170 ;
  assign n3173 = ~n3171 & ~n3172 ;
  assign n3174 = n2592 & n3173 ;
  assign n3175 = ~n3168 & ~n3174 ;
  assign n3176 = n3167 & n3173 ;
  assign n3177 = ~n3167 & ~n3173 ;
  assign n3178 = ~n3176 & ~n3177 ;
  assign n3179 = n3175 & n3178 ;
  assign n3180 = ~n3158 & n3179 ;
  assign n3181 = n2911 & n2926 ;
  assign n3182 = n2937 & n2954 ;
  assign n3183 = ~n3181 & ~n3182 ;
  assign n3184 = n2965 & n2980 ;
  assign n3185 = ~n2965 & ~n2980 ;
  assign n3186 = ~n2990 & ~n3005 ;
  assign n3187 = ~n3185 & ~n3186 ;
  assign n3188 = ~n3184 & ~n3187 ;
  assign n3189 = n3183 & n3188 ;
  assign n3190 = ~n2937 & ~n2954 ;
  assign n3191 = ~n2911 & ~n2926 ;
  assign n3192 = ~n3182 & n3191 ;
  assign n3193 = ~n3190 & ~n3192 ;
  assign n3194 = ~n3189 & n3193 ;
  assign n3195 = n2678 & n2692 ;
  assign n3196 = n2702 & n2719 ;
  assign n3197 = ~n3195 & ~n3196 ;
  assign n3198 = n2823 & ~n2830 ;
  assign n3199 = n2800 & ~n2814 ;
  assign n3200 = ~n3198 & ~n3199 ;
  assign n3201 = ~n2800 & n2814 ;
  assign n3202 = ~n2777 & n2791 ;
  assign n3203 = ~n3201 & ~n3202 ;
  assign n3204 = ~n3200 & n3203 ;
  assign n3205 = ~n2849 & n2858 ;
  assign n3206 = n2866 & ~n2880 ;
  assign n3207 = n2777 & ~n2791 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = ~n3205 & n3208 ;
  assign n3210 = ~n3204 & n3209 ;
  assign n3211 = n2849 & ~n2858 ;
  assign n3212 = ~n2866 & n2880 ;
  assign n3213 = ~n3211 & ~n3212 ;
  assign n3214 = ~n3205 & ~n3213 ;
  assign n3215 = ~n3210 & ~n3214 ;
  assign n3216 = n2730 & n2745 ;
  assign n3217 = n2755 & n2768 ;
  assign n3218 = ~n3216 & ~n3217 ;
  assign n3219 = ~n3215 & n3218 ;
  assign n3220 = ~n2730 & ~n2745 ;
  assign n3221 = ~n2755 & ~n2768 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = ~n3216 & ~n3222 ;
  assign n3224 = ~n3219 & ~n3223 ;
  assign n3225 = n3197 & ~n3224 ;
  assign n3226 = ~n2678 & ~n2692 ;
  assign n3227 = ~n2702 & ~n2719 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = ~n3195 & ~n3228 ;
  assign n3230 = ~n3225 & ~n3229 ;
  assign n3231 = n2990 & n3005 ;
  assign n3232 = ~n3184 & ~n3231 ;
  assign n3233 = n3183 & n3232 ;
  assign n3234 = ~n3230 & n3233 ;
  assign n3235 = n3194 & ~n3234 ;
  assign n3236 = n2579 & n2588 ;
  assign n3237 = n2604 & n2613 ;
  assign n3238 = ~n3236 & ~n3237 ;
  assign n3239 = n2630 & n2640 ;
  assign n3240 = n2657 & n2666 ;
  assign n3241 = ~n3239 & ~n3240 ;
  assign n3242 = n3238 & n3241 ;
  assign n3243 = n3036 & n3046 ;
  assign n3244 = n3056 & n3071 ;
  assign n3245 = ~n3243 & ~n3244 ;
  assign n3246 = n3082 & n3095 ;
  assign n3247 = n3105 & n3118 ;
  assign n3248 = ~n3246 & ~n3247 ;
  assign n3249 = n3245 & n3248 ;
  assign n3250 = n3242 & n3249 ;
  assign n3251 = ~n3235 & n3250 ;
  assign n3252 = ~n3082 & ~n3095 ;
  assign n3253 = ~n3105 & ~n3118 ;
  assign n3254 = ~n3252 & ~n3253 ;
  assign n3255 = ~n3246 & ~n3254 ;
  assign n3256 = n3245 & n3255 ;
  assign n3257 = ~n3036 & ~n3046 ;
  assign n3258 = ~n3056 & ~n3071 ;
  assign n3259 = ~n3243 & n3258 ;
  assign n3260 = ~n3257 & ~n3259 ;
  assign n3261 = ~n3256 & n3260 ;
  assign n3262 = n3242 & ~n3261 ;
  assign n3263 = ~n2630 & ~n2640 ;
  assign n3264 = ~n2657 & ~n2666 ;
  assign n3265 = ~n3263 & ~n3264 ;
  assign n3266 = ~n3240 & ~n3265 ;
  assign n3267 = n3238 & n3266 ;
  assign n3268 = ~n2579 & ~n2588 ;
  assign n3269 = ~n2604 & ~n2613 ;
  assign n3270 = ~n3268 & ~n3269 ;
  assign n3271 = ~n3236 & ~n3270 ;
  assign n3272 = ~n3267 & ~n3271 ;
  assign n3273 = ~n3262 & n3272 ;
  assign n3274 = ~n3251 & n3273 ;
  assign n3275 = n2315 & n2328 ;
  assign n3276 = n2376 & n2385 ;
  assign n3277 = ~n3275 & ~n3276 ;
  assign n3278 = n2424 & n2433 ;
  assign n3279 = n2452 & n2461 ;
  assign n3280 = ~n3278 & ~n3279 ;
  assign n3281 = n3277 & n3280 ;
  assign n3282 = n2498 & n2507 ;
  assign n3283 = n2471 & n2484 ;
  assign n3284 = ~n3282 & ~n3283 ;
  assign n3285 = n2522 & n2531 ;
  assign n3286 = n2541 & n2551 ;
  assign n3287 = ~n3285 & ~n3286 ;
  assign n3288 = n3284 & n3287 ;
  assign n3289 = n3281 & n3288 ;
  assign n3290 = ~n3274 & n3289 ;
  assign n3291 = ~n2522 & ~n2531 ;
  assign n3292 = ~n2541 & ~n2551 ;
  assign n3293 = ~n3291 & ~n3292 ;
  assign n3294 = ~n3285 & ~n3293 ;
  assign n3295 = n3284 & n3294 ;
  assign n3296 = ~n2471 & ~n2484 ;
  assign n3297 = ~n2498 & ~n2507 ;
  assign n3298 = ~n3283 & n3297 ;
  assign n3299 = ~n3296 & ~n3298 ;
  assign n3300 = ~n3295 & n3299 ;
  assign n3301 = n3281 & ~n3300 ;
  assign n3302 = ~n2424 & ~n2433 ;
  assign n3303 = ~n2452 & ~n2461 ;
  assign n3304 = ~n3302 & ~n3303 ;
  assign n3305 = ~n3278 & ~n3304 ;
  assign n3306 = n3277 & n3305 ;
  assign n3307 = ~n2315 & ~n2328 ;
  assign n3308 = ~n2376 & ~n2385 ;
  assign n3309 = ~n3307 & ~n3308 ;
  assign n3310 = ~n3275 & ~n3309 ;
  assign n3311 = ~n3306 & ~n3310 ;
  assign n3312 = ~n3301 & n3311 ;
  assign n3313 = ~n3290 & n3312 ;
  assign n3314 = ~n2244 & n3313 ;
  assign n3315 = n2244 & ~n3313 ;
  assign n3316 = ~n3314 & ~n3315 ;
  assign n3317 = n2033 & n3316 ;
  assign n3318 = ~n2034 & ~n3317 ;
  assign n3319 = ~n3175 & ~n3176 ;
  assign n3320 = ~n3318 & n3319 ;
  assign n3321 = n2050 & ~n2328 ;
  assign n3326 = \P2_reg2_reg[31]/NET0131  & n2208 ;
  assign n3324 = \P2_reg0_reg[31]/NET0131  & n2210 ;
  assign n3325 = \P2_reg1_reg[31]/NET0131  & n2206 ;
  assign n3327 = ~n3324 & ~n3325 ;
  assign n3328 = ~n3326 & n3327 ;
  assign n3329 = ~n2238 & n3328 ;
  assign n3330 = ~n2823 & ~n3329 ;
  assign n3331 = ~n2800 & n3330 ;
  assign n3332 = ~n2777 & n3331 ;
  assign n3333 = ~n2866 & n3332 ;
  assign n3334 = ~n2858 & n3333 ;
  assign n3335 = ~n2702 & ~n2730 ;
  assign n3336 = ~n2755 & n3335 ;
  assign n3337 = n3334 & n3336 ;
  assign n3338 = ~n2678 & ~n2990 ;
  assign n3339 = n3337 & n3338 ;
  assign n3340 = ~n2911 & ~n2937 ;
  assign n3341 = ~n2965 & n3340 ;
  assign n3342 = n3339 & n3341 ;
  assign n3343 = ~n3082 & ~n3105 ;
  assign n3344 = n3342 & n3343 ;
  assign n3346 = ~n2613 & ~n3056 ;
  assign n3347 = ~n2666 & n3346 ;
  assign n3345 = ~n2640 & ~n3046 ;
  assign n3348 = ~n2588 & n3345 ;
  assign n3349 = n3347 & n3348 ;
  assign n3350 = ~n2551 & n3349 ;
  assign n3351 = ~n2507 & ~n2531 ;
  assign n3352 = n3350 & n3351 ;
  assign n3353 = ~n2484 & n3352 ;
  assign n3354 = ~n2461 & n3353 ;
  assign n3355 = n3344 & n3354 ;
  assign n3322 = ~n2385 & ~n2433 ;
  assign n3323 = ~n2328 & n3322 ;
  assign n3356 = ~n2241 & n3323 ;
  assign n3357 = n3355 & n3356 ;
  assign n3360 = \P2_reg1_reg[30]/NET0131  & n2206 ;
  assign n3358 = \P2_reg0_reg[30]/NET0131  & n2210 ;
  assign n3359 = \P2_reg2_reg[30]/NET0131  & n2208 ;
  assign n3361 = ~n3358 & ~n3359 ;
  assign n3362 = ~n3360 & n3361 ;
  assign n3363 = ~n2238 & n3362 ;
  assign n3364 = ~n3357 & n3363 ;
  assign n3365 = n3357 & ~n3363 ;
  assign n3366 = \P2_B_reg/NET0131  & n2043 ;
  assign n3367 = ~n2050 & ~n3366 ;
  assign n3368 = ~n3365 & n3367 ;
  assign n3369 = ~n3364 & n3368 ;
  assign n3370 = ~n3321 & ~n3369 ;
  assign n3371 = ~n2592 & ~n3161 ;
  assign n3372 = n3167 & n3371 ;
  assign n3373 = n3173 & n3372 ;
  assign n3374 = ~n3370 & n3373 ;
  assign n3375 = n3161 & n3177 ;
  assign n3376 = n2191 & n3375 ;
  assign n3377 = n2814 & n2830 ;
  assign n3378 = n2791 & n3377 ;
  assign n3379 = n2880 & n3378 ;
  assign n3380 = n2849 & n3379 ;
  assign n3381 = ~n2768 & n3380 ;
  assign n3382 = ~n2745 & n3381 ;
  assign n3383 = ~n2719 & n3382 ;
  assign n3384 = ~n2692 & n3383 ;
  assign n3385 = ~n2980 & ~n3005 ;
  assign n3386 = ~n2926 & n3385 ;
  assign n3387 = n3384 & n3386 ;
  assign n3388 = ~n2954 & ~n3118 ;
  assign n3389 = n3387 & n3388 ;
  assign n3390 = ~n2579 & ~n2630 ;
  assign n3391 = ~n2657 & n3390 ;
  assign n3392 = ~n2604 & n3391 ;
  assign n3393 = ~n2541 & n3392 ;
  assign n3394 = ~n2498 & ~n2522 ;
  assign n3395 = n3393 & n3394 ;
  assign n3396 = n3389 & n3395 ;
  assign n3397 = ~n3036 & ~n3095 ;
  assign n3398 = ~n3071 & n3397 ;
  assign n3399 = ~n2452 & n3398 ;
  assign n3400 = ~n2471 & n3399 ;
  assign n3401 = ~n2376 & ~n2424 ;
  assign n3402 = n3400 & n3401 ;
  assign n3403 = n3396 & n3402 ;
  assign n3404 = ~n2315 & n3403 ;
  assign n3405 = n2191 & ~n3404 ;
  assign n3406 = ~n2191 & n3404 ;
  assign n3407 = ~n3405 & ~n3406 ;
  assign n3408 = ~n3167 & n3371 ;
  assign n3409 = ~n3173 & n3408 ;
  assign n3410 = n3407 & n3409 ;
  assign n3411 = ~n3376 & ~n3410 ;
  assign n3412 = ~n3374 & n3411 ;
  assign n3413 = n2033 & ~n3412 ;
  assign n3414 = n2592 & ~n3161 ;
  assign n3415 = n3177 & n3414 ;
  assign n3416 = n2237 & n3415 ;
  assign n3417 = ~n2033 & n3373 ;
  assign n3418 = n3176 & ~n3371 ;
  assign n3419 = n2033 & ~n3418 ;
  assign n3420 = n3177 & ~n3414 ;
  assign n3421 = ~n3418 & ~n3420 ;
  assign n3422 = ~n3419 & ~n3421 ;
  assign n3423 = ~n3417 & ~n3422 ;
  assign n3424 = \P2_reg2_reg[29]/NET0131  & ~n3423 ;
  assign n3425 = ~n3416 & ~n3424 ;
  assign n3426 = ~n3413 & n3425 ;
  assign n3427 = ~n3320 & n3426 ;
  assign n3428 = ~n3180 & n3427 ;
  assign n3429 = n2017 & ~n3428 ;
  assign n3430 = ~n1984 & n2016 ;
  assign n3431 = \P2_reg2_reg[29]/NET0131  & n3430 ;
  assign n3432 = ~n3429 & ~n3431 ;
  assign n3433 = \P1_state_reg[0]/NET0131  & ~n3432 ;
  assign n3434 = \P1_state_reg[0]/NET0131  & ~n1984 ;
  assign n3435 = \P2_reg2_reg[29]/NET0131  & ~n3434 ;
  assign n3436 = ~n3433 & ~n3435 ;
  assign n3438 = \P1_B_reg/NET0131  & ~n1944 ;
  assign n3439 = ~\P1_B_reg/NET0131  & n1944 ;
  assign n3440 = ~n3438 & ~n3439 ;
  assign n3441 = ~n1939 & ~n1949 ;
  assign n3442 = ~n3440 & n3441 ;
  assign n3437 = \P1_d_reg[0]/NET0131  & ~n1939 ;
  assign n3443 = n1939 & n1944 ;
  assign n3444 = ~n3437 & ~n3443 ;
  assign n3445 = ~n3442 & n3444 ;
  assign n3446 = \P1_d_reg[1]/NET0131  & ~n1939 ;
  assign n3447 = n1939 & n1949 ;
  assign n3448 = ~n3446 & ~n3447 ;
  assign n3449 = ~n3442 & n3448 ;
  assign n3450 = ~n3445 & ~n3449 ;
  assign n3451 = n1642 & ~n3450 ;
  assign n3452 = n1138 & n1151 ;
  assign n3453 = n1115 & n1128 ;
  assign n3454 = ~n3452 & ~n3453 ;
  assign n3455 = ~n1189 & ~n1202 ;
  assign n3456 = ~n1747 & n3455 ;
  assign n3457 = ~n1748 & ~n3456 ;
  assign n3458 = n3454 & ~n3457 ;
  assign n3459 = ~n1138 & ~n1151 ;
  assign n3460 = ~n1115 & ~n1128 ;
  assign n3461 = ~n3459 & ~n3460 ;
  assign n3462 = ~n3453 & ~n3461 ;
  assign n3463 = ~n3458 & ~n3462 ;
  assign n3464 = n1222 & n1238 ;
  assign n3465 = ~n1741 & ~n3464 ;
  assign n3467 = ~n1390 & ~n1397 ;
  assign n3468 = n1367 & n1381 ;
  assign n3469 = n3467 & ~n3468 ;
  assign n3470 = ~n1367 & ~n1381 ;
  assign n3471 = ~n3469 & ~n3470 ;
  assign n3472 = n1344 & n1358 ;
  assign n3473 = ~n1744 & ~n3472 ;
  assign n3474 = ~n3471 & n3473 ;
  assign n3475 = ~n1344 & ~n1358 ;
  assign n3476 = ~n1745 & ~n3475 ;
  assign n3477 = ~n1744 & ~n3476 ;
  assign n3478 = ~n3474 & ~n3477 ;
  assign n3466 = n1274 & n1288 ;
  assign n3479 = ~n1752 & ~n3466 ;
  assign n3480 = ~n3478 & n3479 ;
  assign n3481 = ~n1274 & ~n1288 ;
  assign n3482 = ~n1751 & ~n3481 ;
  assign n3483 = ~n3466 & ~n3482 ;
  assign n3484 = ~n3480 & ~n3483 ;
  assign n3485 = n3465 & ~n3484 ;
  assign n3486 = ~n1222 & ~n1238 ;
  assign n3487 = ~n1741 & n3486 ;
  assign n3488 = ~n1742 & ~n3487 ;
  assign n3489 = ~n3485 & n3488 ;
  assign n3490 = n1189 & n1202 ;
  assign n3491 = ~n1747 & ~n3490 ;
  assign n3492 = n3454 & n3491 ;
  assign n3493 = ~n3489 & n3492 ;
  assign n3494 = n3463 & ~n3493 ;
  assign n3495 = n785 & n796 ;
  assign n3496 = n829 & n838 ;
  assign n3497 = ~n3495 & ~n3496 ;
  assign n3498 = n638 & n692 ;
  assign n3499 = ~n1798 & ~n3498 ;
  assign n3500 = n3497 & n3499 ;
  assign n3501 = n1026 & n1040 ;
  assign n3502 = ~n1763 & ~n3501 ;
  assign n3503 = n1051 & n1064 ;
  assign n3504 = ~n1761 & ~n3503 ;
  assign n3505 = n3502 & n3504 ;
  assign n3506 = n3500 & n3505 ;
  assign n3507 = ~n3494 & n3506 ;
  assign n3508 = ~n1051 & ~n1064 ;
  assign n3509 = ~n1760 & ~n3508 ;
  assign n3510 = ~n3503 & ~n3509 ;
  assign n3511 = n3502 & n3510 ;
  assign n3512 = ~n1026 & ~n1040 ;
  assign n3513 = ~n1763 & n3512 ;
  assign n3514 = ~n1764 & ~n3513 ;
  assign n3515 = ~n3511 & n3514 ;
  assign n3516 = n3500 & ~n3515 ;
  assign n3517 = ~n785 & ~n796 ;
  assign n3518 = ~n829 & ~n838 ;
  assign n3519 = ~n3495 & n3518 ;
  assign n3520 = ~n3517 & ~n3519 ;
  assign n3521 = n3499 & ~n3520 ;
  assign n3522 = ~n638 & ~n692 ;
  assign n3523 = n1797 & ~n3498 ;
  assign n3524 = ~n3522 & ~n3523 ;
  assign n3525 = ~n3521 & n3524 ;
  assign n3526 = ~n3516 & n3525 ;
  assign n3527 = ~n3507 & n3526 ;
  assign n3528 = ~n1770 & ~n1789 ;
  assign n3529 = ~n1767 & ~n1781 ;
  assign n3530 = n3528 & n3529 ;
  assign n3531 = ~n1777 & ~n1794 ;
  assign n3532 = ~n1775 & ~n1784 ;
  assign n3533 = n3531 & n3532 ;
  assign n3534 = n3530 & n3533 ;
  assign n3535 = ~n3527 & n3534 ;
  assign n3540 = n1774 & ~n1784 ;
  assign n3541 = ~n1785 & ~n3540 ;
  assign n3542 = n3531 & ~n3541 ;
  assign n3543 = n1778 & ~n1794 ;
  assign n3544 = ~n1795 & ~n3543 ;
  assign n3545 = ~n3542 & n3544 ;
  assign n3546 = n3530 & ~n3545 ;
  assign n3536 = ~n1767 & n1782 ;
  assign n3537 = ~n1768 & ~n3536 ;
  assign n3538 = ~n1771 & n3537 ;
  assign n3539 = n3528 & ~n3538 ;
  assign n3547 = ~n1788 & ~n3539 ;
  assign n3548 = ~n3546 & n3547 ;
  assign n3549 = ~n3535 & n3548 ;
  assign n3550 = n1793 & n3549 ;
  assign n3551 = ~n1793 & ~n3549 ;
  assign n3552 = ~n3550 & ~n3551 ;
  assign n3553 = n3450 & ~n3552 ;
  assign n3554 = ~n3451 & ~n3553 ;
  assign n3555 = ~n499 & ~n1911 ;
  assign n3556 = ~n1735 & ~n1897 ;
  assign n3557 = n3555 & n3556 ;
  assign n3558 = ~n3554 & n3557 ;
  assign n3559 = n1211 & ~n1423 ;
  assign n3560 = n1106 & n1429 ;
  assign n3561 = ~n3559 & n3560 ;
  assign n3562 = ~n1103 & n1429 ;
  assign n3563 = n847 & ~n3562 ;
  assign n3564 = ~n3561 & n3563 ;
  assign n3565 = n1426 & n1573 ;
  assign n3566 = ~n3564 & n3565 ;
  assign n3567 = ~n982 & n1573 ;
  assign n3568 = n1583 & ~n3567 ;
  assign n3569 = ~n3566 & n3568 ;
  assign n3570 = n1793 & ~n3569 ;
  assign n3571 = ~n1793 & n3569 ;
  assign n3572 = ~n3570 & ~n3571 ;
  assign n3573 = n3450 & ~n3572 ;
  assign n3574 = ~n3451 & ~n3573 ;
  assign n3575 = ~n1897 & ~n3555 ;
  assign n3576 = ~n3574 & n3575 ;
  assign n3577 = ~n1390 & ~n1677 ;
  assign n3578 = ~n1367 & n3577 ;
  assign n3579 = ~n1344 & n3578 ;
  assign n3580 = ~n1322 & n3579 ;
  assign n3581 = ~n1298 & n3580 ;
  assign n3582 = ~n1162 & ~n1189 ;
  assign n3583 = ~n1222 & ~n1248 ;
  assign n3584 = ~n1274 & n3583 ;
  assign n3585 = n3582 & n3584 ;
  assign n3586 = n3581 & n3585 ;
  assign n3587 = ~n1138 & n3586 ;
  assign n3588 = ~n1026 & ~n1051 ;
  assign n3589 = ~n999 & ~n1075 ;
  assign n3590 = ~n1115 & n3589 ;
  assign n3591 = n3588 & n3590 ;
  assign n3592 = n3587 & n3591 ;
  assign n3593 = ~n838 & n3592 ;
  assign n3594 = ~n692 & ~n973 ;
  assign n3595 = ~n887 & ~n949 ;
  assign n3596 = n3594 & n3595 ;
  assign n3597 = ~n921 & n3596 ;
  assign n3598 = ~n1542 & ~n1570 ;
  assign n3599 = n3597 & n3598 ;
  assign n3600 = ~n1478 & ~n1510 ;
  assign n3601 = n3599 & n3600 ;
  assign n3602 = ~n752 & ~n796 ;
  assign n3603 = ~n1646 & n3602 ;
  assign n3604 = n3601 & n3603 ;
  assign n3605 = n3593 & n3604 ;
  assign n3606 = ~n1618 & ~n3605 ;
  assign n3607 = n1618 & n3605 ;
  assign n3608 = ~n3606 & ~n3607 ;
  assign n3609 = ~n536 & ~n3608 ;
  assign n3610 = n536 & ~n1510 ;
  assign n3611 = ~n3609 & ~n3610 ;
  assign n3612 = n3450 & ~n3611 ;
  assign n3613 = ~n3451 & ~n3612 ;
  assign n3614 = n1898 & ~n3613 ;
  assign n3620 = n743 & n829 ;
  assign n3621 = n785 & n3620 ;
  assign n3622 = ~n875 & ~n939 ;
  assign n3623 = n638 & n3622 ;
  assign n3624 = ~n964 & n3623 ;
  assign n3625 = n3621 & n3624 ;
  assign n3626 = n1381 & n1397 ;
  assign n3627 = n1358 & n3626 ;
  assign n3628 = n1336 & n3627 ;
  assign n3629 = n1313 & n3628 ;
  assign n3630 = n1288 & n3629 ;
  assign n3631 = n1238 & n1263 ;
  assign n3632 = n3630 & n3631 ;
  assign n3633 = n1178 & n1202 ;
  assign n3634 = n3632 & n3633 ;
  assign n3635 = n1128 & n1151 ;
  assign n3636 = n3634 & n3635 ;
  assign n3637 = n1015 & n1040 ;
  assign n3638 = n1064 & n1094 ;
  assign n3639 = n3637 & n3638 ;
  assign n3640 = n3636 & n3639 ;
  assign n3641 = n3625 & n3640 ;
  assign n3642 = ~n911 & ~n1561 ;
  assign n3643 = ~n1463 & ~n1533 ;
  assign n3644 = n3642 & n3643 ;
  assign n3645 = ~n1500 & n3644 ;
  assign n3646 = n3641 & n3645 ;
  assign n3647 = ~n1637 & n3646 ;
  assign n3648 = n1637 & ~n3646 ;
  assign n3649 = ~n3647 & ~n3648 ;
  assign n3650 = n1731 & n1735 ;
  assign n3651 = n3649 & n3650 ;
  assign n3652 = n3450 & n3651 ;
  assign n3615 = ~n1731 & n1897 ;
  assign n3616 = ~n1734 & n1735 ;
  assign n3617 = ~n3450 & n3616 ;
  assign n3618 = ~n3615 & ~n3617 ;
  assign n3619 = n1642 & ~n3618 ;
  assign n3653 = ~n1736 & ~n3450 ;
  assign n3654 = ~n1731 & n1735 ;
  assign n3655 = ~n3653 & n3654 ;
  assign n3656 = n1637 & n3655 ;
  assign n3657 = ~n3619 & ~n3656 ;
  assign n3658 = ~n3652 & n3657 ;
  assign n3659 = ~n3614 & n3658 ;
  assign n3660 = ~n3576 & n3659 ;
  assign n3661 = ~n3558 & n3660 ;
  assign n3662 = ~n1933 & ~n1951 ;
  assign n3663 = ~n3661 & n3662 ;
  assign n3664 = ~n1933 & n1951 ;
  assign n3665 = n1642 & n3664 ;
  assign n3666 = ~n3663 & ~n3665 ;
  assign n3667 = \P1_state_reg[0]/NET0131  & ~n3666 ;
  assign n3668 = \P1_reg3_reg[28]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n3669 = n1642 & n1934 ;
  assign n3670 = ~n3668 & ~n3669 ;
  assign n3671 = ~n3667 & n3670 ;
  assign n3672 = n3445 & ~n3449 ;
  assign n3673 = \P1_reg2_reg[28]/NET0131  & ~n3672 ;
  assign n3674 = ~n3552 & n3672 ;
  assign n3675 = ~n3673 & ~n3674 ;
  assign n3676 = n3557 & ~n3675 ;
  assign n3677 = ~n3572 & n3672 ;
  assign n3678 = ~n3673 & ~n3677 ;
  assign n3679 = n3575 & ~n3678 ;
  assign n3680 = ~n3611 & n3672 ;
  assign n3681 = ~n3673 & ~n3680 ;
  assign n3682 = n1898 & ~n3681 ;
  assign n3687 = n3649 & n3672 ;
  assign n3688 = ~n3673 & ~n3687 ;
  assign n3689 = n3650 & ~n3688 ;
  assign n3683 = n498 & n1735 ;
  assign n3691 = n1637 & n3683 ;
  assign n3692 = n3672 & n3691 ;
  assign n3684 = ~n3672 & n3683 ;
  assign n3685 = ~n3615 & ~n3684 ;
  assign n3686 = \P1_reg2_reg[28]/NET0131  & ~n3685 ;
  assign n3690 = n1642 & n1736 ;
  assign n3693 = ~n3686 & ~n3690 ;
  assign n3694 = ~n3692 & n3693 ;
  assign n3695 = ~n3689 & n3694 ;
  assign n3696 = ~n3682 & n3695 ;
  assign n3697 = ~n3679 & n3696 ;
  assign n3698 = ~n3676 & n3697 ;
  assign n3699 = n3662 & ~n3698 ;
  assign n3700 = \P1_reg2_reg[28]/NET0131  & n3664 ;
  assign n3701 = ~n3699 & ~n3700 ;
  assign n3702 = \P1_state_reg[0]/NET0131  & ~n3701 ;
  assign n3703 = \P1_state_reg[0]/NET0131  & ~n1933 ;
  assign n3704 = \P1_reg2_reg[28]/NET0131  & ~n3703 ;
  assign n3705 = ~n3702 & ~n3704 ;
  assign n3706 = \P1_reg2_reg[29]/NET0131  & ~n3703 ;
  assign n3707 = \P1_reg2_reg[29]/NET0131  & n3664 ;
  assign n3708 = \P1_reg2_reg[29]/NET0131  & ~n3672 ;
  assign n3709 = n536 & ~n1646 ;
  assign n3710 = ~n838 & n3602 ;
  assign n3711 = n3592 & n3710 ;
  assign n3712 = n3601 & n3711 ;
  assign n3713 = ~n1646 & n3712 ;
  assign n3714 = ~n1618 & n3713 ;
  assign n3715 = n1702 & ~n3714 ;
  assign n3716 = ~n1702 & n3714 ;
  assign n3717 = \P1_B_reg/NET0131  & ~n527 ;
  assign n3718 = ~n536 & ~n3717 ;
  assign n3719 = ~n3716 & n3718 ;
  assign n3720 = ~n3715 & n3719 ;
  assign n3721 = ~n3709 & ~n3720 ;
  assign n3722 = n3672 & ~n3721 ;
  assign n3723 = ~n3708 & ~n3722 ;
  assign n3724 = n1898 & ~n3723 ;
  assign n3806 = ~n693 & ~n984 ;
  assign n3807 = ~n753 & ~n797 ;
  assign n3808 = n3806 & n3807 ;
  assign n3809 = ~n1041 & ~n1065 ;
  assign n3810 = ~n1016 & ~n1427 ;
  assign n3811 = n3809 & n3810 ;
  assign n3812 = n3808 & n3811 ;
  assign n3813 = ~n1104 & ~n1129 ;
  assign n3814 = ~n1152 & ~n1861 ;
  assign n3815 = n3813 & n3814 ;
  assign n3816 = ~n1104 & n1208 ;
  assign n3817 = ~n1095 & ~n3816 ;
  assign n3818 = ~n3815 & n3817 ;
  assign n3819 = ~n1399 & n1870 ;
  assign n3820 = ~n1314 & n1360 ;
  assign n3821 = ~n3819 & n3820 ;
  assign n3822 = ~n1314 & ~n1873 ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3824 = ~n1264 & ~n1420 ;
  assign n3825 = ~n1239 & ~n1289 ;
  assign n3826 = n3824 & n3825 ;
  assign n3827 = ~n3823 & n3826 ;
  assign n3828 = ~n1239 & ~n1867 ;
  assign n3829 = n3824 & n3828 ;
  assign n3830 = ~n1203 & ~n1414 ;
  assign n3831 = ~n1420 & ~n3830 ;
  assign n3832 = ~n3829 & ~n3831 ;
  assign n3833 = ~n3827 & n3832 ;
  assign n3834 = ~n1152 & ~n1179 ;
  assign n3835 = n3813 & n3834 ;
  assign n3836 = ~n3833 & n3835 ;
  assign n3837 = n3818 & ~n3836 ;
  assign n3838 = n3812 & ~n3837 ;
  assign n3839 = ~n1041 & ~n1857 ;
  assign n3840 = n3810 & n3839 ;
  assign n3841 = ~n839 & ~n1100 ;
  assign n3842 = ~n1427 & ~n3841 ;
  assign n3843 = ~n3840 & ~n3842 ;
  assign n3844 = n3808 & ~n3843 ;
  assign n3845 = ~n753 & ~n1851 ;
  assign n3846 = n3806 & n3845 ;
  assign n3847 = ~n844 & ~n974 ;
  assign n3848 = ~n984 & ~n3847 ;
  assign n3849 = ~n3846 & ~n3848 ;
  assign n3850 = ~n3844 & n3849 ;
  assign n3851 = ~n3838 & n3850 ;
  assign n3852 = ~n888 & ~n950 ;
  assign n3853 = ~n922 & ~n1571 ;
  assign n3854 = n3852 & n3853 ;
  assign n3855 = ~n1479 & ~n1543 ;
  assign n3856 = ~n1511 & ~n1647 ;
  assign n3857 = n3855 & n3856 ;
  assign n3858 = n3854 & n3857 ;
  assign n3859 = ~n3851 & n3858 ;
  assign n3860 = ~n888 & ~n986 ;
  assign n3861 = n3853 & n3860 ;
  assign n3862 = ~n978 & ~n1578 ;
  assign n3863 = ~n1571 & ~n3862 ;
  assign n3864 = ~n3861 & ~n3863 ;
  assign n3865 = n3857 & ~n3864 ;
  assign n3866 = ~n1479 & ~n1845 ;
  assign n3867 = ~n1575 & ~n3866 ;
  assign n3868 = n3856 & ~n3867 ;
  assign n3869 = ~n1710 & ~n3868 ;
  assign n3870 = ~n3865 & n3869 ;
  assign n3871 = ~n3859 & n3870 ;
  assign n3872 = ~n1780 & n3871 ;
  assign n3873 = n1780 & ~n3871 ;
  assign n3874 = ~n3872 & ~n3873 ;
  assign n3875 = n3672 & n3874 ;
  assign n3876 = ~n3708 & ~n3875 ;
  assign n3877 = n3575 & ~n3876 ;
  assign n3725 = ~n1747 & ~n3452 ;
  assign n3726 = ~n1761 & ~n3453 ;
  assign n3727 = n3725 & n3726 ;
  assign n3728 = ~n3470 & ~n3475 ;
  assign n3729 = ~n3469 & n3728 ;
  assign n3730 = n3473 & ~n3729 ;
  assign n3731 = ~n1745 & ~n1751 ;
  assign n3732 = ~n3730 & n3731 ;
  assign n3733 = ~n1752 & ~n3732 ;
  assign n3734 = ~n1741 & ~n3490 ;
  assign n3735 = ~n3464 & ~n3466 ;
  assign n3736 = n3734 & n3735 ;
  assign n3737 = n3733 & n3736 ;
  assign n3738 = n3727 & n3737 ;
  assign n3739 = ~n3481 & ~n3486 ;
  assign n3740 = ~n3464 & ~n3739 ;
  assign n3741 = n3734 & n3740 ;
  assign n3742 = n1742 & ~n3490 ;
  assign n3743 = ~n3455 & ~n3742 ;
  assign n3744 = ~n3741 & n3743 ;
  assign n3745 = n3727 & ~n3744 ;
  assign n3746 = ~n1748 & ~n3459 ;
  assign n3747 = ~n3452 & ~n3746 ;
  assign n3748 = n3726 & n3747 ;
  assign n3749 = ~n1761 & n3460 ;
  assign n3750 = ~n1760 & ~n3749 ;
  assign n3751 = ~n3748 & n3750 ;
  assign n3752 = ~n3745 & n3751 ;
  assign n3753 = ~n3738 & n3752 ;
  assign n3754 = ~n1775 & ~n3498 ;
  assign n3755 = ~n1798 & ~n3495 ;
  assign n3756 = n3754 & n3755 ;
  assign n3757 = ~n3501 & ~n3503 ;
  assign n3758 = ~n1763 & ~n3496 ;
  assign n3759 = n3757 & n3758 ;
  assign n3760 = n3756 & n3759 ;
  assign n3761 = ~n3753 & n3760 ;
  assign n3762 = ~n3501 & n3508 ;
  assign n3763 = ~n3512 & ~n3762 ;
  assign n3764 = n3758 & ~n3763 ;
  assign n3765 = ~n1764 & ~n3518 ;
  assign n3766 = ~n3496 & ~n3765 ;
  assign n3767 = ~n3764 & ~n3766 ;
  assign n3768 = n3756 & ~n3767 ;
  assign n3769 = ~n1798 & n3517 ;
  assign n3770 = ~n1797 & ~n3769 ;
  assign n3771 = n3754 & ~n3770 ;
  assign n3772 = ~n1775 & n3522 ;
  assign n3773 = ~n1774 & ~n3772 ;
  assign n3774 = ~n3771 & n3773 ;
  assign n3775 = ~n3768 & n3774 ;
  assign n3776 = ~n3761 & n3775 ;
  assign n3778 = ~n1789 & ~n1791 ;
  assign n3777 = ~n1767 & ~n1770 ;
  assign n3779 = ~n1777 & ~n1784 ;
  assign n3780 = ~n1781 & ~n1794 ;
  assign n3781 = n3779 & n3780 ;
  assign n3782 = n3777 & n3781 ;
  assign n3783 = n3778 & n3782 ;
  assign n3784 = ~n3776 & n3783 ;
  assign n3785 = ~n1777 & n1785 ;
  assign n3786 = ~n1778 & ~n3785 ;
  assign n3787 = n3780 & ~n3786 ;
  assign n3788 = ~n1781 & n1795 ;
  assign n3789 = ~n1782 & ~n3788 ;
  assign n3790 = ~n3787 & n3789 ;
  assign n3791 = n3777 & ~n3790 ;
  assign n3792 = n1768 & ~n1770 ;
  assign n3793 = ~n1771 & ~n3792 ;
  assign n3794 = ~n3791 & n3793 ;
  assign n3795 = n3778 & ~n3794 ;
  assign n3796 = n1788 & ~n1791 ;
  assign n3797 = ~n1792 & ~n3796 ;
  assign n3798 = ~n3795 & n3797 ;
  assign n3799 = ~n3784 & n3798 ;
  assign n3800 = n1780 & ~n3799 ;
  assign n3801 = ~n1780 & n3799 ;
  assign n3802 = ~n3800 & ~n3801 ;
  assign n3803 = n3672 & ~n3802 ;
  assign n3804 = ~n3708 & ~n3803 ;
  assign n3805 = n3557 & ~n3804 ;
  assign n3878 = n1607 & ~n3647 ;
  assign n3879 = ~n1607 & n3647 ;
  assign n3880 = ~n3878 & ~n3879 ;
  assign n3881 = n3672 & n3880 ;
  assign n3882 = ~n3708 & ~n3881 ;
  assign n3883 = n3650 & ~n3882 ;
  assign n3884 = n1607 & n3683 ;
  assign n3885 = n3672 & n3884 ;
  assign n3886 = \P1_reg2_reg[29]/NET0131  & ~n3685 ;
  assign n3887 = n1612 & n1736 ;
  assign n3888 = ~n3886 & ~n3887 ;
  assign n3889 = ~n3885 & n3888 ;
  assign n3890 = ~n3883 & n3889 ;
  assign n3891 = ~n3805 & n3890 ;
  assign n3892 = ~n3877 & n3891 ;
  assign n3893 = ~n3724 & n3892 ;
  assign n3894 = n3662 & ~n3893 ;
  assign n3895 = ~n3707 & ~n3894 ;
  assign n3896 = \P1_state_reg[0]/NET0131  & ~n3895 ;
  assign n3897 = ~n3706 & ~n3896 ;
  assign n3898 = \P1_reg0_reg[29]/NET0131  & ~n3703 ;
  assign n3899 = \P1_reg0_reg[29]/NET0131  & n3664 ;
  assign n3900 = n3445 & n3449 ;
  assign n3901 = \P1_reg0_reg[29]/NET0131  & ~n3900 ;
  assign n3902 = ~n3721 & n3900 ;
  assign n3903 = ~n3901 & ~n3902 ;
  assign n3904 = n1898 & ~n3903 ;
  assign n3908 = ~n3802 & n3900 ;
  assign n3909 = ~n3901 & ~n3908 ;
  assign n3910 = n3557 & ~n3909 ;
  assign n3905 = n3874 & n3900 ;
  assign n3906 = ~n3901 & ~n3905 ;
  assign n3907 = n3575 & ~n3906 ;
  assign n3911 = n3880 & n3900 ;
  assign n3912 = ~n3901 & ~n3911 ;
  assign n3913 = n3650 & ~n3912 ;
  assign n3914 = n3884 & n3900 ;
  assign n3915 = ~n1736 & ~n3615 ;
  assign n3916 = n3683 & ~n3900 ;
  assign n3917 = n3915 & ~n3916 ;
  assign n3918 = \P1_reg0_reg[29]/NET0131  & ~n3917 ;
  assign n3919 = ~n3914 & ~n3918 ;
  assign n3920 = ~n3913 & n3919 ;
  assign n3921 = ~n3907 & n3920 ;
  assign n3922 = ~n3910 & n3921 ;
  assign n3923 = ~n3904 & n3922 ;
  assign n3924 = n3662 & ~n3923 ;
  assign n3925 = ~n3899 & ~n3924 ;
  assign n3926 = \P1_state_reg[0]/NET0131  & ~n3925 ;
  assign n3927 = ~n3898 & ~n3926 ;
  assign n3929 = n2043 & n2050 ;
  assign n3928 = ~n2016 & n3176 ;
  assign n3930 = n3371 & n3928 ;
  assign n3931 = n3929 & n3930 ;
  assign n3932 = ~n1984 & ~n3931 ;
  assign n3933 = \P1_state_reg[0]/NET0131  & ~n3932 ;
  assign n3934 = \P2_B_reg/NET0131  & ~n3933 ;
  assign n3935 = \P1_state_reg[0]/NET0131  & n1984 ;
  assign n3981 = ~n2242 & ~n3275 ;
  assign n3936 = ~\P1_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n3937 = ~n2054 & ~n2056 ;
  assign n3938 = ~n2057 & n3937 ;
  assign n3939 = ~n3936 & n3938 ;
  assign n3940 = n2334 & n3939 ;
  assign n3941 = ~n2492 & n3940 ;
  assign n3945 = ~n2333 & n3939 ;
  assign n3942 = ~n2165 & n3937 ;
  assign n3943 = ~n2053 & ~n3942 ;
  assign n3944 = ~n3936 & ~n3943 ;
  assign n3946 = \P1_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n3947 = ~n3944 & ~n3946 ;
  assign n3948 = ~n3945 & n3947 ;
  assign n3949 = ~n3941 & n3948 ;
  assign n3951 = ~\si[31]_pad  & n3949 ;
  assign n3950 = \si[31]_pad  & ~n3949 ;
  assign n3952 = n542 & ~n3950 ;
  assign n3953 = ~n3951 & n3952 ;
  assign n3954 = \P1_datao_reg[31]/NET0131  & n3953 ;
  assign n3955 = ~\P1_datao_reg[31]/NET0131  & ~n3953 ;
  assign n3956 = ~n3954 & ~n3955 ;
  assign n3957 = ~n2051 & n3956 ;
  assign n3959 = ~n3329 & ~n3957 ;
  assign n3960 = \P1_datao_reg[30]/NET0131  & ~n542 ;
  assign n3961 = ~n3936 & ~n3946 ;
  assign n3963 = ~n2058 & n3938 ;
  assign n3966 = n2392 & n3963 ;
  assign n3967 = ~n2516 & n3966 ;
  assign n3964 = ~n2391 & n3963 ;
  assign n3965 = ~n2247 & n3938 ;
  assign n3962 = ~n2054 & n2163 ;
  assign n3968 = ~n2053 & ~n3962 ;
  assign n3969 = ~n3965 & n3968 ;
  assign n3970 = ~n3964 & n3969 ;
  assign n3971 = ~n3967 & n3970 ;
  assign n3973 = ~n3961 & n3971 ;
  assign n3972 = n3961 & ~n3971 ;
  assign n3974 = n542 & ~n3972 ;
  assign n3975 = ~n3973 & n3974 ;
  assign n3976 = ~n3960 & ~n3975 ;
  assign n3977 = ~n2051 & ~n3976 ;
  assign n4188 = ~n3329 & ~n3363 ;
  assign n4189 = n3977 & ~n4188 ;
  assign n4190 = ~n3959 & ~n4189 ;
  assign n4191 = n3981 & n4190 ;
  assign n3989 = ~n3302 & ~n3308 ;
  assign n3990 = ~n3296 & ~n3303 ;
  assign n4060 = ~n3279 & ~n3990 ;
  assign n4061 = ~n3278 & n4060 ;
  assign n4062 = n3989 & ~n4061 ;
  assign n4063 = ~n3276 & ~n4062 ;
  assign n4049 = ~n3276 & ~n3278 ;
  assign n4050 = ~n3279 & ~n3283 ;
  assign n4070 = n4049 & n4050 ;
  assign n4037 = ~n3282 & ~n3285 ;
  assign n4071 = n3268 & ~n3286 ;
  assign n4072 = ~n3292 & ~n4071 ;
  assign n4073 = n4037 & ~n4072 ;
  assign n4029 = ~n3291 & ~n3297 ;
  assign n4074 = ~n3282 & ~n4029 ;
  assign n4075 = ~n4073 & ~n4074 ;
  assign n4038 = ~n3236 & ~n3286 ;
  assign n4076 = n4037 & n4038 ;
  assign n4042 = ~n3237 & ~n3240 ;
  assign n4032 = ~n3257 & ~n3263 ;
  assign n4077 = ~n3239 & ~n4032 ;
  assign n4078 = n4042 & n4077 ;
  assign n4079 = ~n3264 & ~n3269 ;
  assign n4080 = ~n3237 & ~n4079 ;
  assign n4081 = ~n4078 & ~n4080 ;
  assign n4082 = n4076 & ~n4081 ;
  assign n4083 = n4075 & ~n4082 ;
  assign n4192 = n4070 & ~n4083 ;
  assign n4193 = ~n4063 & ~n4192 ;
  assign n4194 = n4191 & ~n4193 ;
  assign n3993 = ~n3244 & ~n3246 ;
  assign n3994 = ~n3190 & ~n3253 ;
  assign n3995 = ~n3247 & ~n3994 ;
  assign n3996 = n3993 & n3995 ;
  assign n3997 = ~n3252 & ~n3258 ;
  assign n3998 = ~n3244 & ~n3997 ;
  assign n3999 = ~n3996 & ~n3998 ;
  assign n4005 = ~n3182 & ~n3247 ;
  assign n4086 = n3993 & n4005 ;
  assign n4000 = ~n3181 & ~n3184 ;
  assign n4012 = ~n3186 & ~n3226 ;
  assign n4087 = ~n3231 & ~n4012 ;
  assign n4088 = n4000 & n4087 ;
  assign n4011 = ~n3185 & ~n3191 ;
  assign n4089 = ~n3181 & ~n4011 ;
  assign n4090 = ~n4088 & ~n4089 ;
  assign n4091 = n4086 & ~n4090 ;
  assign n4092 = n3999 & ~n4091 ;
  assign n4013 = ~n3196 & ~n3216 ;
  assign n4014 = ~n3205 & ~n3217 ;
  assign n4093 = ~n3200 & ~n3201 ;
  assign n4094 = n3208 & ~n4093 ;
  assign n4095 = n3202 & ~n3206 ;
  assign n4096 = ~n3212 & ~n4095 ;
  assign n4097 = ~n4094 & n4096 ;
  assign n4098 = n4014 & ~n4097 ;
  assign n4099 = n3211 & ~n3217 ;
  assign n4100 = ~n3221 & ~n4099 ;
  assign n4101 = ~n4098 & n4100 ;
  assign n4102 = n4013 & ~n4101 ;
  assign n4103 = ~n3220 & ~n3227 ;
  assign n4104 = ~n3196 & ~n4103 ;
  assign n4105 = ~n4102 & ~n4104 ;
  assign n4198 = n4092 & n4105 ;
  assign n4001 = ~n3195 & ~n3231 ;
  assign n4002 = n3187 & ~n4001 ;
  assign n4003 = n4000 & ~n4002 ;
  assign n4004 = ~n3191 & ~n4003 ;
  assign n4006 = n3254 & ~n4005 ;
  assign n4007 = n3993 & ~n4006 ;
  assign n4008 = ~n3258 & ~n4007 ;
  assign n4009 = ~n4004 & ~n4008 ;
  assign n4010 = n3999 & ~n4009 ;
  assign n4043 = ~n3239 & ~n3243 ;
  assign n4084 = n4042 & n4043 ;
  assign n4200 = ~n4010 & n4084 ;
  assign n4201 = ~n4198 & n4200 ;
  assign n4199 = n4070 & n4076 ;
  assign n4202 = n4191 & n4199 ;
  assign n4203 = n4201 & n4202 ;
  assign n3986 = ~n2243 & ~n3307 ;
  assign n4066 = ~n2242 & ~n3986 ;
  assign n4195 = n4066 & n4190 ;
  assign n3980 = ~n3363 & ~n3977 ;
  assign n4196 = ~n3329 & ~n3980 ;
  assign n4197 = n3957 & ~n4196 ;
  assign n4204 = ~n4195 & ~n4197 ;
  assign n4205 = ~n4203 & n4204 ;
  assign n4206 = ~n4194 & n4205 ;
  assign n4207 = n2592 & ~n4206 ;
  assign n4208 = ~n2592 & n4206 ;
  assign n4209 = ~n4207 & ~n4208 ;
  assign n4223 = n3168 & ~n3173 ;
  assign n4224 = ~n4209 & n4223 ;
  assign n3958 = n3329 & n3957 ;
  assign n3978 = n3363 & n3977 ;
  assign n3979 = ~n3959 & ~n3978 ;
  assign n3982 = ~n2243 & ~n3980 ;
  assign n3983 = ~n3981 & n3982 ;
  assign n3984 = n3979 & ~n3983 ;
  assign n3985 = ~n3958 & ~n3984 ;
  assign n3987 = ~n3958 & ~n3980 ;
  assign n3988 = n3986 & n3987 ;
  assign n3991 = n3989 & n3990 ;
  assign n3992 = n3988 & n3991 ;
  assign n4015 = ~n2823 & n2830 ;
  assign n4016 = ~n3199 & n4015 ;
  assign n4017 = n3203 & ~n4016 ;
  assign n4018 = n3208 & ~n4017 ;
  assign n4019 = n3213 & ~n4018 ;
  assign n4020 = n4014 & ~n4019 ;
  assign n4021 = n3222 & ~n4020 ;
  assign n4022 = n4013 & ~n4021 ;
  assign n4023 = ~n3227 & n4012 ;
  assign n4024 = n4011 & n4023 ;
  assign n4025 = n3994 & n4024 ;
  assign n4026 = n3997 & n4025 ;
  assign n4027 = ~n4022 & n4026 ;
  assign n4028 = ~n4010 & ~n4027 ;
  assign n4030 = n3270 & ~n3292 ;
  assign n4031 = n4029 & n4030 ;
  assign n4033 = ~n3264 & n4032 ;
  assign n4034 = n4031 & n4033 ;
  assign n4035 = ~n4028 & n4034 ;
  assign n4036 = n3992 & n4035 ;
  assign n4055 = ~n3985 & ~n4036 ;
  assign n4039 = n3293 & ~n4038 ;
  assign n4040 = n4037 & ~n4039 ;
  assign n4041 = ~n3297 & ~n4040 ;
  assign n4044 = n3265 & ~n4043 ;
  assign n4045 = n4042 & ~n4044 ;
  assign n4046 = n4031 & ~n4045 ;
  assign n4047 = ~n4041 & ~n4046 ;
  assign n4048 = n3992 & ~n4047 ;
  assign n4051 = n3304 & ~n4050 ;
  assign n4052 = n4049 & ~n4051 ;
  assign n4053 = ~n3308 & n3988 ;
  assign n4054 = ~n4052 & n4053 ;
  assign n4056 = ~n4048 & ~n4054 ;
  assign n4057 = n4055 & n4056 ;
  assign n4214 = ~n2592 & n4057 ;
  assign n4213 = n2592 & ~n4057 ;
  assign n4215 = ~n3161 & n3167 ;
  assign n4216 = ~n3173 & n4215 ;
  assign n4217 = ~n4213 & n4216 ;
  assign n4218 = ~n4214 & n4217 ;
  assign n4085 = n4076 & n4084 ;
  assign n4106 = n4001 & ~n4105 ;
  assign n4107 = n4000 & n4106 ;
  assign n4108 = n4086 & n4107 ;
  assign n4109 = n4092 & ~n4108 ;
  assign n4110 = n4085 & ~n4109 ;
  assign n4111 = n4083 & ~n4110 ;
  assign n4064 = n3979 & n3981 ;
  assign n4112 = n4064 & n4070 ;
  assign n4113 = ~n4111 & n4112 ;
  assign n4065 = n4063 & n4064 ;
  assign n4067 = ~n3978 & n4066 ;
  assign n4068 = n3987 & ~n4067 ;
  assign n4069 = ~n3959 & ~n4068 ;
  assign n4114 = ~n4065 & ~n4069 ;
  assign n4115 = ~n4113 & n4114 ;
  assign n4219 = ~\P2_B_reg/NET0131  & n4115 ;
  assign n4220 = ~n3161 & ~n3167 ;
  assign n4221 = n3174 & n4220 ;
  assign n4222 = ~n4219 & n4221 ;
  assign n4227 = ~n4218 & ~n4222 ;
  assign n4228 = ~n4224 & n4227 ;
  assign n4210 = ~\P2_B_reg/NET0131  & n4209 ;
  assign n4211 = n3161 & n3176 ;
  assign n4212 = ~n4210 & n4211 ;
  assign n4058 = ~\P2_B_reg/NET0131  & ~n4057 ;
  assign n4059 = n3176 & ~n4058 ;
  assign n4116 = n3177 & ~n4115 ;
  assign n4117 = ~n4059 & ~n4116 ;
  assign n4118 = n3414 & ~n4117 ;
  assign n4128 = ~n2981 & ~n3010 ;
  assign n4127 = ~n3006 & ~n3011 ;
  assign n4130 = ~n2746 & ~n2891 ;
  assign n4133 = ~n3206 & ~n3212 ;
  assign n4147 = ~n4130 & n4133 ;
  assign n4134 = ~n3202 & ~n3207 ;
  assign n4141 = ~n3205 & ~n3211 ;
  assign n4148 = n4134 & n4141 ;
  assign n4149 = n4147 & n4148 ;
  assign n4153 = ~n4127 & n4149 ;
  assign n4154 = ~n4128 & n4153 ;
  assign n4157 = n3248 & n4154 ;
  assign n4131 = ~n3047 & ~n3129 ;
  assign n4158 = n3254 & ~n4131 ;
  assign n4159 = n4157 & n4158 ;
  assign n4120 = ~n3072 & ~n3130 ;
  assign n4142 = ~n2955 & ~n3015 ;
  assign n4139 = ~n2927 & ~n3016 ;
  assign n4121 = ~n2720 & ~n2897 ;
  assign n4129 = ~n3217 & ~n3221 ;
  assign n4146 = ~n4015 & n4129 ;
  assign n4150 = ~n4121 & n4146 ;
  assign n4123 = ~n2693 & ~n2896 ;
  assign n4124 = ~n3199 & ~n3201 ;
  assign n4125 = ~n3198 & n4124 ;
  assign n4151 = ~n4123 & n4125 ;
  assign n4152 = n4150 & n4151 ;
  assign n4155 = ~n4139 & n4152 ;
  assign n4156 = ~n4142 & n4155 ;
  assign n4160 = ~n4120 & n4156 ;
  assign n4164 = n4159 & n4160 ;
  assign n4126 = ~n2614 & ~n3141 ;
  assign n4144 = ~n2508 & ~n2557 ;
  assign n4165 = ~n4126 & ~n4144 ;
  assign n4166 = n4164 & n4165 ;
  assign n4122 = ~n2532 & ~n2533 ;
  assign n4132 = ~n2641 & ~n3136 ;
  assign n4138 = ~n2552 & ~n3147 ;
  assign n4161 = ~n4132 & ~n4138 ;
  assign n4140 = ~n2589 & ~n3140 ;
  assign n4145 = ~n2667 & ~n3135 ;
  assign n4162 = ~n4140 & ~n4145 ;
  assign n4163 = n4161 & n4162 ;
  assign n4167 = ~n4122 & n4163 ;
  assign n4170 = n4166 & n4167 ;
  assign n4135 = ~n2434 & ~n2563 ;
  assign n4171 = n2244 & ~n4135 ;
  assign n4172 = n4170 & n4171 ;
  assign n4143 = ~n2386 & ~n2562 ;
  assign n4136 = ~n2485 & ~n2556 ;
  assign n4137 = ~n2462 & ~n2564 ;
  assign n4168 = ~n4136 & ~n4137 ;
  assign n4169 = ~n4143 & n4168 ;
  assign n4173 = n3979 & n4169 ;
  assign n4119 = ~n2329 & ~n2567 ;
  assign n4174 = n3987 & ~n4119 ;
  assign n4175 = n4173 & n4174 ;
  assign n4176 = n4172 & n4175 ;
  assign n4177 = n2592 & ~n4176 ;
  assign n4178 = ~n2592 & n4176 ;
  assign n4179 = ~n4177 & ~n4178 ;
  assign n4180 = n3161 & ~n4179 ;
  assign n4181 = \P2_B_reg/NET0131  & n3173 ;
  assign n4182 = ~n3414 & n4181 ;
  assign n4183 = ~n4180 & ~n4182 ;
  assign n4184 = ~n3167 & ~n4183 ;
  assign n4185 = n3408 & n4115 ;
  assign n4186 = ~\P2_B_reg/NET0131  & n4057 ;
  assign n4187 = n3373 & ~n4186 ;
  assign n4225 = ~n4185 & ~n4187 ;
  assign n4226 = ~n4184 & n4225 ;
  assign n4229 = ~n4118 & n4226 ;
  assign n4230 = ~n4212 & n4229 ;
  assign n4231 = n4228 & n4230 ;
  assign n4232 = n3935 & ~n4231 ;
  assign n4233 = ~n3934 & ~n4232 ;
  assign n4234 = \P1_reg1_reg[29]/NET0131  & ~n3703 ;
  assign n4235 = \P1_reg1_reg[29]/NET0131  & n3664 ;
  assign n4236 = ~n3445 & n3449 ;
  assign n4237 = \P1_reg1_reg[29]/NET0131  & ~n4236 ;
  assign n4238 = ~n3721 & n4236 ;
  assign n4239 = ~n4237 & ~n4238 ;
  assign n4240 = n1898 & ~n4239 ;
  assign n4244 = n3874 & n4236 ;
  assign n4245 = ~n4237 & ~n4244 ;
  assign n4246 = n3575 & ~n4245 ;
  assign n4241 = ~n3802 & n4236 ;
  assign n4242 = ~n4237 & ~n4241 ;
  assign n4243 = n3557 & ~n4242 ;
  assign n4247 = n3880 & n4236 ;
  assign n4248 = ~n4237 & ~n4247 ;
  assign n4249 = n3650 & ~n4248 ;
  assign n4250 = n3884 & n4236 ;
  assign n4251 = n3683 & ~n4236 ;
  assign n4252 = n3915 & ~n4251 ;
  assign n4253 = \P1_reg1_reg[29]/NET0131  & ~n4252 ;
  assign n4254 = ~n4250 & ~n4253 ;
  assign n4255 = ~n4249 & n4254 ;
  assign n4256 = ~n4243 & n4255 ;
  assign n4257 = ~n4246 & n4256 ;
  assign n4258 = ~n4240 & n4257 ;
  assign n4259 = n3662 & ~n4258 ;
  assign n4260 = ~n4235 & ~n4259 ;
  assign n4261 = \P1_state_reg[0]/NET0131  & ~n4260 ;
  assign n4262 = ~n4234 & ~n4261 ;
  assign n4266 = n3406 & ~n3977 ;
  assign n4268 = ~n3957 & n4266 ;
  assign n4267 = n3957 & ~n4266 ;
  assign n4269 = n3409 & ~n4267 ;
  assign n4270 = ~n4268 & n4269 ;
  assign n4263 = n3375 & n3957 ;
  assign n4264 = ~n3329 & n3373 ;
  assign n4265 = n3368 & n4264 ;
  assign n4271 = ~n4263 & ~n4265 ;
  assign n4272 = ~n4270 & n4271 ;
  assign n4273 = n2033 & ~n4272 ;
  assign n4274 = ~n3416 & ~n4273 ;
  assign n4275 = \P1_state_reg[0]/NET0131  & n2017 ;
  assign n4276 = ~n4274 & n4275 ;
  assign n4277 = ~n3415 & ~n3419 ;
  assign n4278 = n4275 & ~n4277 ;
  assign n4279 = \P2_reg2_reg[31]/NET0131  & ~n4278 ;
  assign n4280 = ~n4276 & ~n4279 ;
  assign n4283 = n1563 & n3664 ;
  assign n4284 = n1563 & ~n3450 ;
  assign n4307 = n3493 & n3506 ;
  assign n4308 = ~n3463 & n3505 ;
  assign n4309 = n3515 & ~n4308 ;
  assign n4310 = n3500 & ~n4309 ;
  assign n4311 = n3525 & ~n4310 ;
  assign n4312 = ~n4307 & n4311 ;
  assign n4313 = n3533 & ~n4312 ;
  assign n4314 = n3545 & ~n4313 ;
  assign n4315 = n1783 & n4314 ;
  assign n4316 = ~n1783 & ~n4314 ;
  assign n4317 = ~n4315 & ~n4316 ;
  assign n4318 = n3450 & ~n4317 ;
  assign n4319 = ~n4284 & ~n4318 ;
  assign n4320 = n3557 & ~n4319 ;
  assign n4285 = n3597 & n3711 ;
  assign n4286 = ~n1570 & n4285 ;
  assign n4287 = n1542 & ~n4286 ;
  assign n4288 = n3599 & n3711 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4290 = ~n536 & ~n4289 ;
  assign n4291 = n536 & n921 ;
  assign n4292 = ~n4290 & ~n4291 ;
  assign n4293 = n3450 & n4292 ;
  assign n4294 = ~n4284 & ~n4293 ;
  assign n4295 = n1898 & ~n4294 ;
  assign n4322 = ~n1213 & n1429 ;
  assign n4323 = n847 & ~n4322 ;
  assign n4324 = n1426 & ~n4323 ;
  assign n4321 = n1424 & n1430 ;
  assign n4325 = n982 & ~n4321 ;
  assign n4326 = ~n4324 & n4325 ;
  assign n4327 = n1783 & ~n4326 ;
  assign n4328 = ~n1783 & n4326 ;
  assign n4329 = ~n4327 & ~n4328 ;
  assign n4330 = n3450 & ~n4329 ;
  assign n4331 = ~n4284 & ~n4330 ;
  assign n4332 = n3575 & ~n4331 ;
  assign n4297 = n3641 & n3642 ;
  assign n4298 = n910 & n3641 ;
  assign n4299 = n1561 & ~n4298 ;
  assign n4300 = ~n4297 & ~n4299 ;
  assign n4301 = n3450 & n4300 ;
  assign n4302 = ~n4284 & ~n4301 ;
  assign n4303 = n3650 & ~n4302 ;
  assign n4296 = n1561 & n3655 ;
  assign n4304 = ~n3450 & n3683 ;
  assign n4305 = ~n3615 & ~n4304 ;
  assign n4306 = n1563 & ~n4305 ;
  assign n4333 = ~n4296 & ~n4306 ;
  assign n4334 = ~n4303 & n4333 ;
  assign n4335 = ~n4332 & n4334 ;
  assign n4336 = ~n4295 & n4335 ;
  assign n4337 = ~n4320 & n4336 ;
  assign n4338 = n3662 & ~n4337 ;
  assign n4339 = ~n4283 & ~n4338 ;
  assign n4340 = \P1_state_reg[0]/NET0131  & ~n4339 ;
  assign n4281 = \P1_reg3_reg[24]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4282 = n1563 & n1934 ;
  assign n4341 = ~n4281 & ~n4282 ;
  assign n4342 = ~n4340 & n4341 ;
  assign n4343 = \P2_reg2_reg[27]/NET0131  & ~n2033 ;
  assign n4344 = n3280 & n3284 ;
  assign n4345 = n3197 & n3232 ;
  assign n4346 = ~n3224 & n4345 ;
  assign n4347 = n3229 & n3232 ;
  assign n4348 = ~n3188 & ~n4347 ;
  assign n4349 = ~n4346 & n4348 ;
  assign n4350 = n3183 & n3248 ;
  assign n4351 = ~n4349 & n4350 ;
  assign n4352 = ~n3193 & n3248 ;
  assign n4353 = ~n3255 & ~n4352 ;
  assign n4354 = ~n4351 & n4353 ;
  assign n4355 = n3241 & n3245 ;
  assign n4356 = ~n4354 & n4355 ;
  assign n4357 = n3241 & ~n3260 ;
  assign n4358 = ~n3266 & ~n4357 ;
  assign n4359 = ~n4356 & n4358 ;
  assign n4360 = n3238 & n3287 ;
  assign n4361 = ~n4359 & n4360 ;
  assign n4362 = n4344 & n4361 ;
  assign n4364 = n3271 & n3287 ;
  assign n4365 = ~n3294 & ~n4364 ;
  assign n4366 = n4344 & ~n4365 ;
  assign n4363 = n3280 & ~n3299 ;
  assign n4367 = ~n3305 & ~n4363 ;
  assign n4368 = ~n4366 & n4367 ;
  assign n4369 = ~n4362 & n4368 ;
  assign n4370 = n4143 & ~n4369 ;
  assign n4371 = ~n4143 & n4369 ;
  assign n4372 = ~n4370 & ~n4371 ;
  assign n4373 = n2033 & ~n4372 ;
  assign n4374 = ~n4343 & ~n4373 ;
  assign n4375 = n3319 & ~n4374 ;
  assign n4376 = ~n3143 & n3148 ;
  assign n4377 = n2554 & ~n4376 ;
  assign n4378 = ~n2462 & ~n2485 ;
  assign n4379 = ~n2508 & n4378 ;
  assign n4380 = ~n4377 & n4379 ;
  assign n4381 = ~n2462 & ~n2559 ;
  assign n4382 = n2565 & ~n4381 ;
  assign n4383 = ~n4380 & n4382 ;
  assign n4384 = ~n2434 & ~n4383 ;
  assign n4385 = n2770 & ~n2888 ;
  assign n4386 = n2894 & ~n4385 ;
  assign n4387 = n2721 & n3007 ;
  assign n4388 = ~n4386 & n4387 ;
  assign n4389 = n2899 & n3007 ;
  assign n4390 = n3013 & ~n4389 ;
  assign n4391 = ~n4388 & n4390 ;
  assign n4392 = n2668 & n3073 ;
  assign n4393 = n2956 & n3120 ;
  assign n4394 = n4392 & n4393 ;
  assign n4395 = ~n4391 & n4394 ;
  assign n4396 = n3018 & n3120 ;
  assign n4397 = ~n3127 & ~n4396 ;
  assign n4398 = n4392 & ~n4397 ;
  assign n4399 = n2668 & ~n3132 ;
  assign n4400 = ~n3138 & ~n4399 ;
  assign n4401 = ~n4398 & n4400 ;
  assign n4402 = ~n4395 & n4401 ;
  assign n4403 = n2615 & n3148 ;
  assign n4404 = ~n2434 & n4379 ;
  assign n4405 = n4403 & n4404 ;
  assign n4406 = ~n4402 & n4405 ;
  assign n4407 = ~n4384 & ~n4406 ;
  assign n4408 = n4143 & n4407 ;
  assign n4409 = ~n4143 & ~n4407 ;
  assign n4410 = ~n4408 & ~n4409 ;
  assign n4411 = n2033 & ~n4410 ;
  assign n4412 = ~n4343 & ~n4411 ;
  assign n4413 = n3179 & ~n4412 ;
  assign n4414 = n2050 & ~n2433 ;
  assign n4415 = ~n2433 & n3355 ;
  assign n4416 = ~n2385 & n4415 ;
  assign n4417 = n2328 & ~n4416 ;
  assign n4418 = n3323 & n3355 ;
  assign n4419 = ~n2050 & ~n4418 ;
  assign n4420 = ~n4417 & n4419 ;
  assign n4421 = ~n4414 & ~n4420 ;
  assign n4422 = n3373 & ~n4421 ;
  assign n4423 = n2376 & n3375 ;
  assign n4424 = n3396 & n3400 ;
  assign n4425 = ~n2424 & n4424 ;
  assign n4426 = n2376 & ~n4425 ;
  assign n4427 = ~n3403 & ~n4426 ;
  assign n4428 = n3409 & n4427 ;
  assign n4429 = ~n4423 & ~n4428 ;
  assign n4430 = ~n4422 & n4429 ;
  assign n4431 = n2033 & ~n4430 ;
  assign n4432 = n2381 & n3415 ;
  assign n4433 = ~n3375 & ~n3418 ;
  assign n4434 = ~n3419 & ~n4433 ;
  assign n4435 = ~n2033 & n3409 ;
  assign n4436 = ~n4434 & ~n4435 ;
  assign n4437 = ~n3417 & n4436 ;
  assign n4438 = \P2_reg2_reg[27]/NET0131  & ~n4437 ;
  assign n4439 = ~n4432 & ~n4438 ;
  assign n4440 = ~n4431 & n4439 ;
  assign n4441 = ~n4413 & n4440 ;
  assign n4442 = ~n4375 & n4441 ;
  assign n4443 = n2017 & ~n4442 ;
  assign n4444 = \P2_reg2_reg[27]/NET0131  & n3430 ;
  assign n4445 = ~n4443 & ~n4444 ;
  assign n4446 = \P1_state_reg[0]/NET0131  & ~n4445 ;
  assign n4447 = \P2_reg2_reg[27]/NET0131  & ~n3434 ;
  assign n4448 = ~n4446 & ~n4447 ;
  assign n4449 = \P1_reg2_reg[26]/NET0131  & ~n3703 ;
  assign n4450 = \P1_reg2_reg[26]/NET0131  & n3664 ;
  assign n4451 = \P1_reg2_reg[26]/NET0131  & ~n3672 ;
  assign n4452 = n1102 & n1428 ;
  assign n4453 = ~n841 & ~n4452 ;
  assign n4454 = ~n1407 & n1412 ;
  assign n4455 = n1265 & n1421 ;
  assign n4456 = ~n4454 & n4455 ;
  assign n4457 = n1417 & n1421 ;
  assign n4458 = ~n1205 & ~n4457 ;
  assign n4459 = ~n4456 & n4458 ;
  assign n4460 = n1105 & n1153 ;
  assign n4461 = ~n4459 & n4460 ;
  assign n4462 = n1105 & n1210 ;
  assign n4463 = ~n1097 & ~n4462 ;
  assign n4464 = ~n4461 & n4463 ;
  assign n4465 = n1042 & n1428 ;
  assign n4466 = ~n4464 & n4465 ;
  assign n4467 = n4453 & ~n4466 ;
  assign n4468 = n923 & n1572 ;
  assign n4469 = n754 & n985 ;
  assign n4470 = n4468 & n4469 ;
  assign n4471 = ~n4467 & n4470 ;
  assign n4473 = n846 & n985 ;
  assign n4474 = ~n976 & ~n4473 ;
  assign n4475 = n4468 & ~n4474 ;
  assign n4472 = n981 & n1572 ;
  assign n4476 = n1580 & ~n4472 ;
  assign n4477 = ~n4475 & n4476 ;
  assign n4478 = ~n4471 & n4477 ;
  assign n4479 = n1772 & ~n4478 ;
  assign n4480 = ~n1772 & n4478 ;
  assign n4481 = ~n4479 & ~n4480 ;
  assign n4482 = n3672 & ~n4481 ;
  assign n4483 = ~n4451 & ~n4482 ;
  assign n4484 = n3575 & ~n4483 ;
  assign n4519 = n536 & ~n1542 ;
  assign n4520 = ~n1478 & n4288 ;
  assign n4521 = n1510 & ~n4520 ;
  assign n4522 = ~n536 & ~n3712 ;
  assign n4523 = ~n4521 & n4522 ;
  assign n4524 = ~n4519 & ~n4523 ;
  assign n4525 = n3672 & ~n4524 ;
  assign n4526 = ~n4451 & ~n4525 ;
  assign n4527 = n1898 & ~n4526 ;
  assign n4485 = n3529 & n3531 ;
  assign n4486 = ~n3524 & n3532 ;
  assign n4487 = n3541 & ~n4486 ;
  assign n4488 = n3499 & n3532 ;
  assign n4489 = n3497 & n3502 ;
  assign n4490 = n3462 & n3504 ;
  assign n4491 = ~n3510 & ~n4490 ;
  assign n4492 = n4489 & ~n4491 ;
  assign n4493 = n3497 & ~n3514 ;
  assign n4494 = n3520 & ~n4493 ;
  assign n4495 = ~n4492 & n4494 ;
  assign n4496 = n4488 & ~n4495 ;
  assign n4497 = n4487 & ~n4496 ;
  assign n4498 = n4485 & ~n4497 ;
  assign n4500 = n3465 & n3491 ;
  assign n4501 = ~n3484 & n4500 ;
  assign n4502 = ~n3488 & n3491 ;
  assign n4503 = n3457 & ~n4502 ;
  assign n4504 = ~n4501 & n4503 ;
  assign n4505 = n3454 & n3504 ;
  assign n4506 = ~n4504 & n4505 ;
  assign n4507 = n4485 & n4488 ;
  assign n4508 = n4489 & n4507 ;
  assign n4509 = n4506 & n4508 ;
  assign n4499 = n3529 & ~n3544 ;
  assign n4510 = n3537 & ~n4499 ;
  assign n4511 = ~n4509 & n4510 ;
  assign n4512 = ~n4498 & n4511 ;
  assign n4513 = n1772 & n4512 ;
  assign n4514 = ~n1772 & ~n4512 ;
  assign n4515 = ~n4513 & ~n4514 ;
  assign n4516 = n3672 & ~n4515 ;
  assign n4517 = ~n4451 & ~n4516 ;
  assign n4518 = n3557 & ~n4517 ;
  assign n4528 = ~n1533 & n4297 ;
  assign n4529 = n1463 & ~n4528 ;
  assign n4530 = ~n1463 & n4528 ;
  assign n4531 = ~n4529 & ~n4530 ;
  assign n4532 = n3672 & n4531 ;
  assign n4533 = ~n4451 & ~n4532 ;
  assign n4534 = n3650 & ~n4533 ;
  assign n4537 = n1463 & n3683 ;
  assign n4538 = n3672 & n4537 ;
  assign n4535 = \P1_reg2_reg[26]/NET0131  & ~n3685 ;
  assign n4536 = n1474 & n1736 ;
  assign n4539 = ~n4535 & ~n4536 ;
  assign n4540 = ~n4538 & n4539 ;
  assign n4541 = ~n4534 & n4540 ;
  assign n4542 = ~n4518 & n4541 ;
  assign n4543 = ~n4527 & n4542 ;
  assign n4544 = ~n4484 & n4543 ;
  assign n4545 = n3662 & ~n4544 ;
  assign n4546 = ~n4450 & ~n4545 ;
  assign n4547 = \P1_state_reg[0]/NET0131  & ~n4546 ;
  assign n4548 = ~n4449 & ~n4547 ;
  assign n4549 = n1538 & n3664 ;
  assign n4550 = n1538 & ~n3450 ;
  assign n4552 = ~n3737 & n3744 ;
  assign n4553 = n3727 & n3759 ;
  assign n4554 = ~n4552 & n4553 ;
  assign n4551 = ~n3751 & n3759 ;
  assign n4555 = n3767 & ~n4551 ;
  assign n4556 = ~n4554 & n4555 ;
  assign n4557 = n3756 & ~n4556 ;
  assign n4558 = n3774 & ~n4557 ;
  assign n4559 = n3781 & ~n4558 ;
  assign n4560 = n3790 & ~n4559 ;
  assign n4561 = n1769 & n4560 ;
  assign n4562 = ~n1769 & ~n4560 ;
  assign n4563 = ~n4561 & ~n4562 ;
  assign n4564 = n3450 & ~n4563 ;
  assign n4565 = ~n4550 & ~n4564 ;
  assign n4566 = n3557 & ~n4565 ;
  assign n4567 = n1478 & ~n4288 ;
  assign n4568 = ~n4520 & ~n4567 ;
  assign n4569 = ~n536 & ~n4568 ;
  assign n4570 = n536 & n1570 ;
  assign n4571 = ~n4569 & ~n4570 ;
  assign n4572 = n3450 & n4571 ;
  assign n4573 = ~n4550 & ~n4572 ;
  assign n4574 = n1898 & ~n4573 ;
  assign n4577 = n3811 & ~n3818 ;
  assign n4578 = n3843 & ~n4577 ;
  assign n4579 = n3808 & ~n4578 ;
  assign n4580 = n3849 & ~n4579 ;
  assign n4581 = n3854 & ~n4580 ;
  assign n4575 = n3812 & n3854 ;
  assign n4576 = n3836 & n4575 ;
  assign n4582 = n3864 & ~n4576 ;
  assign n4583 = ~n4581 & n4582 ;
  assign n4584 = n1769 & ~n4583 ;
  assign n4585 = ~n1769 & n4583 ;
  assign n4586 = ~n4584 & ~n4585 ;
  assign n4587 = n3450 & ~n4586 ;
  assign n4588 = ~n4550 & ~n4587 ;
  assign n4589 = n3575 & ~n4588 ;
  assign n4593 = n1533 & ~n4297 ;
  assign n4594 = ~n4528 & ~n4593 ;
  assign n4595 = n3650 & n4594 ;
  assign n4596 = n3450 & n4595 ;
  assign n4590 = ~n3450 & n3650 ;
  assign n4591 = n4305 & ~n4590 ;
  assign n4592 = n1538 & ~n4591 ;
  assign n4597 = n1533 & n3655 ;
  assign n4598 = ~n4592 & ~n4597 ;
  assign n4599 = ~n4596 & n4598 ;
  assign n4600 = ~n4589 & n4599 ;
  assign n4601 = ~n4574 & n4600 ;
  assign n4602 = ~n4566 & n4601 ;
  assign n4603 = n3662 & ~n4602 ;
  assign n4604 = ~n4549 & ~n4603 ;
  assign n4605 = \P1_state_reg[0]/NET0131  & ~n4604 ;
  assign n4606 = \P1_reg3_reg[25]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4607 = n1538 & n1934 ;
  assign n4608 = ~n4606 & ~n4607 ;
  assign n4609 = ~n4605 & n4608 ;
  assign n4610 = n2027 & n2032 ;
  assign n4611 = \P2_reg0_reg[29]/NET0131  & ~n4610 ;
  assign n4612 = ~n3156 & n4610 ;
  assign n4613 = ~n4611 & ~n4612 ;
  assign n4614 = n3179 & ~n4613 ;
  assign n4615 = n3316 & n4610 ;
  assign n4616 = ~n4611 & ~n4615 ;
  assign n4617 = n3319 & ~n4616 ;
  assign n4618 = ~n3412 & n4610 ;
  assign n4619 = ~n3415 & ~n3418 ;
  assign n4620 = n3420 & ~n4610 ;
  assign n4621 = n4619 & ~n4620 ;
  assign n4622 = n3373 & ~n4610 ;
  assign n4623 = n4621 & ~n4622 ;
  assign n4624 = \P2_reg0_reg[29]/NET0131  & ~n4623 ;
  assign n4625 = ~n4618 & ~n4624 ;
  assign n4626 = ~n4617 & n4625 ;
  assign n4627 = ~n4614 & n4626 ;
  assign n4628 = n2017 & ~n4627 ;
  assign n4629 = \P2_reg0_reg[29]/NET0131  & n3430 ;
  assign n4630 = ~n4628 & ~n4629 ;
  assign n4631 = \P1_state_reg[0]/NET0131  & ~n4630 ;
  assign n4632 = \P2_reg0_reg[29]/NET0131  & ~n3434 ;
  assign n4633 = ~n4631 & ~n4632 ;
  assign n4634 = \P1_reg2_reg[24]/NET0131  & ~n3703 ;
  assign n4635 = \P1_reg2_reg[24]/NET0131  & n3664 ;
  assign n4636 = \P1_reg2_reg[24]/NET0131  & ~n3672 ;
  assign n4647 = n3672 & ~n4317 ;
  assign n4648 = ~n4636 & ~n4647 ;
  assign n4649 = n3557 & ~n4648 ;
  assign n4637 = n3672 & n4292 ;
  assign n4638 = ~n4636 & ~n4637 ;
  assign n4639 = n1898 & ~n4638 ;
  assign n4650 = n3672 & ~n4329 ;
  assign n4651 = ~n4636 & ~n4650 ;
  assign n4652 = n3575 & ~n4651 ;
  assign n4641 = n3672 & n4300 ;
  assign n4642 = ~n4636 & ~n4641 ;
  assign n4643 = n3650 & ~n4642 ;
  assign n4645 = n1561 & n3683 ;
  assign n4646 = n3672 & n4645 ;
  assign n4640 = \P1_reg2_reg[24]/NET0131  & ~n3685 ;
  assign n4644 = n1563 & n1736 ;
  assign n4653 = ~n4640 & ~n4644 ;
  assign n4654 = ~n4646 & n4653 ;
  assign n4655 = ~n4643 & n4654 ;
  assign n4656 = ~n4652 & n4655 ;
  assign n4657 = ~n4639 & n4656 ;
  assign n4658 = ~n4649 & n4657 ;
  assign n4659 = n3662 & ~n4658 ;
  assign n4660 = ~n4635 & ~n4659 ;
  assign n4661 = \P1_state_reg[0]/NET0131  & ~n4660 ;
  assign n4662 = ~n4634 & ~n4661 ;
  assign n4663 = ~n2027 & n2032 ;
  assign n4664 = \P2_reg1_reg[29]/NET0131  & ~n4663 ;
  assign n4665 = ~n3156 & n4663 ;
  assign n4666 = ~n4664 & ~n4665 ;
  assign n4667 = n3179 & ~n4666 ;
  assign n4668 = n3316 & n4663 ;
  assign n4669 = ~n4664 & ~n4668 ;
  assign n4670 = n3319 & ~n4669 ;
  assign n4671 = ~n3370 & n4663 ;
  assign n4672 = ~n4664 & ~n4671 ;
  assign n4673 = n3373 & ~n4672 ;
  assign n4674 = n3407 & n4663 ;
  assign n4675 = ~n4664 & ~n4674 ;
  assign n4676 = n3409 & ~n4675 ;
  assign n4677 = \P2_reg1_reg[29]/NET0131  & ~n4619 ;
  assign n4678 = n2191 & n4663 ;
  assign n4679 = ~n4664 & ~n4678 ;
  assign n4680 = n3375 & ~n4679 ;
  assign n4681 = ~n4677 & ~n4680 ;
  assign n4682 = ~n4676 & n4681 ;
  assign n4683 = ~n4673 & n4682 ;
  assign n4684 = ~n4670 & n4683 ;
  assign n4685 = ~n4667 & n4684 ;
  assign n4686 = n2017 & ~n4685 ;
  assign n4687 = \P2_reg1_reg[29]/NET0131  & n3430 ;
  assign n4688 = ~n4686 & ~n4687 ;
  assign n4689 = \P1_state_reg[0]/NET0131  & ~n4688 ;
  assign n4690 = \P2_reg1_reg[29]/NET0131  & ~n3434 ;
  assign n4691 = ~n4689 & ~n4690 ;
  assign n4692 = \P1_reg0_reg[28]/NET0131  & ~n3703 ;
  assign n4693 = \P1_reg0_reg[28]/NET0131  & ~n3900 ;
  assign n4694 = ~n3552 & n3900 ;
  assign n4695 = ~n4693 & ~n4694 ;
  assign n4696 = n3557 & ~n4695 ;
  assign n4697 = ~n3572 & n3900 ;
  assign n4698 = ~n4693 & ~n4697 ;
  assign n4699 = n3575 & ~n4698 ;
  assign n4700 = n1898 & ~n3611 ;
  assign n4701 = ~n3651 & ~n3691 ;
  assign n4702 = ~n4700 & n4701 ;
  assign n4703 = n3900 & ~n4702 ;
  assign n4704 = n1731 & ~n3556 ;
  assign n4705 = ~n3900 & n4704 ;
  assign n4706 = n3917 & ~n4705 ;
  assign n4707 = \P1_reg0_reg[28]/NET0131  & ~n4706 ;
  assign n4708 = ~n4703 & ~n4707 ;
  assign n4709 = ~n4699 & n4708 ;
  assign n4710 = ~n4696 & n4709 ;
  assign n4711 = n3662 & ~n4710 ;
  assign n4712 = \P1_reg0_reg[28]/NET0131  & n3664 ;
  assign n4713 = ~n4711 & ~n4712 ;
  assign n4714 = \P1_state_reg[0]/NET0131  & ~n4713 ;
  assign n4715 = ~n4692 & ~n4714 ;
  assign n4716 = \P1_reg0_reg[25]/NET0131  & ~n3703 ;
  assign n4717 = \P1_reg0_reg[25]/NET0131  & n3664 ;
  assign n4718 = \P1_reg0_reg[25]/NET0131  & ~n3900 ;
  assign n4719 = n3900 & ~n4563 ;
  assign n4720 = ~n4718 & ~n4719 ;
  assign n4721 = n3557 & ~n4720 ;
  assign n4727 = n3900 & n4571 ;
  assign n4728 = ~n4718 & ~n4727 ;
  assign n4729 = n1898 & ~n4728 ;
  assign n4722 = n3650 & ~n3900 ;
  assign n4723 = n3917 & ~n4722 ;
  assign n4724 = n3575 & ~n3900 ;
  assign n4725 = n4723 & ~n4724 ;
  assign n4726 = \P1_reg0_reg[25]/NET0131  & ~n4725 ;
  assign n4730 = n3575 & ~n4586 ;
  assign n4731 = n1533 & n3683 ;
  assign n4732 = ~n4595 & ~n4731 ;
  assign n4733 = ~n4730 & n4732 ;
  assign n4734 = n3900 & ~n4733 ;
  assign n4735 = ~n4726 & ~n4734 ;
  assign n4736 = ~n4729 & n4735 ;
  assign n4737 = ~n4721 & n4736 ;
  assign n4738 = n3662 & ~n4737 ;
  assign n4739 = ~n4717 & ~n4738 ;
  assign n4740 = \P1_state_reg[0]/NET0131  & ~n4739 ;
  assign n4741 = ~n4716 & ~n4740 ;
  assign n4742 = \P1_reg1_reg[26]/NET0131  & ~n3703 ;
  assign n4743 = \P1_reg1_reg[26]/NET0131  & n3664 ;
  assign n4761 = n4236 & n4481 ;
  assign n4760 = ~\P1_reg1_reg[26]/NET0131  & ~n4236 ;
  assign n4762 = n3575 & ~n4760 ;
  assign n4763 = ~n4761 & n4762 ;
  assign n4746 = n3557 & ~n4515 ;
  assign n4745 = n1898 & ~n4524 ;
  assign n4744 = n3650 & n4531 ;
  assign n4747 = ~n4537 & ~n4744 ;
  assign n4748 = ~n4745 & n4747 ;
  assign n4749 = ~n4746 & n4748 ;
  assign n4750 = n4236 & ~n4749 ;
  assign n4751 = n1898 & ~n4236 ;
  assign n4752 = n3650 & ~n4236 ;
  assign n4753 = n4252 & ~n4752 ;
  assign n4754 = ~n4751 & n4753 ;
  assign n4755 = ~n1735 & n3555 ;
  assign n4756 = ~n4236 & n4755 ;
  assign n4757 = ~n1897 & n4756 ;
  assign n4758 = n4754 & ~n4757 ;
  assign n4759 = \P1_reg1_reg[26]/NET0131  & ~n4758 ;
  assign n4764 = ~n4750 & ~n4759 ;
  assign n4765 = ~n4763 & n4764 ;
  assign n4766 = n3662 & ~n4765 ;
  assign n4767 = ~n4743 & ~n4766 ;
  assign n4768 = \P1_state_reg[0]/NET0131  & ~n4767 ;
  assign n4769 = ~n4742 & ~n4768 ;
  assign n4770 = \P1_reg1_reg[28]/NET0131  & ~n3703 ;
  assign n4771 = \P1_reg1_reg[28]/NET0131  & ~n4236 ;
  assign n4772 = ~n3552 & n4236 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4774 = n3557 & ~n4773 ;
  assign n4775 = ~n3572 & n4236 ;
  assign n4776 = ~n4771 & ~n4775 ;
  assign n4777 = n3575 & ~n4776 ;
  assign n4778 = n4236 & ~n4702 ;
  assign n4779 = \P1_reg1_reg[28]/NET0131  & ~n4754 ;
  assign n4780 = ~n4778 & ~n4779 ;
  assign n4781 = ~n4777 & n4780 ;
  assign n4782 = ~n4774 & n4781 ;
  assign n4783 = n3662 & ~n4782 ;
  assign n4784 = \P1_reg1_reg[28]/NET0131  & n3664 ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4786 = \P1_state_reg[0]/NET0131  & ~n4785 ;
  assign n4787 = ~n4770 & ~n4786 ;
  assign n4789 = n834 & n3664 ;
  assign n4791 = n834 & ~n3450 ;
  assign n4792 = ~n3494 & n3505 ;
  assign n4793 = n3515 & ~n4792 ;
  assign n4794 = n1787 & n4793 ;
  assign n4795 = ~n1787 & ~n4793 ;
  assign n4796 = ~n4794 & ~n4795 ;
  assign n4797 = n3450 & n4796 ;
  assign n4798 = ~n4791 & ~n4797 ;
  assign n4799 = n3557 & ~n4798 ;
  assign n4800 = n796 & ~n3593 ;
  assign n4801 = ~n796 & n3593 ;
  assign n4802 = ~n4800 & ~n4801 ;
  assign n4803 = ~n536 & ~n4802 ;
  assign n4804 = n536 & n999 ;
  assign n4805 = ~n4803 & ~n4804 ;
  assign n4806 = n3450 & n4805 ;
  assign n4807 = ~n4791 & ~n4806 ;
  assign n4808 = n1898 & ~n4807 ;
  assign n4810 = ~n829 & ~n3640 ;
  assign n4809 = n829 & n3640 ;
  assign n4811 = n3650 & ~n4809 ;
  assign n4812 = ~n4810 & n4811 ;
  assign n4814 = n1425 & ~n1787 ;
  assign n4813 = ~n1425 & n1787 ;
  assign n4815 = n3575 & ~n4813 ;
  assign n4816 = ~n4814 & n4815 ;
  assign n4817 = ~n4812 & ~n4816 ;
  assign n4818 = n3450 & ~n4817 ;
  assign n4790 = ~n829 & n3655 ;
  assign n4819 = ~n3450 & n3575 ;
  assign n4820 = n4591 & ~n4819 ;
  assign n4821 = n834 & ~n4820 ;
  assign n4822 = ~n4790 & ~n4821 ;
  assign n4823 = ~n4818 & n4822 ;
  assign n4824 = ~n4808 & n4823 ;
  assign n4825 = ~n4799 & n4824 ;
  assign n4826 = n3662 & ~n4825 ;
  assign n4827 = ~n4789 & ~n4826 ;
  assign n4828 = \P1_state_reg[0]/NET0131  & ~n4827 ;
  assign n4788 = n834 & n1934 ;
  assign n4829 = \P1_reg3_reg[16]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4830 = ~n4788 & ~n4829 ;
  assign n4831 = ~n4828 & n4830 ;
  assign n4832 = \P1_reg2_reg[31]/NET0131  & ~n3703 ;
  assign n4833 = \P1_reg2_reg[31]/NET0131  & n3664 ;
  assign n4851 = n1671 & n3683 ;
  assign n4852 = ~n1677 & n1898 ;
  assign n4853 = n3719 & n4852 ;
  assign n4854 = ~n4851 & ~n4853 ;
  assign n4855 = n3672 & ~n4854 ;
  assign n4834 = n1094 & n3635 ;
  assign n4835 = n3634 & n4834 ;
  assign n4836 = n1064 & n4835 ;
  assign n4837 = n1040 & n4836 ;
  assign n4838 = n1015 & n3625 ;
  assign n4839 = n4837 & n4838 ;
  assign n4840 = n3645 & n4839 ;
  assign n4841 = ~n1607 & ~n1696 ;
  assign n4842 = ~n1637 & n4841 ;
  assign n4843 = n4840 & n4842 ;
  assign n4844 = ~n1671 & n4843 ;
  assign n4845 = n1671 & ~n4843 ;
  assign n4846 = ~n4844 & ~n4845 ;
  assign n4847 = n3672 & ~n4846 ;
  assign n4848 = ~\P1_reg2_reg[31]/NET0131  & ~n3672 ;
  assign n4849 = n3650 & ~n4848 ;
  assign n4850 = ~n4847 & n4849 ;
  assign n4856 = ~n1735 & ~n3672 ;
  assign n4857 = n3685 & ~n4856 ;
  assign n4858 = \P1_reg2_reg[31]/NET0131  & ~n4857 ;
  assign n4859 = ~n3887 & ~n4858 ;
  assign n4860 = ~n4850 & n4859 ;
  assign n4861 = ~n4855 & n4860 ;
  assign n4862 = n3662 & ~n4861 ;
  assign n4863 = ~n4833 & ~n4862 ;
  assign n4864 = \P1_state_reg[0]/NET0131  & ~n4863 ;
  assign n4865 = ~n4832 & ~n4864 ;
  assign n4866 = \P2_reg2_reg[25]/NET0131  & ~n3434 ;
  assign n4867 = \P2_reg2_reg[25]/NET0131  & n3430 ;
  assign n4868 = \P2_reg2_reg[25]/NET0131  & ~n2033 ;
  assign n4884 = n3234 & n3250 ;
  assign n4881 = ~n3194 & n3249 ;
  assign n4882 = n3261 & ~n4881 ;
  assign n4883 = n3242 & ~n4882 ;
  assign n4885 = n3272 & ~n4883 ;
  assign n4886 = ~n4884 & n4885 ;
  assign n4887 = n3288 & ~n4886 ;
  assign n4888 = n3300 & ~n4887 ;
  assign n4889 = n4137 & ~n4888 ;
  assign n4890 = ~n4137 & n4888 ;
  assign n4891 = ~n4889 & ~n4890 ;
  assign n4892 = n2033 & ~n4891 ;
  assign n4893 = ~n4868 & ~n4892 ;
  assign n4894 = n3319 & ~n4893 ;
  assign n4869 = ~n3122 & n3133 ;
  assign n4870 = n2669 & n3149 ;
  assign n4871 = ~n4869 & n4870 ;
  assign n4872 = ~n3144 & n3149 ;
  assign n4873 = n2560 & ~n4872 ;
  assign n4874 = ~n4871 & n4873 ;
  assign n4875 = n4137 & n4874 ;
  assign n4876 = ~n4137 & ~n4874 ;
  assign n4877 = ~n4875 & ~n4876 ;
  assign n4878 = n2033 & ~n4877 ;
  assign n4879 = ~n4868 & ~n4878 ;
  assign n4880 = n3179 & ~n4879 ;
  assign n4896 = n2433 & ~n3355 ;
  assign n4897 = ~n4415 & ~n4896 ;
  assign n4898 = ~n2050 & ~n4897 ;
  assign n4899 = n2050 & n2484 ;
  assign n4900 = ~n4898 & ~n4899 ;
  assign n4901 = n2033 & n4900 ;
  assign n4902 = ~n4868 & ~n4901 ;
  assign n4903 = n3373 & ~n4902 ;
  assign n4905 = n2452 & n3375 ;
  assign n4906 = n3396 & n3398 ;
  assign n4907 = ~n2471 & n4906 ;
  assign n4908 = n2452 & ~n4907 ;
  assign n4909 = n3409 & ~n4424 ;
  assign n4910 = ~n4908 & n4909 ;
  assign n4911 = ~n4905 & ~n4910 ;
  assign n4912 = n2033 & ~n4911 ;
  assign n4895 = \P2_reg2_reg[25]/NET0131  & n3422 ;
  assign n4904 = n2457 & n3415 ;
  assign n4913 = ~n4895 & ~n4904 ;
  assign n4914 = ~n4912 & n4913 ;
  assign n4915 = ~n4903 & n4914 ;
  assign n4916 = ~n4880 & n4915 ;
  assign n4917 = ~n4894 & n4916 ;
  assign n4918 = n2017 & ~n4917 ;
  assign n4919 = ~n4867 & ~n4918 ;
  assign n4920 = \P1_state_reg[0]/NET0131  & ~n4919 ;
  assign n4921 = ~n4866 & ~n4920 ;
  assign n4924 = n2457 & n3430 ;
  assign n4925 = ~n2027 & ~n2032 ;
  assign n4926 = n2457 & ~n4925 ;
  assign n4930 = ~n4891 & n4925 ;
  assign n4931 = ~n4926 & ~n4930 ;
  assign n4932 = n3319 & ~n4931 ;
  assign n4927 = ~n4877 & n4925 ;
  assign n4928 = ~n4926 & ~n4927 ;
  assign n4929 = n3179 & ~n4928 ;
  assign n4936 = n4900 & n4925 ;
  assign n4937 = ~n4926 & ~n4936 ;
  assign n4938 = n3373 & ~n4937 ;
  assign n4940 = ~n4911 & n4925 ;
  assign n4933 = ~n3418 & n4925 ;
  assign n4934 = ~n3421 & ~n4933 ;
  assign n4935 = n2457 & n4934 ;
  assign n4939 = n2452 & n3415 ;
  assign n4941 = ~n4935 & ~n4939 ;
  assign n4942 = ~n4940 & n4941 ;
  assign n4943 = ~n4938 & n4942 ;
  assign n4944 = ~n4929 & n4943 ;
  assign n4945 = ~n4932 & n4944 ;
  assign n4946 = n2017 & ~n4945 ;
  assign n4947 = ~n4924 & ~n4946 ;
  assign n4948 = \P1_state_reg[0]/NET0131  & ~n4947 ;
  assign n4922 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[25]/NET0131  ;
  assign n4923 = n2457 & n3935 ;
  assign n4949 = ~n4922 & ~n4923 ;
  assign n4950 = ~n4948 & n4949 ;
  assign n4951 = n1474 & n3664 ;
  assign n4952 = n1474 & ~n3450 ;
  assign n4953 = n3450 & ~n4481 ;
  assign n4954 = ~n4952 & ~n4953 ;
  assign n4955 = n3575 & ~n4954 ;
  assign n4959 = n3450 & ~n4524 ;
  assign n4960 = ~n4952 & ~n4959 ;
  assign n4961 = n1898 & ~n4960 ;
  assign n4956 = n3450 & ~n4515 ;
  assign n4957 = ~n4952 & ~n4956 ;
  assign n4958 = n3557 & ~n4957 ;
  assign n4963 = n3450 & n4744 ;
  assign n4962 = n1474 & ~n4591 ;
  assign n4964 = n1463 & n3655 ;
  assign n4965 = ~n4962 & ~n4964 ;
  assign n4966 = ~n4963 & n4965 ;
  assign n4967 = ~n4958 & n4966 ;
  assign n4968 = ~n4961 & n4967 ;
  assign n4969 = ~n4955 & n4968 ;
  assign n4970 = n3662 & ~n4969 ;
  assign n4971 = ~n4951 & ~n4970 ;
  assign n4972 = \P1_state_reg[0]/NET0131  & ~n4971 ;
  assign n4973 = \P1_reg3_reg[26]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4974 = n1474 & n1934 ;
  assign n4975 = ~n4973 & ~n4974 ;
  assign n4976 = ~n4972 & n4975 ;
  assign n4977 = n1506 & ~n3450 ;
  assign n4978 = ~n3823 & n3825 ;
  assign n4979 = ~n3828 & ~n4978 ;
  assign n4980 = n3824 & n3834 ;
  assign n4981 = ~n4979 & n4980 ;
  assign n4982 = n3831 & n3834 ;
  assign n4983 = ~n3814 & ~n4982 ;
  assign n4984 = ~n4981 & n4983 ;
  assign n4985 = n3809 & n3813 ;
  assign n4986 = ~n4984 & n4985 ;
  assign n4987 = n3809 & ~n3817 ;
  assign n4988 = ~n3839 & ~n4987 ;
  assign n4989 = ~n4986 & n4988 ;
  assign n4990 = n3807 & n3810 ;
  assign n4991 = ~n4989 & n4990 ;
  assign n4992 = n3807 & n3842 ;
  assign n4993 = ~n3845 & ~n4992 ;
  assign n4994 = ~n4991 & n4993 ;
  assign n4995 = n3853 & n3855 ;
  assign n4996 = n3806 & n3852 ;
  assign n4997 = n4995 & n4996 ;
  assign n4998 = ~n4994 & n4997 ;
  assign n5000 = n3848 & n3852 ;
  assign n5001 = ~n3860 & ~n5000 ;
  assign n5002 = n4995 & ~n5001 ;
  assign n4999 = n3855 & n3863 ;
  assign n5003 = ~n3866 & ~n4999 ;
  assign n5004 = ~n5002 & n5003 ;
  assign n5005 = ~n4998 & n5004 ;
  assign n5006 = n1790 & ~n5005 ;
  assign n5007 = ~n1790 & n5005 ;
  assign n5008 = ~n5006 & ~n5007 ;
  assign n5009 = n3450 & ~n5008 ;
  assign n5010 = ~n4977 & ~n5009 ;
  assign n5011 = n3575 & ~n5010 ;
  assign n5048 = n1646 & ~n3712 ;
  assign n5049 = ~n3713 & ~n5048 ;
  assign n5050 = ~n536 & ~n5049 ;
  assign n5051 = n536 & n1478 ;
  assign n5052 = ~n5050 & ~n5051 ;
  assign n5053 = n3450 & n5052 ;
  assign n5054 = ~n4977 & ~n5053 ;
  assign n5055 = n1898 & ~n5054 ;
  assign n5012 = n3777 & n3780 ;
  assign n5013 = n3754 & n3779 ;
  assign n5014 = n5012 & n5013 ;
  assign n5015 = n3733 & n3735 ;
  assign n5016 = ~n3740 & ~n5015 ;
  assign n5017 = n3725 & n3734 ;
  assign n5018 = ~n5016 & n5017 ;
  assign n5019 = n3725 & ~n3743 ;
  assign n5020 = ~n3747 & ~n5019 ;
  assign n5021 = ~n5018 & n5020 ;
  assign n5022 = n3755 & n3758 ;
  assign n5023 = n3726 & n3757 ;
  assign n5024 = n5022 & n5023 ;
  assign n5025 = ~n5021 & n5024 ;
  assign n5026 = n5014 & n5025 ;
  assign n5034 = ~n3773 & n3779 ;
  assign n5035 = n3786 & ~n5034 ;
  assign n5036 = n5012 & ~n5035 ;
  assign n5027 = ~n3750 & n3757 ;
  assign n5028 = n3763 & ~n5027 ;
  assign n5029 = n5022 & ~n5028 ;
  assign n5030 = n3755 & n3766 ;
  assign n5031 = n3770 & ~n5030 ;
  assign n5032 = ~n5029 & n5031 ;
  assign n5033 = n5014 & ~n5032 ;
  assign n5037 = n3777 & ~n3789 ;
  assign n5038 = n3793 & ~n5037 ;
  assign n5039 = ~n5033 & n5038 ;
  assign n5040 = ~n5036 & n5039 ;
  assign n5041 = ~n5026 & n5040 ;
  assign n5042 = n1790 & n5041 ;
  assign n5043 = ~n1790 & ~n5041 ;
  assign n5044 = ~n5042 & ~n5043 ;
  assign n5045 = n3450 & ~n5044 ;
  assign n5046 = ~n4977 & ~n5045 ;
  assign n5047 = n3557 & ~n5046 ;
  assign n5056 = n3644 & n4839 ;
  assign n5057 = n1500 & ~n5056 ;
  assign n5058 = ~n4840 & ~n5057 ;
  assign n5059 = n3450 & n5058 ;
  assign n5060 = ~n4977 & ~n5059 ;
  assign n5061 = n3650 & ~n5060 ;
  assign n5062 = n1506 & ~n4305 ;
  assign n5063 = n1500 & n3655 ;
  assign n5064 = ~n5062 & ~n5063 ;
  assign n5065 = ~n5061 & n5064 ;
  assign n5066 = ~n5047 & n5065 ;
  assign n5067 = ~n5055 & n5066 ;
  assign n5068 = ~n5011 & n5067 ;
  assign n5069 = n3662 & ~n5068 ;
  assign n5070 = n1506 & n3664 ;
  assign n5071 = ~n5069 & ~n5070 ;
  assign n5072 = \P1_state_reg[0]/NET0131  & ~n5071 ;
  assign n5073 = \P1_reg3_reg[27]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5074 = n1506 & n1934 ;
  assign n5075 = ~n5073 & ~n5074 ;
  assign n5076 = ~n5072 & n5075 ;
  assign n5077 = n2381 & ~n4925 ;
  assign n5078 = ~n4372 & n4925 ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5080 = n3319 & ~n5079 ;
  assign n5081 = ~n4410 & n4925 ;
  assign n5082 = ~n5077 & ~n5081 ;
  assign n5083 = n3179 & ~n5082 ;
  assign n5084 = ~n4421 & n4925 ;
  assign n5085 = ~n5077 & ~n5084 ;
  assign n5086 = n3373 & ~n5085 ;
  assign n5087 = n4427 & n4925 ;
  assign n5088 = ~n5077 & ~n5087 ;
  assign n5089 = n3409 & ~n5088 ;
  assign n5090 = ~n4433 & ~n4933 ;
  assign n5091 = n2381 & n5090 ;
  assign n5092 = n3375 & n4925 ;
  assign n5093 = ~n3415 & ~n5092 ;
  assign n5094 = n2376 & ~n5093 ;
  assign n5095 = ~n5091 & ~n5094 ;
  assign n5096 = ~n5089 & n5095 ;
  assign n5097 = ~n5086 & n5096 ;
  assign n5098 = ~n5083 & n5097 ;
  assign n5099 = ~n5080 & n5098 ;
  assign n5100 = n2017 & ~n5099 ;
  assign n5101 = n2381 & n3430 ;
  assign n5102 = ~n5100 & ~n5101 ;
  assign n5103 = \P1_state_reg[0]/NET0131  & ~n5102 ;
  assign n5104 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[27]/NET0131  ;
  assign n5105 = n2381 & n3935 ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = ~n5103 & n5106 ;
  assign n5108 = n2324 & ~n4925 ;
  assign n5109 = n4090 & ~n4107 ;
  assign n5110 = n4084 & n4086 ;
  assign n5111 = ~n5109 & n5110 ;
  assign n5112 = ~n3999 & n4084 ;
  assign n5113 = n4081 & ~n5112 ;
  assign n5114 = ~n5111 & n5113 ;
  assign n5115 = n4199 & ~n5114 ;
  assign n5116 = n4070 & ~n4075 ;
  assign n5117 = ~n4063 & ~n5116 ;
  assign n5118 = ~n5115 & n5117 ;
  assign n5119 = n4119 & ~n5118 ;
  assign n5120 = ~n4119 & n5118 ;
  assign n5121 = ~n5119 & ~n5120 ;
  assign n5122 = n4925 & ~n5121 ;
  assign n5123 = ~n5108 & ~n5122 ;
  assign n5124 = n3319 & ~n5123 ;
  assign n5133 = ~n2792 & ~n2885 ;
  assign n5134 = ~n2834 & n5133 ;
  assign n5135 = ~n2881 & ~n5134 ;
  assign n5136 = ~n2720 & ~n2746 ;
  assign n5137 = ~n2769 & ~n2859 ;
  assign n5138 = n5136 & n5137 ;
  assign n5139 = n5135 & n5138 ;
  assign n5140 = ~n2884 & ~n2892 ;
  assign n5141 = ~n2769 & ~n5140 ;
  assign n5142 = n5136 & n5141 ;
  assign n5143 = ~n2720 & n2891 ;
  assign n5144 = ~n2897 & ~n5143 ;
  assign n5145 = ~n5142 & n5144 ;
  assign n5146 = ~n5139 & n5145 ;
  assign n5147 = ~n2693 & ~n3006 ;
  assign n5148 = ~n2927 & ~n2981 ;
  assign n5149 = n5147 & n5148 ;
  assign n5150 = ~n5146 & n5149 ;
  assign n5151 = ~n2896 & ~n3011 ;
  assign n5152 = ~n3006 & ~n5151 ;
  assign n5153 = n5148 & n5152 ;
  assign n5154 = ~n2927 & n3010 ;
  assign n5155 = ~n3016 & ~n5154 ;
  assign n5156 = ~n5153 & n5155 ;
  assign n5157 = ~n5150 & n5156 ;
  assign n5158 = ~n2955 & ~n3119 ;
  assign n5159 = ~n3072 & ~n3096 ;
  assign n5160 = n5158 & n5159 ;
  assign n5161 = ~n2641 & ~n3047 ;
  assign n5162 = ~n2614 & ~n2667 ;
  assign n5163 = n5161 & n5162 ;
  assign n5164 = n5160 & n5163 ;
  assign n5165 = ~n5157 & n5164 ;
  assign n5166 = ~n3015 & ~n3125 ;
  assign n5167 = ~n3119 & ~n5166 ;
  assign n5168 = n5159 & n5167 ;
  assign n5169 = ~n3072 & n3124 ;
  assign n5170 = ~n3130 & ~n5169 ;
  assign n5171 = ~n5168 & n5170 ;
  assign n5172 = n5163 & ~n5171 ;
  assign n5173 = ~n3129 & ~n3136 ;
  assign n5174 = ~n2641 & ~n5173 ;
  assign n5175 = n5162 & n5174 ;
  assign n5176 = ~n3135 & ~n3141 ;
  assign n5177 = ~n2614 & ~n5176 ;
  assign n5178 = ~n5175 & ~n5177 ;
  assign n5179 = ~n5172 & n5178 ;
  assign n5180 = ~n5165 & n5179 ;
  assign n5181 = ~n2589 & ~n3147 ;
  assign n5182 = ~n2508 & ~n2533 ;
  assign n5183 = n5181 & n5182 ;
  assign n5184 = n2435 & n4378 ;
  assign n5185 = n5183 & n5184 ;
  assign n5186 = ~n5180 & n5185 ;
  assign n5187 = n3140 & ~n3147 ;
  assign n5188 = ~n2552 & ~n5187 ;
  assign n5189 = n5182 & ~n5188 ;
  assign n5190 = ~n2508 & n2532 ;
  assign n5191 = ~n2557 & ~n5190 ;
  assign n5192 = ~n5189 & n5191 ;
  assign n5193 = n5184 & ~n5192 ;
  assign n5194 = ~n2462 & n2556 ;
  assign n5195 = ~n2564 & ~n5194 ;
  assign n5196 = n2435 & ~n5195 ;
  assign n5197 = ~n2386 & n2563 ;
  assign n5198 = ~n2562 & ~n5197 ;
  assign n5199 = ~n5196 & n5198 ;
  assign n5200 = ~n5193 & n5199 ;
  assign n5201 = ~n5186 & n5200 ;
  assign n5202 = n4119 & n5201 ;
  assign n5203 = ~n4119 & ~n5201 ;
  assign n5204 = ~n5202 & ~n5203 ;
  assign n5205 = n4925 & ~n5204 ;
  assign n5206 = ~n5108 & ~n5205 ;
  assign n5207 = n3179 & ~n5206 ;
  assign n5125 = n2241 & ~n4418 ;
  assign n5126 = ~n3357 & ~n5125 ;
  assign n5127 = ~n2050 & ~n5126 ;
  assign n5128 = n2050 & n2385 ;
  assign n5129 = ~n5127 & ~n5128 ;
  assign n5130 = n4925 & n5129 ;
  assign n5131 = ~n5108 & ~n5130 ;
  assign n5132 = n3373 & ~n5131 ;
  assign n5209 = n2315 & ~n3403 ;
  assign n5210 = ~n3404 & ~n5209 ;
  assign n5211 = n4925 & n5210 ;
  assign n5212 = ~n5108 & ~n5211 ;
  assign n5213 = n3409 & ~n5212 ;
  assign n5208 = n2324 & n5090 ;
  assign n5214 = n2315 & ~n5093 ;
  assign n5215 = ~n5208 & ~n5214 ;
  assign n5216 = ~n5213 & n5215 ;
  assign n5217 = ~n5132 & n5216 ;
  assign n5218 = ~n5207 & n5217 ;
  assign n5219 = ~n5124 & n5218 ;
  assign n5220 = n2017 & ~n5219 ;
  assign n5221 = n2324 & n3430 ;
  assign n5222 = ~n5220 & ~n5221 ;
  assign n5223 = \P1_state_reg[0]/NET0131  & ~n5222 ;
  assign n5224 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[28]/NET0131  ;
  assign n5225 = n2324 & n3935 ;
  assign n5226 = ~n5224 & ~n5225 ;
  assign n5227 = ~n5223 & n5226 ;
  assign n5228 = \P2_reg0_reg[25]/NET0131  & ~n3434 ;
  assign n5229 = \P2_reg0_reg[25]/NET0131  & n3430 ;
  assign n5234 = \P2_reg0_reg[25]/NET0131  & ~n4610 ;
  assign n5238 = n4610 & ~n4891 ;
  assign n5239 = ~n5234 & ~n5238 ;
  assign n5240 = n3319 & ~n5239 ;
  assign n5235 = n4610 & ~n4877 ;
  assign n5236 = ~n5234 & ~n5235 ;
  assign n5237 = n3179 & ~n5236 ;
  assign n5230 = n3373 & n4900 ;
  assign n5231 = n4911 & ~n5230 ;
  assign n5232 = n4610 & ~n5231 ;
  assign n5233 = \P2_reg0_reg[25]/NET0131  & ~n4623 ;
  assign n5241 = ~n5232 & ~n5233 ;
  assign n5242 = ~n5237 & n5241 ;
  assign n5243 = ~n5240 & n5242 ;
  assign n5244 = n2017 & ~n5243 ;
  assign n5245 = ~n5229 & ~n5244 ;
  assign n5246 = \P1_state_reg[0]/NET0131  & ~n5245 ;
  assign n5247 = ~n5228 & ~n5246 ;
  assign n5248 = \P2_reg0_reg[27]/NET0131  & ~n4610 ;
  assign n5249 = ~n4372 & n4610 ;
  assign n5250 = ~n5248 & ~n5249 ;
  assign n5251 = n3319 & ~n5250 ;
  assign n5252 = ~n4410 & n4610 ;
  assign n5253 = ~n5248 & ~n5252 ;
  assign n5254 = n3179 & ~n5253 ;
  assign n5255 = n3375 & ~n4610 ;
  assign n5256 = n4619 & ~n5255 ;
  assign n5257 = n3409 & ~n4610 ;
  assign n5258 = n5256 & ~n5257 ;
  assign n5259 = ~n4622 & n5258 ;
  assign n5260 = \P2_reg0_reg[27]/NET0131  & ~n5259 ;
  assign n5261 = ~n4430 & n4610 ;
  assign n5262 = ~n5260 & ~n5261 ;
  assign n5263 = ~n5254 & n5262 ;
  assign n5264 = ~n5251 & n5263 ;
  assign n5265 = n2017 & ~n5264 ;
  assign n5266 = \P2_reg0_reg[27]/NET0131  & n3430 ;
  assign n5267 = ~n5265 & ~n5266 ;
  assign n5268 = \P1_state_reg[0]/NET0131  & ~n5267 ;
  assign n5269 = \P2_reg0_reg[27]/NET0131  & ~n3434 ;
  assign n5270 = ~n5268 & ~n5269 ;
  assign n5271 = \P2_reg0_reg[26]/NET0131  & ~n4610 ;
  assign n5272 = n5135 & n5137 ;
  assign n5273 = ~n5141 & ~n5272 ;
  assign n5274 = n5136 & n5147 ;
  assign n5275 = ~n5273 & n5274 ;
  assign n5276 = ~n5144 & n5147 ;
  assign n5277 = ~n5152 & ~n5276 ;
  assign n5278 = ~n5275 & n5277 ;
  assign n5279 = n5148 & n5158 ;
  assign n5280 = ~n5278 & n5279 ;
  assign n5281 = ~n5155 & n5158 ;
  assign n5282 = ~n5167 & ~n5281 ;
  assign n5283 = ~n5280 & n5282 ;
  assign n5284 = n5159 & n5161 ;
  assign n5285 = ~n5283 & n5284 ;
  assign n5286 = n5161 & ~n5170 ;
  assign n5287 = ~n5174 & ~n5286 ;
  assign n5288 = ~n5285 & n5287 ;
  assign n5289 = n5162 & n5181 ;
  assign n5290 = ~n2533 & n4379 ;
  assign n5291 = n5289 & n5290 ;
  assign n5292 = ~n5288 & n5291 ;
  assign n5294 = n5177 & n5181 ;
  assign n5295 = n5188 & ~n5294 ;
  assign n5296 = n5290 & ~n5295 ;
  assign n5293 = n4378 & ~n5191 ;
  assign n5297 = n5195 & ~n5293 ;
  assign n5298 = ~n5296 & n5297 ;
  assign n5299 = ~n5292 & n5298 ;
  assign n5300 = n4135 & n5299 ;
  assign n5301 = ~n4135 & ~n5299 ;
  assign n5302 = ~n5300 & ~n5301 ;
  assign n5303 = n4610 & ~n5302 ;
  assign n5304 = ~n5271 & ~n5303 ;
  assign n5305 = n3179 & ~n5304 ;
  assign n5306 = ~n4087 & ~n4106 ;
  assign n5307 = n3993 & n4043 ;
  assign n5308 = n4000 & n4005 ;
  assign n5309 = n5307 & n5308 ;
  assign n5310 = ~n5306 & n5309 ;
  assign n5311 = n3998 & n4043 ;
  assign n5312 = ~n4077 & ~n5311 ;
  assign n5313 = n4005 & n4089 ;
  assign n5314 = ~n3995 & ~n5313 ;
  assign n5315 = n5307 & ~n5314 ;
  assign n5316 = n5312 & ~n5315 ;
  assign n5317 = ~n5310 & n5316 ;
  assign n5318 = n4037 & n4050 ;
  assign n5319 = n4038 & n4042 ;
  assign n5320 = n5318 & n5319 ;
  assign n5321 = ~n5317 & n5320 ;
  assign n5323 = n4038 & n4080 ;
  assign n5324 = n4072 & ~n5323 ;
  assign n5325 = n5318 & ~n5324 ;
  assign n5322 = n4050 & n4074 ;
  assign n5326 = ~n4060 & ~n5322 ;
  assign n5327 = ~n5325 & n5326 ;
  assign n5328 = ~n5321 & n5327 ;
  assign n5329 = n4135 & ~n5328 ;
  assign n5330 = ~n4135 & n5328 ;
  assign n5331 = ~n5329 & ~n5330 ;
  assign n5332 = n4610 & ~n5331 ;
  assign n5333 = ~n5271 & ~n5332 ;
  assign n5334 = n3319 & ~n5333 ;
  assign n5335 = n2385 & ~n4415 ;
  assign n5336 = ~n4416 & ~n5335 ;
  assign n5337 = ~n2050 & ~n5336 ;
  assign n5338 = n2050 & n2461 ;
  assign n5339 = ~n5337 & ~n5338 ;
  assign n5340 = n3373 & n5339 ;
  assign n5341 = n2424 & n3375 ;
  assign n5342 = n2424 & ~n4424 ;
  assign n5343 = n3409 & ~n4425 ;
  assign n5344 = ~n5342 & n5343 ;
  assign n5345 = ~n5341 & ~n5344 ;
  assign n5346 = ~n5340 & n5345 ;
  assign n5347 = n4610 & ~n5346 ;
  assign n5348 = \P2_reg0_reg[26]/NET0131  & ~n5259 ;
  assign n5349 = ~n5347 & ~n5348 ;
  assign n5350 = ~n5334 & n5349 ;
  assign n5351 = ~n5305 & n5350 ;
  assign n5352 = n2017 & ~n5351 ;
  assign n5353 = \P2_reg0_reg[26]/NET0131  & n3430 ;
  assign n5354 = ~n5352 & ~n5353 ;
  assign n5355 = \P1_state_reg[0]/NET0131  & ~n5354 ;
  assign n5356 = \P2_reg0_reg[26]/NET0131  & ~n3434 ;
  assign n5357 = ~n5355 & ~n5356 ;
  assign n5358 = \P2_reg0_reg[28]/NET0131  & ~n4610 ;
  assign n5359 = n4610 & ~n5121 ;
  assign n5360 = ~n5358 & ~n5359 ;
  assign n5361 = n3319 & ~n5360 ;
  assign n5365 = n4610 & n5129 ;
  assign n5366 = ~n5358 & ~n5365 ;
  assign n5367 = n3373 & ~n5366 ;
  assign n5362 = n4610 & ~n5204 ;
  assign n5363 = ~n5358 & ~n5362 ;
  assign n5364 = n3179 & ~n5363 ;
  assign n5369 = n4610 & n5210 ;
  assign n5370 = ~n5358 & ~n5369 ;
  assign n5371 = n3409 & ~n5370 ;
  assign n5368 = \P2_reg0_reg[28]/NET0131  & ~n5256 ;
  assign n5372 = n2315 & n3375 ;
  assign n5373 = n4610 & n5372 ;
  assign n5374 = ~n5368 & ~n5373 ;
  assign n5375 = ~n5371 & n5374 ;
  assign n5376 = ~n5364 & n5375 ;
  assign n5377 = ~n5367 & n5376 ;
  assign n5378 = ~n5361 & n5377 ;
  assign n5379 = n2017 & ~n5378 ;
  assign n5380 = \P2_reg0_reg[28]/NET0131  & n3430 ;
  assign n5381 = ~n5379 & ~n5380 ;
  assign n5382 = \P1_state_reg[0]/NET0131  & ~n5381 ;
  assign n5383 = \P2_reg0_reg[28]/NET0131  & ~n3434 ;
  assign n5384 = ~n5382 & ~n5383 ;
  assign n5385 = n4275 & n4610 ;
  assign n5386 = ~n4272 & n5385 ;
  assign n5387 = ~n3178 & ~n3371 ;
  assign n5388 = ~n4610 & ~n5387 ;
  assign n5389 = n4275 & ~n5388 ;
  assign n5390 = n5256 & n5389 ;
  assign n5391 = \P2_reg0_reg[31]/NET0131  & ~n5390 ;
  assign n5392 = ~n5386 & ~n5391 ;
  assign n5393 = \P1_reg2_reg[20]/NET0131  & ~n3703 ;
  assign n5394 = \P1_reg2_reg[20]/NET0131  & n3664 ;
  assign n5396 = \P1_reg2_reg[20]/NET0131  & ~n3672 ;
  assign n5407 = n1776 & ~n3527 ;
  assign n5408 = ~n1776 & n3527 ;
  assign n5409 = ~n5407 & ~n5408 ;
  assign n5410 = n3672 & n5409 ;
  assign n5411 = ~n5396 & ~n5410 ;
  assign n5412 = n3557 & ~n5411 ;
  assign n5397 = n3594 & n3711 ;
  assign n5398 = n949 & ~n5397 ;
  assign n5399 = ~n949 & n5397 ;
  assign n5400 = ~n5398 & ~n5399 ;
  assign n5401 = ~n536 & ~n5400 ;
  assign n5402 = n536 & n692 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = n3672 & n5403 ;
  assign n5405 = ~n5396 & ~n5404 ;
  assign n5406 = n1898 & ~n5405 ;
  assign n5414 = n1776 & ~n3564 ;
  assign n5415 = ~n1776 & n3564 ;
  assign n5416 = ~n5414 & ~n5415 ;
  assign n5417 = n3575 & ~n5416 ;
  assign n5413 = n964 & n3683 ;
  assign n5418 = n3621 & n3640 ;
  assign n5419 = n638 & n5418 ;
  assign n5421 = ~n964 & n5419 ;
  assign n5420 = n964 & ~n5419 ;
  assign n5422 = n3650 & ~n5420 ;
  assign n5423 = ~n5421 & n5422 ;
  assign n5424 = ~n5413 & ~n5423 ;
  assign n5425 = ~n5417 & n5424 ;
  assign n5426 = n3672 & ~n5425 ;
  assign n5395 = n969 & n1736 ;
  assign n5427 = n3616 & ~n3672 ;
  assign n5428 = ~n3615 & ~n5427 ;
  assign n5429 = n3575 & ~n3672 ;
  assign n5430 = n5428 & ~n5429 ;
  assign n5431 = \P1_reg2_reg[20]/NET0131  & ~n5430 ;
  assign n5432 = ~n5395 & ~n5431 ;
  assign n5433 = ~n5426 & n5432 ;
  assign n5434 = ~n5406 & n5433 ;
  assign n5435 = ~n5412 & n5434 ;
  assign n5436 = n3662 & ~n5435 ;
  assign n5437 = ~n5394 & ~n5436 ;
  assign n5438 = \P1_state_reg[0]/NET0131  & ~n5437 ;
  assign n5439 = ~n5393 & ~n5438 ;
  assign n5440 = \P1_reg2_reg[25]/NET0131  & ~n3703 ;
  assign n5441 = \P1_reg2_reg[25]/NET0131  & n3664 ;
  assign n5442 = \P1_reg2_reg[25]/NET0131  & ~n3672 ;
  assign n5443 = n3672 & ~n4563 ;
  assign n5444 = ~n5442 & ~n5443 ;
  assign n5445 = n3557 & ~n5444 ;
  assign n5447 = n3672 & n4571 ;
  assign n5448 = ~n5442 & ~n5447 ;
  assign n5449 = n1898 & ~n5448 ;
  assign n5446 = n3672 & ~n4733 ;
  assign n5450 = n1538 & n1736 ;
  assign n5451 = n3650 & ~n3672 ;
  assign n5452 = n3685 & ~n5451 ;
  assign n5453 = ~n5429 & n5452 ;
  assign n5454 = \P1_reg2_reg[25]/NET0131  & ~n5453 ;
  assign n5455 = ~n5450 & ~n5454 ;
  assign n5456 = ~n5446 & n5455 ;
  assign n5457 = ~n5449 & n5456 ;
  assign n5458 = ~n5445 & n5457 ;
  assign n5459 = n3662 & ~n5458 ;
  assign n5460 = ~n5441 & ~n5459 ;
  assign n5461 = \P1_state_reg[0]/NET0131  & ~n5460 ;
  assign n5462 = ~n5440 & ~n5461 ;
  assign n5463 = \P1_reg2_reg[27]/NET0131  & ~n3672 ;
  assign n5464 = n3672 & ~n5008 ;
  assign n5465 = ~n5463 & ~n5464 ;
  assign n5466 = n3575 & ~n5465 ;
  assign n5470 = n3672 & n5052 ;
  assign n5471 = ~n5463 & ~n5470 ;
  assign n5472 = n1898 & ~n5471 ;
  assign n5467 = n3672 & ~n5044 ;
  assign n5468 = ~n5463 & ~n5467 ;
  assign n5469 = n3557 & ~n5468 ;
  assign n5473 = n3672 & n5058 ;
  assign n5474 = ~n5463 & ~n5473 ;
  assign n5475 = n3650 & ~n5474 ;
  assign n5478 = n1500 & n3683 ;
  assign n5479 = n3672 & n5478 ;
  assign n5476 = \P1_reg2_reg[27]/NET0131  & ~n3685 ;
  assign n5477 = n1506 & n1736 ;
  assign n5480 = ~n5476 & ~n5477 ;
  assign n5481 = ~n5479 & n5480 ;
  assign n5482 = ~n5475 & n5481 ;
  assign n5483 = ~n5469 & n5482 ;
  assign n5484 = ~n5472 & n5483 ;
  assign n5485 = ~n5466 & n5484 ;
  assign n5486 = n3662 & ~n5485 ;
  assign n5487 = \P1_reg2_reg[27]/NET0131  & n3664 ;
  assign n5488 = ~n5486 & ~n5487 ;
  assign n5489 = \P1_state_reg[0]/NET0131  & ~n5488 ;
  assign n5490 = \P1_reg2_reg[27]/NET0131  & ~n3703 ;
  assign n5491 = ~n5489 & ~n5490 ;
  assign n5492 = \P2_reg1_reg[24]/NET0131  & ~n3434 ;
  assign n5493 = \P2_reg1_reg[24]/NET0131  & n3430 ;
  assign n5513 = \P2_reg1_reg[24]/NET0131  & ~n4663 ;
  assign n5527 = ~n5156 & n5160 ;
  assign n5528 = n5171 & ~n5527 ;
  assign n5529 = n5163 & ~n5528 ;
  assign n5526 = n5150 & n5164 ;
  assign n5530 = n5178 & ~n5526 ;
  assign n5531 = ~n5529 & n5530 ;
  assign n5532 = n5183 & ~n5531 ;
  assign n5533 = n5192 & ~n5532 ;
  assign n5534 = n4136 & n5533 ;
  assign n5535 = ~n4136 & ~n5533 ;
  assign n5536 = ~n5534 & ~n5535 ;
  assign n5537 = n4663 & ~n5536 ;
  assign n5538 = ~n5513 & ~n5537 ;
  assign n5539 = n3179 & ~n5538 ;
  assign n5517 = n4085 & n4108 ;
  assign n5514 = n4084 & ~n4092 ;
  assign n5515 = n4081 & ~n5514 ;
  assign n5516 = n4076 & ~n5515 ;
  assign n5518 = n4075 & ~n5516 ;
  assign n5519 = ~n5517 & n5518 ;
  assign n5520 = n4136 & ~n5519 ;
  assign n5521 = ~n4136 & n5519 ;
  assign n5522 = ~n5520 & ~n5521 ;
  assign n5523 = n4663 & ~n5522 ;
  assign n5524 = ~n5513 & ~n5523 ;
  assign n5525 = n3319 & ~n5524 ;
  assign n5494 = n2471 & n3375 ;
  assign n5495 = n3344 & n3353 ;
  assign n5496 = n2461 & ~n5495 ;
  assign n5497 = ~n3355 & ~n5496 ;
  assign n5498 = ~n2050 & ~n5497 ;
  assign n5499 = n2050 & n2507 ;
  assign n5500 = n3373 & ~n5499 ;
  assign n5501 = ~n5498 & n5500 ;
  assign n5502 = n2471 & ~n4906 ;
  assign n5503 = n3409 & ~n4907 ;
  assign n5504 = ~n5502 & n5503 ;
  assign n5505 = ~n5501 & ~n5504 ;
  assign n5506 = ~n5494 & n5505 ;
  assign n5507 = n4663 & ~n5506 ;
  assign n5508 = n3420 & ~n4663 ;
  assign n5509 = n4619 & ~n5508 ;
  assign n5510 = n3373 & ~n4663 ;
  assign n5511 = n5509 & ~n5510 ;
  assign n5512 = \P2_reg1_reg[24]/NET0131  & ~n5511 ;
  assign n5540 = ~n5507 & ~n5512 ;
  assign n5541 = ~n5525 & n5540 ;
  assign n5542 = ~n5539 & n5541 ;
  assign n5543 = n2017 & ~n5542 ;
  assign n5544 = ~n5493 & ~n5543 ;
  assign n5545 = \P1_state_reg[0]/NET0131  & ~n5544 ;
  assign n5546 = ~n5492 & ~n5545 ;
  assign n5547 = \P2_reg1_reg[26]/NET0131  & ~n3434 ;
  assign n5548 = \P2_reg1_reg[26]/NET0131  & ~n4663 ;
  assign n5549 = n4663 & ~n5302 ;
  assign n5550 = ~n5548 & ~n5549 ;
  assign n5551 = n3179 & ~n5550 ;
  assign n5552 = n4663 & ~n5331 ;
  assign n5553 = ~n5548 & ~n5552 ;
  assign n5554 = n3319 & ~n5553 ;
  assign n5555 = n4663 & ~n5346 ;
  assign n5556 = \P2_reg1_reg[26]/NET0131  & ~n5511 ;
  assign n5557 = ~n5555 & ~n5556 ;
  assign n5558 = ~n5554 & n5557 ;
  assign n5559 = ~n5551 & n5558 ;
  assign n5560 = n2017 & ~n5559 ;
  assign n5561 = \P2_reg1_reg[26]/NET0131  & n3430 ;
  assign n5562 = ~n5560 & ~n5561 ;
  assign n5563 = \P1_state_reg[0]/NET0131  & ~n5562 ;
  assign n5564 = ~n5547 & ~n5563 ;
  assign n5565 = n3375 & ~n4663 ;
  assign n5566 = n4619 & ~n5565 ;
  assign n5567 = ~n4663 & ~n5387 ;
  assign n5568 = n5566 & ~n5567 ;
  assign n5569 = n4275 & n5568 ;
  assign n5570 = \P2_reg1_reg[27]/NET0131  & ~n5569 ;
  assign n5571 = n2017 & n4663 ;
  assign n5572 = \P1_state_reg[0]/NET0131  & n5571 ;
  assign n5574 = n3319 & ~n4372 ;
  assign n5573 = n3179 & ~n4410 ;
  assign n5575 = n4430 & ~n5573 ;
  assign n5576 = ~n5574 & n5575 ;
  assign n5577 = n5572 & ~n5576 ;
  assign n5578 = ~n5570 & ~n5577 ;
  assign n5579 = \P2_reg1_reg[28]/NET0131  & ~n4663 ;
  assign n5580 = n4663 & ~n5121 ;
  assign n5581 = ~n5579 & ~n5580 ;
  assign n5582 = n3319 & ~n5581 ;
  assign n5586 = n4663 & n5129 ;
  assign n5587 = ~n5579 & ~n5586 ;
  assign n5588 = n3373 & ~n5587 ;
  assign n5583 = n4663 & ~n5204 ;
  assign n5584 = ~n5579 & ~n5583 ;
  assign n5585 = n3179 & ~n5584 ;
  assign n5590 = n4663 & n5210 ;
  assign n5591 = ~n5579 & ~n5590 ;
  assign n5592 = n3409 & ~n5591 ;
  assign n5589 = \P2_reg1_reg[28]/NET0131  & ~n5566 ;
  assign n5593 = n4663 & n5372 ;
  assign n5594 = ~n5589 & ~n5593 ;
  assign n5595 = ~n5592 & n5594 ;
  assign n5596 = ~n5585 & n5595 ;
  assign n5597 = ~n5588 & n5596 ;
  assign n5598 = ~n5582 & n5597 ;
  assign n5599 = n2017 & ~n5598 ;
  assign n5600 = \P2_reg1_reg[28]/NET0131  & n3430 ;
  assign n5601 = ~n5599 & ~n5600 ;
  assign n5602 = \P1_state_reg[0]/NET0131  & ~n5601 ;
  assign n5603 = \P2_reg1_reg[28]/NET0131  & ~n3434 ;
  assign n5604 = ~n5602 & ~n5603 ;
  assign n5605 = ~n3178 & ~n3372 ;
  assign n5606 = ~n4663 & ~n5605 ;
  assign n5607 = n4275 & ~n5606 ;
  assign n5608 = n5509 & n5607 ;
  assign n5609 = \P2_reg1_reg[31]/NET0131  & ~n5608 ;
  assign n5610 = ~n4272 & n5572 ;
  assign n5611 = ~n5609 & ~n5610 ;
  assign n5612 = \P2_reg2_reg[28]/NET0131  & ~n2033 ;
  assign n5613 = n2033 & ~n5121 ;
  assign n5614 = ~n5612 & ~n5613 ;
  assign n5615 = n3319 & ~n5614 ;
  assign n5619 = n2033 & ~n5204 ;
  assign n5620 = ~n5612 & ~n5619 ;
  assign n5621 = n3179 & ~n5620 ;
  assign n5616 = n2033 & n5129 ;
  assign n5617 = ~n5612 & ~n5616 ;
  assign n5618 = n3373 & ~n5617 ;
  assign n5623 = n2033 & n5210 ;
  assign n5624 = ~n5612 & ~n5623 ;
  assign n5625 = n3409 & ~n5624 ;
  assign n5627 = n2033 & n5372 ;
  assign n5622 = \P2_reg2_reg[28]/NET0131  & n4434 ;
  assign n5626 = n2324 & n3415 ;
  assign n5628 = ~n5622 & ~n5626 ;
  assign n5629 = ~n5627 & n5628 ;
  assign n5630 = ~n5625 & n5629 ;
  assign n5631 = ~n5618 & n5630 ;
  assign n5632 = ~n5621 & n5631 ;
  assign n5633 = ~n5615 & n5632 ;
  assign n5634 = n2017 & ~n5633 ;
  assign n5635 = \P2_reg2_reg[28]/NET0131  & n3430 ;
  assign n5636 = ~n5634 & ~n5635 ;
  assign n5637 = \P1_state_reg[0]/NET0131  & ~n5636 ;
  assign n5638 = \P2_reg2_reg[28]/NET0131  & ~n3434 ;
  assign n5639 = ~n5637 & ~n5638 ;
  assign n5640 = \P1_reg0_reg[26]/NET0131  & ~n3703 ;
  assign n5641 = \P1_reg0_reg[26]/NET0131  & n3664 ;
  assign n5647 = n3900 & n4481 ;
  assign n5646 = ~\P1_reg0_reg[26]/NET0131  & ~n3900 ;
  assign n5648 = n3575 & ~n5646 ;
  assign n5649 = ~n5647 & n5648 ;
  assign n5642 = n3900 & ~n4749 ;
  assign n5643 = ~n3900 & n4755 ;
  assign n5644 = n4723 & ~n5643 ;
  assign n5645 = \P1_reg0_reg[26]/NET0131  & ~n5644 ;
  assign n5650 = ~n5642 & ~n5645 ;
  assign n5651 = ~n5649 & n5650 ;
  assign n5652 = n3662 & ~n5651 ;
  assign n5653 = ~n5641 & ~n5652 ;
  assign n5654 = \P1_state_reg[0]/NET0131  & ~n5653 ;
  assign n5655 = ~n5640 & ~n5654 ;
  assign n5656 = \P1_reg0_reg[27]/NET0131  & ~n3900 ;
  assign n5657 = n3900 & ~n5008 ;
  assign n5658 = ~n5656 & ~n5657 ;
  assign n5659 = n3575 & ~n5658 ;
  assign n5663 = n3900 & ~n5044 ;
  assign n5664 = ~n5656 & ~n5663 ;
  assign n5665 = n3557 & ~n5664 ;
  assign n5660 = n3900 & n5052 ;
  assign n5661 = ~n5656 & ~n5660 ;
  assign n5662 = n1898 & ~n5661 ;
  assign n5666 = n3900 & n5058 ;
  assign n5667 = ~n5656 & ~n5666 ;
  assign n5668 = n3650 & ~n5667 ;
  assign n5669 = \P1_reg0_reg[27]/NET0131  & ~n3917 ;
  assign n5670 = n3900 & n5478 ;
  assign n5671 = ~n5669 & ~n5670 ;
  assign n5672 = ~n5668 & n5671 ;
  assign n5673 = ~n5662 & n5672 ;
  assign n5674 = ~n5665 & n5673 ;
  assign n5675 = ~n5659 & n5674 ;
  assign n5676 = n3662 & ~n5675 ;
  assign n5677 = \P1_reg0_reg[27]/NET0131  & n3664 ;
  assign n5678 = ~n5676 & ~n5677 ;
  assign n5679 = \P1_state_reg[0]/NET0131  & ~n5678 ;
  assign n5680 = \P1_reg0_reg[27]/NET0131  & ~n3703 ;
  assign n5681 = ~n5679 & ~n5680 ;
  assign n5682 = \P1_reg1_reg[25]/NET0131  & ~n3703 ;
  assign n5683 = \P1_reg1_reg[25]/NET0131  & n3664 ;
  assign n5684 = \P1_reg1_reg[25]/NET0131  & ~n4236 ;
  assign n5685 = n4236 & ~n4563 ;
  assign n5686 = ~n5684 & ~n5685 ;
  assign n5687 = n3557 & ~n5686 ;
  assign n5688 = n4236 & n4571 ;
  assign n5689 = ~n5684 & ~n5688 ;
  assign n5690 = n1898 & ~n5689 ;
  assign n5691 = n4236 & ~n4586 ;
  assign n5692 = ~n5684 & ~n5691 ;
  assign n5693 = n3575 & ~n5692 ;
  assign n5695 = n4236 & n4594 ;
  assign n5696 = ~n5684 & ~n5695 ;
  assign n5697 = n3650 & ~n5696 ;
  assign n5694 = n4236 & n4731 ;
  assign n5698 = \P1_reg1_reg[25]/NET0131  & ~n4252 ;
  assign n5699 = ~n5694 & ~n5698 ;
  assign n5700 = ~n5697 & n5699 ;
  assign n5701 = ~n5693 & n5700 ;
  assign n5702 = ~n5690 & n5701 ;
  assign n5703 = ~n5687 & n5702 ;
  assign n5704 = n3662 & ~n5703 ;
  assign n5705 = ~n5683 & ~n5704 ;
  assign n5706 = \P1_state_reg[0]/NET0131  & ~n5705 ;
  assign n5707 = ~n5682 & ~n5706 ;
  assign n5708 = \P1_reg1_reg[27]/NET0131  & ~n4236 ;
  assign n5709 = n4236 & ~n5008 ;
  assign n5710 = ~n5708 & ~n5709 ;
  assign n5711 = n3575 & ~n5710 ;
  assign n5715 = n4236 & n5052 ;
  assign n5716 = ~n5708 & ~n5715 ;
  assign n5717 = n1898 & ~n5716 ;
  assign n5712 = n4236 & ~n5044 ;
  assign n5713 = ~n5708 & ~n5712 ;
  assign n5714 = n3557 & ~n5713 ;
  assign n5718 = n4236 & n5058 ;
  assign n5719 = ~n5708 & ~n5718 ;
  assign n5720 = n3650 & ~n5719 ;
  assign n5721 = \P1_reg1_reg[27]/NET0131  & ~n4252 ;
  assign n5722 = n4236 & n5478 ;
  assign n5723 = ~n5721 & ~n5722 ;
  assign n5724 = ~n5720 & n5723 ;
  assign n5725 = ~n5714 & n5724 ;
  assign n5726 = ~n5717 & n5725 ;
  assign n5727 = ~n5711 & n5726 ;
  assign n5728 = n3662 & ~n5727 ;
  assign n5729 = \P1_reg1_reg[27]/NET0131  & n3664 ;
  assign n5730 = ~n5728 & ~n5729 ;
  assign n5731 = \P1_state_reg[0]/NET0131  & ~n5730 ;
  assign n5732 = \P1_reg1_reg[27]/NET0131  & ~n3703 ;
  assign n5733 = ~n5731 & ~n5732 ;
  assign n5735 = n1068 & n3664 ;
  assign n5754 = ~n1762 & n3494 ;
  assign n5753 = n1762 & ~n3494 ;
  assign n5755 = n3557 & ~n5753 ;
  assign n5756 = ~n5754 & n5755 ;
  assign n5738 = ~n1115 & n3587 ;
  assign n5739 = ~n1075 & n5738 ;
  assign n5740 = n1051 & ~n5739 ;
  assign n5741 = ~n1051 & n5739 ;
  assign n5742 = ~n5740 & ~n5741 ;
  assign n5743 = ~n536 & ~n5742 ;
  assign n5737 = n536 & n1115 ;
  assign n5744 = n1898 & ~n5737 ;
  assign n5745 = ~n5743 & n5744 ;
  assign n5747 = n1762 & n3559 ;
  assign n5746 = ~n1762 & ~n3559 ;
  assign n5748 = n3575 & ~n5746 ;
  assign n5749 = ~n5747 & n5748 ;
  assign n5750 = ~n1094 & ~n3636 ;
  assign n5751 = n3650 & ~n4835 ;
  assign n5752 = ~n5750 & n5751 ;
  assign n5757 = ~n5749 & ~n5752 ;
  assign n5758 = ~n5745 & n5757 ;
  assign n5759 = ~n5756 & n5758 ;
  assign n5760 = n3450 & ~n5759 ;
  assign n5736 = ~n1094 & n3655 ;
  assign n5761 = ~n1731 & ~n3556 ;
  assign n5762 = ~n3450 & ~n5761 ;
  assign n5763 = n4305 & ~n5762 ;
  assign n5764 = n1068 & ~n5763 ;
  assign n5765 = ~n5736 & ~n5764 ;
  assign n5766 = ~n5760 & n5765 ;
  assign n5767 = n3662 & ~n5766 ;
  assign n5768 = ~n5735 & ~n5767 ;
  assign n5769 = \P1_state_reg[0]/NET0131  & ~n5768 ;
  assign n5734 = \P1_reg3_reg[12]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5770 = n1068 & n1934 ;
  assign n5771 = ~n5734 & ~n5770 ;
  assign n5772 = ~n5769 & n5771 ;
  assign n5775 = n748 & n3664 ;
  assign n5777 = n748 & ~n3450 ;
  assign n5787 = n1799 & ~n4467 ;
  assign n5788 = ~n1799 & n4467 ;
  assign n5789 = ~n5787 & ~n5788 ;
  assign n5790 = n3450 & ~n5789 ;
  assign n5791 = ~n5777 & ~n5790 ;
  assign n5792 = n3575 & ~n5791 ;
  assign n5778 = n4491 & ~n4506 ;
  assign n5779 = n4489 & ~n5778 ;
  assign n5780 = n4494 & ~n5779 ;
  assign n5781 = n1799 & ~n5780 ;
  assign n5782 = ~n1799 & n5780 ;
  assign n5783 = ~n5781 & ~n5782 ;
  assign n5784 = n3450 & n5783 ;
  assign n5785 = ~n5777 & ~n5784 ;
  assign n5786 = n3557 & ~n5785 ;
  assign n5793 = ~n692 & n3711 ;
  assign n5794 = n692 & ~n3711 ;
  assign n5795 = ~n5793 & ~n5794 ;
  assign n5796 = ~n536 & ~n5795 ;
  assign n5797 = n536 & n796 ;
  assign n5798 = ~n5796 & ~n5797 ;
  assign n5799 = n3450 & n5798 ;
  assign n5800 = ~n5777 & ~n5799 ;
  assign n5801 = n1898 & ~n5800 ;
  assign n5802 = n785 & n4809 ;
  assign n5803 = ~n743 & ~n5802 ;
  assign n5804 = n3650 & ~n5418 ;
  assign n5805 = ~n5803 & n5804 ;
  assign n5806 = n3450 & n5805 ;
  assign n5776 = n748 & ~n3618 ;
  assign n5807 = ~n743 & n3655 ;
  assign n5808 = ~n5776 & ~n5807 ;
  assign n5809 = ~n5806 & n5808 ;
  assign n5810 = ~n5801 & n5809 ;
  assign n5811 = ~n5786 & n5810 ;
  assign n5812 = ~n5792 & n5811 ;
  assign n5813 = n3662 & ~n5812 ;
  assign n5814 = ~n5775 & ~n5813 ;
  assign n5815 = \P1_state_reg[0]/NET0131  & ~n5814 ;
  assign n5773 = \P1_reg3_reg[18]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5774 = n748 & n1934 ;
  assign n5816 = ~n5773 & ~n5774 ;
  assign n5817 = ~n5815 & n5816 ;
  assign n5818 = n2636 & n3430 ;
  assign n5820 = n2636 & ~n4925 ;
  assign n5821 = ~n3056 & n3344 ;
  assign n5822 = n3345 & n5821 ;
  assign n5823 = ~n2666 & n5822 ;
  assign n5824 = n2666 & ~n5822 ;
  assign n5825 = ~n5823 & ~n5824 ;
  assign n5826 = ~n2050 & ~n5825 ;
  assign n5827 = n2050 & n3046 ;
  assign n5828 = ~n5826 & ~n5827 ;
  assign n5829 = n4925 & n5828 ;
  assign n5830 = ~n5820 & ~n5829 ;
  assign n5831 = n3373 & ~n5830 ;
  assign n5838 = ~n3235 & n3249 ;
  assign n5839 = n3261 & ~n5838 ;
  assign n5840 = n4132 & n5839 ;
  assign n5841 = ~n4132 & ~n5839 ;
  assign n5842 = ~n5840 & ~n5841 ;
  assign n5843 = n4925 & n5842 ;
  assign n5844 = ~n5820 & ~n5843 ;
  assign n5845 = n3319 & ~n5844 ;
  assign n5832 = n4132 & n4869 ;
  assign n5833 = ~n4132 & ~n4869 ;
  assign n5834 = ~n5832 & ~n5833 ;
  assign n5835 = n4925 & ~n5834 ;
  assign n5836 = ~n5820 & ~n5835 ;
  assign n5837 = n3179 & ~n5836 ;
  assign n5846 = n3389 & n3398 ;
  assign n5847 = ~n2630 & n5846 ;
  assign n5848 = n2630 & ~n5846 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5850 = n4925 & n5849 ;
  assign n5851 = ~n5820 & ~n5850 ;
  assign n5852 = n3409 & ~n5851 ;
  assign n5819 = n2630 & ~n5093 ;
  assign n5853 = n2636 & n5090 ;
  assign n5854 = ~n5819 & ~n5853 ;
  assign n5855 = ~n5852 & n5854 ;
  assign n5856 = ~n5837 & n5855 ;
  assign n5857 = ~n5845 & n5856 ;
  assign n5858 = ~n5831 & n5857 ;
  assign n5859 = n2017 & ~n5858 ;
  assign n5860 = ~n5818 & ~n5859 ;
  assign n5861 = \P1_state_reg[0]/NET0131  & ~n5860 ;
  assign n5862 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[17]/NET0131  ;
  assign n5863 = n2636 & n3935 ;
  assign n5864 = ~n5862 & ~n5863 ;
  assign n5865 = ~n5861 & n5864 ;
  assign n5866 = n2662 & n3430 ;
  assign n5868 = n2662 & ~n4925 ;
  assign n5869 = n2613 & ~n5823 ;
  assign n5870 = ~n2613 & n5823 ;
  assign n5871 = ~n5869 & ~n5870 ;
  assign n5872 = ~n2050 & ~n5871 ;
  assign n5873 = n2050 & n2640 ;
  assign n5874 = ~n5872 & ~n5873 ;
  assign n5875 = n4925 & n5874 ;
  assign n5876 = ~n5868 & ~n5875 ;
  assign n5877 = n3373 & ~n5876 ;
  assign n5878 = n4145 & ~n5288 ;
  assign n5879 = ~n4145 & n5288 ;
  assign n5880 = ~n5878 & ~n5879 ;
  assign n5881 = n4925 & n5880 ;
  assign n5882 = ~n5868 & ~n5881 ;
  assign n5883 = n3179 & ~n5882 ;
  assign n5884 = n4145 & ~n5317 ;
  assign n5885 = ~n4145 & n5317 ;
  assign n5886 = ~n5884 & ~n5885 ;
  assign n5887 = n4925 & ~n5886 ;
  assign n5888 = ~n5868 & ~n5887 ;
  assign n5889 = n3319 & ~n5888 ;
  assign n5890 = n2657 & ~n5847 ;
  assign n5891 = ~n2657 & n5847 ;
  assign n5892 = ~n5890 & ~n5891 ;
  assign n5893 = n3409 & n5892 ;
  assign n5894 = n4925 & n5893 ;
  assign n5867 = n2662 & n4934 ;
  assign n5895 = n2657 & ~n5093 ;
  assign n5896 = ~n5867 & ~n5895 ;
  assign n5897 = ~n5894 & n5896 ;
  assign n5898 = ~n5889 & n5897 ;
  assign n5899 = ~n5883 & n5898 ;
  assign n5900 = ~n5877 & n5899 ;
  assign n5901 = n2017 & ~n5900 ;
  assign n5902 = ~n5866 & ~n5901 ;
  assign n5903 = \P1_state_reg[0]/NET0131  & ~n5902 ;
  assign n5904 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[18]/NET0131  ;
  assign n5905 = n2662 & n3935 ;
  assign n5906 = ~n5904 & ~n5905 ;
  assign n5907 = ~n5903 & n5906 ;
  assign n5909 = n2609 & n3430 ;
  assign n5929 = n2604 & ~n5891 ;
  assign n5928 = ~n2604 & n5891 ;
  assign n5930 = n3409 & ~n5928 ;
  assign n5931 = ~n5929 & n5930 ;
  assign n5921 = n4126 & n4359 ;
  assign n5920 = ~n4126 & ~n4359 ;
  assign n5922 = n3319 & ~n5920 ;
  assign n5923 = ~n5921 & n5922 ;
  assign n5925 = ~n4126 & n4402 ;
  assign n5924 = n4126 & ~n4402 ;
  assign n5926 = n3179 & ~n5924 ;
  assign n5927 = ~n5925 & n5926 ;
  assign n5932 = ~n5923 & ~n5927 ;
  assign n5933 = ~n5931 & n5932 ;
  assign n5934 = n4925 & ~n5933 ;
  assign n5910 = n2050 & ~n2666 ;
  assign n5912 = n2588 & ~n5870 ;
  assign n5911 = n3344 & n3349 ;
  assign n5913 = ~n2050 & ~n5911 ;
  assign n5914 = ~n5912 & n5913 ;
  assign n5915 = ~n5910 & ~n5914 ;
  assign n5916 = n4925 & n5915 ;
  assign n5917 = ~n2609 & ~n4925 ;
  assign n5918 = n3373 & ~n5917 ;
  assign n5919 = ~n5916 & n5918 ;
  assign n5935 = ~n3179 & ~n3319 ;
  assign n5936 = ~n4925 & ~n5935 ;
  assign n5937 = ~n4934 & ~n5936 ;
  assign n5938 = n2609 & ~n5937 ;
  assign n5939 = n2604 & ~n5093 ;
  assign n5940 = ~n5938 & ~n5939 ;
  assign n5941 = ~n5919 & n5940 ;
  assign n5942 = ~n5934 & n5941 ;
  assign n5943 = n2017 & ~n5942 ;
  assign n5944 = ~n5909 & ~n5943 ;
  assign n5945 = \P1_state_reg[0]/NET0131  & ~n5944 ;
  assign n5908 = n2609 & n3935 ;
  assign n5946 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[19]/NET0131  ;
  assign n5947 = ~n5908 & ~n5946 ;
  assign n5948 = ~n5945 & n5947 ;
  assign n5949 = \P1_reg2_reg[17]/NET0131  & ~n3703 ;
  assign n5950 = \P1_reg2_reg[17]/NET0131  & n3664 ;
  assign n5951 = \P1_reg2_reg[17]/NET0131  & ~n3672 ;
  assign n5965 = n752 & ~n4801 ;
  assign n5966 = ~n3711 & ~n5965 ;
  assign n5967 = ~n536 & ~n5966 ;
  assign n5968 = n536 & n838 ;
  assign n5969 = ~n5967 & ~n5968 ;
  assign n5970 = n3672 & n5969 ;
  assign n5971 = ~n5951 & ~n5970 ;
  assign n5972 = n1898 & ~n5971 ;
  assign n5952 = n3811 & ~n3837 ;
  assign n5953 = n3843 & ~n5952 ;
  assign n5954 = n1773 & n5953 ;
  assign n5955 = ~n1773 & ~n5953 ;
  assign n5956 = ~n5954 & ~n5955 ;
  assign n5957 = n3672 & ~n5956 ;
  assign n5958 = ~n5951 & ~n5957 ;
  assign n5959 = n3575 & ~n5958 ;
  assign n5974 = n1773 & ~n4556 ;
  assign n5975 = ~n1773 & n4556 ;
  assign n5976 = ~n5974 & ~n5975 ;
  assign n5977 = n3672 & ~n5976 ;
  assign n5978 = ~n5951 & ~n5977 ;
  assign n5979 = n3557 & ~n5978 ;
  assign n5960 = ~n785 & ~n4809 ;
  assign n5961 = ~n5802 & ~n5960 ;
  assign n5962 = n3672 & n5961 ;
  assign n5963 = ~n5951 & ~n5962 ;
  assign n5964 = n3650 & ~n5963 ;
  assign n5981 = ~n785 & n3683 ;
  assign n5982 = n3672 & n5981 ;
  assign n5973 = \P1_reg2_reg[17]/NET0131  & ~n3685 ;
  assign n5980 = n792 & n1736 ;
  assign n5983 = ~n5973 & ~n5980 ;
  assign n5984 = ~n5982 & n5983 ;
  assign n5985 = ~n5964 & n5984 ;
  assign n5986 = ~n5979 & n5985 ;
  assign n5987 = ~n5959 & n5986 ;
  assign n5988 = ~n5972 & n5987 ;
  assign n5989 = n3662 & ~n5988 ;
  assign n5990 = ~n5950 & ~n5989 ;
  assign n5991 = \P1_state_reg[0]/NET0131  & ~n5990 ;
  assign n5992 = ~n5949 & ~n5991 ;
  assign n5995 = n969 & n3664 ;
  assign n5997 = n969 & ~n3450 ;
  assign n6001 = n3450 & n5409 ;
  assign n6002 = ~n5997 & ~n6001 ;
  assign n6003 = n3557 & ~n6002 ;
  assign n5998 = n3450 & n5403 ;
  assign n5999 = ~n5997 & ~n5998 ;
  assign n6000 = n1898 & ~n5999 ;
  assign n6004 = n3450 & ~n5416 ;
  assign n6005 = ~n5997 & ~n6004 ;
  assign n6006 = n3575 & ~n6005 ;
  assign n6007 = n3450 & n5423 ;
  assign n5996 = n969 & ~n3618 ;
  assign n6008 = n964 & n3655 ;
  assign n6009 = ~n5996 & ~n6008 ;
  assign n6010 = ~n6007 & n6009 ;
  assign n6011 = ~n6006 & n6010 ;
  assign n6012 = ~n6000 & n6011 ;
  assign n6013 = ~n6003 & n6012 ;
  assign n6014 = n3662 & ~n6013 ;
  assign n6015 = ~n5995 & ~n6014 ;
  assign n6016 = \P1_state_reg[0]/NET0131  & ~n6015 ;
  assign n5993 = \P1_reg3_reg[20]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5994 = n969 & n1934 ;
  assign n6017 = ~n5993 & ~n5994 ;
  assign n6018 = ~n6016 & n6017 ;
  assign n6019 = \P2_reg0_reg[22]/NET0131  & ~n3434 ;
  assign n6020 = \P2_reg0_reg[22]/NET0131  & n3430 ;
  assign n6021 = \P2_reg0_reg[22]/NET0131  & ~n4610 ;
  assign n6022 = ~n5288 & n5289 ;
  assign n6023 = n5295 & ~n6022 ;
  assign n6024 = n4122 & n6023 ;
  assign n6025 = ~n4122 & ~n6023 ;
  assign n6026 = ~n6024 & ~n6025 ;
  assign n6027 = n4610 & ~n6026 ;
  assign n6028 = ~n6021 & ~n6027 ;
  assign n6029 = n3179 & ~n6028 ;
  assign n6030 = ~n5306 & n5308 ;
  assign n6031 = n5314 & ~n6030 ;
  assign n6032 = n5307 & n5319 ;
  assign n6033 = ~n6031 & n6032 ;
  assign n6034 = ~n5312 & n5319 ;
  assign n6035 = n5324 & ~n6034 ;
  assign n6036 = ~n6033 & n6035 ;
  assign n6037 = n4122 & ~n6036 ;
  assign n6038 = ~n4122 & n6036 ;
  assign n6039 = ~n6037 & ~n6038 ;
  assign n6040 = n4610 & ~n6039 ;
  assign n6041 = ~n6021 & ~n6040 ;
  assign n6042 = n3319 & ~n6041 ;
  assign n6044 = n2050 & ~n2551 ;
  assign n6045 = n3344 & n3352 ;
  assign n6046 = n3344 & n3350 ;
  assign n6047 = ~n2531 & n6046 ;
  assign n6048 = ~n2050 & ~n2507 ;
  assign n6049 = ~n6047 & ~n6048 ;
  assign n6050 = ~n6045 & ~n6049 ;
  assign n6051 = ~n6044 & ~n6050 ;
  assign n6052 = n3373 & ~n6051 ;
  assign n6043 = n2522 & n3375 ;
  assign n6053 = n3393 & n5846 ;
  assign n6055 = ~n2522 & n6053 ;
  assign n6054 = n2522 & ~n6053 ;
  assign n6056 = n3409 & ~n6054 ;
  assign n6057 = ~n6055 & n6056 ;
  assign n6058 = ~n6043 & ~n6057 ;
  assign n6059 = ~n6052 & n6058 ;
  assign n6060 = n4610 & ~n6059 ;
  assign n6061 = \P2_reg0_reg[22]/NET0131  & ~n5259 ;
  assign n6062 = ~n6060 & ~n6061 ;
  assign n6063 = ~n6042 & n6062 ;
  assign n6064 = ~n6029 & n6063 ;
  assign n6065 = n2017 & ~n6064 ;
  assign n6066 = ~n6020 & ~n6065 ;
  assign n6067 = \P1_state_reg[0]/NET0131  & ~n6066 ;
  assign n6068 = ~n6019 & ~n6067 ;
  assign n6069 = n3555 & n4856 ;
  assign n6070 = ~n1951 & n3703 ;
  assign n6071 = ~n6069 & n6070 ;
  assign n6072 = n5430 & n6071 ;
  assign n6073 = \P1_reg2_reg[16]/NET0131  & ~n6072 ;
  assign n6074 = n834 & n1736 ;
  assign n6076 = n3557 & n4796 ;
  assign n6077 = n1898 & n4805 ;
  assign n6075 = ~n829 & n3683 ;
  assign n6078 = n4817 & ~n6075 ;
  assign n6079 = ~n6077 & n6078 ;
  assign n6080 = ~n6076 & n6079 ;
  assign n6081 = n3672 & ~n6080 ;
  assign n6082 = ~n6074 & ~n6081 ;
  assign n6083 = n6070 & ~n6082 ;
  assign n6084 = ~n6073 & ~n6083 ;
  assign n6085 = \P2_reg0_reg[24]/NET0131  & ~n3434 ;
  assign n6086 = \P2_reg0_reg[24]/NET0131  & n3430 ;
  assign n6089 = \P2_reg0_reg[24]/NET0131  & ~n4610 ;
  assign n6093 = n4610 & ~n5536 ;
  assign n6094 = ~n6089 & ~n6093 ;
  assign n6095 = n3179 & ~n6094 ;
  assign n6090 = n4610 & ~n5522 ;
  assign n6091 = ~n6089 & ~n6090 ;
  assign n6092 = n3319 & ~n6091 ;
  assign n6087 = n4610 & ~n5506 ;
  assign n6088 = \P2_reg0_reg[24]/NET0131  & ~n5259 ;
  assign n6096 = ~n6087 & ~n6088 ;
  assign n6097 = ~n6092 & n6096 ;
  assign n6098 = ~n6095 & n6097 ;
  assign n6099 = n2017 & ~n6098 ;
  assign n6100 = ~n6086 & ~n6099 ;
  assign n6101 = \P1_state_reg[0]/NET0131  & ~n6100 ;
  assign n6102 = ~n6085 & ~n6101 ;
  assign n6103 = \P2_reg1_reg[25]/NET0131  & ~n3434 ;
  assign n6104 = \P2_reg1_reg[25]/NET0131  & n3430 ;
  assign n6105 = \P2_reg1_reg[25]/NET0131  & ~n4663 ;
  assign n6109 = n4663 & ~n4891 ;
  assign n6110 = ~n6105 & ~n6109 ;
  assign n6111 = n3319 & ~n6110 ;
  assign n6106 = n4663 & ~n4877 ;
  assign n6107 = ~n6105 & ~n6106 ;
  assign n6108 = n3179 & ~n6107 ;
  assign n6113 = n4663 & n4900 ;
  assign n6114 = ~n6105 & ~n6113 ;
  assign n6115 = n3373 & ~n6114 ;
  assign n6112 = \P2_reg1_reg[25]/NET0131  & ~n5509 ;
  assign n6116 = n4663 & ~n4911 ;
  assign n6117 = ~n6112 & ~n6116 ;
  assign n6118 = ~n6115 & n6117 ;
  assign n6119 = ~n6108 & n6118 ;
  assign n6120 = ~n6111 & n6119 ;
  assign n6121 = n2017 & ~n6120 ;
  assign n6122 = ~n6104 & ~n6121 ;
  assign n6123 = \P1_state_reg[0]/NET0131  & ~n6122 ;
  assign n6124 = ~n6103 & ~n6123 ;
  assign n6125 = \P2_reg2_reg[24]/NET0131  & ~n3434 ;
  assign n6126 = \P2_reg2_reg[24]/NET0131  & n3430 ;
  assign n6127 = \P2_reg2_reg[24]/NET0131  & ~n2033 ;
  assign n6131 = n2033 & ~n5536 ;
  assign n6132 = ~n6127 & ~n6131 ;
  assign n6133 = n3179 & ~n6132 ;
  assign n6128 = n2033 & ~n5522 ;
  assign n6129 = ~n6127 & ~n6128 ;
  assign n6130 = n3319 & ~n6129 ;
  assign n6135 = n2033 & ~n5506 ;
  assign n6134 = n2480 & n3415 ;
  assign n6136 = \P2_reg2_reg[24]/NET0131  & ~n4437 ;
  assign n6137 = ~n6134 & ~n6136 ;
  assign n6138 = ~n6135 & n6137 ;
  assign n6139 = ~n6130 & n6138 ;
  assign n6140 = ~n6133 & n6139 ;
  assign n6141 = n2017 & ~n6140 ;
  assign n6142 = ~n6126 & ~n6141 ;
  assign n6143 = \P1_state_reg[0]/NET0131  & ~n6142 ;
  assign n6144 = ~n6125 & ~n6143 ;
  assign n6145 = \P2_reg2_reg[26]/NET0131  & ~n2033 ;
  assign n6146 = n2033 & ~n5302 ;
  assign n6147 = ~n6145 & ~n6146 ;
  assign n6148 = n3179 & ~n6147 ;
  assign n6149 = n2033 & ~n5331 ;
  assign n6150 = ~n6145 & ~n6149 ;
  assign n6151 = n3319 & ~n6150 ;
  assign n6152 = n2033 & ~n5346 ;
  assign n6153 = n2429 & n3415 ;
  assign n6154 = \P2_reg2_reg[26]/NET0131  & ~n4437 ;
  assign n6155 = ~n6153 & ~n6154 ;
  assign n6156 = ~n6152 & n6155 ;
  assign n6157 = ~n6151 & n6156 ;
  assign n6158 = ~n6148 & n6157 ;
  assign n6159 = n2017 & ~n6158 ;
  assign n6160 = \P2_reg2_reg[26]/NET0131  & n3430 ;
  assign n6161 = ~n6159 & ~n6160 ;
  assign n6162 = \P1_state_reg[0]/NET0131  & ~n6161 ;
  assign n6163 = \P2_reg2_reg[26]/NET0131  & ~n3434 ;
  assign n6164 = ~n6162 & ~n6163 ;
  assign n6165 = n3616 & ~n3900 ;
  assign n6166 = n3915 & ~n4724 ;
  assign n6167 = ~n6165 & n6166 ;
  assign n6168 = ~n5643 & n6167 ;
  assign n6169 = n6070 & n6168 ;
  assign n6170 = \P1_reg0_reg[16]/NET0131  & ~n6169 ;
  assign n6171 = n3900 & n6070 ;
  assign n6172 = ~n6080 & n6171 ;
  assign n6173 = ~n6170 & ~n6172 ;
  assign n6174 = \P1_reg0_reg[21]/NET0131  & ~n3703 ;
  assign n6175 = \P1_reg0_reg[21]/NET0131  & n3664 ;
  assign n6176 = ~n3900 & ~n5761 ;
  assign n6177 = n3917 & ~n6176 ;
  assign n6178 = \P1_reg0_reg[21]/NET0131  & ~n6177 ;
  assign n6179 = n887 & ~n5399 ;
  assign n6180 = n3596 & n3711 ;
  assign n6181 = ~n6179 & ~n6180 ;
  assign n6182 = ~n536 & ~n6181 ;
  assign n6183 = n536 & n973 ;
  assign n6184 = ~n6182 & ~n6183 ;
  assign n6185 = n1898 & n6184 ;
  assign n6186 = n939 & ~n5421 ;
  assign n6187 = ~n939 & n5421 ;
  assign n6188 = ~n6186 & ~n6187 ;
  assign n6189 = n3650 & n6188 ;
  assign n6190 = n939 & n3683 ;
  assign n6192 = n1786 & ~n3776 ;
  assign n6191 = ~n1786 & n3776 ;
  assign n6193 = n3557 & ~n6191 ;
  assign n6194 = ~n6192 & n6193 ;
  assign n6196 = ~n1786 & ~n3851 ;
  assign n6195 = n1786 & n3851 ;
  assign n6197 = n3575 & ~n6195 ;
  assign n6198 = ~n6196 & n6197 ;
  assign n6199 = ~n6194 & ~n6198 ;
  assign n6200 = ~n6190 & n6199 ;
  assign n6201 = ~n6189 & n6200 ;
  assign n6202 = ~n6185 & n6201 ;
  assign n6203 = n3900 & ~n6202 ;
  assign n6204 = ~n6178 & ~n6203 ;
  assign n6205 = n3662 & ~n6204 ;
  assign n6206 = ~n6175 & ~n6205 ;
  assign n6207 = \P1_state_reg[0]/NET0131  & ~n6206 ;
  assign n6208 = ~n6174 & ~n6207 ;
  assign n6209 = \P1_reg0_reg[24]/NET0131  & ~n3703 ;
  assign n6210 = \P1_reg0_reg[24]/NET0131  & n3664 ;
  assign n6211 = \P1_reg0_reg[24]/NET0131  & ~n3900 ;
  assign n6220 = n3900 & ~n4317 ;
  assign n6221 = ~n6211 & ~n6220 ;
  assign n6222 = n3557 & ~n6221 ;
  assign n6212 = n3900 & n4292 ;
  assign n6213 = ~n6211 & ~n6212 ;
  assign n6214 = n1898 & ~n6213 ;
  assign n6223 = n3900 & ~n4329 ;
  assign n6224 = ~n6211 & ~n6223 ;
  assign n6225 = n3575 & ~n6224 ;
  assign n6216 = n3900 & n4300 ;
  assign n6217 = ~n6211 & ~n6216 ;
  assign n6218 = n3650 & ~n6217 ;
  assign n6215 = \P1_reg0_reg[24]/NET0131  & ~n3917 ;
  assign n6219 = n3900 & n4645 ;
  assign n6226 = ~n6215 & ~n6219 ;
  assign n6227 = ~n6218 & n6226 ;
  assign n6228 = ~n6225 & n6227 ;
  assign n6229 = ~n6214 & n6228 ;
  assign n6230 = ~n6222 & n6229 ;
  assign n6231 = n3662 & ~n6230 ;
  assign n6232 = ~n6210 & ~n6231 ;
  assign n6233 = \P1_state_reg[0]/NET0131  & ~n6232 ;
  assign n6234 = ~n6209 & ~n6233 ;
  assign n6235 = n3650 & n4846 ;
  assign n6236 = n4854 & ~n6235 ;
  assign n6237 = n6171 & ~n6236 ;
  assign n6238 = n3915 & n6171 ;
  assign n6239 = \P1_reg0_reg[31]/NET0131  & ~n6238 ;
  assign n6240 = ~n6237 & ~n6239 ;
  assign n6241 = n3575 & ~n4236 ;
  assign n6242 = n4753 & ~n6241 ;
  assign n6243 = ~n4756 & n6242 ;
  assign n6244 = n6070 & n6243 ;
  assign n6245 = \P1_reg1_reg[16]/NET0131  & ~n6244 ;
  assign n6246 = n4236 & n6070 ;
  assign n6247 = ~n6080 & n6246 ;
  assign n6248 = ~n6245 & ~n6247 ;
  assign n6249 = \P1_reg1_reg[17]/NET0131  & ~n3703 ;
  assign n6250 = \P1_reg1_reg[17]/NET0131  & n3664 ;
  assign n6251 = n1898 & n5969 ;
  assign n6253 = n3575 & ~n5956 ;
  assign n6254 = n3650 & n5961 ;
  assign n6252 = n3557 & ~n5976 ;
  assign n6255 = ~n5981 & ~n6252 ;
  assign n6256 = ~n6254 & n6255 ;
  assign n6257 = ~n6253 & n6256 ;
  assign n6258 = ~n6251 & n6257 ;
  assign n6259 = n4236 & ~n6258 ;
  assign n6260 = \P1_reg1_reg[17]/NET0131  & ~n6243 ;
  assign n6261 = ~n6259 & ~n6260 ;
  assign n6262 = n3662 & ~n6261 ;
  assign n6263 = ~n6250 & ~n6262 ;
  assign n6264 = \P1_state_reg[0]/NET0131  & ~n6263 ;
  assign n6265 = ~n6249 & ~n6264 ;
  assign n6266 = \P1_reg1_reg[21]/NET0131  & ~n3703 ;
  assign n6267 = \P1_reg1_reg[21]/NET0131  & n3664 ;
  assign n6270 = n4236 & ~n6184 ;
  assign n6269 = ~\P1_reg1_reg[21]/NET0131  & ~n4236 ;
  assign n6271 = n1898 & ~n6269 ;
  assign n6272 = ~n6270 & n6271 ;
  assign n6268 = n4236 & ~n6201 ;
  assign n6273 = n3556 & ~n4236 ;
  assign n6274 = n1732 & ~n4236 ;
  assign n6275 = ~n6273 & ~n6274 ;
  assign n6276 = n4252 & n6275 ;
  assign n6277 = \P1_reg1_reg[21]/NET0131  & ~n6276 ;
  assign n6278 = ~n6268 & ~n6277 ;
  assign n6279 = ~n6272 & n6278 ;
  assign n6280 = n3662 & ~n6279 ;
  assign n6281 = ~n6267 & ~n6280 ;
  assign n6282 = \P1_state_reg[0]/NET0131  & ~n6281 ;
  assign n6283 = ~n6266 & ~n6282 ;
  assign n6284 = \P1_reg1_reg[24]/NET0131  & ~n3703 ;
  assign n6285 = \P1_reg1_reg[24]/NET0131  & n3664 ;
  assign n6286 = \P1_reg1_reg[24]/NET0131  & ~n4236 ;
  assign n6295 = n4236 & ~n4317 ;
  assign n6296 = ~n6286 & ~n6295 ;
  assign n6297 = n3557 & ~n6296 ;
  assign n6287 = n4236 & n4292 ;
  assign n6288 = ~n6286 & ~n6287 ;
  assign n6289 = n1898 & ~n6288 ;
  assign n6298 = n4236 & ~n4329 ;
  assign n6299 = ~n6286 & ~n6298 ;
  assign n6300 = n3575 & ~n6299 ;
  assign n6291 = n4236 & n4300 ;
  assign n6292 = ~n6286 & ~n6291 ;
  assign n6293 = n3650 & ~n6292 ;
  assign n6290 = n4236 & n4645 ;
  assign n6294 = \P1_reg1_reg[24]/NET0131  & ~n4252 ;
  assign n6301 = ~n6290 & ~n6294 ;
  assign n6302 = ~n6293 & n6301 ;
  assign n6303 = ~n6300 & n6302 ;
  assign n6304 = ~n6289 & n6303 ;
  assign n6305 = ~n6297 & n6304 ;
  assign n6306 = n3662 & ~n6305 ;
  assign n6307 = ~n6285 & ~n6306 ;
  assign n6308 = \P1_state_reg[0]/NET0131  & ~n6307 ;
  assign n6309 = ~n6284 & ~n6308 ;
  assign n6310 = ~n6236 & n6246 ;
  assign n6311 = n3915 & n6246 ;
  assign n6312 = \P1_reg1_reg[31]/NET0131  & ~n6311 ;
  assign n6313 = ~n6310 & ~n6312 ;
  assign n6315 = n792 & n3664 ;
  assign n6317 = n792 & ~n3450 ;
  assign n6318 = n3450 & n5969 ;
  assign n6319 = ~n6317 & ~n6318 ;
  assign n6320 = n1898 & ~n6319 ;
  assign n6321 = n3450 & ~n5956 ;
  assign n6322 = ~n6317 & ~n6321 ;
  assign n6323 = n3575 & ~n6322 ;
  assign n6324 = n3450 & ~n5976 ;
  assign n6325 = ~n6317 & ~n6324 ;
  assign n6326 = n3557 & ~n6325 ;
  assign n6327 = n3450 & n6254 ;
  assign n6316 = n792 & ~n3618 ;
  assign n6328 = ~n785 & n3655 ;
  assign n6329 = ~n6316 & ~n6328 ;
  assign n6330 = ~n6327 & n6329 ;
  assign n6331 = ~n6326 & n6330 ;
  assign n6332 = ~n6323 & n6331 ;
  assign n6333 = ~n6320 & n6332 ;
  assign n6334 = n3662 & ~n6333 ;
  assign n6335 = ~n6315 & ~n6334 ;
  assign n6336 = \P1_state_reg[0]/NET0131  & ~n6335 ;
  assign n6314 = n792 & n1934 ;
  assign n6337 = \P1_reg3_reg[17]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6338 = ~n6314 & ~n6337 ;
  assign n6339 = ~n6336 & n6338 ;
  assign n6342 = n688 & n3664 ;
  assign n6344 = n688 & ~n3450 ;
  assign n6351 = n973 & ~n5793 ;
  assign n6352 = ~n5397 & ~n6351 ;
  assign n6353 = ~n536 & ~n6352 ;
  assign n6354 = n536 & n752 ;
  assign n6355 = ~n6353 & ~n6354 ;
  assign n6356 = n3450 & n6355 ;
  assign n6357 = ~n6344 & ~n6356 ;
  assign n6358 = n1898 & ~n6357 ;
  assign n6345 = n1800 & ~n4994 ;
  assign n6346 = ~n1800 & n4994 ;
  assign n6347 = ~n6345 & ~n6346 ;
  assign n6348 = n3450 & n6347 ;
  assign n6349 = ~n6344 & ~n6348 ;
  assign n6350 = n3575 & ~n6349 ;
  assign n6359 = ~n5025 & n5032 ;
  assign n6360 = n1800 & n6359 ;
  assign n6361 = ~n1800 & ~n6359 ;
  assign n6362 = ~n6360 & ~n6361 ;
  assign n6363 = n3450 & n6362 ;
  assign n6364 = ~n6344 & ~n6363 ;
  assign n6365 = n3557 & ~n6364 ;
  assign n6366 = n1015 & n3621 ;
  assign n6367 = n4837 & n6366 ;
  assign n6368 = ~n638 & ~n6367 ;
  assign n6369 = ~n5419 & ~n6368 ;
  assign n6370 = n3650 & n6369 ;
  assign n6371 = n3450 & n6370 ;
  assign n6343 = n688 & ~n3618 ;
  assign n6372 = ~n638 & n3655 ;
  assign n6373 = ~n6343 & ~n6372 ;
  assign n6374 = ~n6371 & n6373 ;
  assign n6375 = ~n6365 & n6374 ;
  assign n6376 = ~n6350 & n6375 ;
  assign n6377 = ~n6358 & n6376 ;
  assign n6378 = n3662 & ~n6377 ;
  assign n6379 = ~n6342 & ~n6378 ;
  assign n6380 = \P1_state_reg[0]/NET0131  & ~n6379 ;
  assign n6340 = n688 & n1934 ;
  assign n6341 = \P1_reg3_reg[19]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6381 = ~n6340 & ~n6341 ;
  assign n6382 = ~n6380 & n6381 ;
  assign n6385 = n2931 & ~n4925 ;
  assign n6386 = n4142 & ~n5109 ;
  assign n6387 = ~n4142 & n5109 ;
  assign n6388 = ~n6386 & ~n6387 ;
  assign n6389 = n4925 & ~n6388 ;
  assign n6390 = ~n6385 & ~n6389 ;
  assign n6391 = n3319 & ~n6390 ;
  assign n6392 = ~n3105 & n3342 ;
  assign n6393 = n3105 & ~n3342 ;
  assign n6394 = ~n6392 & ~n6393 ;
  assign n6395 = ~n2050 & ~n6394 ;
  assign n6396 = n2050 & n2911 ;
  assign n6397 = ~n6395 & ~n6396 ;
  assign n6398 = n4925 & n6397 ;
  assign n6399 = ~n6385 & ~n6398 ;
  assign n6400 = n3373 & ~n6399 ;
  assign n6401 = n4142 & ~n5157 ;
  assign n6402 = ~n4142 & n5157 ;
  assign n6403 = ~n6401 & ~n6402 ;
  assign n6404 = n4925 & n6403 ;
  assign n6405 = ~n6385 & ~n6404 ;
  assign n6406 = n3179 & ~n6405 ;
  assign n6407 = n2954 & ~n3387 ;
  assign n6408 = ~n2954 & n3387 ;
  assign n6409 = n3409 & ~n6408 ;
  assign n6410 = ~n6407 & n6409 ;
  assign n6411 = n4925 & n6410 ;
  assign n6384 = n2931 & n4934 ;
  assign n6412 = n2954 & ~n5093 ;
  assign n6413 = ~n6384 & ~n6412 ;
  assign n6414 = ~n6411 & n6413 ;
  assign n6415 = ~n6406 & n6414 ;
  assign n6416 = ~n6400 & n6415 ;
  assign n6417 = ~n6391 & n6416 ;
  assign n6418 = n2017 & ~n6417 ;
  assign n6419 = n2931 & n3430 ;
  assign n6420 = ~n6418 & ~n6419 ;
  assign n6421 = \P1_state_reg[0]/NET0131  & ~n6420 ;
  assign n6383 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[12]/NET0131  ;
  assign n6422 = n2931 & n3935 ;
  assign n6423 = ~n6383 & ~n6422 ;
  assign n6424 = ~n6421 & n6423 ;
  assign n6427 = n3042 & n3430 ;
  assign n6429 = n3042 & ~n4925 ;
  assign n6430 = ~n3046 & n5821 ;
  assign n6431 = n2640 & ~n6430 ;
  assign n6432 = ~n5822 & ~n6431 ;
  assign n6433 = ~n2050 & ~n6432 ;
  assign n6434 = n2050 & n3056 ;
  assign n6435 = ~n6433 & ~n6434 ;
  assign n6436 = n4925 & n6435 ;
  assign n6437 = ~n6429 & ~n6436 ;
  assign n6438 = n3373 & ~n6437 ;
  assign n6447 = ~n4109 & n4131 ;
  assign n6448 = n4109 & ~n4131 ;
  assign n6449 = ~n6447 & ~n6448 ;
  assign n6450 = n4925 & ~n6449 ;
  assign n6451 = ~n6429 & ~n6450 ;
  assign n6452 = n3319 & ~n6451 ;
  assign n6453 = ~n3095 & n3389 ;
  assign n6454 = ~n3071 & n6453 ;
  assign n6455 = n3036 & ~n6454 ;
  assign n6456 = ~n5846 & ~n6455 ;
  assign n6457 = n4925 & n6456 ;
  assign n6458 = ~n6429 & ~n6457 ;
  assign n6459 = n3409 & ~n6458 ;
  assign n6439 = ~n5157 & n5160 ;
  assign n6440 = n5171 & ~n6439 ;
  assign n6441 = n4131 & n6440 ;
  assign n6442 = ~n4131 & ~n6440 ;
  assign n6443 = ~n6441 & ~n6442 ;
  assign n6444 = n4925 & ~n6443 ;
  assign n6445 = ~n6429 & ~n6444 ;
  assign n6446 = n3179 & ~n6445 ;
  assign n6428 = n3036 & ~n5093 ;
  assign n6460 = n3042 & n5090 ;
  assign n6461 = ~n6428 & ~n6460 ;
  assign n6462 = ~n6446 & n6461 ;
  assign n6463 = ~n6459 & n6462 ;
  assign n6464 = ~n6452 & n6463 ;
  assign n6465 = ~n6438 & n6464 ;
  assign n6466 = n2017 & ~n6465 ;
  assign n6467 = ~n6427 & ~n6466 ;
  assign n6468 = \P1_state_reg[0]/NET0131  & ~n6467 ;
  assign n6425 = n3042 & n3935 ;
  assign n6426 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[16]/NET0131  ;
  assign n6469 = ~n6425 & ~n6426 ;
  assign n6470 = ~n6468 & n6469 ;
  assign n6472 = n1158 & n3664 ;
  assign n6474 = n1158 & ~n3450 ;
  assign n6475 = n1138 & ~n3586 ;
  assign n6476 = ~n3587 & ~n6475 ;
  assign n6477 = ~n536 & ~n6476 ;
  assign n6478 = n536 & n1189 ;
  assign n6479 = ~n6477 & ~n6478 ;
  assign n6480 = n3450 & n6479 ;
  assign n6481 = ~n6474 & ~n6480 ;
  assign n6482 = n1898 & ~n6481 ;
  assign n6483 = n1749 & ~n4552 ;
  assign n6484 = ~n1749 & n4552 ;
  assign n6485 = ~n6483 & ~n6484 ;
  assign n6486 = n3450 & n6485 ;
  assign n6487 = ~n6474 & ~n6486 ;
  assign n6488 = n3557 & ~n6487 ;
  assign n6489 = n1749 & ~n3833 ;
  assign n6490 = ~n1749 & n3833 ;
  assign n6491 = ~n6489 & ~n6490 ;
  assign n6492 = n3450 & ~n6491 ;
  assign n6493 = ~n6474 & ~n6492 ;
  assign n6494 = n3575 & ~n6493 ;
  assign n6495 = n1202 & n3632 ;
  assign n6496 = ~n1178 & ~n6495 ;
  assign n6497 = ~n3634 & n3650 ;
  assign n6498 = ~n6496 & n6497 ;
  assign n6499 = n3450 & n6498 ;
  assign n6473 = n1158 & ~n3618 ;
  assign n6500 = ~n1178 & n3655 ;
  assign n6501 = ~n6473 & ~n6500 ;
  assign n6502 = ~n6499 & n6501 ;
  assign n6503 = ~n6494 & n6502 ;
  assign n6504 = ~n6488 & n6503 ;
  assign n6505 = ~n6482 & n6504 ;
  assign n6506 = n3662 & ~n6505 ;
  assign n6507 = ~n6472 & ~n6506 ;
  assign n6508 = \P1_state_reg[0]/NET0131  & ~n6507 ;
  assign n6471 = \P1_reg3_reg[9]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6509 = n1158 & n1934 ;
  assign n6510 = ~n6471 & ~n6509 ;
  assign n6511 = ~n6508 & n6510 ;
  assign n6512 = \P2_reg2_reg[18]/NET0131  & ~n3434 ;
  assign n6513 = \P2_reg2_reg[18]/NET0131  & n3430 ;
  assign n6515 = \P2_reg2_reg[18]/NET0131  & ~n2033 ;
  assign n6516 = n2033 & n5874 ;
  assign n6517 = ~n6515 & ~n6516 ;
  assign n6518 = n3373 & ~n6517 ;
  assign n6519 = n2033 & n5880 ;
  assign n6520 = ~n6515 & ~n6519 ;
  assign n6521 = n3179 & ~n6520 ;
  assign n6522 = n2033 & ~n5886 ;
  assign n6523 = ~n6515 & ~n6522 ;
  assign n6524 = n3319 & ~n6523 ;
  assign n6525 = n2033 & n5892 ;
  assign n6526 = ~n6515 & ~n6525 ;
  assign n6527 = n3409 & ~n6526 ;
  assign n6528 = n2033 & n2657 ;
  assign n6529 = ~n6515 & ~n6528 ;
  assign n6530 = n3375 & ~n6529 ;
  assign n6514 = n2662 & n3415 ;
  assign n6531 = \P2_reg2_reg[18]/NET0131  & n3418 ;
  assign n6532 = ~n6514 & ~n6531 ;
  assign n6533 = ~n6530 & n6532 ;
  assign n6534 = ~n6527 & n6533 ;
  assign n6535 = ~n6524 & n6534 ;
  assign n6536 = ~n6521 & n6535 ;
  assign n6537 = ~n6518 & n6536 ;
  assign n6538 = n2017 & ~n6537 ;
  assign n6539 = ~n6513 & ~n6538 ;
  assign n6540 = \P1_state_reg[0]/NET0131  & ~n6539 ;
  assign n6541 = ~n6512 & ~n6540 ;
  assign n6542 = n945 & n3664 ;
  assign n6546 = ~n6189 & n6199 ;
  assign n6547 = ~n6185 & n6546 ;
  assign n6548 = n3450 & ~n6547 ;
  assign n6543 = n939 & n3655 ;
  assign n6544 = ~n3615 & ~n3653 ;
  assign n6545 = n945 & ~n6544 ;
  assign n6549 = ~n6543 & ~n6545 ;
  assign n6550 = ~n6548 & n6549 ;
  assign n6551 = n3662 & ~n6550 ;
  assign n6552 = ~n6542 & ~n6551 ;
  assign n6553 = \P1_state_reg[0]/NET0131  & ~n6552 ;
  assign n6554 = n945 & n1934 ;
  assign n6555 = \P1_reg3_reg[21]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6556 = ~n6554 & ~n6555 ;
  assign n6557 = ~n6553 & n6556 ;
  assign n6558 = n883 & n3664 ;
  assign n6559 = n883 & ~n3450 ;
  assign n6560 = n4488 & ~n5780 ;
  assign n6561 = n4487 & ~n6560 ;
  assign n6562 = n1779 & n6561 ;
  assign n6563 = ~n1779 & ~n6561 ;
  assign n6564 = ~n6562 & ~n6563 ;
  assign n6565 = n3450 & ~n6564 ;
  assign n6566 = ~n6559 & ~n6565 ;
  assign n6567 = n3557 & ~n6566 ;
  assign n6568 = n4466 & n4469 ;
  assign n6569 = ~n4453 & n4469 ;
  assign n6570 = n4474 & ~n6569 ;
  assign n6571 = ~n6568 & n6570 ;
  assign n6572 = n1779 & ~n6571 ;
  assign n6573 = ~n1779 & n6571 ;
  assign n6574 = ~n6572 & ~n6573 ;
  assign n6575 = n3450 & ~n6574 ;
  assign n6576 = ~n6559 & ~n6575 ;
  assign n6577 = n3575 & ~n6576 ;
  assign n6579 = n536 & ~n949 ;
  assign n6580 = n921 & ~n6180 ;
  assign n6581 = ~n536 & ~n4285 ;
  assign n6582 = ~n6580 & n6581 ;
  assign n6583 = ~n6579 & ~n6582 ;
  assign n6584 = n1898 & ~n6583 ;
  assign n6585 = n875 & ~n6187 ;
  assign n6586 = ~n3641 & n3650 ;
  assign n6587 = ~n6585 & n6586 ;
  assign n6588 = ~n6584 & ~n6587 ;
  assign n6589 = n3450 & ~n6588 ;
  assign n6578 = n875 & n3655 ;
  assign n6590 = n1898 & ~n3450 ;
  assign n6591 = n4591 & ~n6590 ;
  assign n6592 = n883 & ~n6591 ;
  assign n6593 = ~n6578 & ~n6592 ;
  assign n6594 = ~n6589 & n6593 ;
  assign n6595 = ~n6577 & n6594 ;
  assign n6596 = ~n6567 & n6595 ;
  assign n6597 = n3662 & ~n6596 ;
  assign n6598 = ~n6558 & ~n6597 ;
  assign n6599 = \P1_state_reg[0]/NET0131  & ~n6598 ;
  assign n6600 = \P1_reg3_reg[22]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6601 = n883 & n1934 ;
  assign n6602 = ~n6600 & ~n6601 ;
  assign n6603 = ~n6599 & n6602 ;
  assign n6604 = n2527 & n3430 ;
  assign n6605 = n2527 & ~n4925 ;
  assign n6606 = n4925 & ~n6026 ;
  assign n6607 = ~n6605 & ~n6606 ;
  assign n6608 = n3179 & ~n6607 ;
  assign n6609 = n4925 & ~n6039 ;
  assign n6610 = ~n6605 & ~n6609 ;
  assign n6611 = n3319 & ~n6610 ;
  assign n6613 = n4925 & ~n6051 ;
  assign n6614 = ~n6605 & ~n6613 ;
  assign n6615 = n3373 & ~n6614 ;
  assign n6616 = n4925 & n6057 ;
  assign n6612 = n2527 & n4934 ;
  assign n6617 = n2522 & ~n5093 ;
  assign n6618 = ~n6612 & ~n6617 ;
  assign n6619 = ~n6616 & n6618 ;
  assign n6620 = ~n6615 & n6619 ;
  assign n6621 = ~n6611 & n6620 ;
  assign n6622 = ~n6608 & n6621 ;
  assign n6623 = n2017 & ~n6622 ;
  assign n6624 = ~n6604 & ~n6623 ;
  assign n6625 = \P1_state_reg[0]/NET0131  & ~n6624 ;
  assign n6626 = n2527 & n3935 ;
  assign n6627 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[22]/NET0131  ;
  assign n6628 = ~n6626 & ~n6627 ;
  assign n6629 = ~n6625 & n6628 ;
  assign n6630 = \P1_reg2_reg[12]/NET0131  & ~n6072 ;
  assign n6631 = n1068 & n1736 ;
  assign n6632 = ~n1094 & n3683 ;
  assign n6633 = n5759 & ~n6632 ;
  assign n6634 = n3672 & ~n6633 ;
  assign n6635 = ~n6631 & ~n6634 ;
  assign n6636 = n6070 & ~n6635 ;
  assign n6637 = ~n6630 & ~n6636 ;
  assign n6638 = \P1_reg2_reg[18]/NET0131  & ~n3703 ;
  assign n6639 = \P1_reg2_reg[18]/NET0131  & n3664 ;
  assign n6643 = \P1_reg2_reg[18]/NET0131  & ~n3672 ;
  assign n6647 = n3672 & ~n5789 ;
  assign n6648 = ~n6643 & ~n6647 ;
  assign n6649 = n3575 & ~n6648 ;
  assign n6644 = n3672 & n5783 ;
  assign n6645 = ~n6643 & ~n6644 ;
  assign n6646 = n3557 & ~n6645 ;
  assign n6650 = n3672 & n5798 ;
  assign n6651 = ~n6643 & ~n6650 ;
  assign n6652 = n1898 & ~n6651 ;
  assign n6640 = ~n743 & n3683 ;
  assign n6641 = ~n5805 & ~n6640 ;
  assign n6642 = n3672 & ~n6641 ;
  assign n6653 = \P1_reg2_reg[18]/NET0131  & ~n5452 ;
  assign n6654 = n748 & n1736 ;
  assign n6655 = ~n6653 & ~n6654 ;
  assign n6656 = ~n6642 & n6655 ;
  assign n6657 = ~n6652 & n6656 ;
  assign n6658 = ~n6646 & n6657 ;
  assign n6659 = ~n6649 & n6658 ;
  assign n6660 = n3662 & ~n6659 ;
  assign n6661 = ~n6639 & ~n6660 ;
  assign n6662 = \P1_state_reg[0]/NET0131  & ~n6661 ;
  assign n6663 = ~n6638 & ~n6662 ;
  assign n6664 = \P1_reg2_reg[21]/NET0131  & ~n3703 ;
  assign n6665 = \P1_reg2_reg[21]/NET0131  & n3664 ;
  assign n6666 = ~n6185 & n6200 ;
  assign n6667 = n3672 & ~n6666 ;
  assign n6670 = n3672 & ~n6188 ;
  assign n6671 = ~\P1_reg2_reg[21]/NET0131  & ~n3672 ;
  assign n6672 = n3650 & ~n6671 ;
  assign n6673 = ~n6670 & n6672 ;
  assign n6668 = n945 & n1736 ;
  assign n6669 = \P1_reg2_reg[21]/NET0131  & ~n4857 ;
  assign n6674 = ~n6668 & ~n6669 ;
  assign n6675 = ~n6673 & n6674 ;
  assign n6676 = ~n6667 & n6675 ;
  assign n6677 = n3662 & ~n6676 ;
  assign n6678 = ~n6665 & ~n6677 ;
  assign n6679 = \P1_state_reg[0]/NET0131  & ~n6678 ;
  assign n6680 = ~n6664 & ~n6679 ;
  assign n6681 = \P1_reg2_reg[22]/NET0131  & ~n3703 ;
  assign n6682 = \P1_reg2_reg[22]/NET0131  & n3664 ;
  assign n6683 = \P1_reg2_reg[22]/NET0131  & ~n3672 ;
  assign n6684 = n3672 & ~n6564 ;
  assign n6685 = ~n6683 & ~n6684 ;
  assign n6686 = n3557 & ~n6685 ;
  assign n6687 = n3672 & ~n6574 ;
  assign n6688 = ~n6683 & ~n6687 ;
  assign n6689 = n3575 & ~n6688 ;
  assign n6690 = n875 & n3683 ;
  assign n6691 = n6588 & ~n6690 ;
  assign n6692 = n3672 & ~n6691 ;
  assign n6693 = ~n3672 & n4704 ;
  assign n6694 = n3685 & ~n6693 ;
  assign n6695 = \P1_reg2_reg[22]/NET0131  & ~n6694 ;
  assign n6696 = n883 & n1736 ;
  assign n6697 = ~n6695 & ~n6696 ;
  assign n6698 = ~n6692 & n6697 ;
  assign n6699 = ~n6689 & n6698 ;
  assign n6700 = ~n6686 & n6699 ;
  assign n6701 = n3662 & ~n6700 ;
  assign n6702 = ~n6682 & ~n6701 ;
  assign n6703 = \P1_state_reg[0]/NET0131  & ~n6702 ;
  assign n6704 = ~n6681 & ~n6703 ;
  assign n6706 = n3373 & n5828 ;
  assign n6708 = n3179 & ~n5834 ;
  assign n6707 = n3319 & n5842 ;
  assign n6705 = n3409 & n5849 ;
  assign n6709 = n2630 & n3375 ;
  assign n6710 = ~n6705 & ~n6709 ;
  assign n6711 = ~n6707 & n6710 ;
  assign n6712 = ~n6708 & n6711 ;
  assign n6713 = ~n6706 & n6712 ;
  assign n6714 = n5572 & ~n6713 ;
  assign n6718 = n3319 & ~n4663 ;
  assign n6719 = n5509 & ~n6718 ;
  assign n6715 = n3175 & ~n3177 ;
  assign n6716 = ~n4663 & n6715 ;
  assign n6717 = ~n3176 & n6716 ;
  assign n6720 = ~n5510 & ~n6717 ;
  assign n6721 = n6719 & n6720 ;
  assign n6722 = n4275 & n6721 ;
  assign n6723 = \P2_reg1_reg[17]/NET0131  & ~n6722 ;
  assign n6724 = ~n6714 & ~n6723 ;
  assign n6725 = \P2_reg1_reg[18]/NET0131  & ~n3434 ;
  assign n6726 = \P2_reg1_reg[18]/NET0131  & n3430 ;
  assign n6732 = \P2_reg1_reg[18]/NET0131  & ~n4663 ;
  assign n6733 = n4663 & n5874 ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6735 = n3373 & ~n6734 ;
  assign n6736 = n4663 & n5880 ;
  assign n6737 = ~n6732 & ~n6736 ;
  assign n6738 = n3179 & ~n6737 ;
  assign n6728 = n3319 & ~n5886 ;
  assign n6727 = n2657 & n3375 ;
  assign n6729 = ~n5893 & ~n6727 ;
  assign n6730 = ~n6728 & n6729 ;
  assign n6731 = n4663 & ~n6730 ;
  assign n6739 = \P2_reg1_reg[18]/NET0131  & ~n6719 ;
  assign n6740 = ~n6731 & ~n6739 ;
  assign n6741 = ~n6738 & n6740 ;
  assign n6742 = ~n6735 & n6741 ;
  assign n6743 = n2017 & ~n6742 ;
  assign n6744 = ~n6726 & ~n6743 ;
  assign n6745 = \P1_state_reg[0]/NET0131  & ~n6744 ;
  assign n6746 = ~n6725 & ~n6745 ;
  assign n6747 = ~n2016 & ~n6716 ;
  assign n6748 = n6719 & n6747 ;
  assign n6749 = n3434 & n6748 ;
  assign n6750 = \P2_reg1_reg[19]/NET0131  & ~n6749 ;
  assign n6752 = n3373 & ~n5915 ;
  assign n6751 = n2604 & n3375 ;
  assign n6753 = n5933 & ~n6751 ;
  assign n6754 = ~n6752 & n6753 ;
  assign n6755 = n5572 & ~n6754 ;
  assign n6756 = ~n6750 & ~n6755 ;
  assign n6757 = \P2_reg1_reg[22]/NET0131  & ~n3434 ;
  assign n6758 = \P2_reg1_reg[22]/NET0131  & n3430 ;
  assign n6759 = \P2_reg1_reg[22]/NET0131  & ~n4663 ;
  assign n6760 = n4663 & ~n6026 ;
  assign n6761 = ~n6759 & ~n6760 ;
  assign n6762 = n3179 & ~n6761 ;
  assign n6763 = n4663 & ~n6039 ;
  assign n6764 = ~n6759 & ~n6763 ;
  assign n6765 = n3319 & ~n6764 ;
  assign n6766 = n4663 & ~n6059 ;
  assign n6767 = \P2_reg1_reg[22]/NET0131  & ~n5511 ;
  assign n6768 = ~n6766 & ~n6767 ;
  assign n6769 = ~n6765 & n6768 ;
  assign n6770 = ~n6762 & n6769 ;
  assign n6771 = n2017 & ~n6770 ;
  assign n6772 = ~n6758 & ~n6771 ;
  assign n6773 = \P1_state_reg[0]/NET0131  & ~n6772 ;
  assign n6774 = ~n6757 & ~n6773 ;
  assign n6775 = \P1_reg0_reg[12]/NET0131  & ~n6169 ;
  assign n6776 = n6171 & ~n6633 ;
  assign n6777 = ~n6775 & ~n6776 ;
  assign n6780 = ~n1696 & n3879 ;
  assign n6779 = n1696 & ~n3879 ;
  assign n6781 = n3650 & ~n6779 ;
  assign n6782 = ~n6780 & n6781 ;
  assign n6778 = n1696 & n3683 ;
  assign n6783 = ~n4853 & ~n6778 ;
  assign n6784 = ~n6782 & n6783 ;
  assign n6785 = n3672 & ~n6784 ;
  assign n6786 = ~n3887 & ~n6785 ;
  assign n6787 = n6070 & ~n6786 ;
  assign n6788 = ~n1736 & ~n3672 ;
  assign n6789 = ~n3615 & n6070 ;
  assign n6790 = ~n6788 & n6789 ;
  assign n6791 = \P1_reg2_reg[30]/NET0131  & ~n6790 ;
  assign n6792 = ~n6787 & ~n6791 ;
  assign n6793 = ~n2033 & n3179 ;
  assign n6794 = ~n2033 & n3319 ;
  assign n6795 = ~n6793 & ~n6794 ;
  assign n6796 = n4437 & n6795 ;
  assign n6797 = n4275 & n6796 ;
  assign n6798 = \P2_reg2_reg[17]/NET0131  & ~n6797 ;
  assign n6799 = n2033 & ~n6713 ;
  assign n6800 = n2636 & n3415 ;
  assign n6801 = ~n6799 & ~n6800 ;
  assign n6802 = n4275 & ~n6801 ;
  assign n6803 = ~n6798 & ~n6802 ;
  assign n6804 = n2033 & ~n6754 ;
  assign n6805 = n2609 & n3415 ;
  assign n6806 = ~n6804 & ~n6805 ;
  assign n6807 = n4275 & ~n6806 ;
  assign n6808 = ~n2033 & ~n5387 ;
  assign n6809 = n4275 & ~n6808 ;
  assign n6810 = ~n4434 & n6809 ;
  assign n6811 = \P2_reg2_reg[19]/NET0131  & ~n6810 ;
  assign n6812 = ~n6807 & ~n6811 ;
  assign n6813 = \P2_reg2_reg[20]/NET0131  & ~n3434 ;
  assign n6814 = \P2_reg2_reg[20]/NET0131  & n3430 ;
  assign n6816 = \P2_reg2_reg[20]/NET0131  & ~n2033 ;
  assign n6823 = n4140 & n5114 ;
  assign n6824 = ~n4140 & ~n5114 ;
  assign n6825 = ~n6823 & ~n6824 ;
  assign n6826 = n2033 & n6825 ;
  assign n6827 = ~n6816 & ~n6826 ;
  assign n6828 = n3319 & ~n6827 ;
  assign n6817 = n3392 & n5846 ;
  assign n6818 = n2579 & ~n5928 ;
  assign n6819 = ~n6817 & ~n6818 ;
  assign n6820 = n2033 & n6819 ;
  assign n6821 = ~n6816 & ~n6820 ;
  assign n6822 = n3409 & ~n6821 ;
  assign n6829 = n2551 & ~n5911 ;
  assign n6830 = ~n6046 & ~n6829 ;
  assign n6831 = ~n2050 & ~n6830 ;
  assign n6832 = n2050 & n2613 ;
  assign n6833 = ~n6831 & ~n6832 ;
  assign n6834 = n2033 & n6833 ;
  assign n6835 = ~n6816 & ~n6834 ;
  assign n6836 = n3373 & ~n6835 ;
  assign n6837 = n2579 & n3375 ;
  assign n6839 = ~n4140 & n5180 ;
  assign n6838 = n4140 & ~n5180 ;
  assign n6840 = n3179 & ~n6838 ;
  assign n6841 = ~n6839 & n6840 ;
  assign n6842 = ~n6837 & ~n6841 ;
  assign n6843 = n2033 & ~n6842 ;
  assign n6815 = n2584 & n3415 ;
  assign n6844 = ~n4434 & ~n6793 ;
  assign n6845 = \P2_reg2_reg[20]/NET0131  & ~n6844 ;
  assign n6846 = ~n6815 & ~n6845 ;
  assign n6847 = ~n6843 & n6846 ;
  assign n6848 = ~n6836 & n6847 ;
  assign n6849 = ~n6822 & n6848 ;
  assign n6850 = ~n6828 & n6849 ;
  assign n6851 = n2017 & ~n6850 ;
  assign n6852 = ~n6814 & ~n6851 ;
  assign n6853 = \P1_state_reg[0]/NET0131  & ~n6852 ;
  assign n6854 = ~n6813 & ~n6853 ;
  assign n6856 = \P1_reg0_reg[17]/NET0131  & ~n3900 ;
  assign n6857 = n5969 & n6171 ;
  assign n6858 = ~n6856 & ~n6857 ;
  assign n6859 = n1898 & ~n6858 ;
  assign n6855 = n6171 & ~n6257 ;
  assign n6860 = ~n4724 & n6070 ;
  assign n6861 = ~n1897 & n5643 ;
  assign n6862 = n6860 & ~n6861 ;
  assign n6863 = n4723 & n6862 ;
  assign n6864 = \P1_reg0_reg[17]/NET0131  & ~n6863 ;
  assign n6865 = ~n6855 & ~n6864 ;
  assign n6866 = ~n6859 & n6865 ;
  assign n6867 = \P1_reg0_reg[20]/NET0131  & ~n3703 ;
  assign n6869 = n1898 & n5403 ;
  assign n6868 = n3557 & n5409 ;
  assign n6870 = n5425 & ~n6868 ;
  assign n6871 = ~n6869 & n6870 ;
  assign n6872 = n3662 & n3900 ;
  assign n6873 = ~n6871 & n6872 ;
  assign n6874 = ~n1951 & n6168 ;
  assign n6875 = \P1_reg0_reg[20]/NET0131  & ~n1933 ;
  assign n6876 = ~n6874 & n6875 ;
  assign n6877 = ~n6873 & ~n6876 ;
  assign n6878 = \P1_state_reg[0]/NET0131  & ~n6877 ;
  assign n6879 = ~n6867 & ~n6878 ;
  assign n6880 = \P1_reg0_reg[30]/NET0131  & ~n6238 ;
  assign n6881 = n6171 & ~n6784 ;
  assign n6882 = ~n6880 & ~n6881 ;
  assign n6883 = \P1_reg1_reg[12]/NET0131  & ~n6244 ;
  assign n6884 = n6246 & ~n6633 ;
  assign n6885 = ~n6883 & ~n6884 ;
  assign n6886 = \P1_reg1_reg[20]/NET0131  & ~n3703 ;
  assign n6887 = \P1_reg1_reg[20]/NET0131  & n3664 ;
  assign n6888 = n3616 & ~n4236 ;
  assign n6889 = n3915 & ~n6888 ;
  assign n6890 = ~n6241 & n6889 ;
  assign n6891 = ~n4756 & n6890 ;
  assign n6892 = \P1_reg1_reg[20]/NET0131  & ~n6891 ;
  assign n6893 = n4236 & ~n6871 ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = n3662 & ~n6894 ;
  assign n6896 = ~n6887 & ~n6895 ;
  assign n6897 = \P1_state_reg[0]/NET0131  & ~n6896 ;
  assign n6898 = ~n6886 & ~n6897 ;
  assign n6899 = n5385 & ~n6713 ;
  assign n6900 = n3319 & ~n4610 ;
  assign n6901 = n4621 & ~n6900 ;
  assign n6902 = ~n4610 & n6715 ;
  assign n6903 = n4275 & ~n6902 ;
  assign n6904 = n6901 & n6903 ;
  assign n6905 = \P2_reg0_reg[17]/NET0131  & ~n6904 ;
  assign n6906 = ~n6899 & ~n6905 ;
  assign n6907 = \P2_reg0_reg[18]/NET0131  & ~n3434 ;
  assign n6908 = \P2_reg0_reg[18]/NET0131  & n3430 ;
  assign n6910 = \P2_reg0_reg[18]/NET0131  & ~n4610 ;
  assign n6911 = n4610 & n5874 ;
  assign n6912 = ~n6910 & ~n6911 ;
  assign n6913 = n3373 & ~n6912 ;
  assign n6914 = n4610 & n5880 ;
  assign n6915 = ~n6910 & ~n6914 ;
  assign n6916 = n3179 & ~n6915 ;
  assign n6909 = n4610 & ~n6730 ;
  assign n6917 = \P2_reg0_reg[18]/NET0131  & ~n6901 ;
  assign n6918 = ~n6909 & ~n6917 ;
  assign n6919 = ~n6916 & n6918 ;
  assign n6920 = ~n6913 & n6919 ;
  assign n6921 = n2017 & ~n6920 ;
  assign n6922 = ~n6908 & ~n6921 ;
  assign n6923 = \P1_state_reg[0]/NET0131  & ~n6922 ;
  assign n6924 = ~n6907 & ~n6923 ;
  assign n6925 = \P1_reg1_reg[30]/NET0131  & ~n6311 ;
  assign n6926 = n6246 & ~n6784 ;
  assign n6927 = ~n6925 & ~n6926 ;
  assign n6928 = n5385 & ~n6754 ;
  assign n6929 = \P2_reg0_reg[19]/NET0131  & ~n6904 ;
  assign n6930 = ~n6928 & ~n6929 ;
  assign n6933 = n1111 & n3664 ;
  assign n6937 = n1111 & ~n3450 ;
  assign n6938 = n1075 & ~n5738 ;
  assign n6939 = ~n5739 & ~n6938 ;
  assign n6940 = ~n536 & ~n6939 ;
  assign n6941 = n536 & n1138 ;
  assign n6942 = ~n6940 & ~n6941 ;
  assign n6943 = n3450 & n6942 ;
  assign n6944 = ~n6937 & ~n6943 ;
  assign n6945 = n1898 & ~n6944 ;
  assign n6946 = n1750 & ~n5021 ;
  assign n6947 = ~n1750 & n5021 ;
  assign n6948 = ~n6946 & ~n6947 ;
  assign n6949 = n3450 & ~n6948 ;
  assign n6950 = ~n6937 & ~n6949 ;
  assign n6951 = n3557 & ~n6950 ;
  assign n6958 = n1750 & ~n4984 ;
  assign n6957 = ~n1750 & n4984 ;
  assign n6959 = n3575 & ~n6957 ;
  assign n6960 = ~n6958 & n6959 ;
  assign n6952 = ~n1128 & n3683 ;
  assign n6953 = n1151 & n3634 ;
  assign n6954 = ~n1128 & ~n6953 ;
  assign n6955 = ~n3636 & n3650 ;
  assign n6956 = ~n6954 & n6955 ;
  assign n6961 = ~n6952 & ~n6956 ;
  assign n6962 = ~n6960 & n6961 ;
  assign n6963 = n3450 & ~n6962 ;
  assign n6934 = ~n1128 & n1736 ;
  assign n6935 = n3618 & ~n4819 ;
  assign n6936 = n1111 & ~n6935 ;
  assign n6964 = ~n6934 & ~n6936 ;
  assign n6965 = ~n6963 & n6964 ;
  assign n6966 = ~n6951 & n6965 ;
  assign n6967 = ~n6945 & n6966 ;
  assign n6968 = n3662 & ~n6967 ;
  assign n6969 = ~n6933 & ~n6968 ;
  assign n6970 = \P1_state_reg[0]/NET0131  & ~n6969 ;
  assign n6931 = \P1_reg3_reg[11]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6932 = n1111 & n1934 ;
  assign n6971 = ~n6931 & ~n6932 ;
  assign n6972 = ~n6970 & n6971 ;
  assign n6975 = n1132 & n3664 ;
  assign n6982 = n1132 & ~n3450 ;
  assign n6983 = n1115 & ~n3587 ;
  assign n6984 = ~n5738 & ~n6983 ;
  assign n6985 = ~n536 & ~n6984 ;
  assign n6986 = n536 & n1162 ;
  assign n6987 = ~n6985 & ~n6986 ;
  assign n6988 = n3450 & n6987 ;
  assign n6989 = ~n6982 & ~n6988 ;
  assign n6990 = n1898 & ~n6989 ;
  assign n6997 = n1754 & ~n4504 ;
  assign n6998 = ~n1754 & n4504 ;
  assign n6999 = ~n6997 & ~n6998 ;
  assign n7000 = n3450 & ~n6999 ;
  assign n7001 = ~n6982 & ~n7000 ;
  assign n7002 = n3557 & ~n7001 ;
  assign n6991 = n1754 & ~n4459 ;
  assign n6992 = ~n1754 & n4459 ;
  assign n6993 = ~n6991 & ~n6992 ;
  assign n6994 = n3450 & n6993 ;
  assign n6995 = ~n6982 & ~n6994 ;
  assign n6996 = n3575 & ~n6995 ;
  assign n6976 = ~n1151 & n3683 ;
  assign n6977 = n3650 & ~n6953 ;
  assign n6978 = ~n1151 & ~n3634 ;
  assign n6979 = n6977 & ~n6978 ;
  assign n6980 = ~n6976 & ~n6979 ;
  assign n6981 = n3450 & ~n6980 ;
  assign n7003 = ~n1151 & n1736 ;
  assign n7004 = n1132 & ~n3618 ;
  assign n7005 = ~n7003 & ~n7004 ;
  assign n7006 = ~n6981 & n7005 ;
  assign n7007 = ~n6996 & n7006 ;
  assign n7008 = ~n7002 & n7007 ;
  assign n7009 = ~n6990 & n7008 ;
  assign n7010 = n3662 & ~n7009 ;
  assign n7011 = ~n6975 & ~n7010 ;
  assign n7012 = \P1_state_reg[0]/NET0131  & ~n7011 ;
  assign n6973 = \P1_reg3_reg[10]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6974 = n1132 & n1934 ;
  assign n7013 = ~n6973 & ~n6974 ;
  assign n7014 = ~n7012 & n7013 ;
  assign n7016 = n1021 & n3664 ;
  assign n7036 = n3588 & n5739 ;
  assign n7037 = n999 & ~n7036 ;
  assign n7038 = ~n3592 & ~n7037 ;
  assign n7039 = ~n536 & ~n7038 ;
  assign n7040 = n536 & n1051 ;
  assign n7041 = ~n7039 & ~n7040 ;
  assign n7042 = n3450 & ~n7041 ;
  assign n7035 = ~n1021 & ~n3450 ;
  assign n7043 = n1898 & ~n7035 ;
  assign n7044 = ~n7042 & n7043 ;
  assign n7026 = ~n1756 & n4464 ;
  assign n7025 = n1756 & ~n4464 ;
  assign n7027 = n3575 & ~n7025 ;
  assign n7028 = ~n7026 & n7027 ;
  assign n7018 = ~n1040 & ~n4836 ;
  assign n7019 = n3650 & ~n4837 ;
  assign n7020 = ~n7018 & n7019 ;
  assign n7022 = ~n1756 & ~n5778 ;
  assign n7021 = n1756 & n5778 ;
  assign n7023 = n3557 & ~n7021 ;
  assign n7024 = ~n7022 & n7023 ;
  assign n7029 = ~n7020 & ~n7024 ;
  assign n7030 = ~n7028 & n7029 ;
  assign n7031 = n3450 & ~n7030 ;
  assign n7017 = ~n1040 & n3655 ;
  assign n7032 = ~n3450 & n3556 ;
  assign n7033 = n4591 & ~n7032 ;
  assign n7034 = n1021 & ~n7033 ;
  assign n7045 = ~n7017 & ~n7034 ;
  assign n7046 = ~n7031 & n7045 ;
  assign n7047 = ~n7044 & n7046 ;
  assign n7048 = n3662 & ~n7047 ;
  assign n7049 = ~n7016 & ~n7048 ;
  assign n7050 = \P1_state_reg[0]/NET0131  & ~n7049 ;
  assign n7015 = \P1_reg3_reg[14]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7051 = n1021 & n1934 ;
  assign n7052 = ~n7015 & ~n7051 ;
  assign n7053 = ~n7050 & n7052 ;
  assign n7056 = n994 & n3664 ;
  assign n7058 = n994 & ~n3450 ;
  assign n7059 = ~n5021 & n5023 ;
  assign n7060 = n5028 & ~n7059 ;
  assign n7061 = n1765 & ~n7060 ;
  assign n7062 = ~n1765 & n7060 ;
  assign n7063 = ~n7061 & ~n7062 ;
  assign n7064 = n3450 & n7063 ;
  assign n7065 = ~n7058 & ~n7064 ;
  assign n7066 = n3557 & ~n7065 ;
  assign n7075 = n1765 & ~n4989 ;
  assign n7076 = ~n1765 & n4989 ;
  assign n7077 = ~n7075 & ~n7076 ;
  assign n7078 = n3450 & ~n7077 ;
  assign n7079 = ~n7058 & ~n7078 ;
  assign n7080 = n3575 & ~n7079 ;
  assign n7067 = n838 & ~n3592 ;
  assign n7068 = ~n3593 & ~n7067 ;
  assign n7069 = ~n536 & ~n7068 ;
  assign n7070 = n536 & n1026 ;
  assign n7071 = ~n7069 & ~n7070 ;
  assign n7072 = n3450 & n7071 ;
  assign n7073 = ~n7058 & ~n7072 ;
  assign n7074 = n1898 & ~n7073 ;
  assign n7081 = ~n1015 & ~n4837 ;
  assign n7082 = ~n3640 & ~n7081 ;
  assign n7083 = n3450 & n7082 ;
  assign n7084 = ~n7058 & ~n7083 ;
  assign n7085 = n3650 & ~n7084 ;
  assign n7057 = ~n1015 & n3655 ;
  assign n7086 = n994 & ~n4305 ;
  assign n7087 = ~n7057 & ~n7086 ;
  assign n7088 = ~n7085 & n7087 ;
  assign n7089 = ~n7074 & n7088 ;
  assign n7090 = ~n7080 & n7089 ;
  assign n7091 = ~n7066 & n7090 ;
  assign n7092 = n3662 & ~n7091 ;
  assign n7093 = ~n7056 & ~n7092 ;
  assign n7094 = \P1_state_reg[0]/NET0131  & ~n7093 ;
  assign n7054 = \P1_reg3_reg[15]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7055 = n994 & n1934 ;
  assign n7095 = ~n7054 & ~n7055 ;
  assign n7096 = ~n7094 & n7095 ;
  assign n7099 = n2961 & n3430 ;
  assign n7101 = n2961 & ~n4925 ;
  assign n7108 = ~n2965 & n3339 ;
  assign n7109 = n2911 & ~n7108 ;
  assign n7110 = ~n2911 & n7108 ;
  assign n7111 = ~n7109 & ~n7110 ;
  assign n7112 = ~n2050 & ~n7111 ;
  assign n7113 = n2050 & n2990 ;
  assign n7114 = ~n7112 & ~n7113 ;
  assign n7115 = n4925 & n7114 ;
  assign n7116 = ~n7101 & ~n7115 ;
  assign n7117 = n3373 & ~n7116 ;
  assign n7102 = n4128 & ~n5306 ;
  assign n7103 = ~n4128 & n5306 ;
  assign n7104 = ~n7102 & ~n7103 ;
  assign n7105 = n4925 & ~n7104 ;
  assign n7106 = ~n7101 & ~n7105 ;
  assign n7107 = n3319 & ~n7106 ;
  assign n7118 = n4128 & ~n5278 ;
  assign n7119 = ~n4128 & n5278 ;
  assign n7120 = ~n7118 & ~n7119 ;
  assign n7121 = n4925 & n7120 ;
  assign n7122 = ~n7101 & ~n7121 ;
  assign n7123 = n3179 & ~n7122 ;
  assign n7124 = ~n3005 & n3384 ;
  assign n7126 = n2980 & ~n7124 ;
  assign n7125 = ~n2980 & n7124 ;
  assign n7127 = n3409 & ~n7125 ;
  assign n7128 = ~n7126 & n7127 ;
  assign n7129 = n4925 & n7128 ;
  assign n7100 = n2961 & n4934 ;
  assign n7130 = n2980 & ~n5093 ;
  assign n7131 = ~n7100 & ~n7130 ;
  assign n7132 = ~n7129 & n7131 ;
  assign n7133 = ~n7123 & n7132 ;
  assign n7134 = ~n7107 & n7133 ;
  assign n7135 = ~n7117 & n7134 ;
  assign n7136 = n2017 & ~n7135 ;
  assign n7137 = ~n7099 & ~n7136 ;
  assign n7138 = \P1_state_reg[0]/NET0131  & ~n7137 ;
  assign n7097 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[10]/NET0131  ;
  assign n7098 = n2961 & n3935 ;
  assign n7139 = ~n7097 & ~n7098 ;
  assign n7140 = ~n7138 & n7139 ;
  assign n7143 = n3099 & n3430 ;
  assign n7151 = n3099 & ~n4925 ;
  assign n7152 = n3082 & ~n6392 ;
  assign n7153 = ~n3344 & ~n7152 ;
  assign n7154 = ~n2050 & ~n7153 ;
  assign n7155 = n2050 & n2937 ;
  assign n7156 = ~n7154 & ~n7155 ;
  assign n7157 = n4925 & n7156 ;
  assign n7158 = ~n7151 & ~n7157 ;
  assign n7159 = n3373 & ~n7158 ;
  assign n7160 = ~n3119 & ~n3125 ;
  assign n7168 = ~n3020 & n7160 ;
  assign n7169 = n3020 & ~n7160 ;
  assign n7170 = ~n7168 & ~n7169 ;
  assign n7171 = n4925 & n7170 ;
  assign n7172 = ~n7151 & ~n7171 ;
  assign n7173 = n3179 & ~n7172 ;
  assign n7161 = ~n3235 & n7160 ;
  assign n7162 = n3235 & ~n7160 ;
  assign n7163 = ~n7161 & ~n7162 ;
  assign n7164 = n4925 & ~n7163 ;
  assign n7165 = ~n7151 & ~n7164 ;
  assign n7166 = n3319 & ~n7165 ;
  assign n7145 = ~n3118 & ~n6409 ;
  assign n7146 = n3409 & n6408 ;
  assign n7147 = n3118 & ~n3375 ;
  assign n7148 = ~n7146 & n7147 ;
  assign n7149 = ~n7145 & ~n7148 ;
  assign n7150 = n4925 & n7149 ;
  assign n7144 = n3099 & n4934 ;
  assign n7167 = n3118 & n3415 ;
  assign n7174 = ~n7144 & ~n7167 ;
  assign n7175 = ~n7150 & n7174 ;
  assign n7176 = ~n7166 & n7175 ;
  assign n7177 = ~n7173 & n7176 ;
  assign n7178 = ~n7159 & n7177 ;
  assign n7179 = n2017 & ~n7178 ;
  assign n7180 = ~n7143 & ~n7179 ;
  assign n7181 = \P1_state_reg[0]/NET0131  & ~n7180 ;
  assign n7141 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[13]/NET0131  ;
  assign n7142 = n3099 & n3935 ;
  assign n7182 = ~n7141 & ~n7142 ;
  assign n7183 = ~n7181 & n7182 ;
  assign n7186 = n3051 & n3430 ;
  assign n7188 = n3051 & ~n4925 ;
  assign n7197 = n3046 & ~n5821 ;
  assign n7198 = ~n6430 & ~n7197 ;
  assign n7199 = ~n2050 & ~n7198 ;
  assign n7200 = n2050 & n3082 ;
  assign n7201 = ~n7199 & ~n7200 ;
  assign n7202 = n4925 & n7201 ;
  assign n7203 = ~n7188 & ~n7202 ;
  assign n7204 = n3373 & ~n7203 ;
  assign n7189 = ~n4391 & n4393 ;
  assign n7190 = n4397 & ~n7189 ;
  assign n7191 = n4120 & ~n7190 ;
  assign n7192 = ~n4120 & n7190 ;
  assign n7193 = ~n7191 & ~n7192 ;
  assign n7194 = n4925 & n7193 ;
  assign n7195 = ~n7188 & ~n7194 ;
  assign n7196 = n3179 & ~n7195 ;
  assign n7205 = n4120 & ~n4354 ;
  assign n7206 = ~n4120 & n4354 ;
  assign n7207 = ~n7205 & ~n7206 ;
  assign n7208 = n4925 & ~n7207 ;
  assign n7209 = ~n7188 & ~n7208 ;
  assign n7210 = n3319 & ~n7209 ;
  assign n7211 = n3071 & ~n6453 ;
  assign n7212 = n3409 & ~n6454 ;
  assign n7213 = ~n7211 & n7212 ;
  assign n7214 = n4925 & n7213 ;
  assign n7187 = n3051 & n4934 ;
  assign n7215 = n3071 & ~n5093 ;
  assign n7216 = ~n7187 & ~n7215 ;
  assign n7217 = ~n7214 & n7216 ;
  assign n7218 = ~n7210 & n7217 ;
  assign n7219 = ~n7196 & n7218 ;
  assign n7220 = ~n7204 & n7219 ;
  assign n7221 = n2017 & ~n7220 ;
  assign n7222 = ~n7186 & ~n7221 ;
  assign n7223 = \P1_state_reg[0]/NET0131  & ~n7222 ;
  assign n7184 = n3051 & n3935 ;
  assign n7185 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[15]/NET0131  ;
  assign n7224 = ~n7184 & ~n7185 ;
  assign n7225 = ~n7223 & n7224 ;
  assign n7228 = n2984 & n3430 ;
  assign n7236 = n2984 & ~n4925 ;
  assign n7237 = n2965 & ~n3339 ;
  assign n7238 = ~n7108 & ~n7237 ;
  assign n7239 = ~n2050 & ~n7238 ;
  assign n7240 = n2050 & n2678 ;
  assign n7241 = ~n7239 & ~n7240 ;
  assign n7242 = n4925 & n7241 ;
  assign n7243 = ~n7236 & ~n7242 ;
  assign n7244 = n3373 & ~n7243 ;
  assign n7252 = ~n3230 & n4127 ;
  assign n7253 = n3230 & ~n4127 ;
  assign n7254 = ~n7252 & ~n7253 ;
  assign n7255 = n4925 & ~n7254 ;
  assign n7256 = ~n7236 & ~n7255 ;
  assign n7257 = n3319 & ~n7256 ;
  assign n7245 = ~n2901 & n4127 ;
  assign n7246 = n2901 & ~n4127 ;
  assign n7247 = ~n7245 & ~n7246 ;
  assign n7248 = n4925 & n7247 ;
  assign n7249 = ~n7236 & ~n7248 ;
  assign n7250 = n3179 & ~n7249 ;
  assign n7230 = n3005 & n3375 ;
  assign n7231 = n3005 & ~n3384 ;
  assign n7232 = n3409 & ~n7124 ;
  assign n7233 = ~n7231 & n7232 ;
  assign n7234 = ~n7230 & ~n7233 ;
  assign n7235 = n4925 & ~n7234 ;
  assign n7229 = n2984 & n4934 ;
  assign n7251 = n3005 & n3415 ;
  assign n7258 = ~n7229 & ~n7251 ;
  assign n7259 = ~n7235 & n7258 ;
  assign n7260 = ~n7250 & n7259 ;
  assign n7261 = ~n7257 & n7260 ;
  assign n7262 = ~n7244 & n7261 ;
  assign n7263 = n2017 & ~n7262 ;
  assign n7264 = ~n7228 & ~n7263 ;
  assign n7265 = \P1_state_reg[0]/NET0131  & ~n7264 ;
  assign n7226 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[9]/NET0131  ;
  assign n7227 = n2984 & n3935 ;
  assign n7266 = ~n7226 & ~n7227 ;
  assign n7267 = ~n7265 & n7266 ;
  assign n7270 = n1182 & n3664 ;
  assign n7279 = ~n1274 & n3581 ;
  assign n7280 = ~n1222 & n7279 ;
  assign n7281 = ~n1248 & n7280 ;
  assign n7282 = ~n1189 & n7281 ;
  assign n7283 = ~n536 & ~n1162 ;
  assign n7284 = ~n7282 & ~n7283 ;
  assign n7285 = ~n3586 & ~n7284 ;
  assign n7286 = n536 & ~n1248 ;
  assign n7287 = ~n7285 & ~n7286 ;
  assign n7288 = n1898 & ~n7287 ;
  assign n7289 = ~n1202 & ~n3632 ;
  assign n7290 = n3650 & ~n6495 ;
  assign n7291 = ~n7289 & n7290 ;
  assign n7293 = n1419 & ~n1757 ;
  assign n7292 = ~n1419 & n1757 ;
  assign n7294 = n3575 & ~n7292 ;
  assign n7295 = ~n7293 & n7294 ;
  assign n7296 = ~n7291 & ~n7295 ;
  assign n7297 = ~n7288 & n7296 ;
  assign n7298 = n3450 & ~n7297 ;
  assign n7272 = n1757 & ~n3489 ;
  assign n7273 = ~n1757 & n3489 ;
  assign n7274 = ~n7272 & ~n7273 ;
  assign n7275 = n3450 & n7274 ;
  assign n7276 = ~n1182 & ~n3450 ;
  assign n7277 = n3557 & ~n7276 ;
  assign n7278 = ~n7275 & n7277 ;
  assign n7271 = ~n1202 & n3655 ;
  assign n7299 = ~n6590 & n6935 ;
  assign n7300 = n1182 & ~n7299 ;
  assign n7301 = ~n7271 & ~n7300 ;
  assign n7302 = ~n7278 & n7301 ;
  assign n7303 = ~n7298 & n7302 ;
  assign n7304 = n3662 & ~n7303 ;
  assign n7305 = ~n7270 & ~n7304 ;
  assign n7306 = \P1_state_reg[0]/NET0131  & ~n7305 ;
  assign n7268 = \P1_reg3_reg[8]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7269 = n1182 & n1934 ;
  assign n7307 = ~n7268 & ~n7269 ;
  assign n7308 = ~n7306 & n7307 ;
  assign n7311 = n3409 & n6819 ;
  assign n7310 = n3319 & n6825 ;
  assign n7309 = n3373 & n6833 ;
  assign n7312 = n6842 & ~n7309 ;
  assign n7313 = ~n7310 & n7312 ;
  assign n7314 = ~n7311 & n7313 ;
  assign n7315 = n4925 & ~n7314 ;
  assign n7316 = n2579 & n3415 ;
  assign n7317 = ~n7315 & ~n7316 ;
  assign n7318 = n2017 & ~n7317 ;
  assign n7320 = ~n3415 & ~n4933 ;
  assign n7321 = ~n3319 & n7320 ;
  assign n7319 = n3319 & ~n4925 ;
  assign n7322 = ~n2016 & ~n7319 ;
  assign n7323 = ~n7321 & n7322 ;
  assign n7324 = ~n1984 & n2584 ;
  assign n7325 = ~n7323 & n7324 ;
  assign n7326 = ~n7318 & ~n7325 ;
  assign n7327 = \P1_state_reg[0]/NET0131  & ~n7326 ;
  assign n7328 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[20]/NET0131  ;
  assign n7329 = n2584 & n3935 ;
  assign n7330 = ~n7328 & ~n7329 ;
  assign n7331 = ~n7327 & n7330 ;
  assign n7332 = n917 & ~n3450 ;
  assign n7333 = ~n4994 & n4996 ;
  assign n7334 = n5001 & ~n7333 ;
  assign n7335 = n1796 & n7334 ;
  assign n7336 = ~n1796 & ~n7334 ;
  assign n7337 = ~n7335 & ~n7336 ;
  assign n7338 = n3450 & n7337 ;
  assign n7339 = ~n7332 & ~n7338 ;
  assign n7340 = n3575 & ~n7339 ;
  assign n7341 = n5013 & n5022 ;
  assign n7342 = ~n7060 & n7341 ;
  assign n7343 = n5013 & ~n5031 ;
  assign n7344 = n5035 & ~n7343 ;
  assign n7345 = ~n7342 & n7344 ;
  assign n7346 = n1796 & n7345 ;
  assign n7347 = ~n1796 & ~n7345 ;
  assign n7348 = ~n7346 & ~n7347 ;
  assign n7349 = n3450 & ~n7348 ;
  assign n7350 = ~n7332 & ~n7349 ;
  assign n7351 = n3557 & ~n7350 ;
  assign n7352 = n1570 & ~n4285 ;
  assign n7353 = ~n4286 & ~n7352 ;
  assign n7354 = ~n536 & ~n7353 ;
  assign n7355 = n536 & n887 ;
  assign n7356 = ~n7354 & ~n7355 ;
  assign n7357 = n3450 & n7356 ;
  assign n7358 = ~n7332 & ~n7357 ;
  assign n7359 = n1898 & ~n7358 ;
  assign n7362 = ~n911 & n4839 ;
  assign n7361 = n911 & ~n4839 ;
  assign n7363 = n3650 & ~n7361 ;
  assign n7364 = ~n7362 & n7363 ;
  assign n7365 = n3450 & n7364 ;
  assign n7360 = n917 & ~n3618 ;
  assign n7366 = n911 & n3655 ;
  assign n7367 = ~n7360 & ~n7366 ;
  assign n7368 = ~n7365 & n7367 ;
  assign n7369 = ~n7359 & n7368 ;
  assign n7370 = ~n7351 & n7369 ;
  assign n7371 = ~n7340 & n7370 ;
  assign n7372 = n3662 & ~n7371 ;
  assign n7373 = n917 & n3664 ;
  assign n7374 = ~n7372 & ~n7373 ;
  assign n7375 = \P1_state_reg[0]/NET0131  & ~n7374 ;
  assign n7376 = n917 & n1934 ;
  assign n7377 = \P1_reg3_reg[23]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7378 = ~n7376 & ~n7377 ;
  assign n7379 = ~n7375 & n7378 ;
  assign n7382 = n2547 & n3430 ;
  assign n7384 = n2547 & ~n4925 ;
  assign n7385 = n3146 & n4138 ;
  assign n7386 = ~n3146 & ~n4138 ;
  assign n7387 = ~n7385 & ~n7386 ;
  assign n7388 = n4925 & ~n7387 ;
  assign n7389 = ~n7384 & ~n7388 ;
  assign n7390 = n3179 & ~n7389 ;
  assign n7399 = ~n3274 & n4138 ;
  assign n7400 = n3274 & ~n4138 ;
  assign n7401 = ~n7399 & ~n7400 ;
  assign n7402 = n4925 & ~n7401 ;
  assign n7403 = ~n7384 & ~n7402 ;
  assign n7404 = n3319 & ~n7403 ;
  assign n7391 = n2531 & ~n6046 ;
  assign n7392 = ~n6047 & ~n7391 ;
  assign n7393 = ~n2050 & ~n7392 ;
  assign n7394 = n2050 & n2588 ;
  assign n7395 = ~n7393 & ~n7394 ;
  assign n7396 = n4925 & n7395 ;
  assign n7397 = ~n7384 & ~n7396 ;
  assign n7398 = n3373 & ~n7397 ;
  assign n7405 = n2541 & ~n6817 ;
  assign n7406 = ~n6053 & ~n7405 ;
  assign n7407 = n4925 & n7406 ;
  assign n7408 = ~n7384 & ~n7407 ;
  assign n7409 = n3409 & ~n7408 ;
  assign n7383 = n2541 & ~n5093 ;
  assign n7410 = n2547 & n5090 ;
  assign n7411 = ~n7383 & ~n7410 ;
  assign n7412 = ~n7409 & n7411 ;
  assign n7413 = ~n7398 & n7412 ;
  assign n7414 = ~n7404 & n7413 ;
  assign n7415 = ~n7390 & n7414 ;
  assign n7416 = n2017 & ~n7415 ;
  assign n7417 = ~n7382 & ~n7416 ;
  assign n7418 = \P1_state_reg[0]/NET0131  & ~n7417 ;
  assign n7380 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[21]/NET0131  ;
  assign n7381 = n2547 & n3935 ;
  assign n7419 = ~n7380 & ~n7381 ;
  assign n7420 = ~n7418 & n7419 ;
  assign n7423 = n2503 & n3430 ;
  assign n7424 = n2503 & ~n4925 ;
  assign n7436 = ~n4361 & n4365 ;
  assign n7437 = n4144 & ~n7436 ;
  assign n7438 = ~n4144 & n7436 ;
  assign n7439 = ~n7437 & ~n7438 ;
  assign n7440 = n4925 & ~n7439 ;
  assign n7441 = ~n7424 & ~n7440 ;
  assign n7442 = n3319 & ~n7441 ;
  assign n7425 = n4392 & n4403 ;
  assign n7426 = ~n7190 & n7425 ;
  assign n7427 = ~n4400 & n4403 ;
  assign n7428 = n4377 & ~n7427 ;
  assign n7429 = ~n7426 & n7428 ;
  assign n7430 = n4144 & n7429 ;
  assign n7431 = ~n4144 & ~n7429 ;
  assign n7432 = ~n7430 & ~n7431 ;
  assign n7433 = n4925 & ~n7432 ;
  assign n7434 = ~n7424 & ~n7433 ;
  assign n7435 = n3179 & ~n7434 ;
  assign n7444 = n2484 & ~n6045 ;
  assign n7445 = ~n5495 & ~n7444 ;
  assign n7446 = ~n2050 & ~n7445 ;
  assign n7447 = n2050 & n2531 ;
  assign n7448 = ~n7446 & ~n7447 ;
  assign n7449 = n4925 & n7448 ;
  assign n7450 = ~n7424 & ~n7449 ;
  assign n7451 = n3373 & ~n7450 ;
  assign n7452 = n2498 & ~n6055 ;
  assign n7453 = n3409 & ~n4906 ;
  assign n7454 = ~n7452 & n7453 ;
  assign n7455 = n4925 & n7454 ;
  assign n7443 = n2498 & ~n5093 ;
  assign n7456 = n2503 & n4934 ;
  assign n7457 = ~n7443 & ~n7456 ;
  assign n7458 = ~n7455 & n7457 ;
  assign n7459 = ~n7451 & n7458 ;
  assign n7460 = ~n7435 & n7459 ;
  assign n7461 = ~n7442 & n7460 ;
  assign n7462 = n2017 & ~n7461 ;
  assign n7463 = ~n7423 & ~n7462 ;
  assign n7464 = \P1_state_reg[0]/NET0131  & ~n7463 ;
  assign n7421 = n2503 & n3935 ;
  assign n7422 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[23]/NET0131  ;
  assign n7465 = ~n7421 & ~n7422 ;
  assign n7466 = ~n7464 & n7465 ;
  assign n7467 = \P2_reg0_reg[21]/NET0131  & ~n3434 ;
  assign n7468 = \P2_reg0_reg[21]/NET0131  & n3430 ;
  assign n7470 = \P2_reg0_reg[21]/NET0131  & ~n4610 ;
  assign n7471 = n4610 & ~n7387 ;
  assign n7472 = ~n7470 & ~n7471 ;
  assign n7473 = n3179 & ~n7472 ;
  assign n7477 = n4610 & ~n7401 ;
  assign n7478 = ~n7470 & ~n7477 ;
  assign n7479 = n3319 & ~n7478 ;
  assign n7474 = n4610 & n7395 ;
  assign n7475 = ~n7470 & ~n7474 ;
  assign n7476 = n3373 & ~n7475 ;
  assign n7469 = \P2_reg0_reg[21]/NET0131  & ~n5258 ;
  assign n7480 = n2541 & n3375 ;
  assign n7481 = n3409 & n7406 ;
  assign n7482 = ~n7480 & ~n7481 ;
  assign n7483 = n4610 & ~n7482 ;
  assign n7484 = ~n7469 & ~n7483 ;
  assign n7485 = ~n7476 & n7484 ;
  assign n7486 = ~n7479 & n7485 ;
  assign n7487 = ~n7473 & n7486 ;
  assign n7488 = n2017 & ~n7487 ;
  assign n7489 = ~n7468 & ~n7488 ;
  assign n7490 = \P1_state_reg[0]/NET0131  & ~n7489 ;
  assign n7491 = ~n7467 & ~n7490 ;
  assign n7492 = \P1_reg1_reg[8]/NET0131  & ~n6244 ;
  assign n7493 = n3557 & ~n7274 ;
  assign n7494 = ~n1202 & n3683 ;
  assign n7495 = ~n7493 & ~n7494 ;
  assign n7496 = n7297 & n7495 ;
  assign n7497 = n6246 & ~n7496 ;
  assign n7498 = ~n7492 & ~n7497 ;
  assign n7499 = \P1_reg1_reg[9]/NET0131  & ~n3703 ;
  assign n7500 = \P1_reg1_reg[9]/NET0131  & n3664 ;
  assign n7502 = \P1_reg1_reg[9]/NET0131  & ~n4236 ;
  assign n7511 = n4236 & n6479 ;
  assign n7512 = ~n7502 & ~n7511 ;
  assign n7513 = n1898 & ~n7512 ;
  assign n7503 = n4236 & n6485 ;
  assign n7504 = ~n7502 & ~n7503 ;
  assign n7505 = n3557 & ~n7504 ;
  assign n7501 = \P1_reg1_reg[9]/NET0131  & ~n6242 ;
  assign n7506 = n3575 & ~n6491 ;
  assign n7507 = ~n1178 & n3683 ;
  assign n7508 = ~n6498 & ~n7507 ;
  assign n7509 = ~n7506 & n7508 ;
  assign n7510 = n4236 & ~n7509 ;
  assign n7514 = ~n7501 & ~n7510 ;
  assign n7515 = ~n7505 & n7514 ;
  assign n7516 = ~n7513 & n7515 ;
  assign n7517 = n3662 & ~n7516 ;
  assign n7518 = ~n7500 & ~n7517 ;
  assign n7519 = \P1_state_reg[0]/NET0131  & ~n7518 ;
  assign n7520 = ~n7499 & ~n7519 ;
  assign n7521 = n3375 & n3977 ;
  assign n7522 = ~n4265 & ~n7521 ;
  assign n7523 = n4610 & ~n7522 ;
  assign n7524 = ~n3406 & n3977 ;
  assign n7525 = ~n4266 & ~n7524 ;
  assign n7526 = n4610 & ~n7525 ;
  assign n7527 = ~\P2_reg0_reg[30]/NET0131  & ~n4610 ;
  assign n7528 = n3409 & ~n7527 ;
  assign n7529 = ~n7526 & n7528 ;
  assign n7530 = ~n7523 & ~n7529 ;
  assign n7531 = n4275 & ~n7530 ;
  assign n7532 = ~n4610 & ~n5605 ;
  assign n7533 = n4275 & ~n7532 ;
  assign n7534 = n5256 & n7533 ;
  assign n7535 = \P2_reg0_reg[30]/NET0131  & ~n7534 ;
  assign n7536 = ~n7531 & ~n7535 ;
  assign n7537 = \P1_reg2_reg[19]/NET0131  & ~n3703 ;
  assign n7538 = \P1_reg2_reg[19]/NET0131  & n3664 ;
  assign n7540 = \P1_reg2_reg[19]/NET0131  & ~n3672 ;
  assign n7544 = n3672 & n6355 ;
  assign n7545 = ~n7540 & ~n7544 ;
  assign n7546 = n1898 & ~n7545 ;
  assign n7541 = n3672 & n6347 ;
  assign n7542 = ~n7540 & ~n7541 ;
  assign n7543 = n3575 & ~n7542 ;
  assign n7547 = n3672 & n6362 ;
  assign n7548 = ~n7540 & ~n7547 ;
  assign n7549 = n3557 & ~n7548 ;
  assign n7550 = n3672 & n6369 ;
  assign n7551 = ~n7540 & ~n7550 ;
  assign n7552 = n3650 & ~n7551 ;
  assign n7554 = ~n638 & n3683 ;
  assign n7555 = n3672 & n7554 ;
  assign n7539 = \P1_reg2_reg[19]/NET0131  & ~n3685 ;
  assign n7553 = n688 & n1736 ;
  assign n7556 = ~n7539 & ~n7553 ;
  assign n7557 = ~n7555 & n7556 ;
  assign n7558 = ~n7552 & n7557 ;
  assign n7559 = ~n7549 & n7558 ;
  assign n7560 = ~n7543 & n7559 ;
  assign n7561 = ~n7546 & n7560 ;
  assign n7562 = n3662 & ~n7561 ;
  assign n7563 = ~n7538 & ~n7562 ;
  assign n7564 = \P1_state_reg[0]/NET0131  & ~n7563 ;
  assign n7565 = ~n7537 & ~n7564 ;
  assign n7571 = \P2_reg1_reg[12]/NET0131  & ~n4663 ;
  assign n7572 = n4663 & ~n6388 ;
  assign n7573 = ~n7571 & ~n7572 ;
  assign n7574 = n3319 & ~n7573 ;
  assign n7575 = n4663 & n6397 ;
  assign n7576 = ~n7571 & ~n7575 ;
  assign n7577 = n3373 & ~n7576 ;
  assign n7566 = n3179 & n6403 ;
  assign n7567 = n2954 & n3375 ;
  assign n7568 = ~n6410 & ~n7567 ;
  assign n7569 = ~n7566 & n7568 ;
  assign n7570 = n4663 & ~n7569 ;
  assign n7578 = n5509 & ~n6717 ;
  assign n7579 = \P2_reg1_reg[12]/NET0131  & ~n7578 ;
  assign n7580 = ~n7570 & ~n7579 ;
  assign n7581 = ~n7577 & n7580 ;
  assign n7582 = ~n7574 & n7581 ;
  assign n7583 = n2017 & ~n7582 ;
  assign n7584 = \P2_reg1_reg[12]/NET0131  & n3430 ;
  assign n7585 = ~n7583 & ~n7584 ;
  assign n7586 = \P1_state_reg[0]/NET0131  & ~n7585 ;
  assign n7587 = \P2_reg1_reg[12]/NET0131  & ~n3434 ;
  assign n7588 = ~n7586 & ~n7587 ;
  assign n7589 = \P1_reg2_reg[23]/NET0131  & n3664 ;
  assign n7590 = \P1_reg2_reg[23]/NET0131  & ~n3672 ;
  assign n7591 = n3672 & n7337 ;
  assign n7592 = ~n7590 & ~n7591 ;
  assign n7593 = n3575 & ~n7592 ;
  assign n7594 = n3672 & ~n7348 ;
  assign n7595 = ~n7590 & ~n7594 ;
  assign n7596 = n3557 & ~n7595 ;
  assign n7597 = n1898 & n7356 ;
  assign n7598 = n911 & n3683 ;
  assign n7599 = ~n7364 & ~n7598 ;
  assign n7600 = ~n7597 & n7599 ;
  assign n7601 = n3672 & ~n7600 ;
  assign n7602 = n917 & n1736 ;
  assign n7603 = \P1_reg2_reg[23]/NET0131  & ~n6694 ;
  assign n7604 = ~n7602 & ~n7603 ;
  assign n7605 = ~n7601 & n7604 ;
  assign n7606 = ~n7596 & n7605 ;
  assign n7607 = ~n7593 & n7606 ;
  assign n7608 = n3662 & ~n7607 ;
  assign n7609 = ~n7589 & ~n7608 ;
  assign n7610 = \P1_state_reg[0]/NET0131  & ~n7609 ;
  assign n7611 = \P1_reg2_reg[23]/NET0131  & ~n3703 ;
  assign n7612 = ~n7610 & ~n7611 ;
  assign n7613 = \P2_reg1_reg[16]/NET0131  & ~n3434 ;
  assign n7614 = \P2_reg1_reg[16]/NET0131  & n3430 ;
  assign n7615 = \P2_reg1_reg[16]/NET0131  & ~n6721 ;
  assign n7620 = n3409 & n6456 ;
  assign n7618 = n3036 & n3375 ;
  assign n7619 = n3179 & ~n6443 ;
  assign n7621 = ~n7618 & ~n7619 ;
  assign n7622 = ~n7620 & n7621 ;
  assign n7616 = n3373 & n6435 ;
  assign n7617 = n3319 & ~n6449 ;
  assign n7623 = ~n7616 & ~n7617 ;
  assign n7624 = n7622 & n7623 ;
  assign n7625 = n4663 & ~n7624 ;
  assign n7626 = ~n7615 & ~n7625 ;
  assign n7627 = n2017 & ~n7626 ;
  assign n7628 = ~n7614 & ~n7627 ;
  assign n7629 = \P1_state_reg[0]/NET0131  & ~n7628 ;
  assign n7630 = ~n7613 & ~n7629 ;
  assign n7631 = \P2_reg1_reg[20]/NET0131  & ~n5608 ;
  assign n7632 = n5572 & ~n7314 ;
  assign n7633 = ~n7631 & ~n7632 ;
  assign n7634 = \P2_reg1_reg[21]/NET0131  & ~n3434 ;
  assign n7635 = \P2_reg1_reg[21]/NET0131  & n3430 ;
  assign n7637 = \P2_reg1_reg[21]/NET0131  & ~n4663 ;
  assign n7638 = n4663 & ~n7387 ;
  assign n7639 = ~n7637 & ~n7638 ;
  assign n7640 = n3179 & ~n7639 ;
  assign n7644 = n4663 & ~n7401 ;
  assign n7645 = ~n7637 & ~n7644 ;
  assign n7646 = n3319 & ~n7645 ;
  assign n7641 = n4663 & n7395 ;
  assign n7642 = ~n7637 & ~n7641 ;
  assign n7643 = n3373 & ~n7642 ;
  assign n7636 = \P2_reg1_reg[21]/NET0131  & ~n5509 ;
  assign n7647 = n4663 & ~n7482 ;
  assign n7648 = ~n7636 & ~n7647 ;
  assign n7649 = ~n7643 & n7648 ;
  assign n7650 = ~n7646 & n7649 ;
  assign n7651 = ~n7640 & n7650 ;
  assign n7652 = n2017 & ~n7651 ;
  assign n7653 = ~n7635 & ~n7652 ;
  assign n7654 = \P1_state_reg[0]/NET0131  & ~n7653 ;
  assign n7655 = ~n7634 & ~n7654 ;
  assign n7656 = n3409 & n7525 ;
  assign n7657 = n7522 & ~n7656 ;
  assign n7658 = n5572 & ~n7657 ;
  assign n7659 = \P2_reg1_reg[30]/NET0131  & ~n5569 ;
  assign n7660 = ~n7658 & ~n7659 ;
  assign n7661 = \P2_reg2_reg[12]/NET0131  & ~n3434 ;
  assign n7663 = \P2_reg2_reg[12]/NET0131  & ~n2033 ;
  assign n7664 = n2033 & ~n6388 ;
  assign n7665 = ~n7663 & ~n7664 ;
  assign n7666 = n3319 & ~n7665 ;
  assign n7667 = n2033 & n6397 ;
  assign n7668 = ~n7663 & ~n7667 ;
  assign n7669 = n3373 & ~n7668 ;
  assign n7670 = n2033 & ~n7569 ;
  assign n7662 = n2931 & n3415 ;
  assign n7671 = n4436 & ~n6793 ;
  assign n7672 = \P2_reg2_reg[12]/NET0131  & ~n7671 ;
  assign n7673 = ~n7662 & ~n7672 ;
  assign n7674 = ~n7670 & n7673 ;
  assign n7675 = ~n7669 & n7674 ;
  assign n7676 = ~n7666 & n7675 ;
  assign n7677 = n2017 & ~n7676 ;
  assign n7678 = \P2_reg2_reg[12]/NET0131  & n3430 ;
  assign n7679 = ~n7677 & ~n7678 ;
  assign n7680 = \P1_state_reg[0]/NET0131  & ~n7679 ;
  assign n7681 = ~n7661 & ~n7680 ;
  assign n7682 = \P2_reg2_reg[16]/NET0131  & ~n3434 ;
  assign n7683 = \P2_reg2_reg[16]/NET0131  & n3430 ;
  assign n7685 = n2033 & ~n7624 ;
  assign n7684 = \P2_reg2_reg[16]/NET0131  & ~n6796 ;
  assign n7686 = n3042 & n3415 ;
  assign n7687 = ~n7684 & ~n7686 ;
  assign n7688 = ~n7685 & n7687 ;
  assign n7689 = n2017 & ~n7688 ;
  assign n7690 = ~n7683 & ~n7689 ;
  assign n7691 = \P1_state_reg[0]/NET0131  & ~n7690 ;
  assign n7692 = ~n7682 & ~n7691 ;
  assign n7693 = n1182 & n1736 ;
  assign n7694 = n3672 & ~n7496 ;
  assign n7695 = ~n7693 & ~n7694 ;
  assign n7696 = n6070 & ~n7695 ;
  assign n7697 = ~n3672 & ~n5761 ;
  assign n7698 = n3685 & ~n7697 ;
  assign n7699 = n6070 & n7698 ;
  assign n7700 = \P1_reg2_reg[8]/NET0131  & ~n7699 ;
  assign n7701 = ~n7696 & ~n7700 ;
  assign n7702 = \P2_reg2_reg[21]/NET0131  & ~n3434 ;
  assign n7703 = \P2_reg2_reg[21]/NET0131  & n3430 ;
  assign n7705 = \P2_reg2_reg[21]/NET0131  & ~n2033 ;
  assign n7706 = n2033 & ~n7387 ;
  assign n7707 = ~n7705 & ~n7706 ;
  assign n7708 = n3179 & ~n7707 ;
  assign n7714 = n2033 & ~n7401 ;
  assign n7715 = ~n7705 & ~n7714 ;
  assign n7716 = n3319 & ~n7715 ;
  assign n7709 = n2033 & n7395 ;
  assign n7710 = ~n7705 & ~n7709 ;
  assign n7711 = n3373 & ~n7710 ;
  assign n7713 = n2033 & ~n7482 ;
  assign n7704 = n2547 & n3415 ;
  assign n7712 = \P2_reg2_reg[21]/NET0131  & ~n4436 ;
  assign n7717 = ~n7704 & ~n7712 ;
  assign n7718 = ~n7713 & n7717 ;
  assign n7719 = ~n7711 & n7718 ;
  assign n7720 = ~n7716 & n7719 ;
  assign n7721 = ~n7708 & n7720 ;
  assign n7722 = n2017 & ~n7721 ;
  assign n7723 = ~n7703 & ~n7722 ;
  assign n7724 = \P1_state_reg[0]/NET0131  & ~n7723 ;
  assign n7725 = ~n7702 & ~n7724 ;
  assign n7726 = \P2_reg2_reg[23]/NET0131  & ~n3434 ;
  assign n7727 = \P2_reg2_reg[23]/NET0131  & n3430 ;
  assign n7728 = \P2_reg2_reg[23]/NET0131  & ~n2033 ;
  assign n7732 = n2033 & ~n7439 ;
  assign n7733 = ~n7728 & ~n7732 ;
  assign n7734 = n3319 & ~n7733 ;
  assign n7729 = n2033 & ~n7432 ;
  assign n7730 = ~n7728 & ~n7729 ;
  assign n7731 = n3179 & ~n7730 ;
  assign n7736 = n2033 & n7448 ;
  assign n7737 = ~n7728 & ~n7736 ;
  assign n7738 = n3373 & ~n7737 ;
  assign n7739 = n2498 & n3375 ;
  assign n7740 = ~n7454 & ~n7739 ;
  assign n7741 = n2033 & ~n7740 ;
  assign n7735 = n2503 & n3415 ;
  assign n7742 = \P2_reg2_reg[23]/NET0131  & ~n4436 ;
  assign n7743 = ~n7735 & ~n7742 ;
  assign n7744 = ~n7741 & n7743 ;
  assign n7745 = ~n7738 & n7744 ;
  assign n7746 = ~n7731 & n7745 ;
  assign n7747 = ~n7734 & n7746 ;
  assign n7748 = n2017 & ~n7747 ;
  assign n7749 = ~n7727 & ~n7748 ;
  assign n7750 = \P1_state_reg[0]/NET0131  & ~n7749 ;
  assign n7751 = ~n7726 & ~n7750 ;
  assign n7752 = \P2_reg2_reg[30]/NET0131  & ~n3434 ;
  assign n7753 = \P2_reg2_reg[30]/NET0131  & n3430 ;
  assign n7754 = \P2_reg2_reg[30]/NET0131  & ~n3415 ;
  assign n7755 = ~n2033 & ~n7754 ;
  assign n7756 = \P2_reg2_reg[30]/NET0131  & ~n3419 ;
  assign n7757 = n7657 & ~n7756 ;
  assign n7758 = ~n7755 & ~n7757 ;
  assign n7759 = ~n3416 & ~n7758 ;
  assign n7760 = n2017 & ~n7759 ;
  assign n7761 = ~n7753 & ~n7760 ;
  assign n7762 = \P1_state_reg[0]/NET0131  & ~n7761 ;
  assign n7763 = ~n7752 & ~n7762 ;
  assign n7764 = \P1_reg0_reg[18]/NET0131  & ~n3703 ;
  assign n7765 = \P1_reg0_reg[18]/NET0131  & n3664 ;
  assign n7767 = \P1_reg0_reg[18]/NET0131  & ~n3900 ;
  assign n7771 = n3900 & ~n5789 ;
  assign n7772 = ~n7767 & ~n7771 ;
  assign n7773 = n3575 & ~n7772 ;
  assign n7768 = n3900 & n5783 ;
  assign n7769 = ~n7767 & ~n7768 ;
  assign n7770 = n3557 & ~n7769 ;
  assign n7774 = n3900 & n5798 ;
  assign n7775 = ~n7767 & ~n7774 ;
  assign n7776 = n1898 & ~n7775 ;
  assign n7766 = \P1_reg0_reg[18]/NET0131  & ~n4723 ;
  assign n7777 = n3900 & ~n6641 ;
  assign n7778 = ~n7766 & ~n7777 ;
  assign n7779 = ~n7776 & n7778 ;
  assign n7780 = ~n7770 & n7779 ;
  assign n7781 = ~n7773 & n7780 ;
  assign n7782 = n3662 & ~n7781 ;
  assign n7783 = ~n7765 & ~n7782 ;
  assign n7784 = \P1_state_reg[0]/NET0131  & ~n7783 ;
  assign n7785 = ~n7764 & ~n7784 ;
  assign n7786 = \P1_reg0_reg[19]/NET0131  & ~n3703 ;
  assign n7787 = \P1_reg0_reg[19]/NET0131  & n3664 ;
  assign n7789 = \P1_reg0_reg[19]/NET0131  & ~n3900 ;
  assign n7793 = n3900 & n6355 ;
  assign n7794 = ~n7789 & ~n7793 ;
  assign n7795 = n1898 & ~n7794 ;
  assign n7790 = n3900 & n6347 ;
  assign n7791 = ~n7789 & ~n7790 ;
  assign n7792 = n3575 & ~n7791 ;
  assign n7798 = n3900 & n6362 ;
  assign n7799 = ~n7789 & ~n7798 ;
  assign n7800 = n3557 & ~n7799 ;
  assign n7788 = \P1_reg0_reg[19]/NET0131  & ~n4723 ;
  assign n7796 = ~n6370 & ~n7554 ;
  assign n7797 = n3900 & ~n7796 ;
  assign n7801 = ~n7788 & ~n7797 ;
  assign n7802 = ~n7800 & n7801 ;
  assign n7803 = ~n7792 & n7802 ;
  assign n7804 = ~n7795 & n7803 ;
  assign n7805 = n3662 & ~n7804 ;
  assign n7806 = ~n7787 & ~n7805 ;
  assign n7807 = \P1_state_reg[0]/NET0131  & ~n7806 ;
  assign n7808 = ~n7786 & ~n7807 ;
  assign n7812 = \P1_reg0_reg[22]/NET0131  & ~n3900 ;
  assign n7813 = n6171 & ~n6564 ;
  assign n7814 = ~n7812 & ~n7813 ;
  assign n7815 = n3557 & ~n7814 ;
  assign n7809 = n3575 & ~n6574 ;
  assign n7810 = n6691 & ~n7809 ;
  assign n7811 = n6171 & ~n7810 ;
  assign n7816 = n4706 & n6860 ;
  assign n7817 = \P1_reg0_reg[22]/NET0131  & ~n7816 ;
  assign n7818 = ~n7811 & ~n7817 ;
  assign n7819 = ~n7815 & n7818 ;
  assign n7820 = \P1_reg0_reg[23]/NET0131  & ~n3900 ;
  assign n7821 = n3900 & n7337 ;
  assign n7822 = ~n7820 & ~n7821 ;
  assign n7823 = n3575 & ~n7822 ;
  assign n7824 = n3900 & ~n7348 ;
  assign n7825 = ~n7820 & ~n7824 ;
  assign n7826 = n3557 & ~n7825 ;
  assign n7827 = n3900 & ~n7600 ;
  assign n7828 = \P1_reg0_reg[23]/NET0131  & ~n4706 ;
  assign n7829 = ~n7827 & ~n7828 ;
  assign n7830 = ~n7826 & n7829 ;
  assign n7831 = ~n7823 & n7830 ;
  assign n7832 = n3662 & ~n7831 ;
  assign n7833 = \P1_reg0_reg[23]/NET0131  & n3664 ;
  assign n7834 = ~n7832 & ~n7833 ;
  assign n7835 = \P1_state_reg[0]/NET0131  & ~n7834 ;
  assign n7836 = \P1_reg0_reg[23]/NET0131  & ~n3703 ;
  assign n7837 = ~n7835 & ~n7836 ;
  assign n7838 = \P1_reg0_reg[8]/NET0131  & ~n6238 ;
  assign n7839 = n6171 & ~n7496 ;
  assign n7840 = ~n7838 & ~n7839 ;
  assign n7841 = \P1_reg0_reg[9]/NET0131  & ~n3703 ;
  assign n7842 = \P1_reg0_reg[9]/NET0131  & n3664 ;
  assign n7844 = \P1_reg0_reg[9]/NET0131  & ~n3900 ;
  assign n7849 = n3900 & n6479 ;
  assign n7850 = ~n7844 & ~n7849 ;
  assign n7851 = n1898 & ~n7850 ;
  assign n7845 = n3900 & n6485 ;
  assign n7846 = ~n7844 & ~n7845 ;
  assign n7847 = n3557 & ~n7846 ;
  assign n7843 = \P1_reg0_reg[9]/NET0131  & ~n4725 ;
  assign n7848 = n3900 & ~n7509 ;
  assign n7852 = ~n7843 & ~n7848 ;
  assign n7853 = ~n7847 & n7852 ;
  assign n7854 = ~n7851 & n7853 ;
  assign n7855 = n3662 & ~n7854 ;
  assign n7856 = ~n7842 & ~n7855 ;
  assign n7857 = \P1_state_reg[0]/NET0131  & ~n7856 ;
  assign n7858 = ~n7841 & ~n7857 ;
  assign n7859 = \P1_reg1_reg[18]/NET0131  & ~n3703 ;
  assign n7860 = \P1_reg1_reg[18]/NET0131  & n3664 ;
  assign n7862 = \P1_reg1_reg[18]/NET0131  & ~n4236 ;
  assign n7866 = n4236 & ~n5789 ;
  assign n7867 = ~n7862 & ~n7866 ;
  assign n7868 = n3575 & ~n7867 ;
  assign n7863 = n4236 & n5783 ;
  assign n7864 = ~n7862 & ~n7863 ;
  assign n7865 = n3557 & ~n7864 ;
  assign n7869 = n4236 & n5798 ;
  assign n7870 = ~n7862 & ~n7869 ;
  assign n7871 = n1898 & ~n7870 ;
  assign n7861 = \P1_reg1_reg[18]/NET0131  & ~n4753 ;
  assign n7872 = n4236 & ~n6641 ;
  assign n7873 = ~n7861 & ~n7872 ;
  assign n7874 = ~n7871 & n7873 ;
  assign n7875 = ~n7865 & n7874 ;
  assign n7876 = ~n7868 & n7875 ;
  assign n7877 = n3662 & ~n7876 ;
  assign n7878 = ~n7860 & ~n7877 ;
  assign n7879 = \P1_state_reg[0]/NET0131  & ~n7878 ;
  assign n7880 = ~n7859 & ~n7879 ;
  assign n7881 = \P1_reg1_reg[19]/NET0131  & ~n3703 ;
  assign n7882 = \P1_reg1_reg[19]/NET0131  & n3664 ;
  assign n7884 = \P1_reg1_reg[19]/NET0131  & ~n4236 ;
  assign n7888 = n4236 & n6355 ;
  assign n7889 = ~n7884 & ~n7888 ;
  assign n7890 = n1898 & ~n7889 ;
  assign n7885 = n4236 & n6347 ;
  assign n7886 = ~n7884 & ~n7885 ;
  assign n7887 = n3575 & ~n7886 ;
  assign n7892 = n4236 & n6362 ;
  assign n7893 = ~n7884 & ~n7892 ;
  assign n7894 = n3557 & ~n7893 ;
  assign n7883 = \P1_reg1_reg[19]/NET0131  & ~n4753 ;
  assign n7891 = n4236 & ~n7796 ;
  assign n7895 = ~n7883 & ~n7891 ;
  assign n7896 = ~n7894 & n7895 ;
  assign n7897 = ~n7887 & n7896 ;
  assign n7898 = ~n7890 & n7897 ;
  assign n7899 = n3662 & ~n7898 ;
  assign n7900 = ~n7882 & ~n7899 ;
  assign n7901 = \P1_state_reg[0]/NET0131  & ~n7900 ;
  assign n7902 = ~n7881 & ~n7901 ;
  assign n7904 = \P1_reg1_reg[22]/NET0131  & ~n4236 ;
  assign n7905 = n6246 & ~n6564 ;
  assign n7906 = ~n7904 & ~n7905 ;
  assign n7907 = n3557 & ~n7906 ;
  assign n7903 = n6246 & ~n7810 ;
  assign n7908 = n4753 & n6070 ;
  assign n7909 = ~n6241 & n7908 ;
  assign n7910 = ~n4751 & n7909 ;
  assign n7911 = \P1_reg1_reg[22]/NET0131  & ~n7910 ;
  assign n7912 = ~n7903 & ~n7911 ;
  assign n7913 = ~n7907 & n7912 ;
  assign n7914 = \P1_reg1_reg[23]/NET0131  & ~n3703 ;
  assign n7915 = \P1_reg1_reg[23]/NET0131  & ~n4236 ;
  assign n7916 = n4236 & n7337 ;
  assign n7917 = ~n7915 & ~n7916 ;
  assign n7918 = n3575 & ~n7917 ;
  assign n7919 = n4236 & ~n7348 ;
  assign n7920 = ~n7915 & ~n7919 ;
  assign n7921 = n3557 & ~n7920 ;
  assign n7922 = n4236 & ~n7600 ;
  assign n7923 = ~n4751 & n6889 ;
  assign n7924 = \P1_reg1_reg[23]/NET0131  & ~n7923 ;
  assign n7925 = ~n7922 & ~n7924 ;
  assign n7926 = ~n7921 & n7925 ;
  assign n7927 = ~n7918 & n7926 ;
  assign n7928 = n3662 & ~n7927 ;
  assign n7929 = \P1_reg1_reg[23]/NET0131  & n3664 ;
  assign n7930 = ~n7928 & ~n7929 ;
  assign n7931 = \P1_state_reg[0]/NET0131  & ~n7930 ;
  assign n7932 = ~n7914 & ~n7931 ;
  assign n7933 = \P2_reg0_reg[12]/NET0131  & ~n3434 ;
  assign n7935 = \P2_reg0_reg[12]/NET0131  & ~n4610 ;
  assign n7936 = n4610 & ~n6388 ;
  assign n7937 = ~n7935 & ~n7936 ;
  assign n7938 = n3319 & ~n7937 ;
  assign n7939 = n4610 & n6397 ;
  assign n7940 = ~n7935 & ~n7939 ;
  assign n7941 = n3373 & ~n7940 ;
  assign n7942 = n4610 & n6403 ;
  assign n7943 = ~n7935 & ~n7942 ;
  assign n7944 = n3179 & ~n7943 ;
  assign n7945 = n4610 & ~n6407 ;
  assign n7946 = ~n6408 & n7945 ;
  assign n7947 = ~n7935 & ~n7946 ;
  assign n7948 = n3409 & ~n7947 ;
  assign n7934 = \P2_reg0_reg[12]/NET0131  & ~n4619 ;
  assign n7949 = n2954 & n4610 ;
  assign n7950 = ~n7935 & ~n7949 ;
  assign n7951 = n3375 & ~n7950 ;
  assign n7952 = ~n7934 & ~n7951 ;
  assign n7953 = ~n7948 & n7952 ;
  assign n7954 = ~n7944 & n7953 ;
  assign n7955 = ~n7941 & n7954 ;
  assign n7956 = ~n7938 & n7955 ;
  assign n7957 = n2017 & ~n7956 ;
  assign n7958 = \P2_reg0_reg[12]/NET0131  & n3430 ;
  assign n7959 = ~n7957 & ~n7958 ;
  assign n7960 = \P1_state_reg[0]/NET0131  & ~n7959 ;
  assign n7961 = ~n7933 & ~n7960 ;
  assign n7962 = \P2_reg0_reg[16]/NET0131  & ~n3434 ;
  assign n7963 = \P2_reg0_reg[16]/NET0131  & n3430 ;
  assign n7965 = \P2_reg0_reg[16]/NET0131  & ~n4610 ;
  assign n7972 = n4610 & n6435 ;
  assign n7973 = ~n7965 & ~n7972 ;
  assign n7974 = n3373 & ~n7973 ;
  assign n7966 = n4610 & ~n6449 ;
  assign n7967 = ~n7965 & ~n7966 ;
  assign n7968 = n3319 & ~n7967 ;
  assign n7964 = n4610 & ~n7622 ;
  assign n7969 = n3179 & ~n4610 ;
  assign n7970 = n5258 & ~n7969 ;
  assign n7971 = \P2_reg0_reg[16]/NET0131  & ~n7970 ;
  assign n7975 = ~n7964 & ~n7971 ;
  assign n7976 = ~n7968 & n7975 ;
  assign n7977 = ~n7974 & n7976 ;
  assign n7978 = n2017 & ~n7977 ;
  assign n7979 = ~n7963 & ~n7978 ;
  assign n7980 = \P1_state_reg[0]/NET0131  & ~n7979 ;
  assign n7981 = ~n7962 & ~n7980 ;
  assign n7982 = ~n5257 & n7534 ;
  assign n7983 = \P2_reg0_reg[20]/NET0131  & ~n7982 ;
  assign n7984 = n5385 & ~n7314 ;
  assign n7985 = ~n7983 & ~n7984 ;
  assign n7987 = n1045 & n3664 ;
  assign n8005 = n1026 & ~n5741 ;
  assign n8006 = ~n7036 & ~n8005 ;
  assign n8007 = ~n536 & ~n8006 ;
  assign n8008 = n536 & n1075 ;
  assign n8009 = ~n8007 & ~n8008 ;
  assign n8010 = n3450 & ~n8009 ;
  assign n8004 = ~n1045 & ~n3450 ;
  assign n8011 = n1898 & ~n8004 ;
  assign n8012 = ~n8010 & n8011 ;
  assign n7997 = ~n1766 & n3837 ;
  assign n7996 = n1766 & ~n3837 ;
  assign n7998 = n3575 & ~n7996 ;
  assign n7999 = ~n7997 & n7998 ;
  assign n7989 = ~n1064 & ~n4835 ;
  assign n7990 = n3650 & ~n4836 ;
  assign n7991 = ~n7989 & n7990 ;
  assign n7993 = ~n1766 & ~n3753 ;
  assign n7992 = n1766 & n3753 ;
  assign n7994 = n3557 & ~n7992 ;
  assign n7995 = ~n7993 & n7994 ;
  assign n8000 = ~n7991 & ~n7995 ;
  assign n8001 = ~n7999 & n8000 ;
  assign n8002 = n3450 & ~n8001 ;
  assign n7988 = ~n1064 & n3655 ;
  assign n8003 = n1045 & ~n7033 ;
  assign n8013 = ~n7988 & ~n8003 ;
  assign n8014 = ~n8002 & n8013 ;
  assign n8015 = ~n8012 & n8014 ;
  assign n8016 = n3662 & ~n8015 ;
  assign n8017 = ~n7987 & ~n8016 ;
  assign n8018 = \P1_state_reg[0]/NET0131  & ~n8017 ;
  assign n7986 = n1045 & n1934 ;
  assign n8019 = \P1_reg3_reg[13]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8020 = ~n7986 & ~n8019 ;
  assign n8021 = ~n8018 & n8020 ;
  assign n8023 = n2905 & n3430 ;
  assign n8025 = n2905 & ~n4925 ;
  assign n8026 = n2937 & ~n7110 ;
  assign n8027 = ~n3342 & ~n8026 ;
  assign n8028 = ~n2050 & ~n8027 ;
  assign n8029 = n2050 & n2965 ;
  assign n8030 = ~n8028 & ~n8029 ;
  assign n8031 = n4925 & n8030 ;
  assign n8032 = ~n8025 & ~n8031 ;
  assign n8033 = n3373 & ~n8032 ;
  assign n8034 = n4139 & ~n4391 ;
  assign n8035 = ~n4139 & n4391 ;
  assign n8036 = ~n8034 & ~n8035 ;
  assign n8037 = n4925 & n8036 ;
  assign n8038 = ~n8025 & ~n8037 ;
  assign n8039 = n3179 & ~n8038 ;
  assign n8044 = n4139 & ~n4349 ;
  assign n8045 = ~n4139 & n4349 ;
  assign n8046 = ~n8044 & ~n8045 ;
  assign n8047 = n4925 & ~n8046 ;
  assign n8048 = ~n8025 & ~n8047 ;
  assign n8049 = n3319 & ~n8048 ;
  assign n8040 = n2926 & ~n7125 ;
  assign n8041 = ~n3387 & n3409 ;
  assign n8042 = ~n8040 & n8041 ;
  assign n8043 = n4925 & n8042 ;
  assign n8024 = n2905 & n4934 ;
  assign n8050 = n2926 & ~n5093 ;
  assign n8051 = ~n8024 & ~n8050 ;
  assign n8052 = ~n8043 & n8051 ;
  assign n8053 = ~n8049 & n8052 ;
  assign n8054 = ~n8039 & n8053 ;
  assign n8055 = ~n8033 & n8054 ;
  assign n8056 = n2017 & ~n8055 ;
  assign n8057 = ~n8023 & ~n8056 ;
  assign n8058 = \P1_state_reg[0]/NET0131  & ~n8057 ;
  assign n8022 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[11]/NET0131  ;
  assign n8059 = n2905 & n3935 ;
  assign n8060 = ~n8022 & ~n8059 ;
  assign n8061 = ~n8058 & n8060 ;
  assign n8064 = n3077 & n3430 ;
  assign n8066 = n3077 & ~n4925 ;
  assign n8067 = ~n3096 & ~n3124 ;
  assign n8068 = n6031 & n8067 ;
  assign n8069 = ~n6031 & ~n8067 ;
  assign n8070 = ~n8068 & ~n8069 ;
  assign n8071 = n4925 & n8070 ;
  assign n8072 = ~n8066 & ~n8071 ;
  assign n8073 = n3319 & ~n8072 ;
  assign n8080 = n3056 & ~n3344 ;
  assign n8081 = ~n5821 & ~n8080 ;
  assign n8082 = ~n2050 & ~n8081 ;
  assign n8083 = n2050 & n3105 ;
  assign n8084 = ~n8082 & ~n8083 ;
  assign n8085 = n4925 & n8084 ;
  assign n8086 = ~n8066 & ~n8085 ;
  assign n8087 = n3373 & ~n8086 ;
  assign n8074 = n5283 & n8067 ;
  assign n8075 = ~n5283 & ~n8067 ;
  assign n8076 = ~n8074 & ~n8075 ;
  assign n8077 = n4925 & ~n8076 ;
  assign n8078 = ~n8066 & ~n8077 ;
  assign n8079 = n3179 & ~n8078 ;
  assign n8088 = n3095 & ~n3389 ;
  assign n8089 = n3409 & ~n6453 ;
  assign n8090 = ~n8088 & n8089 ;
  assign n8091 = n4925 & n8090 ;
  assign n8065 = n3077 & n4934 ;
  assign n8092 = n3095 & ~n5093 ;
  assign n8093 = ~n8065 & ~n8092 ;
  assign n8094 = ~n8091 & n8093 ;
  assign n8095 = ~n8079 & n8094 ;
  assign n8096 = ~n8087 & n8095 ;
  assign n8097 = ~n8073 & n8096 ;
  assign n8098 = n2017 & ~n8097 ;
  assign n8099 = ~n8064 & ~n8098 ;
  assign n8100 = \P1_state_reg[0]/NET0131  & ~n8099 ;
  assign n8062 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[14]/NET0131  ;
  assign n8063 = n3077 & n3935 ;
  assign n8101 = ~n8062 & ~n8063 ;
  assign n8102 = ~n8100 & n8101 ;
  assign n8103 = n1291 & n3664 ;
  assign n8104 = n1274 & ~n3581 ;
  assign n8105 = ~n7279 & ~n8104 ;
  assign n8106 = ~n536 & ~n8105 ;
  assign n8107 = n536 & n1322 ;
  assign n8108 = ~n8106 & ~n8107 ;
  assign n8127 = n3450 & ~n8108 ;
  assign n8128 = n1898 & ~n8127 ;
  assign n8129 = n3618 & ~n7032 ;
  assign n8130 = ~n8128 & n8129 ;
  assign n8131 = n1291 & ~n8130 ;
  assign n8109 = n1898 & n8108 ;
  assign n8119 = n1406 & n1753 ;
  assign n8118 = ~n1406 & ~n1753 ;
  assign n8120 = n3575 & ~n8118 ;
  assign n8121 = ~n8119 & n8120 ;
  assign n8115 = ~n1753 & n3478 ;
  assign n8114 = n1753 & ~n3478 ;
  assign n8116 = n3557 & ~n8114 ;
  assign n8117 = ~n8115 & n8116 ;
  assign n8110 = ~n1313 & n3683 ;
  assign n8111 = ~n1313 & ~n3628 ;
  assign n8112 = ~n3629 & n3650 ;
  assign n8113 = ~n8111 & n8112 ;
  assign n8122 = ~n8110 & ~n8113 ;
  assign n8123 = ~n8117 & n8122 ;
  assign n8124 = ~n8121 & n8123 ;
  assign n8125 = ~n8109 & n8124 ;
  assign n8126 = n3450 & ~n8125 ;
  assign n8132 = ~n1313 & n1736 ;
  assign n8133 = ~n8126 & ~n8132 ;
  assign n8134 = ~n8131 & n8133 ;
  assign n8135 = n3662 & ~n8134 ;
  assign n8136 = ~n8103 & ~n8135 ;
  assign n8137 = \P1_state_reg[0]/NET0131  & ~n8136 ;
  assign n8138 = \P1_state_reg[0]/NET0131  & ~n1291 ;
  assign n8139 = ~\P1_reg3_reg[4]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8140 = ~n8138 & ~n8139 ;
  assign n8141 = ~n3703 & n8140 ;
  assign n8142 = ~n8137 & ~n8141 ;
  assign n8145 = n2674 & n3430 ;
  assign n8147 = n2674 & ~n4925 ;
  assign n8154 = n2050 & ~n2702 ;
  assign n8155 = ~n2678 & n3337 ;
  assign n8156 = n2990 & ~n8155 ;
  assign n8157 = ~n2050 & ~n3339 ;
  assign n8158 = ~n8156 & n8157 ;
  assign n8159 = ~n8154 & ~n8158 ;
  assign n8160 = n4925 & ~n8159 ;
  assign n8161 = ~n8147 & ~n8160 ;
  assign n8162 = n3373 & ~n8161 ;
  assign n8148 = n4105 & n4123 ;
  assign n8149 = ~n4105 & ~n4123 ;
  assign n8150 = ~n8148 & ~n8149 ;
  assign n8151 = n4925 & n8150 ;
  assign n8152 = ~n8147 & ~n8151 ;
  assign n8153 = n3319 & ~n8152 ;
  assign n8163 = n4123 & n5146 ;
  assign n8164 = ~n4123 & ~n5146 ;
  assign n8165 = ~n8163 & ~n8164 ;
  assign n8166 = n4925 & ~n8165 ;
  assign n8167 = ~n8147 & ~n8166 ;
  assign n8168 = n3179 & ~n8167 ;
  assign n8169 = n2692 & ~n3383 ;
  assign n8170 = ~n3384 & n3409 ;
  assign n8171 = ~n8169 & n8170 ;
  assign n8172 = n4925 & n8171 ;
  assign n8146 = n2674 & n4934 ;
  assign n8173 = n2692 & ~n5093 ;
  assign n8174 = ~n8146 & ~n8173 ;
  assign n8175 = ~n8172 & n8174 ;
  assign n8176 = ~n8168 & n8175 ;
  assign n8177 = ~n8153 & n8176 ;
  assign n8178 = ~n8162 & n8177 ;
  assign n8179 = n2017 & ~n8178 ;
  assign n8180 = ~n8145 & ~n8179 ;
  assign n8181 = \P1_state_reg[0]/NET0131  & ~n8180 ;
  assign n8143 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[8]/NET0131  ;
  assign n8144 = n2674 & n3935 ;
  assign n8182 = ~n8143 & ~n8144 ;
  assign n8183 = ~n8181 & n8182 ;
  assign n8185 = n1270 & n3664 ;
  assign n8186 = n1222 & ~n7279 ;
  assign n8187 = ~n7280 & ~n8186 ;
  assign n8188 = ~n536 & ~n8187 ;
  assign n8189 = n536 & n1298 ;
  assign n8190 = ~n8188 & ~n8189 ;
  assign n8209 = n3450 & ~n8190 ;
  assign n8210 = n1898 & ~n8209 ;
  assign n8211 = n8129 & ~n8210 ;
  assign n8212 = n1270 & ~n8211 ;
  assign n8191 = n1898 & n8190 ;
  assign n8201 = ~n1758 & n3733 ;
  assign n8200 = n1758 & ~n3733 ;
  assign n8202 = n3557 & ~n8200 ;
  assign n8203 = ~n8201 & n8202 ;
  assign n8197 = ~n1758 & n3823 ;
  assign n8196 = n1758 & ~n3823 ;
  assign n8198 = n3575 & ~n8196 ;
  assign n8199 = ~n8197 & n8198 ;
  assign n8192 = ~n1288 & n3683 ;
  assign n8193 = ~n1288 & ~n3629 ;
  assign n8194 = ~n3630 & n3650 ;
  assign n8195 = ~n8193 & n8194 ;
  assign n8204 = ~n8192 & ~n8195 ;
  assign n8205 = ~n8199 & n8204 ;
  assign n8206 = ~n8203 & n8205 ;
  assign n8207 = ~n8191 & n8206 ;
  assign n8208 = n3450 & ~n8207 ;
  assign n8213 = ~n1288 & n1736 ;
  assign n8214 = ~n8208 & ~n8213 ;
  assign n8215 = ~n8212 & n8214 ;
  assign n8216 = n3662 & ~n8215 ;
  assign n8217 = ~n8185 & ~n8216 ;
  assign n8218 = \P1_state_reg[0]/NET0131  & ~n8217 ;
  assign n8184 = \P1_reg3_reg[5]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8219 = n1270 & n1934 ;
  assign n8220 = ~n8184 & ~n8219 ;
  assign n8221 = ~n8218 & n8220 ;
  assign n8222 = \P2_reg0_reg[23]/NET0131  & ~n3434 ;
  assign n8223 = \P2_reg0_reg[23]/NET0131  & n3430 ;
  assign n8224 = \P2_reg0_reg[23]/NET0131  & ~n4610 ;
  assign n8228 = n4610 & ~n7439 ;
  assign n8229 = ~n8224 & ~n8228 ;
  assign n8230 = n3319 & ~n8229 ;
  assign n8225 = n4610 & ~n7432 ;
  assign n8226 = ~n8224 & ~n8225 ;
  assign n8227 = n3179 & ~n8226 ;
  assign n8232 = n4610 & n7448 ;
  assign n8233 = ~n8224 & ~n8232 ;
  assign n8234 = n3373 & ~n8233 ;
  assign n8231 = \P2_reg0_reg[23]/NET0131  & ~n5258 ;
  assign n8235 = n4610 & ~n7740 ;
  assign n8236 = ~n8231 & ~n8235 ;
  assign n8237 = ~n8234 & n8236 ;
  assign n8238 = ~n8227 & n8237 ;
  assign n8239 = ~n8230 & n8238 ;
  assign n8240 = n2017 & ~n8239 ;
  assign n8241 = ~n8223 & ~n8240 ;
  assign n8242 = \P1_state_reg[0]/NET0131  & ~n8241 ;
  assign n8243 = ~n8222 & ~n8242 ;
  assign n8244 = \P1_reg2_reg[10]/NET0131  & ~n3703 ;
  assign n8245 = \P1_reg2_reg[10]/NET0131  & n3664 ;
  assign n8247 = \P1_reg2_reg[10]/NET0131  & ~n3672 ;
  assign n8248 = n3672 & n6987 ;
  assign n8249 = ~n8247 & ~n8248 ;
  assign n8250 = n1898 & ~n8249 ;
  assign n8254 = n3672 & ~n6999 ;
  assign n8255 = ~n8247 & ~n8254 ;
  assign n8256 = n3557 & ~n8255 ;
  assign n8251 = n3672 & n6993 ;
  assign n8252 = ~n8247 & ~n8251 ;
  assign n8253 = n3575 & ~n8252 ;
  assign n8246 = n3672 & ~n6980 ;
  assign n8257 = n1132 & n1736 ;
  assign n8258 = \P1_reg2_reg[10]/NET0131  & ~n5428 ;
  assign n8259 = ~n8257 & ~n8258 ;
  assign n8260 = ~n8246 & n8259 ;
  assign n8261 = ~n8253 & n8260 ;
  assign n8262 = ~n8256 & n8261 ;
  assign n8263 = ~n8250 & n8262 ;
  assign n8264 = n3662 & ~n8263 ;
  assign n8265 = ~n8245 & ~n8264 ;
  assign n8266 = \P1_state_reg[0]/NET0131  & ~n8265 ;
  assign n8267 = ~n8244 & ~n8266 ;
  assign n8268 = \P1_reg2_reg[11]/NET0131  & ~n3703 ;
  assign n8269 = \P1_reg2_reg[11]/NET0131  & n3664 ;
  assign n8271 = \P1_reg2_reg[11]/NET0131  & ~n3672 ;
  assign n8282 = n3672 & n6942 ;
  assign n8283 = ~n8271 & ~n8282 ;
  assign n8284 = n1898 & ~n8283 ;
  assign n8272 = n3672 & ~n6948 ;
  assign n8273 = ~n8271 & ~n8272 ;
  assign n8274 = n3557 & ~n8273 ;
  assign n8275 = n1128 & n6977 ;
  assign n8276 = ~n498 & ~n6953 ;
  assign n8277 = ~n1128 & n3616 ;
  assign n8278 = ~n8276 & n8277 ;
  assign n8279 = ~n8275 & ~n8278 ;
  assign n8280 = ~n6960 & n8279 ;
  assign n8281 = n3672 & ~n8280 ;
  assign n8270 = \P1_reg2_reg[11]/NET0131  & ~n5430 ;
  assign n8285 = n1111 & n1736 ;
  assign n8286 = ~n8270 & ~n8285 ;
  assign n8287 = ~n8281 & n8286 ;
  assign n8288 = ~n8274 & n8287 ;
  assign n8289 = ~n8284 & n8288 ;
  assign n8290 = n3662 & ~n8289 ;
  assign n8291 = ~n8269 & ~n8290 ;
  assign n8292 = \P1_state_reg[0]/NET0131  & ~n8291 ;
  assign n8293 = ~n8268 & ~n8292 ;
  assign n8294 = \P1_reg2_reg[13]/NET0131  & ~n7699 ;
  assign n8295 = n1045 & n1736 ;
  assign n8296 = n1898 & n8009 ;
  assign n8297 = ~n1064 & n3683 ;
  assign n8298 = n8001 & ~n8297 ;
  assign n8299 = ~n8296 & n8298 ;
  assign n8300 = n3672 & ~n8299 ;
  assign n8301 = ~n8295 & ~n8300 ;
  assign n8302 = n6070 & ~n8301 ;
  assign n8303 = ~n8294 & ~n8302 ;
  assign n8304 = \P1_reg2_reg[14]/NET0131  & ~n3703 ;
  assign n8305 = \P1_reg2_reg[14]/NET0131  & n3664 ;
  assign n8307 = ~n1040 & n3683 ;
  assign n8308 = n7030 & ~n8307 ;
  assign n8309 = n1898 & n7041 ;
  assign n8310 = n8308 & ~n8309 ;
  assign n8311 = n3672 & ~n8310 ;
  assign n8306 = \P1_reg2_reg[14]/NET0131  & ~n7698 ;
  assign n8312 = n1021 & n1736 ;
  assign n8313 = ~n8306 & ~n8312 ;
  assign n8314 = ~n8311 & n8313 ;
  assign n8315 = n3662 & ~n8314 ;
  assign n8316 = ~n8305 & ~n8315 ;
  assign n8317 = \P1_state_reg[0]/NET0131  & ~n8316 ;
  assign n8318 = ~n8304 & ~n8317 ;
  assign n8319 = \P1_reg2_reg[15]/NET0131  & ~n3703 ;
  assign n8320 = \P1_reg2_reg[15]/NET0131  & n3664 ;
  assign n8322 = \P1_reg2_reg[15]/NET0131  & ~n3672 ;
  assign n8323 = n3672 & n7063 ;
  assign n8324 = ~n8322 & ~n8323 ;
  assign n8325 = n3557 & ~n8324 ;
  assign n8329 = n3672 & ~n7077 ;
  assign n8330 = ~n8322 & ~n8329 ;
  assign n8331 = n3575 & ~n8330 ;
  assign n8326 = n3672 & n7071 ;
  assign n8327 = ~n8322 & ~n8326 ;
  assign n8328 = n1898 & ~n8327 ;
  assign n8332 = n3672 & n7082 ;
  assign n8333 = ~n8322 & ~n8332 ;
  assign n8334 = n3650 & ~n8333 ;
  assign n8336 = ~n1015 & n3683 ;
  assign n8337 = n3672 & n8336 ;
  assign n8321 = \P1_reg2_reg[15]/NET0131  & ~n3685 ;
  assign n8335 = n994 & n1736 ;
  assign n8338 = ~n8321 & ~n8335 ;
  assign n8339 = ~n8337 & n8338 ;
  assign n8340 = ~n8334 & n8339 ;
  assign n8341 = ~n8328 & n8340 ;
  assign n8342 = ~n8331 & n8341 ;
  assign n8343 = ~n8325 & n8342 ;
  assign n8344 = n3662 & ~n8343 ;
  assign n8345 = ~n8320 & ~n8344 ;
  assign n8346 = \P1_state_reg[0]/NET0131  & ~n8345 ;
  assign n8347 = ~n8319 & ~n8346 ;
  assign n8348 = \P2_reg0_reg[9]/NET0131  & ~n3434 ;
  assign n8349 = \P2_reg0_reg[9]/NET0131  & n3430 ;
  assign n8351 = \P2_reg0_reg[9]/NET0131  & ~n4610 ;
  assign n8352 = n4610 & n7241 ;
  assign n8353 = ~n8351 & ~n8352 ;
  assign n8354 = n3373 & ~n8353 ;
  assign n8358 = n4610 & ~n7254 ;
  assign n8359 = ~n8351 & ~n8358 ;
  assign n8360 = n3319 & ~n8359 ;
  assign n8355 = n4610 & n7247 ;
  assign n8356 = ~n8351 & ~n8355 ;
  assign n8357 = n3179 & ~n8356 ;
  assign n8350 = n4610 & ~n7234 ;
  assign n8361 = \P2_reg0_reg[9]/NET0131  & ~n4621 ;
  assign n8362 = ~n8350 & ~n8361 ;
  assign n8363 = ~n8357 & n8362 ;
  assign n8364 = ~n8360 & n8363 ;
  assign n8365 = ~n8354 & n8364 ;
  assign n8366 = n2017 & ~n8365 ;
  assign n8367 = ~n8349 & ~n8366 ;
  assign n8368 = \P1_state_reg[0]/NET0131  & ~n8367 ;
  assign n8369 = ~n8348 & ~n8368 ;
  assign n8370 = \P2_reg1_reg[10]/NET0131  & ~n3434 ;
  assign n8371 = \P2_reg1_reg[10]/NET0131  & n3430 ;
  assign n8373 = \P2_reg1_reg[10]/NET0131  & ~n4663 ;
  assign n8377 = n4663 & n7114 ;
  assign n8378 = ~n8373 & ~n8377 ;
  assign n8379 = n3373 & ~n8378 ;
  assign n8374 = n4663 & ~n7104 ;
  assign n8375 = ~n8373 & ~n8374 ;
  assign n8376 = n3319 & ~n8375 ;
  assign n8380 = n4663 & n7120 ;
  assign n8381 = ~n8373 & ~n8380 ;
  assign n8382 = n3179 & ~n8381 ;
  assign n8372 = \P2_reg1_reg[10]/NET0131  & ~n5509 ;
  assign n8383 = n2980 & n3375 ;
  assign n8384 = ~n7128 & ~n8383 ;
  assign n8385 = n4663 & ~n8384 ;
  assign n8386 = ~n8372 & ~n8385 ;
  assign n8387 = ~n8382 & n8386 ;
  assign n8388 = ~n8376 & n8387 ;
  assign n8389 = ~n8379 & n8388 ;
  assign n8390 = n2017 & ~n8389 ;
  assign n8391 = ~n8371 & ~n8390 ;
  assign n8392 = \P1_state_reg[0]/NET0131  & ~n8391 ;
  assign n8393 = ~n8370 & ~n8392 ;
  assign n8394 = \P2_reg1_reg[13]/NET0131  & ~n3434 ;
  assign n8395 = \P2_reg1_reg[13]/NET0131  & n3430 ;
  assign n8397 = \P2_reg1_reg[13]/NET0131  & ~n4663 ;
  assign n8398 = n4663 & n7156 ;
  assign n8399 = ~n8397 & ~n8398 ;
  assign n8400 = n3373 & ~n8399 ;
  assign n8404 = n4663 & n7170 ;
  assign n8405 = ~n8397 & ~n8404 ;
  assign n8406 = n3179 & ~n8405 ;
  assign n8401 = n4663 & ~n7163 ;
  assign n8402 = ~n8397 & ~n8401 ;
  assign n8403 = n3319 & ~n8402 ;
  assign n8396 = n4663 & n7149 ;
  assign n8407 = \P2_reg1_reg[13]/NET0131  & ~n5509 ;
  assign n8408 = ~n8396 & ~n8407 ;
  assign n8409 = ~n8403 & n8408 ;
  assign n8410 = ~n8406 & n8409 ;
  assign n8411 = ~n8400 & n8410 ;
  assign n8412 = n2017 & ~n8411 ;
  assign n8413 = ~n8395 & ~n8412 ;
  assign n8414 = \P1_state_reg[0]/NET0131  & ~n8413 ;
  assign n8415 = ~n8394 & ~n8414 ;
  assign n8416 = \P2_reg1_reg[15]/NET0131  & ~n3434 ;
  assign n8417 = \P2_reg1_reg[15]/NET0131  & n3430 ;
  assign n8424 = \P2_reg1_reg[15]/NET0131  & ~n4663 ;
  assign n8428 = n4663 & n7201 ;
  assign n8429 = ~n8424 & ~n8428 ;
  assign n8430 = n3373 & ~n8429 ;
  assign n8425 = n4663 & n7193 ;
  assign n8426 = ~n8424 & ~n8425 ;
  assign n8427 = n3179 & ~n8426 ;
  assign n8418 = n3071 & n3375 ;
  assign n8419 = ~n7213 & ~n8418 ;
  assign n8420 = n3319 & ~n7207 ;
  assign n8421 = n8419 & ~n8420 ;
  assign n8422 = n4663 & ~n8421 ;
  assign n8423 = \P2_reg1_reg[15]/NET0131  & ~n6719 ;
  assign n8431 = ~n8422 & ~n8423 ;
  assign n8432 = ~n8427 & n8431 ;
  assign n8433 = ~n8430 & n8432 ;
  assign n8434 = n2017 & ~n8433 ;
  assign n8435 = ~n8417 & ~n8434 ;
  assign n8436 = \P1_state_reg[0]/NET0131  & ~n8435 ;
  assign n8437 = ~n8416 & ~n8436 ;
  assign n8438 = \P2_reg1_reg[23]/NET0131  & ~n3434 ;
  assign n8439 = \P2_reg1_reg[23]/NET0131  & n3430 ;
  assign n8440 = \P2_reg1_reg[23]/NET0131  & ~n4663 ;
  assign n8444 = n4663 & ~n7439 ;
  assign n8445 = ~n8440 & ~n8444 ;
  assign n8446 = n3319 & ~n8445 ;
  assign n8441 = n4663 & ~n7432 ;
  assign n8442 = ~n8440 & ~n8441 ;
  assign n8443 = n3179 & ~n8442 ;
  assign n8448 = n4663 & n7448 ;
  assign n8449 = ~n8440 & ~n8448 ;
  assign n8450 = n3373 & ~n8449 ;
  assign n8447 = \P2_reg1_reg[23]/NET0131  & ~n5509 ;
  assign n8451 = n4663 & ~n7740 ;
  assign n8452 = ~n8447 & ~n8451 ;
  assign n8453 = ~n8450 & n8452 ;
  assign n8454 = ~n8443 & n8453 ;
  assign n8455 = ~n8446 & n8454 ;
  assign n8456 = n2017 & ~n8455 ;
  assign n8457 = ~n8439 & ~n8456 ;
  assign n8458 = \P1_state_reg[0]/NET0131  & ~n8457 ;
  assign n8459 = ~n8438 & ~n8458 ;
  assign n8460 = \P2_reg1_reg[9]/NET0131  & ~n3434 ;
  assign n8461 = \P2_reg1_reg[9]/NET0131  & n3430 ;
  assign n8463 = \P2_reg1_reg[9]/NET0131  & ~n4663 ;
  assign n8464 = n4663 & n7241 ;
  assign n8465 = ~n8463 & ~n8464 ;
  assign n8466 = n3373 & ~n8465 ;
  assign n8470 = n4663 & ~n7254 ;
  assign n8471 = ~n8463 & ~n8470 ;
  assign n8472 = n3319 & ~n8471 ;
  assign n8467 = n4663 & n7247 ;
  assign n8468 = ~n8463 & ~n8467 ;
  assign n8469 = n3179 & ~n8468 ;
  assign n8462 = n4663 & ~n7234 ;
  assign n8473 = \P2_reg1_reg[9]/NET0131  & ~n5509 ;
  assign n8474 = ~n8462 & ~n8473 ;
  assign n8475 = ~n8469 & n8474 ;
  assign n8476 = ~n8472 & n8475 ;
  assign n8477 = ~n8466 & n8476 ;
  assign n8478 = n2017 & ~n8477 ;
  assign n8479 = ~n8461 & ~n8478 ;
  assign n8480 = \P1_state_reg[0]/NET0131  & ~n8479 ;
  assign n8481 = ~n8460 & ~n8480 ;
  assign n8482 = \P2_reg2_reg[10]/NET0131  & ~n3434 ;
  assign n8483 = \P2_reg2_reg[10]/NET0131  & n3430 ;
  assign n8485 = \P2_reg2_reg[10]/NET0131  & ~n2033 ;
  assign n8489 = n2033 & n7114 ;
  assign n8490 = ~n8485 & ~n8489 ;
  assign n8491 = n3373 & ~n8490 ;
  assign n8486 = n2033 & ~n7104 ;
  assign n8487 = ~n8485 & ~n8486 ;
  assign n8488 = n3319 & ~n8487 ;
  assign n8494 = n2033 & n7120 ;
  assign n8495 = ~n8485 & ~n8494 ;
  assign n8496 = n3179 & ~n8495 ;
  assign n8493 = n2033 & ~n8384 ;
  assign n8484 = n2961 & n3415 ;
  assign n8492 = \P2_reg2_reg[10]/NET0131  & ~n4436 ;
  assign n8497 = ~n8484 & ~n8492 ;
  assign n8498 = ~n8493 & n8497 ;
  assign n8499 = ~n8496 & n8498 ;
  assign n8500 = ~n8488 & n8499 ;
  assign n8501 = ~n8491 & n8500 ;
  assign n8502 = n2017 & ~n8501 ;
  assign n8503 = ~n8483 & ~n8502 ;
  assign n8504 = \P1_state_reg[0]/NET0131  & ~n8503 ;
  assign n8505 = ~n8482 & ~n8504 ;
  assign n8506 = \P2_reg2_reg[13]/NET0131  & ~n3434 ;
  assign n8507 = \P2_reg2_reg[13]/NET0131  & n3430 ;
  assign n8510 = \P2_reg2_reg[13]/NET0131  & ~n2033 ;
  assign n8511 = n2033 & n7156 ;
  assign n8512 = ~n8510 & ~n8511 ;
  assign n8513 = n3373 & ~n8512 ;
  assign n8518 = n2033 & n7170 ;
  assign n8519 = ~n8510 & ~n8518 ;
  assign n8520 = n3179 & ~n8519 ;
  assign n8514 = n2033 & ~n7163 ;
  assign n8515 = ~n8510 & ~n8514 ;
  assign n8516 = n3319 & ~n8515 ;
  assign n8509 = n2033 & n7149 ;
  assign n8508 = \P2_reg2_reg[13]/NET0131  & n3422 ;
  assign n8517 = n3099 & n3415 ;
  assign n8521 = ~n8508 & ~n8517 ;
  assign n8522 = ~n8509 & n8521 ;
  assign n8523 = ~n8516 & n8522 ;
  assign n8524 = ~n8520 & n8523 ;
  assign n8525 = ~n8513 & n8524 ;
  assign n8526 = n2017 & ~n8525 ;
  assign n8527 = ~n8507 & ~n8526 ;
  assign n8528 = \P1_state_reg[0]/NET0131  & ~n8527 ;
  assign n8529 = ~n8506 & ~n8528 ;
  assign n8530 = \P2_reg2_reg[15]/NET0131  & ~n3434 ;
  assign n8531 = \P2_reg2_reg[15]/NET0131  & n3430 ;
  assign n8533 = \P2_reg2_reg[15]/NET0131  & ~n2033 ;
  assign n8537 = n2033 & n7201 ;
  assign n8538 = ~n8533 & ~n8537 ;
  assign n8539 = n3373 & ~n8538 ;
  assign n8534 = n2033 & n7193 ;
  assign n8535 = ~n8533 & ~n8534 ;
  assign n8536 = n3179 & ~n8535 ;
  assign n8543 = n2033 & ~n8419 ;
  assign n8540 = n2033 & ~n7207 ;
  assign n8541 = ~n8533 & ~n8540 ;
  assign n8542 = n3319 & ~n8541 ;
  assign n8532 = n3051 & n3415 ;
  assign n8544 = \P2_reg2_reg[15]/NET0131  & ~n4436 ;
  assign n8545 = ~n8532 & ~n8544 ;
  assign n8546 = ~n8542 & n8545 ;
  assign n8547 = ~n8543 & n8546 ;
  assign n8548 = ~n8536 & n8547 ;
  assign n8549 = ~n8539 & n8548 ;
  assign n8550 = n2017 & ~n8549 ;
  assign n8551 = ~n8531 & ~n8550 ;
  assign n8552 = \P1_state_reg[0]/NET0131  & ~n8551 ;
  assign n8553 = ~n8530 & ~n8552 ;
  assign n8554 = \P1_reg2_reg[9]/NET0131  & ~n3703 ;
  assign n8555 = \P1_reg2_reg[9]/NET0131  & n3664 ;
  assign n8557 = \P1_reg2_reg[9]/NET0131  & ~n3672 ;
  assign n8558 = n3672 & n6479 ;
  assign n8559 = ~n8557 & ~n8558 ;
  assign n8560 = n1898 & ~n8559 ;
  assign n8564 = n3672 & n6485 ;
  assign n8565 = ~n8557 & ~n8564 ;
  assign n8566 = n3557 & ~n8565 ;
  assign n8561 = n3672 & ~n6491 ;
  assign n8562 = ~n8557 & ~n8561 ;
  assign n8563 = n3575 & ~n8562 ;
  assign n8568 = n1178 & n7290 ;
  assign n8569 = ~n498 & ~n6495 ;
  assign n8570 = ~n1178 & n3616 ;
  assign n8571 = ~n8569 & n8570 ;
  assign n8572 = ~n8568 & ~n8571 ;
  assign n8573 = n3672 & ~n8572 ;
  assign n8556 = \P1_reg2_reg[9]/NET0131  & ~n5428 ;
  assign n8567 = n1158 & n1736 ;
  assign n8574 = ~n8556 & ~n8567 ;
  assign n8575 = ~n8573 & n8574 ;
  assign n8576 = ~n8563 & n8575 ;
  assign n8577 = ~n8566 & n8576 ;
  assign n8578 = ~n8560 & n8577 ;
  assign n8579 = n3662 & ~n8578 ;
  assign n8580 = ~n8555 & ~n8579 ;
  assign n8581 = \P1_state_reg[0]/NET0131  & ~n8580 ;
  assign n8582 = ~n8554 & ~n8581 ;
  assign n8583 = \P2_reg2_reg[9]/NET0131  & ~n3434 ;
  assign n8584 = \P2_reg2_reg[9]/NET0131  & n3430 ;
  assign n8587 = \P2_reg2_reg[9]/NET0131  & ~n2033 ;
  assign n8588 = n2033 & n7241 ;
  assign n8589 = ~n8587 & ~n8588 ;
  assign n8590 = n3373 & ~n8589 ;
  assign n8595 = n2033 & ~n7254 ;
  assign n8596 = ~n8587 & ~n8595 ;
  assign n8597 = n3319 & ~n8596 ;
  assign n8591 = n2033 & n7247 ;
  assign n8592 = ~n8587 & ~n8591 ;
  assign n8593 = n3179 & ~n8592 ;
  assign n8586 = n2033 & ~n7234 ;
  assign n8585 = \P2_reg2_reg[9]/NET0131  & n3422 ;
  assign n8594 = n2984 & n3415 ;
  assign n8598 = ~n8585 & ~n8594 ;
  assign n8599 = ~n8586 & n8598 ;
  assign n8600 = ~n8593 & n8599 ;
  assign n8601 = ~n8597 & n8600 ;
  assign n8602 = ~n8590 & n8601 ;
  assign n8603 = n2017 & ~n8602 ;
  assign n8604 = ~n8584 & ~n8603 ;
  assign n8605 = \P1_state_reg[0]/NET0131  & ~n8604 ;
  assign n8606 = ~n8583 & ~n8605 ;
  assign n8607 = \P1_reg0_reg[15]/NET0131  & ~n3703 ;
  assign n8608 = \P1_reg0_reg[15]/NET0131  & n3664 ;
  assign n8610 = \P1_reg0_reg[15]/NET0131  & ~n3900 ;
  assign n8611 = n3900 & n7063 ;
  assign n8612 = ~n8610 & ~n8611 ;
  assign n8613 = n3557 & ~n8612 ;
  assign n8617 = n3900 & ~n7077 ;
  assign n8618 = ~n8610 & ~n8617 ;
  assign n8619 = n3575 & ~n8618 ;
  assign n8614 = n3900 & n7071 ;
  assign n8615 = ~n8610 & ~n8614 ;
  assign n8616 = n1898 & ~n8615 ;
  assign n8620 = n3900 & n7082 ;
  assign n8621 = ~n8610 & ~n8620 ;
  assign n8622 = n3650 & ~n8621 ;
  assign n8609 = n3900 & n8336 ;
  assign n8623 = \P1_reg0_reg[15]/NET0131  & ~n3917 ;
  assign n8624 = ~n8609 & ~n8623 ;
  assign n8625 = ~n8622 & n8624 ;
  assign n8626 = ~n8616 & n8625 ;
  assign n8627 = ~n8619 & n8626 ;
  assign n8628 = ~n8613 & n8627 ;
  assign n8629 = n3662 & ~n8628 ;
  assign n8630 = ~n8608 & ~n8629 ;
  assign n8631 = \P1_state_reg[0]/NET0131  & ~n8630 ;
  assign n8632 = ~n8607 & ~n8631 ;
  assign n8633 = \P1_reg1_reg[15]/NET0131  & ~n3703 ;
  assign n8634 = \P1_reg1_reg[15]/NET0131  & n3664 ;
  assign n8636 = \P1_reg1_reg[15]/NET0131  & ~n4236 ;
  assign n8637 = n4236 & n7063 ;
  assign n8638 = ~n8636 & ~n8637 ;
  assign n8639 = n3557 & ~n8638 ;
  assign n8643 = n4236 & ~n7077 ;
  assign n8644 = ~n8636 & ~n8643 ;
  assign n8645 = n3575 & ~n8644 ;
  assign n8640 = n4236 & n7071 ;
  assign n8641 = ~n8636 & ~n8640 ;
  assign n8642 = n1898 & ~n8641 ;
  assign n8646 = n4236 & n7082 ;
  assign n8647 = ~n8636 & ~n8646 ;
  assign n8648 = n3650 & ~n8647 ;
  assign n8635 = \P1_reg1_reg[15]/NET0131  & ~n4252 ;
  assign n8649 = n4236 & n8336 ;
  assign n8650 = ~n8635 & ~n8649 ;
  assign n8651 = ~n8648 & n8650 ;
  assign n8652 = ~n8642 & n8651 ;
  assign n8653 = ~n8645 & n8652 ;
  assign n8654 = ~n8639 & n8653 ;
  assign n8655 = n3662 & ~n8654 ;
  assign n8656 = ~n8634 & ~n8655 ;
  assign n8657 = \P1_state_reg[0]/NET0131  & ~n8656 ;
  assign n8658 = ~n8633 & ~n8657 ;
  assign n8659 = \P2_reg0_reg[10]/NET0131  & ~n3434 ;
  assign n8660 = \P2_reg0_reg[10]/NET0131  & n3430 ;
  assign n8662 = \P2_reg0_reg[10]/NET0131  & ~n4610 ;
  assign n8666 = n4610 & n7114 ;
  assign n8667 = ~n8662 & ~n8666 ;
  assign n8668 = n3373 & ~n8667 ;
  assign n8663 = n4610 & ~n7104 ;
  assign n8664 = ~n8662 & ~n8663 ;
  assign n8665 = n3319 & ~n8664 ;
  assign n8669 = n4610 & n7120 ;
  assign n8670 = ~n8662 & ~n8669 ;
  assign n8671 = n3179 & ~n8670 ;
  assign n8661 = n4610 & ~n8384 ;
  assign n8672 = \P2_reg0_reg[10]/NET0131  & ~n4621 ;
  assign n8673 = ~n8661 & ~n8672 ;
  assign n8674 = ~n8671 & n8673 ;
  assign n8675 = ~n8665 & n8674 ;
  assign n8676 = ~n8668 & n8675 ;
  assign n8677 = n2017 & ~n8676 ;
  assign n8678 = ~n8660 & ~n8677 ;
  assign n8679 = \P1_state_reg[0]/NET0131  & ~n8678 ;
  assign n8680 = ~n8659 & ~n8679 ;
  assign n8681 = \P2_reg0_reg[13]/NET0131  & ~n3434 ;
  assign n8682 = \P2_reg0_reg[13]/NET0131  & n3430 ;
  assign n8684 = \P2_reg0_reg[13]/NET0131  & ~n4610 ;
  assign n8685 = n4610 & n7156 ;
  assign n8686 = ~n8684 & ~n8685 ;
  assign n8687 = n3373 & ~n8686 ;
  assign n8691 = n4610 & n7170 ;
  assign n8692 = ~n8684 & ~n8691 ;
  assign n8693 = n3179 & ~n8692 ;
  assign n8688 = n4610 & ~n7163 ;
  assign n8689 = ~n8684 & ~n8688 ;
  assign n8690 = n3319 & ~n8689 ;
  assign n8683 = \P2_reg0_reg[13]/NET0131  & ~n4621 ;
  assign n8694 = n4610 & n7149 ;
  assign n8695 = ~n8683 & ~n8694 ;
  assign n8696 = ~n8690 & n8695 ;
  assign n8697 = ~n8693 & n8696 ;
  assign n8698 = ~n8687 & n8697 ;
  assign n8699 = n2017 & ~n8698 ;
  assign n8700 = ~n8682 & ~n8699 ;
  assign n8701 = \P1_state_reg[0]/NET0131  & ~n8700 ;
  assign n8702 = ~n8681 & ~n8701 ;
  assign n8703 = \P2_reg0_reg[15]/NET0131  & ~n3434 ;
  assign n8704 = \P2_reg0_reg[15]/NET0131  & n3430 ;
  assign n8707 = \P2_reg0_reg[15]/NET0131  & ~n4610 ;
  assign n8711 = n4610 & n7201 ;
  assign n8712 = ~n8707 & ~n8711 ;
  assign n8713 = n3373 & ~n8712 ;
  assign n8708 = n4610 & n7193 ;
  assign n8709 = ~n8707 & ~n8708 ;
  assign n8710 = n3179 & ~n8709 ;
  assign n8705 = \P2_reg0_reg[15]/NET0131  & ~n6901 ;
  assign n8706 = n4610 & ~n8421 ;
  assign n8714 = ~n8705 & ~n8706 ;
  assign n8715 = ~n8710 & n8714 ;
  assign n8716 = ~n8713 & n8715 ;
  assign n8717 = n2017 & ~n8716 ;
  assign n8718 = ~n8704 & ~n8717 ;
  assign n8719 = \P1_state_reg[0]/NET0131  & ~n8718 ;
  assign n8720 = ~n8703 & ~n8719 ;
  assign n8721 = n6070 & n6891 ;
  assign n8722 = \P1_reg1_reg[4]/NET0131  & ~n8721 ;
  assign n8723 = n6246 & ~n8125 ;
  assign n8724 = ~n8722 & ~n8723 ;
  assign n8726 = ~\P1_reg3_reg[3]/NET0131  & n3664 ;
  assign n8746 = n1298 & ~n3580 ;
  assign n8747 = ~n3581 & ~n8746 ;
  assign n8748 = ~n536 & ~n8747 ;
  assign n8749 = n536 & n1344 ;
  assign n8750 = ~n8748 & ~n8749 ;
  assign n8751 = n3450 & ~n8750 ;
  assign n8745 = \P1_reg3_reg[3]/NET0131  & ~n3450 ;
  assign n8752 = n1898 & ~n8745 ;
  assign n8753 = ~n8751 & n8752 ;
  assign n8735 = ~n1745 & n3730 ;
  assign n8733 = ~n3472 & ~n3729 ;
  assign n8734 = ~n1746 & ~n8733 ;
  assign n8736 = n3557 & ~n8734 ;
  assign n8737 = ~n8735 & n8736 ;
  assign n8728 = ~n1359 & ~n3819 ;
  assign n8730 = n1746 & ~n8728 ;
  assign n8729 = ~n1746 & n8728 ;
  assign n8731 = n3575 & ~n8729 ;
  assign n8732 = ~n8730 & n8731 ;
  assign n8738 = ~n1336 & ~n3627 ;
  assign n8739 = ~n3628 & n3650 ;
  assign n8740 = ~n8738 & n8739 ;
  assign n8741 = ~n8732 & ~n8740 ;
  assign n8742 = ~n8737 & n8741 ;
  assign n8743 = n3450 & ~n8742 ;
  assign n8727 = ~n1336 & n3655 ;
  assign n8744 = ~\P1_reg3_reg[3]/NET0131  & ~n8129 ;
  assign n8754 = ~n8727 & ~n8744 ;
  assign n8755 = ~n8743 & n8754 ;
  assign n8756 = ~n8753 & n8755 ;
  assign n8757 = n3662 & ~n8756 ;
  assign n8758 = ~n8726 & ~n8757 ;
  assign n8759 = \P1_state_reg[0]/NET0131  & ~n8758 ;
  assign n8725 = \P1_reg3_reg[3]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8760 = ~\P1_reg3_reg[3]/NET0131  & n1934 ;
  assign n8761 = ~n8725 & ~n8760 ;
  assign n8762 = ~n8759 & n8761 ;
  assign n8764 = n2853 & n3430 ;
  assign n8766 = n2755 & ~n3334 ;
  assign n8767 = ~n2755 & n3334 ;
  assign n8768 = ~n8766 & ~n8767 ;
  assign n8769 = ~n2050 & ~n8768 ;
  assign n8770 = n2050 & n2866 ;
  assign n8771 = ~n8769 & ~n8770 ;
  assign n8772 = n4925 & ~n8771 ;
  assign n8773 = ~n2853 & ~n4925 ;
  assign n8774 = n3373 & ~n8773 ;
  assign n8775 = ~n8772 & n8774 ;
  assign n8784 = ~n4141 & n5135 ;
  assign n8783 = n4141 & ~n5135 ;
  assign n8785 = n3179 & ~n8783 ;
  assign n8786 = ~n8784 & n8785 ;
  assign n8776 = ~n2849 & ~n3379 ;
  assign n8777 = ~n3380 & n3409 ;
  assign n8778 = ~n8776 & n8777 ;
  assign n8780 = n4097 & ~n4141 ;
  assign n8779 = ~n4097 & n4141 ;
  assign n8781 = n3319 & ~n8779 ;
  assign n8782 = ~n8780 & n8781 ;
  assign n8787 = ~n8778 & ~n8782 ;
  assign n8788 = ~n8786 & n8787 ;
  assign n8789 = n4925 & ~n8788 ;
  assign n8765 = n2853 & ~n5937 ;
  assign n8790 = ~n2849 & ~n5093 ;
  assign n8791 = ~n8765 & ~n8790 ;
  assign n8792 = ~n8789 & n8791 ;
  assign n8793 = ~n8775 & n8792 ;
  assign n8794 = n2017 & ~n8793 ;
  assign n8795 = ~n8764 & ~n8794 ;
  assign n8796 = \P1_state_reg[0]/NET0131  & ~n8795 ;
  assign n8763 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n8797 = n2853 & n3935 ;
  assign n8798 = ~n8763 & ~n8797 ;
  assign n8799 = ~n8796 & n8798 ;
  assign n8802 = n2749 & ~n4925 ;
  assign n8803 = n2730 & ~n8767 ;
  assign n8804 = ~n2730 & n8767 ;
  assign n8805 = ~n8803 & ~n8804 ;
  assign n8806 = ~n2050 & ~n8805 ;
  assign n8807 = n2050 & n2858 ;
  assign n8808 = ~n8806 & ~n8807 ;
  assign n8809 = n4925 & n8808 ;
  assign n8810 = ~n8802 & ~n8809 ;
  assign n8811 = n3373 & ~n8810 ;
  assign n8812 = n2888 & ~n4129 ;
  assign n8813 = ~n2888 & n4129 ;
  assign n8814 = ~n8812 & ~n8813 ;
  assign n8815 = n4925 & ~n8814 ;
  assign n8816 = ~n8802 & ~n8815 ;
  assign n8817 = n3179 & ~n8816 ;
  assign n8818 = n3215 & ~n4129 ;
  assign n8819 = ~n3215 & n4129 ;
  assign n8820 = ~n8818 & ~n8819 ;
  assign n8821 = n4925 & n8820 ;
  assign n8822 = ~n8802 & ~n8821 ;
  assign n8823 = n3319 & ~n8822 ;
  assign n8824 = n2768 & ~n3380 ;
  assign n8825 = ~n3381 & n3409 ;
  assign n8826 = ~n8824 & n8825 ;
  assign n8827 = n4925 & n8826 ;
  assign n8801 = n2749 & n4934 ;
  assign n8828 = n2768 & ~n5093 ;
  assign n8829 = ~n8801 & ~n8828 ;
  assign n8830 = ~n8827 & n8829 ;
  assign n8831 = ~n8823 & n8830 ;
  assign n8832 = ~n8817 & n8831 ;
  assign n8833 = ~n8811 & n8832 ;
  assign n8834 = n2017 & ~n8833 ;
  assign n8835 = n2749 & n3430 ;
  assign n8836 = ~n8834 & ~n8835 ;
  assign n8837 = \P1_state_reg[0]/NET0131  & ~n8836 ;
  assign n8800 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[5]/NET0131  ;
  assign n8838 = n2749 & n3935 ;
  assign n8839 = ~n8800 & ~n8838 ;
  assign n8840 = ~n8837 & n8839 ;
  assign n8843 = n2698 & n3430 ;
  assign n8845 = n2698 & ~n4925 ;
  assign n8852 = n2678 & ~n3337 ;
  assign n8853 = ~n8155 & ~n8852 ;
  assign n8854 = ~n2050 & ~n8853 ;
  assign n8855 = n2050 & n2730 ;
  assign n8856 = ~n8854 & ~n8855 ;
  assign n8857 = n4925 & n8856 ;
  assign n8858 = ~n8845 & ~n8857 ;
  assign n8859 = n3373 & ~n8858 ;
  assign n8846 = n4121 & ~n4386 ;
  assign n8847 = ~n4121 & n4386 ;
  assign n8848 = ~n8846 & ~n8847 ;
  assign n8849 = n4925 & n8848 ;
  assign n8850 = ~n8845 & ~n8849 ;
  assign n8851 = n3179 & ~n8850 ;
  assign n8860 = ~n3224 & n4121 ;
  assign n8861 = n3224 & ~n4121 ;
  assign n8862 = ~n8860 & ~n8861 ;
  assign n8863 = n4925 & ~n8862 ;
  assign n8864 = ~n8845 & ~n8863 ;
  assign n8865 = n3319 & ~n8864 ;
  assign n8866 = n2719 & ~n3382 ;
  assign n8867 = ~n3383 & ~n8866 ;
  assign n8868 = n3409 & n8867 ;
  assign n8869 = n4925 & n8868 ;
  assign n8844 = n2698 & n4934 ;
  assign n8870 = n2719 & ~n5093 ;
  assign n8871 = ~n8844 & ~n8870 ;
  assign n8872 = ~n8869 & n8871 ;
  assign n8873 = ~n8865 & n8872 ;
  assign n8874 = ~n8851 & n8873 ;
  assign n8875 = ~n8859 & n8874 ;
  assign n8876 = n2017 & ~n8875 ;
  assign n8877 = ~n8843 & ~n8876 ;
  assign n8878 = \P1_state_reg[0]/NET0131  & ~n8877 ;
  assign n8841 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[7]/NET0131  ;
  assign n8842 = n2698 & n3935 ;
  assign n8879 = ~n8841 & ~n8842 ;
  assign n8880 = ~n8878 & n8879 ;
  assign n8882 = n1218 & n3664 ;
  assign n8883 = n1248 & ~n7280 ;
  assign n8884 = ~n7281 & ~n8883 ;
  assign n8885 = ~n536 & ~n8884 ;
  assign n8886 = n536 & n1274 ;
  assign n8887 = ~n8885 & ~n8886 ;
  assign n8907 = n3450 & ~n8887 ;
  assign n8908 = n1898 & ~n8907 ;
  assign n8909 = n8129 & ~n8908 ;
  assign n8910 = n1218 & ~n8909 ;
  assign n8888 = n1898 & n8887 ;
  assign n8899 = ~n1740 & ~n3484 ;
  assign n8898 = n1740 & n3484 ;
  assign n8900 = n3557 & ~n8898 ;
  assign n8901 = ~n8899 & n8900 ;
  assign n8895 = ~n1740 & n4454 ;
  assign n8894 = n1740 & ~n4454 ;
  assign n8896 = n3575 & ~n8894 ;
  assign n8897 = ~n8895 & n8896 ;
  assign n8889 = ~n1238 & n3683 ;
  assign n8890 = ~n1238 & ~n3630 ;
  assign n8891 = n1238 & n3630 ;
  assign n8892 = n3650 & ~n8891 ;
  assign n8893 = ~n8890 & n8892 ;
  assign n8902 = ~n8889 & ~n8893 ;
  assign n8903 = ~n8897 & n8902 ;
  assign n8904 = ~n8901 & n8903 ;
  assign n8905 = ~n8888 & n8904 ;
  assign n8906 = n3450 & ~n8905 ;
  assign n8911 = ~n1238 & n1736 ;
  assign n8912 = ~n8906 & ~n8911 ;
  assign n8913 = ~n8910 & n8912 ;
  assign n8914 = n3662 & ~n8913 ;
  assign n8915 = ~n8882 & ~n8914 ;
  assign n8916 = \P1_state_reg[0]/NET0131  & ~n8915 ;
  assign n8881 = \P1_reg3_reg[6]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8917 = n1218 & n1934 ;
  assign n8918 = ~n8881 & ~n8917 ;
  assign n8919 = ~n8916 & n8918 ;
  assign n8921 = n1243 & n3664 ;
  assign n8922 = n1189 & ~n7281 ;
  assign n8923 = ~n7282 & ~n8922 ;
  assign n8924 = ~n536 & ~n8923 ;
  assign n8925 = n536 & n1222 ;
  assign n8926 = ~n8924 & ~n8925 ;
  assign n8927 = n1898 & n8926 ;
  assign n8937 = ~n1743 & n5016 ;
  assign n8936 = n1743 & ~n5016 ;
  assign n8938 = n3557 & ~n8936 ;
  assign n8939 = ~n8937 & n8938 ;
  assign n8929 = n1743 & n4979 ;
  assign n8928 = ~n1743 & ~n4979 ;
  assign n8930 = n3575 & ~n8928 ;
  assign n8931 = ~n8929 & n8930 ;
  assign n8932 = n3650 & n8891 ;
  assign n8933 = ~n3683 & ~n8932 ;
  assign n8934 = ~n1263 & ~n8933 ;
  assign n8935 = n1263 & n8892 ;
  assign n8940 = ~n8934 & ~n8935 ;
  assign n8941 = ~n8931 & n8940 ;
  assign n8942 = ~n8939 & n8941 ;
  assign n8943 = ~n8927 & n8942 ;
  assign n8944 = n3450 & ~n8943 ;
  assign n8945 = ~n6590 & n8129 ;
  assign n8946 = n1243 & ~n8945 ;
  assign n8947 = ~n1263 & n1736 ;
  assign n8948 = ~n8946 & ~n8947 ;
  assign n8949 = ~n8944 & n8948 ;
  assign n8950 = n3662 & ~n8949 ;
  assign n8951 = ~n8921 & ~n8950 ;
  assign n8952 = \P1_state_reg[0]/NET0131  & ~n8951 ;
  assign n8920 = \P1_reg3_reg[7]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8953 = n1243 & n1934 ;
  assign n8954 = ~n8920 & ~n8953 ;
  assign n8955 = ~n8952 & n8954 ;
  assign n8956 = \P2_reg0_reg[4]/NET0131  & ~n3434 ;
  assign n8957 = \P2_reg0_reg[4]/NET0131  & n3430 ;
  assign n8958 = n5258 & ~n6900 ;
  assign n8959 = ~n6902 & n8958 ;
  assign n8960 = \P2_reg0_reg[4]/NET0131  & ~n8959 ;
  assign n8961 = ~n2849 & n3375 ;
  assign n8962 = n3373 & n8771 ;
  assign n8963 = n8788 & ~n8962 ;
  assign n8964 = ~n8961 & n8963 ;
  assign n8965 = n4610 & ~n8964 ;
  assign n8966 = ~n8960 & ~n8965 ;
  assign n8967 = n2017 & ~n8966 ;
  assign n8968 = ~n8957 & ~n8967 ;
  assign n8969 = \P1_state_reg[0]/NET0131  & ~n8968 ;
  assign n8970 = ~n8956 & ~n8969 ;
  assign n8971 = \P2_reg1_reg[4]/NET0131  & ~n3434 ;
  assign n8972 = \P2_reg1_reg[4]/NET0131  & n3430 ;
  assign n8973 = \P2_reg1_reg[4]/NET0131  & ~n6721 ;
  assign n8974 = n4663 & ~n8964 ;
  assign n8975 = ~n8973 & ~n8974 ;
  assign n8976 = n2017 & ~n8975 ;
  assign n8977 = ~n8972 & ~n8976 ;
  assign n8978 = \P1_state_reg[0]/NET0131  & ~n8977 ;
  assign n8979 = ~n8971 & ~n8978 ;
  assign n8980 = ~\P1_reg2_reg[4]/NET0131  & ~n3672 ;
  assign n8981 = n3672 & ~n8108 ;
  assign n8982 = n1898 & ~n8981 ;
  assign n8983 = n3672 & ~n8124 ;
  assign n8984 = n6070 & ~n8983 ;
  assign n8985 = ~n8982 & n8984 ;
  assign n8986 = ~n8980 & ~n8985 ;
  assign n8987 = n1291 & n1736 ;
  assign n8988 = n3556 & ~n3672 ;
  assign n8989 = n5428 & ~n8988 ;
  assign n8990 = \P1_reg2_reg[4]/NET0131  & ~n8989 ;
  assign n8991 = ~n8987 & ~n8990 ;
  assign n8992 = ~n8986 & n8991 ;
  assign n8993 = ~\P1_reg2_reg[4]/NET0131  & ~n6070 ;
  assign n8994 = ~n8992 & ~n8993 ;
  assign n8995 = \P2_reg2_reg[8]/NET0131  & ~n3434 ;
  assign n8996 = \P2_reg2_reg[8]/NET0131  & n3430 ;
  assign n8998 = \P2_reg2_reg[8]/NET0131  & ~n2033 ;
  assign n9002 = n2033 & ~n8159 ;
  assign n9003 = ~n8998 & ~n9002 ;
  assign n9004 = n3373 & ~n9003 ;
  assign n8999 = n2033 & n8150 ;
  assign n9000 = ~n8998 & ~n8999 ;
  assign n9001 = n3319 & ~n9000 ;
  assign n9009 = n2033 & ~n8165 ;
  assign n9010 = ~n8998 & ~n9009 ;
  assign n9011 = n3179 & ~n9010 ;
  assign n9006 = n2692 & n3375 ;
  assign n9007 = ~n8171 & ~n9006 ;
  assign n9008 = n2033 & ~n9007 ;
  assign n8997 = n2674 & n3415 ;
  assign n9005 = \P2_reg2_reg[8]/NET0131  & ~n4436 ;
  assign n9012 = ~n8997 & ~n9005 ;
  assign n9013 = ~n9008 & n9012 ;
  assign n9014 = ~n9011 & n9013 ;
  assign n9015 = ~n9001 & n9014 ;
  assign n9016 = ~n9004 & n9015 ;
  assign n9017 = n2017 & ~n9016 ;
  assign n9018 = ~n8996 & ~n9017 ;
  assign n9019 = \P1_state_reg[0]/NET0131  & ~n9018 ;
  assign n9020 = ~n8995 & ~n9019 ;
  assign n9021 = \P1_reg1_reg[5]/NET0131  & ~n8721 ;
  assign n9022 = n6246 & ~n8207 ;
  assign n9023 = ~n9021 & ~n9022 ;
  assign n9024 = \P2_reg0_reg[8]/NET0131  & ~n3434 ;
  assign n9025 = \P2_reg0_reg[8]/NET0131  & n3430 ;
  assign n9027 = \P2_reg0_reg[8]/NET0131  & ~n4610 ;
  assign n9031 = n4610 & ~n8159 ;
  assign n9032 = ~n9027 & ~n9031 ;
  assign n9033 = n3373 & ~n9032 ;
  assign n9028 = n4610 & n8150 ;
  assign n9029 = ~n9027 & ~n9028 ;
  assign n9030 = n3319 & ~n9029 ;
  assign n9034 = n4610 & ~n8165 ;
  assign n9035 = ~n9027 & ~n9034 ;
  assign n9036 = n3179 & ~n9035 ;
  assign n9026 = \P2_reg0_reg[8]/NET0131  & ~n5258 ;
  assign n9037 = n4610 & ~n9007 ;
  assign n9038 = ~n9026 & ~n9037 ;
  assign n9039 = ~n9036 & n9038 ;
  assign n9040 = ~n9030 & n9039 ;
  assign n9041 = ~n9033 & n9040 ;
  assign n9042 = n2017 & ~n9041 ;
  assign n9043 = ~n9025 & ~n9042 ;
  assign n9044 = \P1_state_reg[0]/NET0131  & ~n9043 ;
  assign n9045 = ~n9024 & ~n9044 ;
  assign n9046 = \P2_reg1_reg[11]/NET0131  & ~n6749 ;
  assign n9048 = n3373 & n8030 ;
  assign n9049 = n3179 & n8036 ;
  assign n9050 = n3319 & ~n8046 ;
  assign n9047 = n2926 & n3375 ;
  assign n9051 = ~n8042 & ~n9047 ;
  assign n9052 = ~n9050 & n9051 ;
  assign n9053 = ~n9049 & n9052 ;
  assign n9054 = ~n9048 & n9053 ;
  assign n9055 = n5572 & ~n9054 ;
  assign n9056 = ~n9046 & ~n9055 ;
  assign n9057 = \P2_reg1_reg[8]/NET0131  & ~n3434 ;
  assign n9058 = \P2_reg1_reg[8]/NET0131  & n3430 ;
  assign n9060 = \P2_reg1_reg[8]/NET0131  & ~n4663 ;
  assign n9064 = n4663 & ~n8159 ;
  assign n9065 = ~n9060 & ~n9064 ;
  assign n9066 = n3373 & ~n9065 ;
  assign n9061 = n4663 & n8150 ;
  assign n9062 = ~n9060 & ~n9061 ;
  assign n9063 = n3319 & ~n9062 ;
  assign n9067 = n4663 & ~n8165 ;
  assign n9068 = ~n9060 & ~n9067 ;
  assign n9069 = n3179 & ~n9068 ;
  assign n9059 = \P2_reg1_reg[8]/NET0131  & ~n5509 ;
  assign n9070 = n4663 & ~n9007 ;
  assign n9071 = ~n9059 & ~n9070 ;
  assign n9072 = ~n9069 & n9071 ;
  assign n9073 = ~n9063 & n9072 ;
  assign n9074 = ~n9066 & n9073 ;
  assign n9075 = n2017 & ~n9074 ;
  assign n9076 = ~n9058 & ~n9075 ;
  assign n9077 = \P1_state_reg[0]/NET0131  & ~n9076 ;
  assign n9078 = ~n9057 & ~n9077 ;
  assign n9079 = \P1_reg0_reg[10]/NET0131  & ~n3703 ;
  assign n9080 = \P1_reg0_reg[10]/NET0131  & n3664 ;
  assign n9082 = \P1_reg0_reg[10]/NET0131  & ~n3900 ;
  assign n9083 = n3900 & n6987 ;
  assign n9084 = ~n9082 & ~n9083 ;
  assign n9085 = n1898 & ~n9084 ;
  assign n9089 = n3900 & n6993 ;
  assign n9090 = ~n9082 & ~n9089 ;
  assign n9091 = n3575 & ~n9090 ;
  assign n9086 = n3900 & ~n6999 ;
  assign n9087 = ~n9082 & ~n9086 ;
  assign n9088 = n3557 & ~n9087 ;
  assign n9081 = \P1_reg0_reg[10]/NET0131  & ~n4723 ;
  assign n9092 = n3900 & ~n6980 ;
  assign n9093 = ~n9081 & ~n9092 ;
  assign n9094 = ~n9088 & n9093 ;
  assign n9095 = ~n9091 & n9094 ;
  assign n9096 = ~n9085 & n9095 ;
  assign n9097 = n3662 & ~n9096 ;
  assign n9098 = ~n9080 & ~n9097 ;
  assign n9099 = \P1_state_reg[0]/NET0131  & ~n9098 ;
  assign n9100 = ~n9079 & ~n9099 ;
  assign n9101 = ~\P1_reg2_reg[5]/NET0131  & ~n3672 ;
  assign n9102 = n3672 & ~n8190 ;
  assign n9103 = n1898 & ~n9102 ;
  assign n9104 = n3672 & ~n8206 ;
  assign n9105 = n6070 & ~n9104 ;
  assign n9106 = ~n9103 & n9105 ;
  assign n9107 = ~n9101 & ~n9106 ;
  assign n9108 = n1270 & n1736 ;
  assign n9109 = \P1_reg2_reg[5]/NET0131  & ~n8989 ;
  assign n9110 = ~n9108 & ~n9109 ;
  assign n9111 = ~n9107 & n9110 ;
  assign n9112 = ~\P1_reg2_reg[5]/NET0131  & ~n6070 ;
  assign n9113 = ~n9111 & ~n9112 ;
  assign n9114 = n2905 & n3415 ;
  assign n9115 = n2033 & ~n9054 ;
  assign n9116 = ~n9114 & ~n9115 ;
  assign n9117 = n4275 & ~n9116 ;
  assign n9118 = \P2_reg2_reg[11]/NET0131  & ~n6797 ;
  assign n9119 = ~n9117 & ~n9118 ;
  assign n9120 = \P2_reg2_reg[14]/NET0131  & ~n3434 ;
  assign n9121 = \P2_reg2_reg[14]/NET0131  & n3430 ;
  assign n9123 = \P2_reg2_reg[14]/NET0131  & ~n2033 ;
  assign n9124 = n2033 & n8070 ;
  assign n9125 = ~n9123 & ~n9124 ;
  assign n9126 = n3319 & ~n9125 ;
  assign n9130 = n2033 & n8084 ;
  assign n9131 = ~n9123 & ~n9130 ;
  assign n9132 = n3373 & ~n9131 ;
  assign n9127 = n2033 & ~n8076 ;
  assign n9128 = ~n9123 & ~n9127 ;
  assign n9129 = n3179 & ~n9128 ;
  assign n9134 = n3095 & n3375 ;
  assign n9135 = ~n8090 & ~n9134 ;
  assign n9136 = n2033 & ~n9135 ;
  assign n9122 = \P2_reg2_reg[14]/NET0131  & ~n4436 ;
  assign n9133 = n3077 & n3415 ;
  assign n9137 = ~n9122 & ~n9133 ;
  assign n9138 = ~n9136 & n9137 ;
  assign n9139 = ~n9129 & n9138 ;
  assign n9140 = ~n9132 & n9139 ;
  assign n9141 = ~n9126 & n9140 ;
  assign n9142 = n2017 & ~n9141 ;
  assign n9143 = ~n9121 & ~n9142 ;
  assign n9144 = \P1_state_reg[0]/NET0131  & ~n9143 ;
  assign n9145 = ~n9120 & ~n9144 ;
  assign n9147 = \P1_reg0_reg[11]/NET0131  & ~n3900 ;
  assign n9148 = n3900 & n6942 ;
  assign n9149 = ~n9147 & ~n9148 ;
  assign n9150 = n1898 & ~n9149 ;
  assign n9151 = n3900 & ~n6948 ;
  assign n9152 = ~n9147 & ~n9151 ;
  assign n9153 = n3557 & ~n9152 ;
  assign n9146 = \P1_reg0_reg[11]/NET0131  & ~n6167 ;
  assign n9154 = n3900 & ~n6962 ;
  assign n9155 = ~n9146 & ~n9154 ;
  assign n9156 = ~n9153 & n9155 ;
  assign n9157 = ~n9150 & n9156 ;
  assign n9158 = n3662 & ~n9157 ;
  assign n9159 = \P1_reg0_reg[11]/NET0131  & n3664 ;
  assign n9160 = ~n9158 & ~n9159 ;
  assign n9161 = \P1_state_reg[0]/NET0131  & ~n9160 ;
  assign n9162 = \P1_reg0_reg[11]/NET0131  & ~n3703 ;
  assign n9163 = ~n9161 & ~n9162 ;
  assign n9164 = \P1_reg0_reg[13]/NET0131  & ~n3703 ;
  assign n9165 = \P1_reg0_reg[13]/NET0131  & n3664 ;
  assign n9166 = \P1_reg0_reg[13]/NET0131  & ~n6177 ;
  assign n9167 = n3900 & ~n8299 ;
  assign n9168 = ~n9166 & ~n9167 ;
  assign n9169 = n3662 & ~n9168 ;
  assign n9170 = ~n9165 & ~n9169 ;
  assign n9171 = \P1_state_reg[0]/NET0131  & ~n9170 ;
  assign n9172 = ~n9164 & ~n9171 ;
  assign n9173 = n6070 & n6177 ;
  assign n9174 = \P1_reg0_reg[14]/NET0131  & ~n9173 ;
  assign n9175 = n6171 & ~n8310 ;
  assign n9176 = ~n9174 & ~n9175 ;
  assign n9177 = \P1_reg0_reg[4]/NET0131  & ~n6169 ;
  assign n9178 = n6171 & ~n8125 ;
  assign n9179 = ~n9177 & ~n9178 ;
  assign n9180 = n6171 & ~n8207 ;
  assign n9181 = \P1_reg0_reg[5]/NET0131  & ~n6169 ;
  assign n9182 = ~n9180 & ~n9181 ;
  assign n9183 = \P1_reg1_reg[10]/NET0131  & ~n3703 ;
  assign n9184 = \P1_reg1_reg[10]/NET0131  & n3664 ;
  assign n9186 = \P1_reg1_reg[10]/NET0131  & ~n4236 ;
  assign n9187 = n4236 & n6987 ;
  assign n9188 = ~n9186 & ~n9187 ;
  assign n9189 = n1898 & ~n9188 ;
  assign n9193 = n4236 & n6993 ;
  assign n9194 = ~n9186 & ~n9193 ;
  assign n9195 = n3575 & ~n9194 ;
  assign n9190 = n4236 & ~n6999 ;
  assign n9191 = ~n9186 & ~n9190 ;
  assign n9192 = n3557 & ~n9191 ;
  assign n9185 = \P1_reg1_reg[10]/NET0131  & ~n6889 ;
  assign n9196 = n4236 & ~n6980 ;
  assign n9197 = ~n9185 & ~n9196 ;
  assign n9198 = ~n9192 & n9197 ;
  assign n9199 = ~n9195 & n9198 ;
  assign n9200 = ~n9189 & n9199 ;
  assign n9201 = n3662 & ~n9200 ;
  assign n9202 = ~n9184 & ~n9201 ;
  assign n9203 = \P1_state_reg[0]/NET0131  & ~n9202 ;
  assign n9204 = ~n9183 & ~n9203 ;
  assign n9205 = \P1_reg1_reg[11]/NET0131  & ~n3703 ;
  assign n9206 = \P1_reg1_reg[11]/NET0131  & n3664 ;
  assign n9208 = \P1_reg1_reg[11]/NET0131  & ~n4236 ;
  assign n9209 = n4236 & n6942 ;
  assign n9210 = ~n9208 & ~n9209 ;
  assign n9211 = n1898 & ~n9210 ;
  assign n9212 = n4236 & ~n6948 ;
  assign n9213 = ~n9208 & ~n9212 ;
  assign n9214 = n3557 & ~n9213 ;
  assign n9207 = \P1_reg1_reg[11]/NET0131  & ~n6890 ;
  assign n9215 = n4236 & ~n6962 ;
  assign n9216 = ~n9207 & ~n9215 ;
  assign n9217 = ~n9214 & n9216 ;
  assign n9218 = ~n9211 & n9217 ;
  assign n9219 = n3662 & ~n9218 ;
  assign n9220 = ~n9206 & ~n9219 ;
  assign n9221 = \P1_state_reg[0]/NET0131  & ~n9220 ;
  assign n9222 = ~n9205 & ~n9221 ;
  assign n9224 = \P1_reg1_reg[13]/NET0131  & ~n4236 ;
  assign n9225 = n6246 & n8009 ;
  assign n9226 = ~n9224 & ~n9225 ;
  assign n9227 = n1898 & ~n9226 ;
  assign n9223 = n6246 & ~n8298 ;
  assign n9228 = ~n4757 & n7909 ;
  assign n9229 = \P1_reg1_reg[13]/NET0131  & ~n9228 ;
  assign n9230 = ~n9223 & ~n9229 ;
  assign n9231 = ~n9227 & n9230 ;
  assign n9233 = \P1_reg1_reg[14]/NET0131  & ~n4236 ;
  assign n9234 = n6246 & n7041 ;
  assign n9235 = ~n9233 & ~n9234 ;
  assign n9236 = n1898 & ~n9235 ;
  assign n9232 = n6246 & ~n8308 ;
  assign n9237 = \P1_reg1_reg[14]/NET0131  & ~n9228 ;
  assign n9238 = ~n9232 & ~n9237 ;
  assign n9239 = ~n9236 & n9238 ;
  assign n9240 = n5385 & ~n9054 ;
  assign n9241 = n4621 & n7533 ;
  assign n9242 = \P2_reg0_reg[11]/NET0131  & ~n9241 ;
  assign n9243 = ~n9240 & ~n9242 ;
  assign n9246 = ~\P2_reg3_reg[3]/NET0131  & ~n4925 ;
  assign n9247 = n2858 & ~n3333 ;
  assign n9248 = ~n3334 & ~n9247 ;
  assign n9249 = ~n2050 & ~n9248 ;
  assign n9250 = n2050 & n2777 ;
  assign n9251 = ~n9249 & ~n9250 ;
  assign n9252 = n4925 & n9251 ;
  assign n9253 = ~n9246 & ~n9252 ;
  assign n9254 = n3373 & ~n9253 ;
  assign n9255 = n2835 & ~n4133 ;
  assign n9256 = ~n2835 & n4133 ;
  assign n9257 = ~n9255 & ~n9256 ;
  assign n9258 = n4925 & ~n9257 ;
  assign n9259 = ~n9246 & ~n9258 ;
  assign n9260 = n3179 & ~n9259 ;
  assign n9261 = ~n3204 & ~n3207 ;
  assign n9262 = ~n4133 & n9261 ;
  assign n9263 = n4133 & ~n9261 ;
  assign n9264 = ~n9262 & ~n9263 ;
  assign n9265 = n4925 & ~n9264 ;
  assign n9266 = ~n9246 & ~n9265 ;
  assign n9267 = n3319 & ~n9266 ;
  assign n9268 = ~n2880 & ~n3378 ;
  assign n9269 = ~n3379 & ~n9268 ;
  assign n9270 = n3409 & n9269 ;
  assign n9271 = n4925 & n9270 ;
  assign n9245 = ~\P2_reg3_reg[3]/NET0131  & n4934 ;
  assign n9272 = ~n2880 & ~n5093 ;
  assign n9273 = ~n9245 & ~n9272 ;
  assign n9274 = ~n9271 & n9273 ;
  assign n9275 = ~n9267 & n9274 ;
  assign n9276 = ~n9260 & n9275 ;
  assign n9277 = ~n9254 & n9276 ;
  assign n9278 = n2017 & ~n9277 ;
  assign n9279 = ~\P2_reg3_reg[3]/NET0131  & n3430 ;
  assign n9280 = ~n9278 & ~n9279 ;
  assign n9281 = \P1_state_reg[0]/NET0131  & ~n9280 ;
  assign n9244 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[3]/NET0131  ;
  assign n9282 = ~\P2_reg3_reg[3]/NET0131  & n3935 ;
  assign n9283 = ~n9244 & ~n9282 ;
  assign n9284 = ~n9281 & n9283 ;
  assign n9287 = n2726 & ~n4925 ;
  assign n9288 = n2050 & ~n2755 ;
  assign n9289 = n2702 & ~n8804 ;
  assign n9290 = ~n2050 & ~n3337 ;
  assign n9291 = ~n9289 & n9290 ;
  assign n9292 = ~n9288 & ~n9291 ;
  assign n9293 = n4925 & ~n9292 ;
  assign n9294 = ~n9287 & ~n9293 ;
  assign n9295 = n3373 & ~n9294 ;
  assign n9296 = n4130 & ~n5273 ;
  assign n9297 = ~n4130 & n5273 ;
  assign n9298 = ~n9296 & ~n9297 ;
  assign n9299 = n4925 & n9298 ;
  assign n9300 = ~n9287 & ~n9299 ;
  assign n9301 = n3179 & ~n9300 ;
  assign n9302 = ~n4101 & n4130 ;
  assign n9303 = n4101 & ~n4130 ;
  assign n9304 = ~n9302 & ~n9303 ;
  assign n9305 = n4925 & ~n9304 ;
  assign n9306 = ~n9287 & ~n9305 ;
  assign n9307 = n3319 & ~n9306 ;
  assign n9308 = n2745 & ~n3381 ;
  assign n9309 = ~n3382 & n3409 ;
  assign n9310 = ~n9308 & n9309 ;
  assign n9311 = n4925 & n9310 ;
  assign n9286 = n2726 & n4934 ;
  assign n9312 = n2745 & ~n5093 ;
  assign n9313 = ~n9286 & ~n9312 ;
  assign n9314 = ~n9311 & n9313 ;
  assign n9315 = ~n9307 & n9314 ;
  assign n9316 = ~n9301 & n9315 ;
  assign n9317 = ~n9295 & n9316 ;
  assign n9318 = n2017 & ~n9317 ;
  assign n9319 = n2726 & n3430 ;
  assign n9320 = ~n9318 & ~n9319 ;
  assign n9321 = \P1_state_reg[0]/NET0131  & ~n9320 ;
  assign n9285 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[6]/NET0131  ;
  assign n9322 = n2726 & n3935 ;
  assign n9323 = ~n9285 & ~n9322 ;
  assign n9324 = ~n9321 & n9323 ;
  assign n9325 = \P2_reg2_reg[5]/NET0131  & ~n3434 ;
  assign n9327 = \P2_reg2_reg[5]/NET0131  & ~n2033 ;
  assign n9328 = n2033 & n8808 ;
  assign n9329 = ~n9327 & ~n9328 ;
  assign n9330 = n3373 & ~n9329 ;
  assign n9331 = n2033 & ~n8814 ;
  assign n9332 = ~n9327 & ~n9331 ;
  assign n9333 = n3179 & ~n9332 ;
  assign n9337 = n3319 & n8820 ;
  assign n9336 = n2768 & n3375 ;
  assign n9338 = ~n8826 & ~n9336 ;
  assign n9339 = ~n9337 & n9338 ;
  assign n9340 = n2033 & ~n9339 ;
  assign n9326 = n2749 & n3415 ;
  assign n9334 = n4436 & ~n6794 ;
  assign n9335 = \P2_reg2_reg[5]/NET0131  & ~n9334 ;
  assign n9341 = ~n9326 & ~n9335 ;
  assign n9342 = ~n9340 & n9341 ;
  assign n9343 = ~n9333 & n9342 ;
  assign n9344 = ~n9330 & n9343 ;
  assign n9345 = n2017 & ~n9344 ;
  assign n9346 = \P2_reg2_reg[5]/NET0131  & n3430 ;
  assign n9347 = ~n9345 & ~n9346 ;
  assign n9348 = \P1_state_reg[0]/NET0131  & ~n9347 ;
  assign n9349 = ~n9325 & ~n9348 ;
  assign n9351 = \P1_reg1_reg[7]/NET0131  & ~n4236 ;
  assign n9352 = n6246 & n8926 ;
  assign n9353 = ~n9351 & ~n9352 ;
  assign n9354 = n1898 & ~n9353 ;
  assign n9350 = n6246 & ~n8942 ;
  assign n9355 = \P1_reg1_reg[7]/NET0131  & ~n9228 ;
  assign n9356 = ~n9350 & ~n9355 ;
  assign n9357 = ~n9354 & n9356 ;
  assign n9358 = \P2_reg0_reg[5]/NET0131  & ~n3434 ;
  assign n9360 = \P2_reg0_reg[5]/NET0131  & ~n4610 ;
  assign n9361 = n4610 & n8808 ;
  assign n9362 = ~n9360 & ~n9361 ;
  assign n9363 = n3373 & ~n9362 ;
  assign n9364 = n4610 & ~n8814 ;
  assign n9365 = ~n9360 & ~n9364 ;
  assign n9366 = n3179 & ~n9365 ;
  assign n9359 = \P2_reg0_reg[5]/NET0131  & ~n8958 ;
  assign n9367 = n4610 & ~n9339 ;
  assign n9368 = ~n9359 & ~n9367 ;
  assign n9369 = ~n9366 & n9368 ;
  assign n9370 = ~n9363 & n9369 ;
  assign n9371 = n2017 & ~n9370 ;
  assign n9372 = \P2_reg0_reg[5]/NET0131  & n3430 ;
  assign n9373 = ~n9371 & ~n9372 ;
  assign n9374 = \P1_state_reg[0]/NET0131  & ~n9373 ;
  assign n9375 = ~n9358 & ~n9374 ;
  assign n9376 = \P2_reg0_reg[7]/NET0131  & ~n3434 ;
  assign n9377 = \P2_reg0_reg[7]/NET0131  & n3430 ;
  assign n9384 = \P2_reg0_reg[7]/NET0131  & ~n4610 ;
  assign n9388 = n4610 & n8856 ;
  assign n9389 = ~n9384 & ~n9388 ;
  assign n9390 = n3373 & ~n9389 ;
  assign n9385 = n4610 & n8848 ;
  assign n9386 = ~n9384 & ~n9385 ;
  assign n9387 = n3179 & ~n9386 ;
  assign n9378 = \P2_reg0_reg[7]/NET0131  & ~n8958 ;
  assign n9380 = n3319 & ~n8862 ;
  assign n9379 = n2719 & n3375 ;
  assign n9381 = ~n8868 & ~n9379 ;
  assign n9382 = ~n9380 & n9381 ;
  assign n9383 = n4610 & ~n9382 ;
  assign n9391 = ~n9378 & ~n9383 ;
  assign n9392 = ~n9387 & n9391 ;
  assign n9393 = ~n9390 & n9392 ;
  assign n9394 = n2017 & ~n9393 ;
  assign n9395 = ~n9377 & ~n9394 ;
  assign n9396 = \P1_state_reg[0]/NET0131  & ~n9395 ;
  assign n9397 = ~n9376 & ~n9396 ;
  assign n9398 = \P2_reg1_reg[14]/NET0131  & ~n3434 ;
  assign n9399 = \P2_reg1_reg[14]/NET0131  & n3430 ;
  assign n9401 = \P2_reg1_reg[14]/NET0131  & ~n4663 ;
  assign n9402 = n4663 & n8070 ;
  assign n9403 = ~n9401 & ~n9402 ;
  assign n9404 = n3319 & ~n9403 ;
  assign n9408 = n4663 & ~n8076 ;
  assign n9409 = ~n9401 & ~n9408 ;
  assign n9410 = n3179 & ~n9409 ;
  assign n9405 = n4663 & n8084 ;
  assign n9406 = ~n9401 & ~n9405 ;
  assign n9407 = n3373 & ~n9406 ;
  assign n9400 = \P2_reg1_reg[14]/NET0131  & ~n5509 ;
  assign n9411 = n4663 & ~n9135 ;
  assign n9412 = ~n9400 & ~n9411 ;
  assign n9413 = ~n9407 & n9412 ;
  assign n9414 = ~n9410 & n9413 ;
  assign n9415 = ~n9404 & n9414 ;
  assign n9416 = n2017 & ~n9415 ;
  assign n9417 = ~n9399 & ~n9416 ;
  assign n9418 = \P1_state_reg[0]/NET0131  & ~n9417 ;
  assign n9419 = ~n9398 & ~n9418 ;
  assign n9420 = \P2_reg1_reg[5]/NET0131  & ~n3434 ;
  assign n9422 = \P2_reg1_reg[5]/NET0131  & ~n4663 ;
  assign n9423 = n4663 & n8808 ;
  assign n9424 = ~n9422 & ~n9423 ;
  assign n9425 = n3373 & ~n9424 ;
  assign n9426 = n4663 & ~n8814 ;
  assign n9427 = ~n9422 & ~n9426 ;
  assign n9428 = n3179 & ~n9427 ;
  assign n9421 = \P2_reg1_reg[5]/NET0131  & ~n6719 ;
  assign n9429 = n4663 & ~n9339 ;
  assign n9430 = ~n9421 & ~n9429 ;
  assign n9431 = ~n9428 & n9430 ;
  assign n9432 = ~n9425 & n9431 ;
  assign n9433 = n2017 & ~n9432 ;
  assign n9434 = \P2_reg1_reg[5]/NET0131  & n3430 ;
  assign n9435 = ~n9433 & ~n9434 ;
  assign n9436 = \P1_state_reg[0]/NET0131  & ~n9435 ;
  assign n9437 = ~n9420 & ~n9436 ;
  assign n9438 = \P1_reg2_reg[3]/NET0131  & ~n3703 ;
  assign n9439 = \P1_reg2_reg[3]/NET0131  & n3664 ;
  assign n9441 = ~n1336 & n3683 ;
  assign n9442 = n8742 & ~n9441 ;
  assign n9443 = n1898 & n8750 ;
  assign n9444 = n9442 & ~n9443 ;
  assign n9445 = n3672 & ~n9444 ;
  assign n9440 = ~\P1_reg3_reg[3]/NET0131  & n1736 ;
  assign n9446 = n1898 & ~n3672 ;
  assign n9447 = n8989 & ~n9446 ;
  assign n9448 = \P1_reg2_reg[3]/NET0131  & ~n9447 ;
  assign n9449 = ~n9440 & ~n9448 ;
  assign n9450 = ~n9445 & n9449 ;
  assign n9451 = n3662 & ~n9450 ;
  assign n9452 = ~n9439 & ~n9451 ;
  assign n9453 = \P1_state_reg[0]/NET0131  & ~n9452 ;
  assign n9454 = ~n9438 & ~n9453 ;
  assign n9455 = \P2_reg1_reg[7]/NET0131  & ~n3434 ;
  assign n9456 = \P2_reg1_reg[7]/NET0131  & n3430 ;
  assign n9459 = \P2_reg1_reg[7]/NET0131  & ~n4663 ;
  assign n9463 = n4663 & n8856 ;
  assign n9464 = ~n9459 & ~n9463 ;
  assign n9465 = n3373 & ~n9464 ;
  assign n9460 = n4663 & n8848 ;
  assign n9461 = ~n9459 & ~n9460 ;
  assign n9462 = n3179 & ~n9461 ;
  assign n9457 = \P2_reg1_reg[7]/NET0131  & ~n6719 ;
  assign n9458 = n4663 & ~n9382 ;
  assign n9466 = ~n9457 & ~n9458 ;
  assign n9467 = ~n9462 & n9466 ;
  assign n9468 = ~n9465 & n9467 ;
  assign n9469 = n2017 & ~n9468 ;
  assign n9470 = ~n9456 & ~n9469 ;
  assign n9471 = \P1_state_reg[0]/NET0131  & ~n9470 ;
  assign n9472 = ~n9455 & ~n9471 ;
  assign n9473 = ~\P1_reg2_reg[6]/NET0131  & ~n3672 ;
  assign n9474 = n3672 & ~n8887 ;
  assign n9475 = n1898 & ~n9474 ;
  assign n9476 = n3672 & ~n8904 ;
  assign n9477 = n6070 & ~n9476 ;
  assign n9478 = ~n9475 & n9477 ;
  assign n9479 = ~n9473 & ~n9478 ;
  assign n9480 = n1218 & n1736 ;
  assign n9481 = \P1_reg2_reg[6]/NET0131  & ~n8989 ;
  assign n9482 = ~n9480 & ~n9481 ;
  assign n9483 = ~n9479 & n9482 ;
  assign n9484 = ~\P1_reg2_reg[6]/NET0131  & ~n6070 ;
  assign n9485 = ~n9483 & ~n9484 ;
  assign n9486 = n1243 & n1736 ;
  assign n9487 = n3672 & ~n8943 ;
  assign n9488 = ~n9486 & ~n9487 ;
  assign n9489 = n6070 & ~n9488 ;
  assign n9490 = \P1_reg2_reg[7]/NET0131  & ~n6072 ;
  assign n9491 = ~n9489 & ~n9490 ;
  assign n9492 = \P2_reg2_reg[4]/NET0131  & ~n3434 ;
  assign n9494 = n2033 & ~n8963 ;
  assign n9498 = n2033 & n2849 ;
  assign n9497 = ~\P2_reg2_reg[4]/NET0131  & ~n2033 ;
  assign n9499 = n3375 & ~n9497 ;
  assign n9500 = ~n9498 & n9499 ;
  assign n9493 = n2853 & n3415 ;
  assign n9495 = ~n3418 & ~n6808 ;
  assign n9496 = \P2_reg2_reg[4]/NET0131  & ~n9495 ;
  assign n9501 = ~n9493 & ~n9496 ;
  assign n9502 = ~n9500 & n9501 ;
  assign n9503 = ~n9494 & n9502 ;
  assign n9504 = n2017 & ~n9503 ;
  assign n9505 = \P2_reg2_reg[4]/NET0131  & n3430 ;
  assign n9506 = ~n9504 & ~n9505 ;
  assign n9507 = \P1_state_reg[0]/NET0131  & ~n9506 ;
  assign n9508 = ~n9492 & ~n9507 ;
  assign n9509 = \P2_reg2_reg[7]/NET0131  & ~n3434 ;
  assign n9510 = \P2_reg2_reg[7]/NET0131  & n3430 ;
  assign n9512 = \P2_reg2_reg[7]/NET0131  & ~n2033 ;
  assign n9516 = n2033 & n8856 ;
  assign n9517 = ~n9512 & ~n9516 ;
  assign n9518 = n3373 & ~n9517 ;
  assign n9513 = n2033 & n8848 ;
  assign n9514 = ~n9512 & ~n9513 ;
  assign n9515 = n3179 & ~n9514 ;
  assign n9519 = n2033 & ~n8862 ;
  assign n9520 = ~n9512 & ~n9519 ;
  assign n9521 = n3319 & ~n9520 ;
  assign n9522 = n2033 & n8867 ;
  assign n9523 = ~n9512 & ~n9522 ;
  assign n9524 = n3409 & ~n9523 ;
  assign n9525 = n2033 & n2719 ;
  assign n9526 = ~n9512 & ~n9525 ;
  assign n9527 = n3375 & ~n9526 ;
  assign n9511 = n2698 & n3415 ;
  assign n9528 = \P2_reg2_reg[7]/NET0131  & n3418 ;
  assign n9529 = ~n9511 & ~n9528 ;
  assign n9530 = ~n9527 & n9529 ;
  assign n9531 = ~n9524 & n9530 ;
  assign n9532 = ~n9521 & n9531 ;
  assign n9533 = ~n9515 & n9532 ;
  assign n9534 = ~n9518 & n9533 ;
  assign n9535 = n2017 & ~n9534 ;
  assign n9536 = ~n9510 & ~n9535 ;
  assign n9537 = \P1_state_reg[0]/NET0131  & ~n9536 ;
  assign n9538 = ~n9509 & ~n9537 ;
  assign n9539 = n6171 & ~n9444 ;
  assign n9540 = \P1_reg0_reg[3]/NET0131  & ~n6238 ;
  assign n9541 = ~n9539 & ~n9540 ;
  assign n9542 = n6171 & ~n8943 ;
  assign n9543 = \P1_reg0_reg[7]/NET0131  & ~n6169 ;
  assign n9544 = ~n9542 & ~n9543 ;
  assign n9545 = \P2_reg0_reg[14]/NET0131  & ~n3434 ;
  assign n9546 = \P2_reg0_reg[14]/NET0131  & n3430 ;
  assign n9548 = \P2_reg0_reg[14]/NET0131  & ~n4610 ;
  assign n9549 = n4610 & n8070 ;
  assign n9550 = ~n9548 & ~n9549 ;
  assign n9551 = n3319 & ~n9550 ;
  assign n9555 = n4610 & ~n8076 ;
  assign n9556 = ~n9548 & ~n9555 ;
  assign n9557 = n3179 & ~n9556 ;
  assign n9552 = n4610 & n8084 ;
  assign n9553 = ~n9548 & ~n9552 ;
  assign n9554 = n3373 & ~n9553 ;
  assign n9547 = n4610 & ~n9135 ;
  assign n9558 = \P2_reg0_reg[14]/NET0131  & ~n4621 ;
  assign n9559 = ~n9547 & ~n9558 ;
  assign n9560 = ~n9554 & n9559 ;
  assign n9561 = ~n9557 & n9560 ;
  assign n9562 = ~n9551 & n9561 ;
  assign n9563 = n2017 & ~n9562 ;
  assign n9564 = ~n9546 & ~n9563 ;
  assign n9565 = \P1_state_reg[0]/NET0131  & ~n9564 ;
  assign n9566 = ~n9545 & ~n9565 ;
  assign n9568 = \P1_reg1_reg[3]/NET0131  & ~n4236 ;
  assign n9569 = n6246 & n8750 ;
  assign n9570 = ~n9568 & ~n9569 ;
  assign n9571 = n1898 & ~n9570 ;
  assign n9567 = n6246 & ~n9442 ;
  assign n9572 = \P1_reg1_reg[3]/NET0131  & ~n9228 ;
  assign n9573 = ~n9567 & ~n9572 ;
  assign n9574 = ~n9571 & n9573 ;
  assign n9575 = n1322 & ~n3579 ;
  assign n9576 = ~n3580 & ~n9575 ;
  assign n9577 = ~n536 & ~n9576 ;
  assign n9578 = n536 & n1367 ;
  assign n9579 = ~n9577 & ~n9578 ;
  assign n9580 = n1898 & n9579 ;
  assign n9590 = ~n1400 & n1759 ;
  assign n9589 = n1400 & ~n1759 ;
  assign n9591 = n3575 & ~n9589 ;
  assign n9592 = ~n9590 & n9591 ;
  assign n9586 = ~n1759 & ~n3471 ;
  assign n9585 = n1759 & n3471 ;
  assign n9587 = n3557 & ~n9585 ;
  assign n9588 = ~n9586 & n9587 ;
  assign n9581 = ~n1358 & n3683 ;
  assign n9582 = ~n1358 & ~n3626 ;
  assign n9583 = ~n3627 & n3650 ;
  assign n9584 = ~n9582 & n9583 ;
  assign n9593 = ~n9581 & ~n9584 ;
  assign n9594 = ~n9588 & n9593 ;
  assign n9595 = ~n9592 & n9594 ;
  assign n9596 = ~n9580 & n9595 ;
  assign n9597 = n3450 & ~n9596 ;
  assign n9598 = ~n1358 & n1736 ;
  assign n9599 = ~n9597 & ~n9598 ;
  assign n9600 = n6070 & ~n9599 ;
  assign n9601 = n3450 & ~n9579 ;
  assign n9602 = n1898 & ~n9601 ;
  assign n9603 = n6070 & n8129 ;
  assign n9604 = ~n9602 & n9603 ;
  assign n9605 = \P1_reg3_reg[2]/NET0131  & ~n9604 ;
  assign n9606 = ~n9600 & ~n9605 ;
  assign n9607 = n6246 & ~n8905 ;
  assign n9608 = ~n1735 & ~n3615 ;
  assign n9609 = ~n4236 & n9608 ;
  assign n9610 = n6070 & ~n9609 ;
  assign n9611 = n6889 & n9610 ;
  assign n9612 = \P1_reg1_reg[6]/NET0131  & ~n9611 ;
  assign n9613 = ~n9607 & ~n9612 ;
  assign n9615 = \P2_reg0_reg[3]/NET0131  & ~n4610 ;
  assign n9616 = n4610 & n9251 ;
  assign n9617 = ~n9615 & ~n9616 ;
  assign n9618 = n3373 & ~n9617 ;
  assign n9619 = n4610 & ~n9257 ;
  assign n9620 = ~n9615 & ~n9619 ;
  assign n9621 = n3179 & ~n9620 ;
  assign n9614 = \P2_reg0_reg[3]/NET0131  & ~n8958 ;
  assign n9623 = n3319 & ~n9264 ;
  assign n9622 = ~n2880 & n3375 ;
  assign n9624 = ~n9270 & ~n9622 ;
  assign n9625 = ~n9623 & n9624 ;
  assign n9626 = n4610 & ~n9625 ;
  assign n9627 = ~n9614 & ~n9626 ;
  assign n9628 = ~n9621 & n9627 ;
  assign n9629 = ~n9618 & n9628 ;
  assign n9630 = n2017 & ~n9629 ;
  assign n9631 = \P2_reg0_reg[3]/NET0131  & n3430 ;
  assign n9632 = ~n9630 & ~n9631 ;
  assign n9633 = \P1_state_reg[0]/NET0131  & ~n9632 ;
  assign n9634 = \P2_reg0_reg[3]/NET0131  & ~n3434 ;
  assign n9635 = ~n9633 & ~n9634 ;
  assign n9636 = \P2_reg1_reg[3]/NET0131  & ~n3434 ;
  assign n9638 = \P2_reg1_reg[3]/NET0131  & ~n4663 ;
  assign n9639 = n4663 & n9251 ;
  assign n9640 = ~n9638 & ~n9639 ;
  assign n9641 = n3373 & ~n9640 ;
  assign n9642 = n4663 & ~n9257 ;
  assign n9643 = ~n9638 & ~n9642 ;
  assign n9644 = n3179 & ~n9643 ;
  assign n9637 = \P2_reg1_reg[3]/NET0131  & ~n6719 ;
  assign n9645 = n4663 & ~n9625 ;
  assign n9646 = ~n9637 & ~n9645 ;
  assign n9647 = ~n9644 & n9646 ;
  assign n9648 = ~n9641 & n9647 ;
  assign n9649 = n2017 & ~n9648 ;
  assign n9650 = \P2_reg1_reg[3]/NET0131  & n3430 ;
  assign n9651 = ~n9649 & ~n9650 ;
  assign n9652 = \P1_state_reg[0]/NET0131  & ~n9651 ;
  assign n9653 = ~n9636 & ~n9652 ;
  assign n9655 = n2033 & n9251 ;
  assign n9656 = \P2_reg2_reg[3]/NET0131  & ~n2033 ;
  assign n9657 = ~n9655 & ~n9656 ;
  assign n9658 = n3373 & ~n9657 ;
  assign n9659 = n2033 & ~n9257 ;
  assign n9660 = ~n9656 & ~n9659 ;
  assign n9661 = n3179 & ~n9660 ;
  assign n9662 = n2033 & ~n9264 ;
  assign n9663 = ~n9656 & ~n9662 ;
  assign n9664 = n3319 & ~n9663 ;
  assign n9665 = n2033 & n9269 ;
  assign n9666 = ~n9656 & ~n9665 ;
  assign n9667 = n3409 & ~n9666 ;
  assign n9668 = n2033 & ~n2880 ;
  assign n9669 = ~n9656 & ~n9668 ;
  assign n9670 = n3375 & ~n9669 ;
  assign n9654 = ~\P2_reg3_reg[3]/NET0131  & n3415 ;
  assign n9671 = \P2_reg2_reg[3]/NET0131  & n3418 ;
  assign n9672 = ~n9654 & ~n9671 ;
  assign n9673 = ~n9670 & n9672 ;
  assign n9674 = ~n9667 & n9673 ;
  assign n9675 = ~n9664 & n9674 ;
  assign n9676 = ~n9661 & n9675 ;
  assign n9677 = ~n9658 & n9676 ;
  assign n9678 = n2017 & ~n9677 ;
  assign n9679 = \P2_reg2_reg[3]/NET0131  & n3430 ;
  assign n9680 = ~n9678 & ~n9679 ;
  assign n9681 = \P1_state_reg[0]/NET0131  & ~n9680 ;
  assign n9682 = \P2_reg2_reg[3]/NET0131  & ~n3434 ;
  assign n9683 = ~n9681 & ~n9682 ;
  assign n9684 = \P2_reg2_reg[6]/NET0131  & ~n3434 ;
  assign n9685 = \P2_reg2_reg[6]/NET0131  & n3430 ;
  assign n9687 = \P2_reg2_reg[6]/NET0131  & ~n2033 ;
  assign n9692 = n2033 & ~n9292 ;
  assign n9693 = ~n9687 & ~n9692 ;
  assign n9694 = n3373 & ~n9693 ;
  assign n9688 = n2033 & n9298 ;
  assign n9689 = ~n9687 & ~n9688 ;
  assign n9690 = n3179 & ~n9689 ;
  assign n9696 = n3319 & ~n9304 ;
  assign n9695 = n2745 & n3375 ;
  assign n9697 = ~n9310 & ~n9695 ;
  assign n9698 = ~n9696 & n9697 ;
  assign n9699 = n2033 & ~n9698 ;
  assign n9686 = n2726 & n3415 ;
  assign n9691 = \P2_reg2_reg[6]/NET0131  & ~n9334 ;
  assign n9700 = ~n9686 & ~n9691 ;
  assign n9701 = ~n9699 & n9700 ;
  assign n9702 = ~n9690 & n9701 ;
  assign n9703 = ~n9694 & n9702 ;
  assign n9704 = n2017 & ~n9703 ;
  assign n9705 = ~n9685 & ~n9704 ;
  assign n9706 = \P1_state_reg[0]/NET0131  & ~n9705 ;
  assign n9707 = ~n9684 & ~n9706 ;
  assign n9708 = \P1_reg0_reg[6]/NET0131  & ~n6169 ;
  assign n9709 = n6171 & ~n8905 ;
  assign n9710 = ~n9708 & ~n9709 ;
  assign n9712 = \P2_reg0_reg[6]/NET0131  & ~n4610 ;
  assign n9713 = n4610 & ~n9292 ;
  assign n9714 = ~n9712 & ~n9713 ;
  assign n9715 = n3373 & ~n9714 ;
  assign n9716 = n4610 & n9298 ;
  assign n9717 = ~n9712 & ~n9716 ;
  assign n9718 = n3179 & ~n9717 ;
  assign n9711 = \P2_reg0_reg[6]/NET0131  & ~n8958 ;
  assign n9719 = n4610 & ~n9698 ;
  assign n9720 = ~n9711 & ~n9719 ;
  assign n9721 = ~n9718 & n9720 ;
  assign n9722 = ~n9715 & n9721 ;
  assign n9723 = n2017 & ~n9722 ;
  assign n9724 = \P2_reg0_reg[6]/NET0131  & n3430 ;
  assign n9725 = ~n9723 & ~n9724 ;
  assign n9726 = \P1_state_reg[0]/NET0131  & ~n9725 ;
  assign n9727 = \P2_reg0_reg[6]/NET0131  & ~n3434 ;
  assign n9728 = ~n9726 & ~n9727 ;
  assign n9729 = ~\P1_reg2_reg[2]/NET0131  & ~n3672 ;
  assign n9730 = n3672 & ~n9579 ;
  assign n9731 = n1898 & ~n9730 ;
  assign n9732 = n3672 & ~n9595 ;
  assign n9733 = n6070 & ~n9732 ;
  assign n9734 = ~n9731 & n9733 ;
  assign n9735 = ~n9729 & ~n9734 ;
  assign n9736 = \P1_reg3_reg[2]/NET0131  & n1736 ;
  assign n9737 = \P1_reg2_reg[2]/NET0131  & ~n8989 ;
  assign n9738 = ~n9736 & ~n9737 ;
  assign n9739 = ~n9735 & n9738 ;
  assign n9740 = ~\P1_reg2_reg[2]/NET0131  & ~n6070 ;
  assign n9741 = ~n9739 & ~n9740 ;
  assign n9743 = \P2_reg1_reg[6]/NET0131  & ~n4663 ;
  assign n9744 = n4663 & ~n9292 ;
  assign n9745 = ~n9743 & ~n9744 ;
  assign n9746 = n3373 & ~n9745 ;
  assign n9747 = n4663 & n9298 ;
  assign n9748 = ~n9743 & ~n9747 ;
  assign n9749 = n3179 & ~n9748 ;
  assign n9742 = \P2_reg1_reg[6]/NET0131  & ~n6719 ;
  assign n9750 = n4663 & ~n9698 ;
  assign n9751 = ~n9742 & ~n9750 ;
  assign n9752 = ~n9749 & n9751 ;
  assign n9753 = ~n9746 & n9752 ;
  assign n9754 = n2017 & ~n9753 ;
  assign n9755 = \P2_reg1_reg[6]/NET0131  & n3430 ;
  assign n9756 = ~n9754 & ~n9755 ;
  assign n9757 = \P1_state_reg[0]/NET0131  & ~n9756 ;
  assign n9758 = \P2_reg1_reg[6]/NET0131  & ~n3434 ;
  assign n9759 = ~n9757 & ~n9758 ;
  assign n9760 = \P1_reg0_reg[2]/NET0131  & ~n6169 ;
  assign n9761 = n6171 & ~n9596 ;
  assign n9762 = ~n9760 & ~n9761 ;
  assign n9763 = n6246 & ~n9596 ;
  assign n9764 = \P1_reg1_reg[2]/NET0131  & ~n8721 ;
  assign n9765 = ~n9763 & ~n9764 ;
  assign n9766 = ~n1381 & n3655 ;
  assign n9767 = n1344 & ~n3578 ;
  assign n9768 = ~n3579 & ~n9767 ;
  assign n9769 = ~n536 & ~n9768 ;
  assign n9770 = n536 & n1390 ;
  assign n9771 = ~n9769 & ~n9770 ;
  assign n9772 = n1898 & n9771 ;
  assign n9781 = n1398 & ~n1755 ;
  assign n9780 = ~n1398 & n1755 ;
  assign n9782 = n3575 & ~n9780 ;
  assign n9783 = ~n9781 & n9782 ;
  assign n9773 = ~n1381 & ~n1397 ;
  assign n9774 = ~n3626 & n3650 ;
  assign n9775 = ~n9773 & n9774 ;
  assign n9777 = ~n1755 & n3467 ;
  assign n9776 = n1755 & ~n3467 ;
  assign n9778 = n3557 & ~n9776 ;
  assign n9779 = ~n9777 & n9778 ;
  assign n9784 = ~n9775 & ~n9779 ;
  assign n9785 = ~n9783 & n9784 ;
  assign n9786 = ~n9772 & n9785 ;
  assign n9787 = n3450 & ~n9786 ;
  assign n9788 = ~n9766 & ~n9787 ;
  assign n9789 = n6070 & ~n9788 ;
  assign n9790 = n6070 & ~n6590 ;
  assign n9791 = n7033 & n9790 ;
  assign n9792 = \P1_reg3_reg[1]/NET0131  & ~n9791 ;
  assign n9793 = ~n9789 & ~n9792 ;
  assign n9794 = ~\P2_reg3_reg[1]/NET0131  & ~n4925 ;
  assign n9795 = n2777 & ~n3331 ;
  assign n9796 = ~n3332 & ~n9795 ;
  assign n9797 = ~n2050 & ~n9796 ;
  assign n9798 = n2050 & n2823 ;
  assign n9799 = ~n9797 & ~n9798 ;
  assign n9800 = n4925 & ~n9799 ;
  assign n9801 = n3373 & ~n9800 ;
  assign n9802 = ~n2814 & ~n2830 ;
  assign n9803 = ~n3377 & ~n9802 ;
  assign n9804 = n3409 & n9803 ;
  assign n9805 = n3198 & ~n4124 ;
  assign n9806 = n3319 & ~n4125 ;
  assign n9807 = ~n9805 & n9806 ;
  assign n9809 = ~n2831 & n4124 ;
  assign n9808 = n2831 & ~n4124 ;
  assign n9810 = n3179 & ~n9808 ;
  assign n9811 = ~n9809 & n9810 ;
  assign n9812 = ~n9807 & ~n9811 ;
  assign n9813 = ~n9804 & n9812 ;
  assign n9814 = n4925 & ~n9813 ;
  assign n9815 = n4275 & ~n9814 ;
  assign n9816 = ~n9801 & n9815 ;
  assign n9817 = ~n9794 & ~n9816 ;
  assign n9818 = ~n2814 & ~n5093 ;
  assign n9819 = ~n9817 & ~n9818 ;
  assign n9820 = n4275 & ~n9819 ;
  assign n9821 = ~\P2_reg3_reg[1]/NET0131  & ~n9820 ;
  assign n9822 = ~n3178 & ~n3408 ;
  assign n9823 = ~n4925 & ~n9822 ;
  assign n9824 = ~n5090 & ~n9823 ;
  assign n9825 = n9819 & n9824 ;
  assign n9826 = ~n9821 & ~n9825 ;
  assign n9827 = ~\P2_reg3_reg[2]/NET0131  & ~n4925 ;
  assign n9828 = n2866 & ~n3332 ;
  assign n9829 = ~n3333 & ~n9828 ;
  assign n9830 = ~n2050 & ~n9829 ;
  assign n9831 = n2050 & n2800 ;
  assign n9832 = ~n9830 & ~n9831 ;
  assign n9833 = n4925 & ~n9832 ;
  assign n9834 = n3373 & ~n9833 ;
  assign n9843 = n2833 & ~n4134 ;
  assign n9842 = ~n2833 & n4134 ;
  assign n9844 = n3179 & ~n9842 ;
  assign n9845 = ~n9843 & n9844 ;
  assign n9835 = ~n2791 & ~n3377 ;
  assign n9836 = ~n3378 & n3409 ;
  assign n9837 = ~n9835 & n9836 ;
  assign n9839 = ~n4093 & n4134 ;
  assign n9838 = n4093 & ~n4134 ;
  assign n9840 = n3319 & ~n9838 ;
  assign n9841 = ~n9839 & n9840 ;
  assign n9846 = ~n9837 & ~n9841 ;
  assign n9847 = ~n9845 & n9846 ;
  assign n9848 = n4925 & ~n9847 ;
  assign n9849 = n4275 & ~n9848 ;
  assign n9850 = ~n9834 & n9849 ;
  assign n9851 = ~n9827 & ~n9850 ;
  assign n9852 = ~n2791 & ~n5093 ;
  assign n9853 = ~n9851 & ~n9852 ;
  assign n9854 = n4275 & ~n9853 ;
  assign n9855 = ~\P2_reg3_reg[2]/NET0131  & ~n9854 ;
  assign n9856 = n9824 & n9853 ;
  assign n9857 = ~n9855 & ~n9856 ;
  assign n9858 = ~n2791 & n3375 ;
  assign n9859 = n9847 & ~n9858 ;
  assign n9860 = n3373 & n9832 ;
  assign n9861 = n9859 & ~n9860 ;
  assign n9862 = n5385 & ~n9861 ;
  assign n9863 = \P2_reg0_reg[2]/NET0131  & ~n7982 ;
  assign n9864 = ~n9862 & ~n9863 ;
  assign n9865 = \P2_reg1_reg[2]/NET0131  & ~n3434 ;
  assign n9866 = \P2_reg1_reg[2]/NET0131  & n3430 ;
  assign n9867 = n4663 & ~n9861 ;
  assign n9868 = \P2_reg1_reg[2]/NET0131  & ~n5568 ;
  assign n9869 = ~n9867 & ~n9868 ;
  assign n9870 = n2017 & ~n9869 ;
  assign n9871 = ~n9866 & ~n9870 ;
  assign n9872 = \P1_state_reg[0]/NET0131  & ~n9871 ;
  assign n9873 = ~n9865 & ~n9872 ;
  assign n9874 = \P1_reg0_reg[1]/NET0131  & ~n3703 ;
  assign n9875 = \P1_reg0_reg[1]/NET0131  & n3664 ;
  assign n9876 = ~n1381 & n3683 ;
  assign n9877 = n9785 & ~n9876 ;
  assign n9878 = ~n9772 & n9877 ;
  assign n9879 = n3900 & ~n9878 ;
  assign n9880 = \P1_reg0_reg[1]/NET0131  & ~n6177 ;
  assign n9881 = ~n9879 & ~n9880 ;
  assign n9882 = n3662 & ~n9881 ;
  assign n9883 = ~n9875 & ~n9882 ;
  assign n9884 = \P1_state_reg[0]/NET0131  & ~n9883 ;
  assign n9885 = ~n9874 & ~n9884 ;
  assign n9887 = \P1_reg1_reg[1]/NET0131  & ~n4236 ;
  assign n9888 = n6246 & n9771 ;
  assign n9889 = ~n9887 & ~n9888 ;
  assign n9890 = n1898 & ~n9889 ;
  assign n9886 = n6246 & ~n9877 ;
  assign n9891 = ~n6273 & n7908 ;
  assign n9892 = \P1_reg1_reg[1]/NET0131  & ~n9891 ;
  assign n9893 = ~n9886 & ~n9892 ;
  assign n9894 = ~n9890 & n9893 ;
  assign n9895 = \P2_reg2_reg[1]/NET0131  & ~n3434 ;
  assign n9896 = \P2_reg2_reg[1]/NET0131  & n3430 ;
  assign n9903 = \P2_reg2_reg[1]/NET0131  & ~n2033 ;
  assign n9904 = n2033 & n9799 ;
  assign n9905 = ~n9903 & ~n9904 ;
  assign n9906 = n3373 & ~n9905 ;
  assign n9900 = ~n2814 & n3375 ;
  assign n9901 = n9812 & ~n9900 ;
  assign n9902 = n2033 & ~n9901 ;
  assign n9907 = n2033 & n9803 ;
  assign n9908 = ~n9903 & ~n9907 ;
  assign n9909 = n3409 & ~n9908 ;
  assign n9897 = \P2_reg3_reg[1]/NET0131  & n3415 ;
  assign n9898 = ~n4434 & n6795 ;
  assign n9899 = \P2_reg2_reg[1]/NET0131  & ~n9898 ;
  assign n9910 = ~n9897 & ~n9899 ;
  assign n9911 = ~n9909 & n9910 ;
  assign n9912 = ~n9902 & n9911 ;
  assign n9913 = ~n9906 & n9912 ;
  assign n9914 = n2017 & ~n9913 ;
  assign n9915 = ~n9896 & ~n9914 ;
  assign n9916 = \P1_state_reg[0]/NET0131  & ~n9915 ;
  assign n9917 = ~n9895 & ~n9916 ;
  assign n9918 = \P1_reg3_reg[1]/NET0131  & n1736 ;
  assign n9919 = n3672 & ~n9878 ;
  assign n9920 = ~n9918 & ~n9919 ;
  assign n9921 = n6070 & ~n9920 ;
  assign n9922 = n3555 & n8988 ;
  assign n9923 = ~n5429 & n6070 ;
  assign n9924 = ~n9922 & n9923 ;
  assign n9925 = n6694 & n9924 ;
  assign n9926 = \P1_reg2_reg[1]/NET0131  & ~n9925 ;
  assign n9927 = ~n9921 & ~n9926 ;
  assign n9928 = \P2_reg1_reg[1]/NET0131  & ~n3434 ;
  assign n9929 = n3373 & n9799 ;
  assign n9930 = ~n9804 & n9901 ;
  assign n9931 = ~n9929 & n9930 ;
  assign n9932 = n5571 & ~n9931 ;
  assign n9933 = \P2_reg1_reg[1]/NET0131  & ~n1984 ;
  assign n9934 = ~n6748 & n9933 ;
  assign n9935 = ~n9932 & ~n9934 ;
  assign n9936 = \P1_state_reg[0]/NET0131  & ~n9935 ;
  assign n9937 = ~n9928 & ~n9936 ;
  assign n9938 = ~\P2_reg2_reg[2]/NET0131  & ~n2033 ;
  assign n9940 = n2033 & ~n9832 ;
  assign n9941 = n3373 & ~n9940 ;
  assign n9939 = n2033 & ~n9859 ;
  assign n9942 = n4275 & ~n9939 ;
  assign n9943 = ~n9941 & n9942 ;
  assign n9944 = ~n9938 & ~n9943 ;
  assign n9945 = \P2_reg3_reg[2]/NET0131  & n3415 ;
  assign n9946 = ~n9944 & ~n9945 ;
  assign n9947 = n4275 & ~n9946 ;
  assign n9948 = ~\P2_reg2_reg[2]/NET0131  & ~n9947 ;
  assign n9949 = ~n3422 & n6795 ;
  assign n9950 = n9946 & n9949 ;
  assign n9951 = ~n9948 & ~n9950 ;
  assign n9953 = \P2_reg0_reg[1]/NET0131  & ~n4610 ;
  assign n9954 = n5385 & n9799 ;
  assign n9955 = ~n9953 & ~n9954 ;
  assign n9956 = n3373 & ~n9955 ;
  assign n9952 = n5385 & ~n9930 ;
  assign n9957 = n4275 & ~n7969 ;
  assign n9958 = n6901 & n9957 ;
  assign n9959 = \P2_reg0_reg[1]/NET0131  & ~n9958 ;
  assign n9960 = ~n9952 & ~n9959 ;
  assign n9961 = ~n9956 & n9960 ;
  assign n9964 = n1367 & ~n3577 ;
  assign n9965 = ~n536 & ~n3578 ;
  assign n9966 = ~n9964 & n9965 ;
  assign n9967 = n1898 & n9966 ;
  assign n9962 = ~n1397 & n3616 ;
  assign n9963 = ~n1739 & n3556 ;
  assign n9968 = ~n9962 & ~n9963 ;
  assign n9969 = ~n9967 & n9968 ;
  assign n9970 = n3450 & ~n9969 ;
  assign n9971 = ~n1397 & n1736 ;
  assign n9972 = ~n9970 & ~n9971 ;
  assign n9973 = n6070 & ~n9972 ;
  assign n9974 = n3450 & ~n9966 ;
  assign n9975 = n1898 & ~n9974 ;
  assign n9976 = n9603 & ~n9975 ;
  assign n9977 = \P1_reg3_reg[0]/NET0131  & ~n9976 ;
  assign n9978 = ~n9973 & ~n9977 ;
  assign n9982 = n2800 & ~n3330 ;
  assign n9983 = ~n2050 & n3373 ;
  assign n9984 = ~n3331 & n9983 ;
  assign n9985 = ~n9982 & n9984 ;
  assign n9979 = ~n2830 & n3420 ;
  assign n9980 = ~n3198 & ~n4015 ;
  assign n9981 = ~n5935 & ~n9980 ;
  assign n9986 = ~n9979 & ~n9981 ;
  assign n9987 = ~n9985 & n9986 ;
  assign n9988 = n4925 & ~n9987 ;
  assign n9989 = ~n2830 & n3415 ;
  assign n9990 = ~n9988 & ~n9989 ;
  assign n9991 = n4275 & ~n9990 ;
  assign n9992 = n4275 & ~n9985 ;
  assign n9993 = ~n7320 & n9992 ;
  assign n9994 = \P2_reg3_reg[0]/NET0131  & ~n9993 ;
  assign n9995 = ~n9991 & ~n9994 ;
  assign n9996 = n3672 & ~n9969 ;
  assign n9997 = \P1_reg3_reg[0]/NET0131  & n1736 ;
  assign n9998 = ~n9996 & ~n9997 ;
  assign n9999 = n6070 & ~n9998 ;
  assign n10000 = n3672 & ~n9966 ;
  assign n10001 = n1898 & ~n10000 ;
  assign n10002 = n6070 & n8989 ;
  assign n10003 = ~n10001 & n10002 ;
  assign n10004 = \P1_reg2_reg[0]/NET0131  & ~n10003 ;
  assign n10005 = ~n9999 & ~n10004 ;
  assign n10006 = n5572 & ~n9987 ;
  assign n10007 = \P2_reg1_reg[0]/NET0131  & ~n6749 ;
  assign n10008 = ~n10006 & ~n10007 ;
  assign n10009 = \P1_reg0_reg[0]/NET0131  & ~n6238 ;
  assign n10010 = n6171 & ~n9969 ;
  assign n10011 = ~n10009 & ~n10010 ;
  assign n10012 = n2033 & ~n9987 ;
  assign n10013 = \P2_reg3_reg[0]/NET0131  & n3415 ;
  assign n10014 = ~n10012 & ~n10013 ;
  assign n10015 = n4275 & ~n10014 ;
  assign n10016 = ~n2033 & ~n5605 ;
  assign n10017 = ~n3422 & ~n10016 ;
  assign n10018 = n9992 & n10017 ;
  assign n10019 = \P2_reg2_reg[0]/NET0131  & ~n10018 ;
  assign n10020 = ~n10015 & ~n10019 ;
  assign n10021 = \P1_reg1_reg[0]/NET0131  & ~n9611 ;
  assign n10022 = n6246 & ~n9969 ;
  assign n10023 = ~n10021 & ~n10022 ;
  assign n10024 = n5385 & ~n9987 ;
  assign n10025 = ~n4622 & n9958 ;
  assign n10026 = \P2_reg0_reg[0]/NET0131  & ~n10025 ;
  assign n10027 = ~n10024 & ~n10026 ;
  assign n10028 = \P1_state_reg[0]/NET0131  & ~n1949 ;
  assign n10029 = ~\P1_state_reg[0]/NET0131  & n1532 ;
  assign n10030 = ~n10028 & ~n10029 ;
  assign n10031 = ~\P1_state_reg[0]/NET0131  & ~n1499 ;
  assign n10032 = \P1_state_reg[0]/NET0131  & ~n527 ;
  assign n10033 = ~n10031 & ~n10032 ;
  assign n10034 = ~\P1_state_reg[0]/NET0131  & ~n2451 ;
  assign n10035 = \P1_state_reg[0]/NET0131  & ~n1994 ;
  assign n10036 = ~n10034 & ~n10035 ;
  assign n10037 = ~\P1_state_reg[0]/NET0131  & ~n2375 ;
  assign n10038 = \P1_state_reg[0]/NET0131  & n2043 ;
  assign n10039 = ~n10037 & ~n10038 ;
  assign n10040 = ~\P1_state_reg[0]/NET0131  & ~n1462 ;
  assign n10041 = \P1_state_reg[0]/NET0131  & ~n1939 ;
  assign n10042 = ~n10040 & ~n10041 ;
  assign n10043 = ~\P1_state_reg[0]/NET0131  & ~n2423 ;
  assign n10044 = \P1_state_reg[0]/NET0131  & ~n2014 ;
  assign n10045 = ~n10043 & ~n10044 ;
  assign n10046 = ~\P1_state_reg[0]/NET0131  & ~n2470 ;
  assign n10047 = \P1_state_reg[0]/NET0131  & n2007 ;
  assign n10048 = ~n10046 & ~n10047 ;
  assign n10049 = \P1_state_reg[0]/NET0131  & ~n2970 ;
  assign n10050 = ~\P1_state_reg[0]/NET0131  & n2978 ;
  assign n10051 = ~n10049 & ~n10050 ;
  assign n10052 = \P1_state_reg[0]/NET0131  & ~n2916 ;
  assign n10053 = ~\P1_state_reg[0]/NET0131  & n2924 ;
  assign n10054 = ~n10052 & ~n10053 ;
  assign n10055 = \P1_state_reg[0]/NET0131  & ~n2943 ;
  assign n10056 = ~\P1_state_reg[0]/NET0131  & n2952 ;
  assign n10057 = ~n10055 & ~n10056 ;
  assign n10058 = ~\P1_state_reg[0]/NET0131  & ~n3116 ;
  assign n10059 = \P1_state_reg[0]/NET0131  & ~n3108 ;
  assign n10060 = ~n10058 & ~n10059 ;
  assign n10061 = ~\P1_state_reg[0]/NET0131  & ~n3093 ;
  assign n10062 = \P1_state_reg[0]/NET0131  & n3085 ;
  assign n10063 = ~n10061 & ~n10062 ;
  assign n10064 = \P1_state_reg[0]/NET0131  & ~n3061 ;
  assign n10065 = ~\P1_state_reg[0]/NET0131  & n3069 ;
  assign n10066 = ~n10064 & ~n10065 ;
  assign n10067 = \P1_state_reg[0]/NET0131  & ~n3026 ;
  assign n10068 = ~\P1_state_reg[0]/NET0131  & n3034 ;
  assign n10069 = ~n10067 & ~n10068 ;
  assign n10070 = ~\P1_state_reg[0]/NET0131  & ~n2628 ;
  assign n10071 = \P1_state_reg[0]/NET0131  & n2619 ;
  assign n10072 = ~n10070 & ~n10071 ;
  assign n10073 = \P1_state_reg[0]/NET0131  & ~n2647 ;
  assign n10074 = ~\P1_state_reg[0]/NET0131  & n2655 ;
  assign n10075 = ~n10073 & ~n10074 ;
  assign n10076 = ~\P1_state_reg[0]/NET0131  & ~n2602 ;
  assign n10077 = \P1_state_reg[0]/NET0131  & n2592 ;
  assign n10078 = ~n10076 & ~n10077 ;
  assign n10079 = \P1_state_reg[0]/NET0131  & ~n2812 ;
  assign n10080 = ~\P1_state_reg[0]/NET0131  & n2807 ;
  assign n10081 = ~n10079 & ~n10080 ;
  assign n10082 = \P1_state_reg[0]/NET0131  & ~n3161 ;
  assign n10083 = ~\P1_state_reg[0]/NET0131  & n2578 ;
  assign n10084 = ~n10082 & ~n10083 ;
  assign n10085 = \P1_state_reg[0]/NET0131  & ~n3167 ;
  assign n10086 = ~\P1_state_reg[0]/NET0131  & n2540 ;
  assign n10087 = ~n10085 & ~n10086 ;
  assign n10088 = \P1_state_reg[0]/NET0131  & ~n3173 ;
  assign n10089 = ~\P1_state_reg[0]/NET0131  & n2521 ;
  assign n10090 = ~n10088 & ~n10089 ;
  assign n10091 = ~\P1_state_reg[0]/NET0131  & ~n2497 ;
  assign n10092 = ~n3935 & ~n10091 ;
  assign n10093 = ~\P1_state_reg[0]/NET0131  & ~n2314 ;
  assign n10094 = \P1_state_reg[0]/NET0131  & n2050 ;
  assign n10095 = ~n10093 & ~n10094 ;
  assign n10096 = \P1_state_reg[0]/NET0131  & ~n2205 ;
  assign n10097 = ~\P1_state_reg[0]/NET0131  & n2190 ;
  assign n10098 = ~n10096 & ~n10097 ;
  assign n10099 = ~\P1_state_reg[0]/NET0131  & ~n2784 ;
  assign n10100 = \P1_state_reg[0]/NET0131  & n2789 ;
  assign n10101 = ~n10099 & ~n10100 ;
  assign n10102 = ~\P1_state_reg[0]/NET0131  & ~n3976 ;
  assign n10103 = \P1_state_reg[0]/NET0131  & n2199 ;
  assign n10104 = ~n10102 & ~n10103 ;
  assign n10105 = ~\P1_state_reg[0]/NET0131  & ~n2878 ;
  assign n10106 = \P1_state_reg[0]/NET0131  & n2870 ;
  assign n10107 = ~n10105 & ~n10106 ;
  assign n10108 = \P1_state_reg[0]/NET0131  & ~n2847 ;
  assign n10109 = ~\P1_state_reg[0]/NET0131  & n2842 ;
  assign n10110 = ~n10108 & ~n10109 ;
  assign n10111 = ~\P1_state_reg[0]/NET0131  & ~n2766 ;
  assign n10112 = \P1_state_reg[0]/NET0131  & ~n2758 ;
  assign n10113 = ~n10111 & ~n10112 ;
  assign n10114 = \P1_state_reg[0]/NET0131  & ~n2735 ;
  assign n10115 = ~\P1_state_reg[0]/NET0131  & n2743 ;
  assign n10116 = ~n10114 & ~n10115 ;
  assign n10117 = \P1_state_reg[0]/NET0131  & ~n2709 ;
  assign n10118 = ~\P1_state_reg[0]/NET0131  & n2717 ;
  assign n10119 = ~n10117 & ~n10118 ;
  assign n10120 = ~\P1_state_reg[0]/NET0131  & ~n2690 ;
  assign n10121 = \P1_state_reg[0]/NET0131  & n2682 ;
  assign n10122 = ~n10120 & ~n10121 ;
  assign n10123 = \P1_state_reg[0]/NET0131  & ~n2995 ;
  assign n10124 = ~\P1_state_reg[0]/NET0131  & n3003 ;
  assign n10125 = ~n10123 & ~n10124 ;
  assign n10126 = ~\P1_state_reg[0]/NET0131  & ~n1145 ;
  assign n10127 = \P1_state_reg[0]/NET0131  & ~n1149 ;
  assign n10128 = ~n10126 & ~n10127 ;
  assign n10129 = ~\P1_state_reg[0]/NET0131  & ~n1122 ;
  assign n10130 = \P1_state_reg[0]/NET0131  & n1126 ;
  assign n10131 = ~n10129 & ~n10130 ;
  assign n10132 = ~\P1_state_reg[0]/NET0131  & ~n1083 ;
  assign n10133 = \P1_state_reg[0]/NET0131  & n1092 ;
  assign n10134 = ~n10132 & ~n10133 ;
  assign n10135 = ~\P1_state_reg[0]/NET0131  & ~n1058 ;
  assign n10136 = \P1_state_reg[0]/NET0131  & n1062 ;
  assign n10137 = ~n10135 & ~n10136 ;
  assign n10138 = ~\P1_state_reg[0]/NET0131  & ~n1033 ;
  assign n10139 = \P1_state_reg[0]/NET0131  & ~n1038 ;
  assign n10140 = ~n10138 & ~n10139 ;
  assign n10141 = ~\P1_state_reg[0]/NET0131  & ~n1006 ;
  assign n10142 = \P1_state_reg[0]/NET0131  & n1013 ;
  assign n10143 = ~n10141 & ~n10142 ;
  assign n10144 = ~\P1_state_reg[0]/NET0131  & ~n823 ;
  assign n10145 = \P1_state_reg[0]/NET0131  & n827 ;
  assign n10146 = ~n10144 & ~n10145 ;
  assign n10147 = ~\P1_state_reg[0]/NET0131  & ~n779 ;
  assign n10148 = \P1_state_reg[0]/NET0131  & n783 ;
  assign n10149 = ~n10147 & ~n10148 ;
  assign n10150 = ~\P1_state_reg[0]/NET0131  & ~n735 ;
  assign n10151 = \P1_state_reg[0]/NET0131  & n741 ;
  assign n10152 = ~n10150 & ~n10151 ;
  assign n10153 = ~\P1_state_reg[0]/NET0131  & ~n635 ;
  assign n10154 = \P1_state_reg[0]/NET0131  & ~n516 ;
  assign n10155 = ~n10153 & ~n10154 ;
  assign n10156 = \P1_state_reg[0]/NET0131  & ~n1371 ;
  assign n10157 = ~\P1_state_reg[0]/NET0131  & n1379 ;
  assign n10158 = ~n10156 & ~n10157 ;
  assign n10159 = \P1_state_reg[0]/NET0131  & ~n498 ;
  assign n10160 = ~\P1_state_reg[0]/NET0131  & n963 ;
  assign n10161 = ~n10159 & ~n10160 ;
  assign n10162 = \P1_state_reg[0]/NET0131  & ~n486 ;
  assign n10163 = ~\P1_state_reg[0]/NET0131  & n938 ;
  assign n10164 = ~n10162 & ~n10163 ;
  assign n10165 = \P1_state_reg[0]/NET0131  & ~n506 ;
  assign n10166 = ~\P1_state_reg[0]/NET0131  & n874 ;
  assign n10167 = ~n10165 & ~n10166 ;
  assign n10168 = ~\P1_state_reg[0]/NET0131  & ~n910 ;
  assign n10169 = ~n1934 & ~n10168 ;
  assign n10170 = \P1_state_reg[0]/NET0131  & ~n1944 ;
  assign n10171 = ~\P1_state_reg[0]/NET0131  & n1560 ;
  assign n10172 = ~n10170 & ~n10171 ;
  assign n10173 = ~\P1_state_reg[0]/NET0131  & ~n1636 ;
  assign n10174 = \P1_state_reg[0]/NET0131  & n536 ;
  assign n10175 = ~n10173 & ~n10174 ;
  assign n10176 = ~\P1_state_reg[0]/NET0131  & ~n1606 ;
  assign n10177 = \P1_state_reg[0]/NET0131  & n662 ;
  assign n10178 = ~n10176 & ~n10177 ;
  assign n10179 = ~\P1_state_reg[0]/NET0131  & ~n1351 ;
  assign n10180 = \P1_state_reg[0]/NET0131  & n1356 ;
  assign n10181 = ~n10179 & ~n10180 ;
  assign n10182 = ~\P1_state_reg[0]/NET0131  & ~n1695 ;
  assign n10183 = \P1_state_reg[0]/NET0131  & n650 ;
  assign n10184 = ~n10182 & ~n10183 ;
  assign n10185 = ~\P1_state_reg[0]/NET0131  & n1670 ;
  assign n10186 = ~\P1_IR_reg[29]/NET0131  & ~\P1_IR_reg[30]/NET0131  ;
  assign n10187 = \P1_IR_reg[31]/NET0131  & \P1_state_reg[0]/NET0131  ;
  assign n10188 = n10186 & n10187 ;
  assign n10189 = n643 & n10188 ;
  assign n10190 = n523 & n10189 ;
  assign n10191 = ~n10185 & ~n10190 ;
  assign n10192 = ~\P1_state_reg[0]/NET0131  & ~n1329 ;
  assign n10193 = \P1_state_reg[0]/NET0131  & n1334 ;
  assign n10194 = ~n10192 & ~n10193 ;
  assign n10195 = \P1_state_reg[0]/NET0131  & n1302 ;
  assign n10196 = ~\P1_state_reg[0]/NET0131  & n1311 ;
  assign n10197 = ~n10195 & ~n10196 ;
  assign n10198 = ~\P1_state_reg[0]/NET0131  & ~n1281 ;
  assign n10199 = \P1_state_reg[0]/NET0131  & ~n1286 ;
  assign n10200 = ~n10198 & ~n10199 ;
  assign n10201 = ~\P1_state_reg[0]/NET0131  & ~n1230 ;
  assign n10202 = \P1_state_reg[0]/NET0131  & n1236 ;
  assign n10203 = ~n10201 & ~n10202 ;
  assign n10204 = ~\P1_state_reg[0]/NET0131  & ~n1255 ;
  assign n10205 = \P1_state_reg[0]/NET0131  & n1261 ;
  assign n10206 = ~n10204 & ~n10205 ;
  assign n10207 = ~\P1_state_reg[0]/NET0131  & ~n1196 ;
  assign n10208 = \P1_state_reg[0]/NET0131  & ~n1200 ;
  assign n10209 = ~n10207 & ~n10208 ;
  assign n10210 = ~\P1_state_reg[0]/NET0131  & ~n1169 ;
  assign n10211 = \P1_state_reg[0]/NET0131  & n1176 ;
  assign n10212 = ~n10210 & ~n10211 ;
  assign n10213 = ~\P1_state_reg[0]/NET0131  & n3956 ;
  assign n10214 = \P1_state_reg[0]/NET0131  & ~\P2_IR_reg[29]/NET0131  ;
  assign n10215 = ~\P2_IR_reg[30]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n10216 = n10214 & n10215 ;
  assign n10217 = n2192 & n10216 ;
  assign n10218 = n2039 & n10217 ;
  assign n10219 = ~n10213 & ~n10218 ;
  assign n10259 = \P2_reg1_reg[6]/NET0131  & n2735 ;
  assign n10260 = ~\P2_reg1_reg[6]/NET0131  & ~n2735 ;
  assign n10261 = ~n10259 & ~n10260 ;
  assign n10262 = \P2_reg1_reg[5]/NET0131  & ~n2758 ;
  assign n10263 = ~\P2_reg1_reg[5]/NET0131  & n2758 ;
  assign n10264 = \P2_reg1_reg[4]/NET0131  & ~n2847 ;
  assign n10265 = ~\P2_reg1_reg[4]/NET0131  & n2847 ;
  assign n10266 = \P2_reg1_reg[3]/NET0131  & n2870 ;
  assign n10267 = ~\P2_reg1_reg[3]/NET0131  & ~n2870 ;
  assign n10268 = \P2_reg1_reg[2]/NET0131  & n2789 ;
  assign n10269 = ~\P2_reg1_reg[2]/NET0131  & ~n2789 ;
  assign n10270 = \P2_reg1_reg[1]/NET0131  & ~n2812 ;
  assign n10271 = ~\P2_reg1_reg[1]/NET0131  & n2812 ;
  assign n10272 = \P2_IR_reg[0]/NET0131  & \P2_reg1_reg[0]/NET0131  ;
  assign n10273 = ~n10271 & n10272 ;
  assign n10274 = ~n10270 & ~n10273 ;
  assign n10275 = ~n10269 & ~n10274 ;
  assign n10276 = ~n10268 & ~n10275 ;
  assign n10277 = ~n10267 & ~n10276 ;
  assign n10278 = ~n10266 & ~n10277 ;
  assign n10279 = ~n10265 & ~n10278 ;
  assign n10280 = ~n10264 & ~n10279 ;
  assign n10281 = ~n10263 & ~n10280 ;
  assign n10282 = ~n10262 & ~n10281 ;
  assign n10284 = ~n10261 & n10282 ;
  assign n10258 = ~n2043 & n2050 ;
  assign n10283 = n10261 & ~n10282 ;
  assign n10285 = n10258 & ~n10283 ;
  assign n10286 = ~n10284 & n10285 ;
  assign n10230 = \P2_reg2_reg[6]/NET0131  & n2735 ;
  assign n10231 = ~\P2_reg2_reg[6]/NET0131  & ~n2735 ;
  assign n10232 = ~n10230 & ~n10231 ;
  assign n10233 = \P2_reg2_reg[5]/NET0131  & ~n2758 ;
  assign n10234 = ~\P2_reg2_reg[5]/NET0131  & n2758 ;
  assign n10235 = \P2_reg2_reg[4]/NET0131  & ~n2847 ;
  assign n10236 = ~\P2_reg2_reg[4]/NET0131  & n2847 ;
  assign n10237 = \P2_reg2_reg[3]/NET0131  & n2870 ;
  assign n10238 = ~\P2_reg2_reg[3]/NET0131  & ~n2870 ;
  assign n10239 = \P2_reg2_reg[2]/NET0131  & n2789 ;
  assign n10240 = ~\P2_reg2_reg[2]/NET0131  & ~n2789 ;
  assign n10241 = \P2_reg2_reg[1]/NET0131  & ~n2812 ;
  assign n10242 = ~\P2_reg2_reg[1]/NET0131  & n2812 ;
  assign n10243 = \P2_IR_reg[0]/NET0131  & \P2_reg2_reg[0]/NET0131  ;
  assign n10244 = ~n10242 & n10243 ;
  assign n10245 = ~n10241 & ~n10244 ;
  assign n10246 = ~n10240 & ~n10245 ;
  assign n10247 = ~n10239 & ~n10246 ;
  assign n10248 = ~n10238 & ~n10247 ;
  assign n10249 = ~n10237 & ~n10248 ;
  assign n10250 = ~n10236 & ~n10249 ;
  assign n10251 = ~n10235 & ~n10250 ;
  assign n10252 = ~n10234 & ~n10251 ;
  assign n10253 = ~n10233 & ~n10252 ;
  assign n10255 = n10232 & ~n10253 ;
  assign n10254 = ~n10232 & n10253 ;
  assign n10256 = n3929 & ~n10254 ;
  assign n10257 = ~n10255 & n10256 ;
  assign n10222 = ~n2043 & ~n3430 ;
  assign n10223 = ~n2050 & n2735 ;
  assign n10224 = ~n10222 & n10223 ;
  assign n10225 = ~n2016 & ~n3176 ;
  assign n10226 = ~n1984 & ~n10225 ;
  assign n10227 = ~n2051 & ~n10226 ;
  assign n10228 = ~n3430 & ~n10227 ;
  assign n10229 = \P2_addr_reg[6]/NET0131  & n10228 ;
  assign n10287 = ~n10224 & ~n10229 ;
  assign n10288 = ~n10257 & n10287 ;
  assign n10289 = ~n10286 & n10288 ;
  assign n10220 = ~n1984 & n3928 ;
  assign n10221 = ~\P2_addr_reg[6]/NET0131  & n10220 ;
  assign n10290 = \P1_state_reg[0]/NET0131  & ~n10221 ;
  assign n10291 = ~n10289 & n10290 ;
  assign n10292 = ~n9285 & ~n10291 ;
  assign n10332 = ~\P2_reg1_reg[12]/NET0131  & ~n2943 ;
  assign n10333 = ~\P2_reg1_reg[11]/NET0131  & ~n2916 ;
  assign n10334 = ~\P2_reg1_reg[10]/NET0131  & ~n2970 ;
  assign n10335 = ~n10333 & ~n10334 ;
  assign n10336 = ~\P2_reg1_reg[9]/NET0131  & ~n2995 ;
  assign n10337 = ~\P2_reg1_reg[8]/NET0131  & ~n2682 ;
  assign n10338 = ~n10259 & n10282 ;
  assign n10339 = ~\P2_reg1_reg[7]/NET0131  & ~n2709 ;
  assign n10340 = ~n10260 & ~n10339 ;
  assign n10341 = ~n10338 & n10340 ;
  assign n10342 = \P2_reg1_reg[7]/NET0131  & n2709 ;
  assign n10343 = \P2_reg1_reg[8]/NET0131  & n2682 ;
  assign n10344 = ~n10342 & ~n10343 ;
  assign n10345 = ~n10341 & n10344 ;
  assign n10346 = ~n10337 & ~n10345 ;
  assign n10347 = ~n10336 & n10346 ;
  assign n10348 = \P2_reg1_reg[9]/NET0131  & n2995 ;
  assign n10349 = \P2_reg1_reg[10]/NET0131  & n2970 ;
  assign n10350 = ~n10348 & ~n10349 ;
  assign n10351 = ~n10347 & n10350 ;
  assign n10352 = n10335 & ~n10351 ;
  assign n10353 = \P2_reg1_reg[12]/NET0131  & n2943 ;
  assign n10354 = \P2_reg1_reg[11]/NET0131  & n2916 ;
  assign n10355 = ~n10353 & ~n10354 ;
  assign n10356 = ~n10352 & n10355 ;
  assign n10357 = ~n10332 & ~n10356 ;
  assign n10358 = \P2_reg1_reg[13]/NET0131  & ~n3108 ;
  assign n10359 = ~\P2_reg1_reg[13]/NET0131  & n3108 ;
  assign n10360 = ~n10358 & ~n10359 ;
  assign n10362 = ~n10357 & ~n10360 ;
  assign n10361 = n10357 & n10360 ;
  assign n10363 = n10258 & ~n10361 ;
  assign n10364 = ~n10362 & n10363 ;
  assign n10299 = \P2_reg2_reg[13]/NET0131  & ~n3108 ;
  assign n10300 = ~\P2_reg2_reg[13]/NET0131  & n3108 ;
  assign n10301 = ~n10299 & ~n10300 ;
  assign n10302 = ~\P2_reg2_reg[12]/NET0131  & ~n2943 ;
  assign n10303 = ~\P2_reg2_reg[11]/NET0131  & ~n2916 ;
  assign n10304 = ~\P2_reg2_reg[10]/NET0131  & ~n2970 ;
  assign n10305 = ~n10303 & ~n10304 ;
  assign n10306 = ~\P2_reg2_reg[9]/NET0131  & ~n2995 ;
  assign n10307 = ~\P2_reg2_reg[8]/NET0131  & ~n2682 ;
  assign n10308 = ~n10230 & n10253 ;
  assign n10309 = ~\P2_reg2_reg[7]/NET0131  & ~n2709 ;
  assign n10310 = ~n10231 & ~n10309 ;
  assign n10311 = ~n10308 & n10310 ;
  assign n10312 = \P2_reg2_reg[7]/NET0131  & n2709 ;
  assign n10313 = \P2_reg2_reg[8]/NET0131  & n2682 ;
  assign n10314 = ~n10312 & ~n10313 ;
  assign n10315 = ~n10311 & n10314 ;
  assign n10316 = ~n10307 & ~n10315 ;
  assign n10317 = ~n10306 & n10316 ;
  assign n10318 = \P2_reg2_reg[9]/NET0131  & n2995 ;
  assign n10319 = \P2_reg2_reg[10]/NET0131  & n2970 ;
  assign n10320 = ~n10318 & ~n10319 ;
  assign n10321 = ~n10317 & n10320 ;
  assign n10322 = n10305 & ~n10321 ;
  assign n10323 = \P2_reg2_reg[11]/NET0131  & n2916 ;
  assign n10324 = \P2_reg2_reg[12]/NET0131  & n2943 ;
  assign n10325 = ~n10323 & ~n10324 ;
  assign n10326 = ~n10322 & n10325 ;
  assign n10327 = ~n10302 & ~n10326 ;
  assign n10329 = ~n10301 & ~n10327 ;
  assign n10328 = n10301 & n10327 ;
  assign n10330 = n3929 & ~n10328 ;
  assign n10331 = ~n10329 & n10330 ;
  assign n10294 = ~\P2_addr_reg[13]/NET0131  & ~n10226 ;
  assign n10295 = n10228 & ~n10294 ;
  assign n10296 = ~n2043 & n10294 ;
  assign n10297 = ~n2050 & ~n3108 ;
  assign n10298 = ~n10296 & n10297 ;
  assign n10365 = ~n10295 & ~n10298 ;
  assign n10366 = ~n10331 & n10365 ;
  assign n10367 = ~n10364 & n10366 ;
  assign n10293 = ~\P2_addr_reg[13]/NET0131  & n10220 ;
  assign n10368 = \P1_state_reg[0]/NET0131  & ~n10293 ;
  assign n10369 = ~n10367 & n10368 ;
  assign n10370 = ~n7141 & ~n10369 ;
  assign n10382 = ~\P2_IR_reg[0]/NET0131  & ~\P2_reg2_reg[0]/NET0131  ;
  assign n10383 = ~n10243 & ~n10382 ;
  assign n10384 = n3929 & n10383 ;
  assign n10377 = n2043 & ~n2050 ;
  assign n10378 = \P2_IR_reg[0]/NET0131  & n10377 ;
  assign n10379 = ~\P2_IR_reg[0]/NET0131  & ~\P2_reg1_reg[0]/NET0131  ;
  assign n10380 = ~n10272 & ~n10379 ;
  assign n10381 = n10258 & n10380 ;
  assign n10385 = ~n10378 & ~n10381 ;
  assign n10386 = ~n10384 & n10385 ;
  assign n10387 = ~n10220 & ~n10386 ;
  assign n10371 = n2051 & ~n3430 ;
  assign n10372 = \P2_addr_reg[0]/NET0131  & n10371 ;
  assign n10373 = n2016 & n2829 ;
  assign n10374 = \P2_addr_reg[0]/NET0131  & n3928 ;
  assign n10375 = ~n10373 & ~n10374 ;
  assign n10376 = ~n1984 & ~n10375 ;
  assign n10388 = ~n10372 & ~n10376 ;
  assign n10389 = ~n10387 & n10388 ;
  assign n10390 = \P1_state_reg[0]/NET0131  & ~n10389 ;
  assign n10391 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[0]/NET0131  ;
  assign n10392 = ~n10390 & ~n10391 ;
  assign n10409 = ~n10304 & ~n10319 ;
  assign n10410 = ~n10311 & ~n10312 ;
  assign n10411 = ~n10307 & ~n10410 ;
  assign n10412 = ~n10313 & ~n10318 ;
  assign n10413 = ~n10411 & n10412 ;
  assign n10414 = ~n10306 & ~n10413 ;
  assign n10416 = n10409 & n10414 ;
  assign n10415 = ~n10409 & ~n10414 ;
  assign n10417 = n3929 & ~n10415 ;
  assign n10418 = ~n10416 & n10417 ;
  assign n10396 = ~n10334 & ~n10349 ;
  assign n10397 = ~n10341 & ~n10342 ;
  assign n10398 = ~n10337 & ~n10397 ;
  assign n10399 = ~n10343 & ~n10348 ;
  assign n10400 = ~n10398 & n10399 ;
  assign n10401 = ~n10336 & ~n10400 ;
  assign n10403 = n10396 & n10401 ;
  assign n10402 = ~n10396 & ~n10401 ;
  assign n10404 = n10258 & ~n10402 ;
  assign n10405 = ~n10403 & n10404 ;
  assign n10394 = ~\P2_addr_reg[10]/NET0131  & ~n10226 ;
  assign n10395 = n10228 & ~n10394 ;
  assign n10406 = ~n2043 & n10394 ;
  assign n10407 = ~n2050 & n2970 ;
  assign n10408 = ~n10406 & n10407 ;
  assign n10419 = ~n10395 & ~n10408 ;
  assign n10420 = ~n10405 & n10419 ;
  assign n10421 = ~n10418 & n10420 ;
  assign n10393 = ~\P2_addr_reg[10]/NET0131  & n10220 ;
  assign n10422 = \P1_state_reg[0]/NET0131  & ~n10393 ;
  assign n10423 = ~n10421 & n10422 ;
  assign n10424 = ~n7097 & ~n10423 ;
  assign n10437 = n10352 & ~n10354 ;
  assign n10434 = ~n10333 & ~n10354 ;
  assign n10435 = ~n10334 & ~n10351 ;
  assign n10436 = ~n10434 & ~n10435 ;
  assign n10438 = n10258 & ~n10436 ;
  assign n10439 = ~n10437 & n10438 ;
  assign n10431 = n10322 & ~n10323 ;
  assign n10428 = ~n10303 & ~n10323 ;
  assign n10429 = ~n10304 & ~n10321 ;
  assign n10430 = ~n10428 & ~n10429 ;
  assign n10432 = n3929 & ~n10430 ;
  assign n10433 = ~n10431 & n10432 ;
  assign n10426 = ~\P2_addr_reg[11]/NET0131  & ~n10226 ;
  assign n10427 = n10228 & ~n10426 ;
  assign n10440 = ~n2043 & n10426 ;
  assign n10441 = ~n2050 & n2916 ;
  assign n10442 = ~n10440 & n10441 ;
  assign n10443 = ~n10427 & ~n10442 ;
  assign n10444 = ~n10433 & n10443 ;
  assign n10445 = ~n10439 & n10444 ;
  assign n10425 = ~\P2_addr_reg[11]/NET0131  & n10220 ;
  assign n10446 = \P1_state_reg[0]/NET0131  & ~n10425 ;
  assign n10447 = ~n10445 & n10446 ;
  assign n10448 = ~n8022 & ~n10447 ;
  assign n10463 = ~n10332 & ~n10353 ;
  assign n10464 = ~n10349 & ~n10401 ;
  assign n10465 = n10335 & ~n10464 ;
  assign n10466 = ~n10354 & ~n10465 ;
  assign n10468 = ~n10463 & n10466 ;
  assign n10467 = n10463 & ~n10466 ;
  assign n10469 = n10258 & ~n10467 ;
  assign n10470 = ~n10468 & n10469 ;
  assign n10455 = ~n10302 & ~n10324 ;
  assign n10456 = ~n10319 & ~n10414 ;
  assign n10457 = n10305 & ~n10456 ;
  assign n10458 = ~n10323 & ~n10457 ;
  assign n10460 = ~n10455 & n10458 ;
  assign n10459 = n10455 & ~n10458 ;
  assign n10461 = n3929 & ~n10459 ;
  assign n10462 = ~n10460 & n10461 ;
  assign n10450 = ~\P2_addr_reg[12]/NET0131  & ~n10226 ;
  assign n10451 = n10228 & ~n10450 ;
  assign n10452 = ~n2043 & n10450 ;
  assign n10453 = ~n2050 & n2943 ;
  assign n10454 = ~n10452 & n10453 ;
  assign n10471 = ~n10451 & ~n10454 ;
  assign n10472 = ~n10462 & n10471 ;
  assign n10473 = ~n10470 & n10472 ;
  assign n10449 = ~\P2_addr_reg[12]/NET0131  & n10220 ;
  assign n10474 = \P1_state_reg[0]/NET0131  & ~n10449 ;
  assign n10475 = ~n10473 & n10474 ;
  assign n10476 = ~n6383 & ~n10475 ;
  assign n10494 = \P2_reg1_reg[14]/NET0131  & n3085 ;
  assign n10495 = ~\P2_reg1_reg[14]/NET0131  & ~n3085 ;
  assign n10496 = ~n10494 & ~n10495 ;
  assign n10497 = ~n10332 & ~n10466 ;
  assign n10498 = ~n10353 & ~n10358 ;
  assign n10499 = ~n10497 & n10498 ;
  assign n10500 = ~n10359 & ~n10499 ;
  assign n10502 = n10496 & n10500 ;
  assign n10501 = ~n10496 & ~n10500 ;
  assign n10503 = n10258 & ~n10501 ;
  assign n10504 = ~n10502 & n10503 ;
  assign n10480 = \P2_reg2_reg[14]/NET0131  & n3085 ;
  assign n10481 = ~\P2_reg2_reg[14]/NET0131  & ~n3085 ;
  assign n10482 = ~n10480 & ~n10481 ;
  assign n10483 = ~n10302 & ~n10458 ;
  assign n10484 = ~n10299 & ~n10324 ;
  assign n10485 = ~n10483 & n10484 ;
  assign n10486 = ~n10300 & ~n10485 ;
  assign n10488 = n10482 & n10486 ;
  assign n10487 = ~n10482 & ~n10486 ;
  assign n10489 = n3929 & ~n10487 ;
  assign n10490 = ~n10488 & n10489 ;
  assign n10478 = ~\P2_addr_reg[14]/NET0131  & ~n10226 ;
  assign n10479 = n10228 & ~n10478 ;
  assign n10491 = ~n2043 & n10478 ;
  assign n10492 = ~n2050 & n3085 ;
  assign n10493 = ~n10491 & n10492 ;
  assign n10505 = ~n10479 & ~n10493 ;
  assign n10506 = ~n10490 & n10505 ;
  assign n10507 = ~n10504 & n10506 ;
  assign n10477 = ~\P2_addr_reg[14]/NET0131  & n10220 ;
  assign n10508 = \P1_state_reg[0]/NET0131  & ~n10477 ;
  assign n10509 = ~n10507 & n10508 ;
  assign n10510 = ~n8062 & ~n10509 ;
  assign n10528 = \P2_reg1_reg[15]/NET0131  & n3061 ;
  assign n10529 = ~\P2_reg1_reg[15]/NET0131  & ~n3061 ;
  assign n10530 = ~n10528 & ~n10529 ;
  assign n10531 = n10357 & ~n10359 ;
  assign n10532 = ~n10358 & ~n10494 ;
  assign n10533 = ~n10531 & n10532 ;
  assign n10534 = ~n10495 & ~n10533 ;
  assign n10536 = n10530 & n10534 ;
  assign n10535 = ~n10530 & ~n10534 ;
  assign n10537 = n10258 & ~n10535 ;
  assign n10538 = ~n10536 & n10537 ;
  assign n10514 = ~\P2_reg2_reg[15]/NET0131  & ~n3061 ;
  assign n10515 = \P2_reg2_reg[15]/NET0131  & n3061 ;
  assign n10516 = ~n10514 & ~n10515 ;
  assign n10517 = ~n10300 & n10327 ;
  assign n10518 = ~n10299 & ~n10480 ;
  assign n10519 = ~n10517 & n10518 ;
  assign n10520 = ~n10481 & ~n10519 ;
  assign n10522 = n10516 & n10520 ;
  assign n10521 = ~n10516 & ~n10520 ;
  assign n10523 = n3929 & ~n10521 ;
  assign n10524 = ~n10522 & n10523 ;
  assign n10512 = ~\P2_addr_reg[15]/NET0131  & ~n10226 ;
  assign n10513 = n10228 & ~n10512 ;
  assign n10525 = ~n2043 & n10512 ;
  assign n10526 = ~n2050 & n3061 ;
  assign n10527 = ~n10525 & n10526 ;
  assign n10539 = ~n10513 & ~n10527 ;
  assign n10540 = ~n10524 & n10539 ;
  assign n10541 = ~n10538 & n10540 ;
  assign n10511 = ~\P2_addr_reg[15]/NET0131  & n10220 ;
  assign n10542 = \P1_state_reg[0]/NET0131  & ~n10511 ;
  assign n10543 = ~n10541 & n10542 ;
  assign n10544 = ~n7185 & ~n10543 ;
  assign n10563 = \P2_reg2_reg[16]/NET0131  & n3026 ;
  assign n10564 = ~\P2_reg2_reg[16]/NET0131  & ~n3026 ;
  assign n10565 = ~n10563 & ~n10564 ;
  assign n10566 = ~n10481 & n10486 ;
  assign n10567 = ~n10480 & ~n10515 ;
  assign n10568 = ~n10566 & n10567 ;
  assign n10569 = ~n10514 & ~n10568 ;
  assign n10571 = ~n10565 & ~n10569 ;
  assign n10570 = n10565 & n10569 ;
  assign n10572 = n3929 & ~n10570 ;
  assign n10573 = ~n10571 & n10572 ;
  assign n10551 = \P2_reg1_reg[16]/NET0131  & n3026 ;
  assign n10552 = ~\P2_reg1_reg[16]/NET0131  & ~n3026 ;
  assign n10553 = ~n10551 & ~n10552 ;
  assign n10554 = ~n10495 & ~n10529 ;
  assign n10555 = n10500 & n10554 ;
  assign n10556 = ~n10494 & ~n10528 ;
  assign n10557 = ~n10529 & ~n10556 ;
  assign n10558 = ~n10555 & ~n10557 ;
  assign n10560 = ~n10553 & n10558 ;
  assign n10559 = n10553 & ~n10558 ;
  assign n10561 = n10258 & ~n10559 ;
  assign n10562 = ~n10560 & n10561 ;
  assign n10546 = ~\P2_addr_reg[16]/NET0131  & ~n10226 ;
  assign n10547 = n10228 & ~n10546 ;
  assign n10548 = ~n2043 & n10546 ;
  assign n10549 = ~n2050 & n3026 ;
  assign n10550 = ~n10548 & n10549 ;
  assign n10574 = ~n10547 & ~n10550 ;
  assign n10575 = ~n10562 & n10574 ;
  assign n10576 = ~n10573 & n10575 ;
  assign n10545 = ~\P2_addr_reg[16]/NET0131  & n10220 ;
  assign n10577 = \P1_state_reg[0]/NET0131  & ~n10545 ;
  assign n10578 = ~n10576 & n10577 ;
  assign n10579 = ~n6426 & ~n10578 ;
  assign n10583 = ~\P2_reg2_reg[17]/NET0131  & ~n2619 ;
  assign n10584 = \P2_reg2_reg[17]/NET0131  & n2619 ;
  assign n10585 = ~n10583 & ~n10584 ;
  assign n10586 = ~n10514 & n10520 ;
  assign n10587 = ~n10515 & ~n10563 ;
  assign n10588 = ~n10586 & n10587 ;
  assign n10589 = ~n10564 & ~n10588 ;
  assign n10591 = n10585 & n10589 ;
  assign n10590 = ~n10585 & ~n10589 ;
  assign n10592 = n3929 & ~n10590 ;
  assign n10593 = ~n10591 & n10592 ;
  assign n10597 = ~\P2_reg1_reg[17]/NET0131  & ~n2619 ;
  assign n10598 = \P2_reg1_reg[17]/NET0131  & n2619 ;
  assign n10599 = ~n10597 & ~n10598 ;
  assign n10600 = ~n10533 & n10554 ;
  assign n10601 = ~n10528 & ~n10551 ;
  assign n10602 = ~n10600 & n10601 ;
  assign n10603 = ~n10552 & ~n10602 ;
  assign n10605 = n10599 & n10603 ;
  assign n10604 = ~n10599 & ~n10603 ;
  assign n10606 = n10258 & ~n10604 ;
  assign n10607 = ~n10605 & n10606 ;
  assign n10581 = ~\P2_addr_reg[17]/NET0131  & ~n10226 ;
  assign n10582 = n10228 & ~n10581 ;
  assign n10594 = ~n2043 & n10581 ;
  assign n10595 = ~n2050 & n2619 ;
  assign n10596 = ~n10594 & n10595 ;
  assign n10608 = ~n10582 & ~n10596 ;
  assign n10609 = ~n10607 & n10608 ;
  assign n10610 = ~n10593 & n10609 ;
  assign n10580 = ~\P2_addr_reg[17]/NET0131  & n10220 ;
  assign n10611 = \P1_state_reg[0]/NET0131  & ~n10580 ;
  assign n10612 = ~n10610 & n10611 ;
  assign n10613 = ~n5862 & ~n10612 ;
  assign n10625 = ~n10241 & ~n10242 ;
  assign n10626 = ~n10243 & ~n10625 ;
  assign n10627 = n10243 & n10625 ;
  assign n10628 = ~n10626 & ~n10627 ;
  assign n10629 = n3929 & n10628 ;
  assign n10619 = ~n2812 & n10377 ;
  assign n10620 = ~n10270 & ~n10271 ;
  assign n10621 = n10272 & n10620 ;
  assign n10622 = ~n10272 & ~n10620 ;
  assign n10623 = ~n10621 & ~n10622 ;
  assign n10624 = n10258 & n10623 ;
  assign n10630 = ~n10619 & ~n10624 ;
  assign n10631 = ~n10629 & n10630 ;
  assign n10632 = ~n10220 & ~n10631 ;
  assign n10614 = \P2_addr_reg[1]/NET0131  & n10371 ;
  assign n10615 = n2016 & n2813 ;
  assign n10616 = \P2_addr_reg[1]/NET0131  & n3928 ;
  assign n10617 = ~n10615 & ~n10616 ;
  assign n10618 = ~n1984 & ~n10617 ;
  assign n10633 = ~n10614 & ~n10618 ;
  assign n10634 = ~n10632 & n10633 ;
  assign n10635 = \P1_state_reg[0]/NET0131  & ~n10634 ;
  assign n10636 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[1]/NET0131  ;
  assign n10637 = ~n10635 & ~n10636 ;
  assign n10649 = ~n10239 & ~n10240 ;
  assign n10650 = n10245 & ~n10649 ;
  assign n10651 = ~n10245 & n10649 ;
  assign n10652 = ~n10650 & ~n10651 ;
  assign n10653 = n3929 & n10652 ;
  assign n10643 = n2789 & n10377 ;
  assign n10644 = ~n10268 & ~n10269 ;
  assign n10645 = ~n10274 & n10644 ;
  assign n10646 = n10274 & ~n10644 ;
  assign n10647 = ~n10645 & ~n10646 ;
  assign n10648 = n10258 & n10647 ;
  assign n10654 = ~n10643 & ~n10648 ;
  assign n10655 = ~n10653 & n10654 ;
  assign n10656 = ~n10220 & ~n10655 ;
  assign n10638 = \P2_addr_reg[2]/NET0131  & n10371 ;
  assign n10639 = n2016 & n2790 ;
  assign n10640 = \P2_addr_reg[2]/NET0131  & n3928 ;
  assign n10641 = ~n10639 & ~n10640 ;
  assign n10642 = ~n1984 & ~n10641 ;
  assign n10657 = ~n10638 & ~n10642 ;
  assign n10658 = ~n10656 & n10657 ;
  assign n10659 = \P1_state_reg[0]/NET0131  & ~n10658 ;
  assign n10660 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[2]/NET0131  ;
  assign n10661 = ~n10659 & ~n10660 ;
  assign n10669 = ~n10237 & ~n10238 ;
  assign n10670 = n10247 & ~n10669 ;
  assign n10671 = ~n10247 & n10669 ;
  assign n10672 = ~n10670 & ~n10671 ;
  assign n10673 = n3929 & n10672 ;
  assign n10663 = n2870 & n10377 ;
  assign n10664 = ~n10266 & ~n10267 ;
  assign n10665 = ~n10276 & n10664 ;
  assign n10666 = n10276 & ~n10664 ;
  assign n10667 = ~n10665 & ~n10666 ;
  assign n10668 = n10258 & n10667 ;
  assign n10674 = ~n10663 & ~n10668 ;
  assign n10675 = ~n10673 & n10674 ;
  assign n10682 = ~n3928 & ~n10675 ;
  assign n10679 = ~n2016 & n2051 ;
  assign n10680 = ~n3928 & ~n10679 ;
  assign n10681 = \P2_addr_reg[3]/NET0131  & ~n10680 ;
  assign n10678 = n2016 & n2871 ;
  assign n10683 = ~n1984 & ~n10678 ;
  assign n10684 = ~n10681 & n10683 ;
  assign n10685 = ~n10682 & n10684 ;
  assign n10662 = \P2_addr_reg[3]/NET0131  & n2051 ;
  assign n10676 = n1984 & ~n10662 ;
  assign n10677 = n10675 & n10676 ;
  assign n10686 = \P1_state_reg[0]/NET0131  & ~n10677 ;
  assign n10687 = ~n10685 & n10686 ;
  assign n10688 = ~n9244 & ~n10687 ;
  assign n10696 = ~n10235 & ~n10236 ;
  assign n10698 = ~n10249 & n10696 ;
  assign n10697 = n10249 & ~n10696 ;
  assign n10699 = n3929 & ~n10697 ;
  assign n10700 = ~n10698 & n10699 ;
  assign n10690 = ~n2847 & n10377 ;
  assign n10691 = ~n10264 & ~n10265 ;
  assign n10693 = ~n10278 & n10691 ;
  assign n10692 = n10278 & ~n10691 ;
  assign n10694 = n10258 & ~n10692 ;
  assign n10695 = ~n10693 & n10694 ;
  assign n10701 = ~n10690 & ~n10695 ;
  assign n10702 = ~n10700 & n10701 ;
  assign n10703 = ~n3928 & ~n10702 ;
  assign n10704 = \P2_addr_reg[4]/NET0131  & ~n10680 ;
  assign n10689 = n2016 & n2848 ;
  assign n10705 = ~n1984 & ~n10689 ;
  assign n10706 = ~n10704 & n10705 ;
  assign n10707 = ~n10703 & n10706 ;
  assign n10708 = \P2_addr_reg[4]/NET0131  & n2051 ;
  assign n10709 = n1984 & ~n10708 ;
  assign n10710 = n10702 & n10709 ;
  assign n10711 = \P1_state_reg[0]/NET0131  & ~n10710 ;
  assign n10712 = ~n10707 & n10711 ;
  assign n10713 = ~n8763 & ~n10712 ;
  assign n10715 = ~n10262 & ~n10263 ;
  assign n10717 = ~n10280 & n10715 ;
  assign n10716 = n10280 & ~n10715 ;
  assign n10718 = n10258 & ~n10716 ;
  assign n10719 = ~n10717 & n10718 ;
  assign n10720 = ~\P2_addr_reg[5]/NET0131  & ~n10226 ;
  assign n10721 = n10228 & ~n10720 ;
  assign n10730 = ~n10719 & ~n10721 ;
  assign n10722 = ~n10233 & ~n10234 ;
  assign n10724 = ~n10251 & n10722 ;
  assign n10723 = n10251 & ~n10722 ;
  assign n10725 = n3929 & ~n10723 ;
  assign n10726 = ~n10724 & n10725 ;
  assign n10727 = ~n2043 & n10720 ;
  assign n10728 = ~n2050 & ~n2758 ;
  assign n10729 = ~n10727 & n10728 ;
  assign n10731 = ~n10726 & ~n10729 ;
  assign n10732 = n10730 & n10731 ;
  assign n10714 = ~\P2_addr_reg[5]/NET0131  & n10220 ;
  assign n10733 = \P1_state_reg[0]/NET0131  & ~n10714 ;
  assign n10734 = ~n10732 & n10733 ;
  assign n10735 = ~n8800 & ~n10734 ;
  assign n10745 = ~n10339 & ~n10342 ;
  assign n10746 = ~n10260 & ~n10338 ;
  assign n10748 = n10745 & n10746 ;
  assign n10747 = ~n10745 & ~n10746 ;
  assign n10749 = n10258 & ~n10747 ;
  assign n10750 = ~n10748 & n10749 ;
  assign n10739 = ~n10309 & ~n10312 ;
  assign n10740 = ~n10231 & ~n10308 ;
  assign n10742 = n10739 & n10740 ;
  assign n10741 = ~n10739 & ~n10740 ;
  assign n10743 = n3929 & ~n10741 ;
  assign n10744 = ~n10742 & n10743 ;
  assign n10737 = ~\P2_addr_reg[7]/NET0131  & ~n10226 ;
  assign n10738 = n10228 & ~n10737 ;
  assign n10751 = ~n2043 & n10737 ;
  assign n10752 = ~n2050 & n2709 ;
  assign n10753 = ~n10751 & n10752 ;
  assign n10754 = ~n10738 & ~n10753 ;
  assign n10755 = ~n10744 & n10754 ;
  assign n10756 = ~n10750 & n10755 ;
  assign n10736 = ~\P2_addr_reg[7]/NET0131  & n10220 ;
  assign n10757 = \P1_state_reg[0]/NET0131  & ~n10736 ;
  assign n10758 = ~n10756 & n10757 ;
  assign n10759 = ~n8841 & ~n10758 ;
  assign n10771 = ~n10307 & ~n10313 ;
  assign n10773 = ~n10410 & n10771 ;
  assign n10772 = n10410 & ~n10771 ;
  assign n10774 = n3929 & ~n10772 ;
  assign n10775 = ~n10773 & n10774 ;
  assign n10766 = ~n10337 & ~n10343 ;
  assign n10768 = ~n10397 & n10766 ;
  assign n10767 = n10397 & ~n10766 ;
  assign n10769 = n10258 & ~n10767 ;
  assign n10770 = ~n10768 & n10769 ;
  assign n10761 = ~\P2_addr_reg[8]/NET0131  & ~n10226 ;
  assign n10762 = n10228 & ~n10761 ;
  assign n10763 = ~n2043 & n10761 ;
  assign n10764 = ~n2050 & n2682 ;
  assign n10765 = ~n10763 & n10764 ;
  assign n10776 = ~n10762 & ~n10765 ;
  assign n10777 = ~n10770 & n10776 ;
  assign n10778 = ~n10775 & n10777 ;
  assign n10760 = ~\P2_addr_reg[8]/NET0131  & n10220 ;
  assign n10779 = \P1_state_reg[0]/NET0131  & ~n10760 ;
  assign n10780 = ~n10778 & n10779 ;
  assign n10781 = ~n8143 & ~n10780 ;
  assign n10793 = ~n10336 & ~n10348 ;
  assign n10795 = ~n10346 & ~n10793 ;
  assign n10794 = n10346 & n10793 ;
  assign n10796 = n10258 & ~n10794 ;
  assign n10797 = ~n10795 & n10796 ;
  assign n10788 = ~n10306 & ~n10318 ;
  assign n10790 = ~n10316 & ~n10788 ;
  assign n10789 = n10316 & n10788 ;
  assign n10791 = n3929 & ~n10789 ;
  assign n10792 = ~n10790 & n10791 ;
  assign n10783 = ~\P2_addr_reg[9]/NET0131  & ~n10226 ;
  assign n10784 = n10228 & ~n10783 ;
  assign n10785 = ~n2043 & n10783 ;
  assign n10786 = ~n2050 & n2995 ;
  assign n10787 = ~n10785 & n10786 ;
  assign n10798 = ~n10784 & ~n10787 ;
  assign n10799 = ~n10792 & n10798 ;
  assign n10800 = ~n10797 & n10799 ;
  assign n10782 = ~\P2_addr_reg[9]/NET0131  & n10220 ;
  assign n10801 = \P1_state_reg[0]/NET0131  & ~n10782 ;
  assign n10802 = ~n10800 & n10801 ;
  assign n10803 = ~n7226 & ~n10802 ;
  assign n10820 = \P2_reg2_reg[18]/NET0131  & n2647 ;
  assign n10821 = ~\P2_reg2_reg[18]/NET0131  & ~n2647 ;
  assign n10822 = ~n10820 & ~n10821 ;
  assign n10823 = ~n10564 & n10569 ;
  assign n10824 = ~n10563 & ~n10584 ;
  assign n10825 = ~n10823 & n10824 ;
  assign n10826 = ~n10583 & ~n10825 ;
  assign n10828 = n10822 & n10826 ;
  assign n10827 = ~n10822 & ~n10826 ;
  assign n10829 = n3929 & ~n10827 ;
  assign n10830 = ~n10828 & n10829 ;
  assign n10804 = \P2_reg1_reg[18]/NET0131  & n2647 ;
  assign n10805 = ~\P2_reg1_reg[18]/NET0131  & ~n2647 ;
  assign n10806 = ~n10804 & ~n10805 ;
  assign n10807 = ~n10552 & ~n10558 ;
  assign n10808 = ~n10551 & ~n10598 ;
  assign n10809 = ~n10807 & n10808 ;
  assign n10810 = ~n10597 & ~n10809 ;
  assign n10812 = n10806 & n10810 ;
  assign n10811 = ~n10806 & ~n10810 ;
  assign n10813 = n10258 & ~n10811 ;
  assign n10814 = ~n10812 & n10813 ;
  assign n10815 = ~\P2_addr_reg[18]/NET0131  & ~n10226 ;
  assign n10816 = n10228 & ~n10815 ;
  assign n10817 = ~n2043 & n10815 ;
  assign n10818 = ~n2050 & n2647 ;
  assign n10819 = ~n10817 & n10818 ;
  assign n10831 = ~n10816 & ~n10819 ;
  assign n10832 = ~n10814 & n10831 ;
  assign n10833 = ~n10830 & n10832 ;
  assign n10834 = ~\P2_addr_reg[18]/NET0131  & n10220 ;
  assign n10835 = \P1_state_reg[0]/NET0131  & ~n10834 ;
  assign n10836 = ~n10833 & n10835 ;
  assign n10837 = ~n5904 & ~n10836 ;
  assign n10854 = ~n10598 & ~n10603 ;
  assign n10855 = ~n10597 & ~n10805 ;
  assign n10856 = ~n10854 & n10855 ;
  assign n10857 = ~n10804 & ~n10856 ;
  assign n10858 = \P2_reg1_reg[19]/NET0131  & ~n10857 ;
  assign n10859 = ~\P2_reg1_reg[19]/NET0131  & n10857 ;
  assign n10860 = ~n10858 & ~n10859 ;
  assign n10862 = ~n2592 & ~n10860 ;
  assign n10861 = n2592 & n10860 ;
  assign n10863 = n10258 & ~n10861 ;
  assign n10864 = ~n10862 & n10863 ;
  assign n10838 = ~n10584 & ~n10589 ;
  assign n10839 = ~n10583 & ~n10821 ;
  assign n10840 = ~n10838 & n10839 ;
  assign n10841 = ~n10820 & ~n10840 ;
  assign n10842 = ~\P2_reg2_reg[19]/NET0131  & ~n2592 ;
  assign n10843 = \P2_reg2_reg[19]/NET0131  & n2592 ;
  assign n10844 = ~n10842 & ~n10843 ;
  assign n10846 = n10841 & ~n10844 ;
  assign n10845 = ~n10841 & n10844 ;
  assign n10847 = n3929 & ~n10845 ;
  assign n10848 = ~n10846 & n10847 ;
  assign n10849 = ~\P2_addr_reg[19]/NET0131  & ~n10226 ;
  assign n10850 = n10228 & ~n10849 ;
  assign n10851 = ~n2043 & n10849 ;
  assign n10852 = ~n2050 & n2592 ;
  assign n10853 = ~n10851 & n10852 ;
  assign n10865 = ~n10850 & ~n10853 ;
  assign n10866 = ~n10848 & n10865 ;
  assign n10867 = ~n10864 & n10866 ;
  assign n10868 = ~\P2_addr_reg[19]/NET0131  & n10220 ;
  assign n10869 = \P1_state_reg[0]/NET0131  & ~n10868 ;
  assign n10870 = ~n10867 & n10869 ;
  assign n10871 = ~n5946 & ~n10870 ;
  assign n10872 = ~\P1_reg3_reg[2]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n10874 = ~\P1_IR_reg[0]/NET0131  & ~\P1_reg2_reg[0]/NET0131  ;
  assign n10875 = \P1_IR_reg[0]/NET0131  & \P1_reg2_reg[0]/NET0131  ;
  assign n10876 = ~n10874 & ~n10875 ;
  assign n10877 = n1936 & n10876 ;
  assign n10878 = n527 & n536 ;
  assign n10879 = \P1_IR_reg[0]/NET0131  & \P1_reg1_reg[0]/NET0131  ;
  assign n10880 = ~\P1_IR_reg[0]/NET0131  & ~\P1_reg1_reg[0]/NET0131  ;
  assign n10881 = ~n10879 & ~n10880 ;
  assign n10882 = n10878 & n10881 ;
  assign n10883 = ~n10877 & ~n10882 ;
  assign n10873 = \P1_IR_reg[0]/NET0131  & ~n536 ;
  assign n10884 = n1951 & ~n10873 ;
  assign n10885 = n10883 & n10884 ;
  assign n10886 = ~\P1_addr_reg[2]/NET0131  & n1897 ;
  assign n10887 = ~n1951 & n10886 ;
  assign n10888 = ~n10885 & ~n10887 ;
  assign n10889 = ~n1933 & ~n10888 ;
  assign n10904 = ~n1897 & ~n1951 ;
  assign n10905 = ~n1933 & ~n10904 ;
  assign n10890 = \P1_addr_reg[2]/NET0131  & n537 ;
  assign n10891 = ~n527 & ~n536 ;
  assign n10892 = n1356 & n10891 ;
  assign n10917 = ~n10890 & ~n10892 ;
  assign n10893 = \P1_reg1_reg[2]/NET0131  & n1356 ;
  assign n10894 = ~\P1_reg1_reg[2]/NET0131  & ~n1356 ;
  assign n10895 = ~n10893 & ~n10894 ;
  assign n10896 = ~\P1_reg1_reg[1]/NET0131  & n1371 ;
  assign n10897 = \P1_reg1_reg[1]/NET0131  & ~n1371 ;
  assign n10898 = ~n10879 & ~n10897 ;
  assign n10899 = ~n10896 & ~n10898 ;
  assign n10900 = n10895 & n10899 ;
  assign n10901 = ~n10895 & ~n10899 ;
  assign n10902 = ~n10900 & ~n10901 ;
  assign n10903 = n10878 & n10902 ;
  assign n10906 = \P1_reg2_reg[2]/NET0131  & n1356 ;
  assign n10907 = ~\P1_reg2_reg[2]/NET0131  & ~n1356 ;
  assign n10908 = ~n10906 & ~n10907 ;
  assign n10909 = ~\P1_reg2_reg[1]/NET0131  & n1371 ;
  assign n10910 = \P1_reg2_reg[1]/NET0131  & ~n1371 ;
  assign n10911 = ~n10875 & ~n10910 ;
  assign n10912 = ~n10909 & ~n10911 ;
  assign n10913 = ~n10908 & ~n10912 ;
  assign n10914 = n10908 & n10912 ;
  assign n10915 = ~n10913 & ~n10914 ;
  assign n10916 = n1936 & n10915 ;
  assign n10918 = ~n10903 & ~n10916 ;
  assign n10919 = n10917 & n10918 ;
  assign n10920 = ~n10905 & n10919 ;
  assign n10921 = ~n10889 & ~n10920 ;
  assign n10922 = \P1_state_reg[0]/NET0131  & ~n10921 ;
  assign n10923 = ~n10872 & ~n10922 ;
  assign n10924 = ~\P1_addr_reg[4]/NET0131  & n1897 ;
  assign n10925 = ~n1951 & n10924 ;
  assign n10926 = ~n10885 & ~n10925 ;
  assign n10927 = ~n1933 & ~n10926 ;
  assign n10928 = n1302 & n10891 ;
  assign n10929 = \P1_addr_reg[4]/NET0131  & n537 ;
  assign n10956 = ~n10928 & ~n10929 ;
  assign n10930 = \P1_reg2_reg[4]/NET0131  & n1302 ;
  assign n10931 = ~\P1_reg2_reg[4]/NET0131  & ~n1302 ;
  assign n10932 = ~n10930 & ~n10931 ;
  assign n10933 = ~\P1_reg2_reg[3]/NET0131  & ~n1334 ;
  assign n10934 = \P1_reg2_reg[3]/NET0131  & n1334 ;
  assign n10935 = ~n10906 & ~n10912 ;
  assign n10936 = ~n10907 & ~n10935 ;
  assign n10937 = ~n10934 & ~n10936 ;
  assign n10938 = ~n10933 & ~n10937 ;
  assign n10939 = n10932 & n10938 ;
  assign n10940 = ~n10932 & ~n10938 ;
  assign n10941 = ~n10939 & ~n10940 ;
  assign n10942 = n1936 & n10941 ;
  assign n10943 = \P1_reg1_reg[4]/NET0131  & n1302 ;
  assign n10944 = ~\P1_reg1_reg[4]/NET0131  & ~n1302 ;
  assign n10945 = ~n10943 & ~n10944 ;
  assign n10946 = ~\P1_reg1_reg[3]/NET0131  & ~n1334 ;
  assign n10947 = \P1_reg1_reg[3]/NET0131  & n1334 ;
  assign n10948 = ~n10893 & ~n10899 ;
  assign n10949 = ~n10894 & ~n10948 ;
  assign n10950 = ~n10947 & ~n10949 ;
  assign n10951 = ~n10946 & ~n10950 ;
  assign n10952 = ~n10945 & ~n10951 ;
  assign n10953 = n10945 & n10951 ;
  assign n10954 = ~n10952 & ~n10953 ;
  assign n10955 = n10878 & n10954 ;
  assign n10957 = ~n10942 & ~n10955 ;
  assign n10958 = n10956 & n10957 ;
  assign n10959 = ~n10905 & n10958 ;
  assign n10960 = ~n10927 & ~n10959 ;
  assign n10961 = \P1_state_reg[0]/NET0131  & ~n10960 ;
  assign n10962 = ~n8139 & ~n10961 ;
  assign n10963 = \P1_state_reg[0]/NET0131  & ~n10227 ;
  assign n10964 = ~n537 & ~n10905 ;
  assign n10965 = \P1_state_reg[0]/NET0131  & ~n10964 ;
  assign n10968 = \P1_state_reg[0]/NET0131  & ~n10905 ;
  assign n10992 = \P1_reg1_reg[8]/NET0131  & ~n1200 ;
  assign n10993 = ~\P1_reg1_reg[8]/NET0131  & n1200 ;
  assign n10994 = ~n10992 & ~n10993 ;
  assign n10995 = \P1_reg1_reg[7]/NET0131  & n1261 ;
  assign n10996 = ~\P1_reg1_reg[7]/NET0131  & ~n1261 ;
  assign n10997 = ~\P1_reg1_reg[6]/NET0131  & ~n1236 ;
  assign n10998 = \P1_reg1_reg[6]/NET0131  & n1236 ;
  assign n10999 = ~\P1_reg1_reg[5]/NET0131  & n1286 ;
  assign n11000 = \P1_reg1_reg[5]/NET0131  & ~n1286 ;
  assign n11001 = ~n10943 & ~n10951 ;
  assign n11002 = ~n10944 & ~n11001 ;
  assign n11003 = ~n11000 & ~n11002 ;
  assign n11004 = ~n10999 & ~n11003 ;
  assign n11005 = ~n10998 & ~n11004 ;
  assign n11006 = ~n10997 & ~n11005 ;
  assign n11007 = ~n10996 & n11006 ;
  assign n11008 = ~n10995 & ~n11007 ;
  assign n11010 = ~n10994 & n11008 ;
  assign n11009 = n10994 & ~n11008 ;
  assign n11011 = n10878 & ~n11009 ;
  assign n11012 = ~n11010 & n11011 ;
  assign n10971 = \P1_reg2_reg[8]/NET0131  & ~n1200 ;
  assign n10972 = ~\P1_reg2_reg[8]/NET0131  & n1200 ;
  assign n10973 = ~n10971 & ~n10972 ;
  assign n10974 = \P1_reg2_reg[7]/NET0131  & n1261 ;
  assign n10975 = ~\P1_reg2_reg[7]/NET0131  & ~n1261 ;
  assign n10976 = ~\P1_reg2_reg[6]/NET0131  & ~n1236 ;
  assign n10977 = \P1_reg2_reg[6]/NET0131  & n1236 ;
  assign n10978 = ~\P1_reg2_reg[5]/NET0131  & n1286 ;
  assign n10979 = \P1_reg2_reg[5]/NET0131  & ~n1286 ;
  assign n10980 = ~n10930 & ~n10938 ;
  assign n10981 = ~n10931 & ~n10980 ;
  assign n10982 = ~n10979 & ~n10981 ;
  assign n10983 = ~n10978 & ~n10982 ;
  assign n10984 = ~n10977 & ~n10983 ;
  assign n10985 = ~n10976 & ~n10984 ;
  assign n10986 = ~n10975 & n10985 ;
  assign n10987 = ~n10974 & ~n10986 ;
  assign n10989 = ~n10973 & n10987 ;
  assign n10988 = n10973 & ~n10987 ;
  assign n10990 = n1936 & ~n10988 ;
  assign n10991 = ~n10989 & n10990 ;
  assign n10969 = ~n1200 & n10891 ;
  assign n10970 = \P1_addr_reg[8]/NET0131  & n537 ;
  assign n11013 = ~n10969 & ~n10970 ;
  assign n11014 = ~n10991 & n11013 ;
  assign n11015 = ~n11012 & n11014 ;
  assign n11016 = n10968 & ~n11015 ;
  assign n10966 = n1897 & n6070 ;
  assign n10967 = \P1_addr_reg[8]/NET0131  & n10966 ;
  assign n11017 = ~n7268 & ~n10967 ;
  assign n11018 = ~n11016 & n11017 ;
  assign n11027 = ~n10976 & ~n10977 ;
  assign n11029 = n10983 & n11027 ;
  assign n11028 = ~n10983 & ~n11027 ;
  assign n11030 = n1936 & ~n11028 ;
  assign n11031 = ~n11029 & n11030 ;
  assign n11021 = ~n10997 & ~n10998 ;
  assign n11023 = n11004 & n11021 ;
  assign n11022 = ~n11004 & ~n11021 ;
  assign n11024 = n10878 & ~n11022 ;
  assign n11025 = ~n11023 & n11024 ;
  assign n11020 = \P1_addr_reg[6]/NET0131  & n537 ;
  assign n11026 = n1236 & n10891 ;
  assign n11032 = ~n11020 & ~n11026 ;
  assign n11033 = ~n11025 & n11032 ;
  assign n11034 = ~n11031 & n11033 ;
  assign n11035 = n10968 & ~n11034 ;
  assign n11019 = \P1_addr_reg[6]/NET0131  & n10966 ;
  assign n11036 = ~n8881 & ~n11019 ;
  assign n11037 = ~n11035 & n11036 ;
  assign n11047 = ~n10995 & n11007 ;
  assign n11045 = ~n10995 & ~n10996 ;
  assign n11046 = ~n11006 & ~n11045 ;
  assign n11048 = n10878 & ~n11046 ;
  assign n11049 = ~n11047 & n11048 ;
  assign n11042 = ~n10974 & n10986 ;
  assign n11040 = ~n10974 & ~n10975 ;
  assign n11041 = ~n10985 & ~n11040 ;
  assign n11043 = n1936 & ~n11041 ;
  assign n11044 = ~n11042 & n11043 ;
  assign n11038 = n1261 & n10891 ;
  assign n11039 = \P1_addr_reg[7]/NET0131  & n537 ;
  assign n11050 = ~n11038 & ~n11039 ;
  assign n11051 = ~n11044 & n11050 ;
  assign n11052 = ~n11049 & n11051 ;
  assign n11055 = ~n1897 & n11052 ;
  assign n11054 = ~\P1_addr_reg[7]/NET0131  & n1897 ;
  assign n11056 = n6070 & ~n11054 ;
  assign n11057 = ~n11055 & n11056 ;
  assign n11053 = n1934 & ~n11052 ;
  assign n11058 = ~n8920 & ~n11053 ;
  assign n11059 = ~n11057 & n11058 ;
  assign n11060 = ~\P1_addr_reg[3]/NET0131  & n1897 ;
  assign n11061 = n6070 & ~n11060 ;
  assign n11062 = ~n1934 & ~n11061 ;
  assign n11063 = ~n537 & ~n10966 ;
  assign n11064 = \P1_addr_reg[3]/NET0131  & ~n11063 ;
  assign n11071 = ~n10933 & ~n10934 ;
  assign n11072 = ~n10936 & ~n11071 ;
  assign n11073 = n10936 & n11071 ;
  assign n11074 = ~n11072 & ~n11073 ;
  assign n11075 = n1936 & n11074 ;
  assign n11065 = ~n10946 & ~n10947 ;
  assign n11066 = ~n10949 & ~n11065 ;
  assign n11067 = n10949 & n11065 ;
  assign n11068 = ~n11066 & ~n11067 ;
  assign n11069 = n10878 & n11068 ;
  assign n11070 = n1334 & n10891 ;
  assign n11076 = ~n11069 & ~n11070 ;
  assign n11077 = ~n11075 & n11076 ;
  assign n11078 = ~n11064 & n11077 ;
  assign n11079 = ~n11062 & ~n11078 ;
  assign n11080 = ~n8725 & ~n11079 ;
  assign n11081 = \P1_reg3_reg[0]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11082 = ~\P1_addr_reg[0]/NET0131  & n1897 ;
  assign n11083 = n6070 & ~n11082 ;
  assign n11084 = ~n1934 & ~n11083 ;
  assign n11086 = \P1_addr_reg[0]/NET0131  & ~n11063 ;
  assign n11085 = ~n527 & n10873 ;
  assign n11087 = n10883 & ~n11085 ;
  assign n11088 = ~n11086 & n11087 ;
  assign n11089 = ~n11084 & ~n11088 ;
  assign n11090 = ~n11081 & ~n11089 ;
  assign n11091 = ~\P1_addr_reg[10]/NET0131  & n1897 ;
  assign n11092 = n6070 & ~n11091 ;
  assign n11093 = ~n1934 & ~n11092 ;
  assign n11109 = \P1_reg1_reg[10]/NET0131  & ~n1149 ;
  assign n11110 = ~\P1_reg1_reg[10]/NET0131  & n1149 ;
  assign n11111 = ~n11109 & ~n11110 ;
  assign n11112 = ~\P1_reg1_reg[9]/NET0131  & ~n1176 ;
  assign n11113 = \P1_reg1_reg[9]/NET0131  & n1176 ;
  assign n11114 = ~n10992 & n11008 ;
  assign n11115 = ~n10993 & ~n11114 ;
  assign n11116 = ~n11113 & ~n11115 ;
  assign n11117 = ~n11112 & ~n11116 ;
  assign n11119 = ~n11111 & ~n11117 ;
  assign n11118 = n11111 & n11117 ;
  assign n11120 = n10878 & ~n11118 ;
  assign n11121 = ~n11119 & n11120 ;
  assign n11096 = \P1_reg2_reg[10]/NET0131  & ~n1149 ;
  assign n11097 = ~\P1_reg2_reg[10]/NET0131  & n1149 ;
  assign n11098 = ~n11096 & ~n11097 ;
  assign n11099 = ~\P1_reg2_reg[9]/NET0131  & ~n1176 ;
  assign n11100 = ~n10972 & ~n10987 ;
  assign n11101 = \P1_reg2_reg[9]/NET0131  & n1176 ;
  assign n11102 = ~n10971 & ~n11101 ;
  assign n11103 = ~n11100 & n11102 ;
  assign n11104 = ~n11099 & ~n11103 ;
  assign n11106 = ~n11098 & ~n11104 ;
  assign n11105 = n11098 & n11104 ;
  assign n11107 = n1936 & ~n11105 ;
  assign n11108 = ~n11106 & n11107 ;
  assign n11094 = \P1_addr_reg[10]/NET0131  & ~n11063 ;
  assign n11095 = ~n1149 & n10891 ;
  assign n11122 = ~n11094 & ~n11095 ;
  assign n11123 = ~n11108 & n11122 ;
  assign n11124 = ~n11121 & n11123 ;
  assign n11125 = ~n11093 & ~n11124 ;
  assign n11126 = ~n6973 & ~n11125 ;
  assign n11143 = ~\P1_reg2_reg[11]/NET0131  & ~n1126 ;
  assign n11144 = \P1_reg2_reg[11]/NET0131  & n1126 ;
  assign n11145 = ~n11143 & ~n11144 ;
  assign n11146 = ~n10971 & ~n10974 ;
  assign n11147 = ~n10986 & n11146 ;
  assign n11148 = ~n10972 & ~n11147 ;
  assign n11149 = ~n11097 & ~n11099 ;
  assign n11150 = n11148 & n11149 ;
  assign n11151 = ~n11097 & n11101 ;
  assign n11152 = ~n11096 & ~n11151 ;
  assign n11153 = ~n11150 & n11152 ;
  assign n11155 = ~n11145 & n11153 ;
  assign n11154 = n11145 & ~n11153 ;
  assign n11156 = n1936 & ~n11154 ;
  assign n11157 = ~n11155 & n11156 ;
  assign n11130 = ~\P1_reg1_reg[11]/NET0131  & ~n1126 ;
  assign n11131 = \P1_reg1_reg[11]/NET0131  & n1126 ;
  assign n11132 = ~n11130 & ~n11131 ;
  assign n11133 = ~n10993 & ~n11110 ;
  assign n11134 = ~n11112 & n11133 ;
  assign n11135 = ~n11114 & n11134 ;
  assign n11136 = ~n11110 & n11113 ;
  assign n11137 = ~n11109 & ~n11136 ;
  assign n11138 = ~n11135 & n11137 ;
  assign n11140 = ~n11132 & n11138 ;
  assign n11139 = n11132 & ~n11138 ;
  assign n11141 = n10878 & ~n11139 ;
  assign n11142 = ~n11140 & n11141 ;
  assign n11128 = \P1_addr_reg[11]/NET0131  & n537 ;
  assign n11129 = n1126 & n10891 ;
  assign n11158 = ~n11128 & ~n11129 ;
  assign n11159 = ~n11142 & n11158 ;
  assign n11160 = ~n11157 & n11159 ;
  assign n11161 = n10968 & ~n11160 ;
  assign n11127 = \P1_addr_reg[11]/NET0131  & n10966 ;
  assign n11162 = ~n6931 & ~n11127 ;
  assign n11163 = ~n11161 & n11162 ;
  assign n11164 = ~\P1_addr_reg[12]/NET0131  & n1897 ;
  assign n11165 = n6070 & ~n11164 ;
  assign n11166 = ~n1934 & ~n11165 ;
  assign n11180 = \P1_reg1_reg[12]/NET0131  & n1092 ;
  assign n11181 = ~\P1_reg1_reg[12]/NET0131  & ~n1092 ;
  assign n11182 = ~n11180 & ~n11181 ;
  assign n11183 = ~n11110 & n11117 ;
  assign n11184 = ~n11109 & ~n11131 ;
  assign n11185 = ~n11183 & n11184 ;
  assign n11186 = ~n11130 & ~n11185 ;
  assign n11188 = ~n11182 & ~n11186 ;
  assign n11187 = n11182 & n11186 ;
  assign n11189 = n10878 & ~n11187 ;
  assign n11190 = ~n11188 & n11189 ;
  assign n11169 = \P1_reg2_reg[12]/NET0131  & n1092 ;
  assign n11170 = ~\P1_reg2_reg[12]/NET0131  & ~n1092 ;
  assign n11171 = ~n11169 & ~n11170 ;
  assign n11172 = ~n11097 & n11104 ;
  assign n11173 = ~n11096 & ~n11144 ;
  assign n11174 = ~n11172 & n11173 ;
  assign n11175 = ~n11143 & ~n11174 ;
  assign n11177 = ~n11171 & ~n11175 ;
  assign n11176 = n11171 & n11175 ;
  assign n11178 = n1936 & ~n11176 ;
  assign n11179 = ~n11177 & n11178 ;
  assign n11167 = n1092 & n10891 ;
  assign n11168 = \P1_addr_reg[12]/NET0131  & ~n11063 ;
  assign n11191 = ~n11167 & ~n11168 ;
  assign n11192 = ~n11179 & n11191 ;
  assign n11193 = ~n11190 & n11192 ;
  assign n11194 = ~n11166 & ~n11193 ;
  assign n11195 = ~n5734 & ~n11194 ;
  assign n11197 = ~\P1_addr_reg[13]/NET0131  & n1897 ;
  assign n11198 = n6070 & ~n11197 ;
  assign n11199 = ~n1934 & ~n11198 ;
  assign n11213 = \P1_reg2_reg[13]/NET0131  & n1062 ;
  assign n11214 = ~\P1_reg2_reg[13]/NET0131  & ~n1062 ;
  assign n11215 = ~n11213 & ~n11214 ;
  assign n11216 = ~n11143 & ~n11153 ;
  assign n11217 = ~n11144 & ~n11169 ;
  assign n11218 = ~n11216 & n11217 ;
  assign n11219 = ~n11170 & ~n11218 ;
  assign n11221 = n11215 & n11219 ;
  assign n11220 = ~n11215 & ~n11219 ;
  assign n11222 = n1936 & ~n11220 ;
  assign n11223 = ~n11221 & n11222 ;
  assign n11202 = ~n11130 & ~n11138 ;
  assign n11203 = ~n11131 & ~n11180 ;
  assign n11204 = ~n11202 & n11203 ;
  assign n11205 = ~n11181 & ~n11204 ;
  assign n11206 = \P1_reg1_reg[13]/NET0131  & n1062 ;
  assign n11207 = ~\P1_reg1_reg[13]/NET0131  & ~n1062 ;
  assign n11208 = ~n11206 & ~n11207 ;
  assign n11210 = n11205 & n11208 ;
  assign n11209 = ~n11205 & ~n11208 ;
  assign n11211 = n10878 & ~n11209 ;
  assign n11212 = ~n11210 & n11211 ;
  assign n11200 = n1062 & n10891 ;
  assign n11201 = \P1_addr_reg[13]/NET0131  & n537 ;
  assign n11224 = ~n11200 & ~n11201 ;
  assign n11225 = ~n11212 & n11224 ;
  assign n11226 = ~n11223 & n11225 ;
  assign n11227 = ~n11199 & ~n11226 ;
  assign n11196 = \P1_addr_reg[13]/NET0131  & n10966 ;
  assign n11228 = ~n8019 & ~n11196 ;
  assign n11229 = ~n11227 & n11228 ;
  assign n11230 = ~\P1_addr_reg[14]/NET0131  & n1897 ;
  assign n11231 = n6070 & ~n11230 ;
  assign n11232 = ~n1934 & ~n11231 ;
  assign n11246 = \P1_reg1_reg[14]/NET0131  & ~n1038 ;
  assign n11247 = ~\P1_reg1_reg[14]/NET0131  & n1038 ;
  assign n11248 = ~n11246 & ~n11247 ;
  assign n11249 = ~n11181 & n11186 ;
  assign n11250 = ~n11180 & ~n11206 ;
  assign n11251 = ~n11249 & n11250 ;
  assign n11252 = ~n11207 & ~n11251 ;
  assign n11254 = ~n11248 & ~n11252 ;
  assign n11253 = n11248 & n11252 ;
  assign n11255 = n10878 & ~n11253 ;
  assign n11256 = ~n11254 & n11255 ;
  assign n11235 = \P1_reg2_reg[14]/NET0131  & ~n1038 ;
  assign n11236 = ~\P1_reg2_reg[14]/NET0131  & n1038 ;
  assign n11237 = ~n11235 & ~n11236 ;
  assign n11238 = ~n11170 & n11175 ;
  assign n11239 = ~n11169 & ~n11213 ;
  assign n11240 = ~n11238 & n11239 ;
  assign n11241 = ~n11214 & ~n11240 ;
  assign n11243 = ~n11237 & ~n11241 ;
  assign n11242 = n11237 & n11241 ;
  assign n11244 = n1936 & ~n11242 ;
  assign n11245 = ~n11243 & n11244 ;
  assign n11233 = ~n1038 & n10891 ;
  assign n11234 = \P1_addr_reg[14]/NET0131  & ~n11063 ;
  assign n11257 = ~n11233 & ~n11234 ;
  assign n11258 = ~n11245 & n11257 ;
  assign n11259 = ~n11256 & n11258 ;
  assign n11260 = ~n11232 & ~n11259 ;
  assign n11261 = ~n7015 & ~n11260 ;
  assign n11263 = ~\P1_addr_reg[16]/NET0131  & n1897 ;
  assign n11264 = n6070 & ~n11263 ;
  assign n11265 = ~n1934 & ~n11264 ;
  assign n11267 = \P1_reg1_reg[16]/NET0131  & n827 ;
  assign n11268 = ~\P1_reg1_reg[16]/NET0131  & ~n827 ;
  assign n11269 = ~n11267 & ~n11268 ;
  assign n11270 = ~\P1_reg1_reg[15]/NET0131  & ~n1013 ;
  assign n11271 = ~n11247 & n11252 ;
  assign n11272 = \P1_reg1_reg[15]/NET0131  & n1013 ;
  assign n11273 = ~n11246 & ~n11272 ;
  assign n11274 = ~n11271 & n11273 ;
  assign n11275 = ~n11270 & ~n11274 ;
  assign n11277 = n11269 & n11275 ;
  assign n11276 = ~n11269 & ~n11275 ;
  assign n11278 = n10878 & ~n11276 ;
  assign n11279 = ~n11277 & n11278 ;
  assign n11281 = \P1_reg2_reg[16]/NET0131  & n827 ;
  assign n11282 = ~\P1_reg2_reg[16]/NET0131  & ~n827 ;
  assign n11283 = ~n11281 & ~n11282 ;
  assign n11284 = ~\P1_reg2_reg[15]/NET0131  & ~n1013 ;
  assign n11285 = ~n11236 & n11241 ;
  assign n11286 = \P1_reg2_reg[15]/NET0131  & n1013 ;
  assign n11287 = ~n11235 & ~n11286 ;
  assign n11288 = ~n11285 & n11287 ;
  assign n11289 = ~n11284 & ~n11288 ;
  assign n11291 = n11283 & n11289 ;
  assign n11290 = ~n11283 & ~n11289 ;
  assign n11292 = n1936 & ~n11290 ;
  assign n11293 = ~n11291 & n11292 ;
  assign n11266 = \P1_addr_reg[16]/NET0131  & n537 ;
  assign n11280 = n827 & n10891 ;
  assign n11294 = ~n11266 & ~n11280 ;
  assign n11295 = ~n11293 & n11294 ;
  assign n11296 = ~n11279 & n11295 ;
  assign n11297 = ~n11265 & ~n11296 ;
  assign n11262 = \P1_addr_reg[16]/NET0131  & n10966 ;
  assign n11298 = ~n4829 & ~n11262 ;
  assign n11299 = ~n11297 & n11298 ;
  assign n11300 = ~\P1_addr_reg[17]/NET0131  & n1897 ;
  assign n11301 = n6070 & ~n11300 ;
  assign n11302 = ~n1934 & ~n11301 ;
  assign n11304 = \P1_reg1_reg[17]/NET0131  & n783 ;
  assign n11305 = ~\P1_reg1_reg[17]/NET0131  & ~n783 ;
  assign n11306 = ~n11304 & ~n11305 ;
  assign n11307 = n11205 & ~n11207 ;
  assign n11308 = ~n11206 & ~n11246 ;
  assign n11309 = ~n11307 & n11308 ;
  assign n11310 = ~n11247 & ~n11309 ;
  assign n11311 = ~n11270 & n11310 ;
  assign n11312 = ~n11267 & ~n11272 ;
  assign n11313 = ~n11311 & n11312 ;
  assign n11314 = ~n11268 & ~n11313 ;
  assign n11316 = n11306 & n11314 ;
  assign n11315 = ~n11306 & ~n11314 ;
  assign n11317 = n10878 & ~n11315 ;
  assign n11318 = ~n11316 & n11317 ;
  assign n11320 = \P1_reg2_reg[17]/NET0131  & n783 ;
  assign n11321 = ~\P1_reg2_reg[17]/NET0131  & ~n783 ;
  assign n11322 = ~n11320 & ~n11321 ;
  assign n11323 = ~n11170 & ~n11214 ;
  assign n11324 = ~n11218 & n11323 ;
  assign n11325 = ~n11213 & ~n11235 ;
  assign n11326 = ~n11324 & n11325 ;
  assign n11327 = ~n11236 & ~n11326 ;
  assign n11328 = ~n11284 & n11327 ;
  assign n11329 = ~n11281 & ~n11286 ;
  assign n11330 = ~n11328 & n11329 ;
  assign n11331 = ~n11282 & ~n11330 ;
  assign n11333 = n11322 & n11331 ;
  assign n11332 = ~n11322 & ~n11331 ;
  assign n11334 = n1936 & ~n11332 ;
  assign n11335 = ~n11333 & n11334 ;
  assign n11303 = n783 & n10891 ;
  assign n11319 = \P1_addr_reg[17]/NET0131  & ~n11063 ;
  assign n11336 = ~n11303 & ~n11319 ;
  assign n11337 = ~n11335 & n11336 ;
  assign n11338 = ~n11318 & n11337 ;
  assign n11339 = ~n11302 & ~n11338 ;
  assign n11340 = ~n6337 & ~n11339 ;
  assign n11341 = ~\P1_addr_reg[18]/NET0131  & n1897 ;
  assign n11342 = n6070 & ~n11341 ;
  assign n11343 = ~n1934 & ~n11342 ;
  assign n11358 = \P1_reg1_reg[18]/NET0131  & n741 ;
  assign n11359 = ~\P1_reg1_reg[18]/NET0131  & ~n741 ;
  assign n11360 = ~n11358 & ~n11359 ;
  assign n11361 = ~n11268 & ~n11305 ;
  assign n11362 = n11275 & n11361 ;
  assign n11363 = n11267 & ~n11305 ;
  assign n11364 = ~n11304 & ~n11363 ;
  assign n11365 = ~n11362 & n11364 ;
  assign n11367 = n11360 & ~n11365 ;
  assign n11366 = ~n11360 & n11365 ;
  assign n11368 = n10878 & ~n11366 ;
  assign n11369 = ~n11367 & n11368 ;
  assign n11346 = \P1_reg2_reg[18]/NET0131  & n741 ;
  assign n11347 = ~\P1_reg2_reg[18]/NET0131  & ~n741 ;
  assign n11348 = ~n11346 & ~n11347 ;
  assign n11349 = ~n11282 & ~n11321 ;
  assign n11350 = n11289 & n11349 ;
  assign n11351 = n11281 & ~n11321 ;
  assign n11352 = ~n11320 & ~n11351 ;
  assign n11353 = ~n11350 & n11352 ;
  assign n11355 = ~n11348 & n11353 ;
  assign n11354 = n11348 & ~n11353 ;
  assign n11356 = n1936 & ~n11354 ;
  assign n11357 = ~n11355 & n11356 ;
  assign n11344 = \P1_addr_reg[18]/NET0131  & n537 ;
  assign n11345 = n741 & n10891 ;
  assign n11370 = ~n11344 & ~n11345 ;
  assign n11371 = ~n11357 & n11370 ;
  assign n11372 = ~n11369 & n11371 ;
  assign n11373 = ~n11343 & ~n11372 ;
  assign n11374 = \P1_addr_reg[18]/NET0131  & n10966 ;
  assign n11375 = ~n5773 & ~n11374 ;
  assign n11376 = ~n11373 & n11375 ;
  assign n11377 = ~\P1_addr_reg[19]/NET0131  & n1897 ;
  assign n11378 = n6070 & ~n11377 ;
  assign n11379 = ~n1934 & ~n11378 ;
  assign n11393 = ~n11304 & ~n11314 ;
  assign n11394 = ~n11305 & ~n11359 ;
  assign n11395 = ~n11393 & n11394 ;
  assign n11396 = ~n11358 & ~n11395 ;
  assign n11397 = \P1_reg1_reg[19]/NET0131  & n516 ;
  assign n11398 = ~\P1_reg1_reg[19]/NET0131  & ~n516 ;
  assign n11399 = ~n11397 & ~n11398 ;
  assign n11401 = ~n11396 & ~n11399 ;
  assign n11400 = n11396 & n11399 ;
  assign n11402 = n10878 & ~n11400 ;
  assign n11403 = ~n11401 & n11402 ;
  assign n11382 = ~n11320 & ~n11331 ;
  assign n11383 = ~n11321 & ~n11347 ;
  assign n11384 = ~n11382 & n11383 ;
  assign n11385 = ~n11346 & ~n11384 ;
  assign n11386 = \P1_reg2_reg[19]/NET0131  & n516 ;
  assign n11387 = ~\P1_reg2_reg[19]/NET0131  & ~n516 ;
  assign n11388 = ~n11386 & ~n11387 ;
  assign n11390 = ~n11385 & ~n11388 ;
  assign n11389 = n11385 & n11388 ;
  assign n11391 = n1936 & ~n11389 ;
  assign n11392 = ~n11390 & n11391 ;
  assign n11380 = \P1_addr_reg[19]/NET0131  & n537 ;
  assign n11381 = ~n516 & n10891 ;
  assign n11404 = ~n11380 & ~n11381 ;
  assign n11405 = ~n11392 & n11404 ;
  assign n11406 = ~n11403 & n11405 ;
  assign n11407 = ~n11379 & ~n11406 ;
  assign n11408 = \P1_addr_reg[19]/NET0131  & n10966 ;
  assign n11409 = ~n6341 & ~n11408 ;
  assign n11410 = ~n11407 & n11409 ;
  assign n11411 = ~\P1_addr_reg[15]/NET0131  & n1897 ;
  assign n11412 = n6070 & ~n11411 ;
  assign n11413 = ~n1934 & ~n11412 ;
  assign n11421 = ~n11270 & ~n11272 ;
  assign n11423 = ~n11310 & ~n11421 ;
  assign n11422 = n11310 & n11421 ;
  assign n11424 = n10878 & ~n11422 ;
  assign n11425 = ~n11423 & n11424 ;
  assign n11416 = ~n11284 & ~n11286 ;
  assign n11418 = ~n11327 & ~n11416 ;
  assign n11417 = n11327 & n11416 ;
  assign n11419 = n1936 & ~n11417 ;
  assign n11420 = ~n11418 & n11419 ;
  assign n11414 = n1013 & n10891 ;
  assign n11415 = \P1_addr_reg[15]/NET0131  & ~n11063 ;
  assign n11426 = ~n11414 & ~n11415 ;
  assign n11427 = ~n11420 & n11426 ;
  assign n11428 = ~n11425 & n11427 ;
  assign n11429 = ~n11413 & ~n11428 ;
  assign n11430 = ~n7054 & ~n11429 ;
  assign n11431 = \P1_reg3_reg[1]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11432 = ~\P1_addr_reg[1]/NET0131  & n1897 ;
  assign n11433 = n6070 & ~n11432 ;
  assign n11434 = ~n1934 & ~n11433 ;
  assign n11435 = \P1_addr_reg[1]/NET0131  & ~n11063 ;
  assign n11442 = ~n10909 & ~n10910 ;
  assign n11443 = ~n10875 & ~n11442 ;
  assign n11444 = n10875 & n11442 ;
  assign n11445 = ~n11443 & ~n11444 ;
  assign n11446 = n1936 & n11445 ;
  assign n11436 = ~n10896 & ~n10897 ;
  assign n11437 = ~n10879 & ~n11436 ;
  assign n11438 = n10879 & n11436 ;
  assign n11439 = ~n11437 & ~n11438 ;
  assign n11440 = n10878 & n11439 ;
  assign n11441 = ~n1371 & n10891 ;
  assign n11447 = ~n11440 & ~n11441 ;
  assign n11448 = ~n11446 & n11447 ;
  assign n11449 = ~n11435 & n11448 ;
  assign n11450 = ~n11434 & ~n11449 ;
  assign n11451 = ~n11431 & ~n11450 ;
  assign n11458 = ~n10999 & ~n11000 ;
  assign n11460 = n11002 & n11458 ;
  assign n11459 = ~n11002 & ~n11458 ;
  assign n11461 = n10878 & ~n11459 ;
  assign n11462 = ~n11460 & n11461 ;
  assign n11452 = ~n1286 & n10891 ;
  assign n11453 = ~n10978 & ~n10979 ;
  assign n11455 = n10981 & n11453 ;
  assign n11454 = ~n10981 & ~n11453 ;
  assign n11456 = n1936 & ~n11454 ;
  assign n11457 = ~n11455 & n11456 ;
  assign n11463 = ~n11452 & ~n11457 ;
  assign n11464 = ~n11462 & n11463 ;
  assign n11465 = n10968 & ~n11464 ;
  assign n11466 = \P1_addr_reg[5]/NET0131  & \P1_state_reg[0]/NET0131  ;
  assign n11467 = ~n3664 & n11466 ;
  assign n11468 = ~n11063 & n11467 ;
  assign n11469 = ~n8184 & ~n11468 ;
  assign n11470 = ~n11465 & n11469 ;
  assign n11472 = ~\P1_addr_reg[9]/NET0131  & n1897 ;
  assign n11473 = n6070 & ~n11472 ;
  assign n11474 = ~n1934 & ~n11473 ;
  assign n11482 = ~n11112 & ~n11113 ;
  assign n11484 = ~n11115 & ~n11482 ;
  assign n11483 = n11115 & n11482 ;
  assign n11485 = n10878 & ~n11483 ;
  assign n11486 = ~n11484 & n11485 ;
  assign n11477 = ~n11099 & ~n11101 ;
  assign n11479 = ~n11148 & ~n11477 ;
  assign n11478 = n11148 & n11477 ;
  assign n11480 = n1936 & ~n11478 ;
  assign n11481 = ~n11479 & n11480 ;
  assign n11475 = \P1_addr_reg[9]/NET0131  & n537 ;
  assign n11476 = n1176 & n10891 ;
  assign n11487 = ~n11475 & ~n11476 ;
  assign n11488 = ~n11481 & n11487 ;
  assign n11489 = ~n11486 & n11488 ;
  assign n11490 = ~n11474 & ~n11489 ;
  assign n11471 = \P1_addr_reg[9]/NET0131  & n10966 ;
  assign n11491 = ~n6471 & ~n11471 ;
  assign n11492 = ~n11490 & n11491 ;
  assign n11493 = \P1_state_reg[0]/NET0131  & n3430 ;
  assign n11494 = \P1_state_reg[0]/NET0131  & n3664 ;
  assign n11497 = n2480 & ~n4925 ;
  assign n11501 = n4925 & ~n5522 ;
  assign n11502 = ~n11497 & ~n11501 ;
  assign n11503 = n3319 & ~n11502 ;
  assign n11498 = n4925 & ~n5536 ;
  assign n11499 = ~n11497 & ~n11498 ;
  assign n11500 = n3179 & ~n11499 ;
  assign n11504 = n4925 & ~n5505 ;
  assign n11496 = n2471 & ~n5093 ;
  assign n11505 = ~n3178 & n3371 ;
  assign n11506 = ~n4925 & n11505 ;
  assign n11507 = ~n5090 & ~n11506 ;
  assign n11508 = n2480 & ~n11507 ;
  assign n11509 = ~n11496 & ~n11508 ;
  assign n11510 = ~n11504 & n11509 ;
  assign n11511 = ~n11500 & n11510 ;
  assign n11512 = ~n11503 & n11511 ;
  assign n11513 = n4275 & ~n11512 ;
  assign n11495 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[24]/NET0131  ;
  assign n11514 = \P1_state_reg[0]/NET0131  & ~n2017 ;
  assign n11515 = n2480 & n11514 ;
  assign n11516 = ~n11495 & ~n11515 ;
  assign n11517 = ~n11513 & n11516 ;
  assign n11520 = n2429 & ~n4925 ;
  assign n11521 = n4925 & ~n5302 ;
  assign n11522 = ~n11520 & ~n11521 ;
  assign n11523 = n3179 & ~n11522 ;
  assign n11524 = n4925 & ~n5331 ;
  assign n11525 = ~n11520 & ~n11524 ;
  assign n11526 = n3319 & ~n11525 ;
  assign n11527 = n4925 & n5339 ;
  assign n11528 = ~n11520 & ~n11527 ;
  assign n11529 = n3373 & ~n11528 ;
  assign n11530 = n4925 & n5344 ;
  assign n11519 = n2424 & ~n5093 ;
  assign n11531 = n2429 & n4934 ;
  assign n11532 = ~n11519 & ~n11531 ;
  assign n11533 = ~n11530 & n11532 ;
  assign n11534 = ~n11529 & n11533 ;
  assign n11535 = ~n11526 & n11534 ;
  assign n11536 = ~n11523 & n11535 ;
  assign n11537 = n4275 & ~n11536 ;
  assign n11518 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[26]/NET0131  ;
  assign n11538 = n2429 & n11514 ;
  assign n11539 = ~n11518 & ~n11538 ;
  assign n11540 = ~n11537 & n11539 ;
  assign n11547 = n3319 & ~n6039 ;
  assign n11548 = n6059 & ~n11547 ;
  assign n11549 = n2033 & ~n11548 ;
  assign n11541 = \P2_reg2_reg[22]/NET0131  & ~n2033 ;
  assign n11546 = n3420 & n11541 ;
  assign n11550 = n2527 & n3415 ;
  assign n11551 = ~n11546 & ~n11550 ;
  assign n11552 = ~n11549 & n11551 ;
  assign n11553 = n4275 & ~n11552 ;
  assign n11542 = n2033 & n4275 ;
  assign n11543 = ~n6026 & n11542 ;
  assign n11544 = ~n11541 & ~n11543 ;
  assign n11545 = n3179 & ~n11544 ;
  assign n11554 = ~n3418 & n4275 ;
  assign n11555 = ~n3417 & n11554 ;
  assign n11556 = ~n6794 & n11555 ;
  assign n11557 = \P2_reg2_reg[22]/NET0131  & ~n11556 ;
  assign n11558 = ~n11545 & ~n11557 ;
  assign n11559 = ~n11553 & n11558 ;
  assign n11560 = ~\P1_rd_reg/NET0131  & ~\P2_rd_reg/NET0131  ;
  assign n11561 = \P1_rd_reg/NET0131  & \P2_rd_reg/NET0131  ;
  assign n11562 = ~n11560 & ~n11561 ;
  assign n11563 = \P1_addr_reg[0]/NET0131  & \P2_addr_reg[0]/NET0131  ;
  assign n11564 = ~\P1_addr_reg[0]/NET0131  & ~\P2_addr_reg[0]/NET0131  ;
  assign n11565 = ~n11563 & ~n11564 ;
  assign n11566 = \P1_addr_reg[10]/NET0131  & \P2_addr_reg[10]/NET0131  ;
  assign n11567 = ~\P1_addr_reg[10]/NET0131  & ~\P2_addr_reg[10]/NET0131  ;
  assign n11568 = ~n11566 & ~n11567 ;
  assign n11569 = ~\P1_addr_reg[9]/NET0131  & ~\P2_addr_reg[9]/NET0131  ;
  assign n11570 = \P1_addr_reg[9]/NET0131  & \P2_addr_reg[9]/NET0131  ;
  assign n11571 = ~\P1_addr_reg[8]/NET0131  & ~\P2_addr_reg[8]/NET0131  ;
  assign n11572 = \P1_addr_reg[8]/NET0131  & \P2_addr_reg[8]/NET0131  ;
  assign n11573 = ~\P1_addr_reg[7]/NET0131  & ~\P2_addr_reg[7]/NET0131  ;
  assign n11574 = \P1_addr_reg[7]/NET0131  & \P2_addr_reg[7]/NET0131  ;
  assign n11575 = ~\P1_addr_reg[6]/NET0131  & ~\P2_addr_reg[6]/NET0131  ;
  assign n11576 = \P1_addr_reg[6]/NET0131  & \P2_addr_reg[6]/NET0131  ;
  assign n11577 = ~\P1_addr_reg[5]/NET0131  & ~\P2_addr_reg[5]/NET0131  ;
  assign n11578 = \P1_addr_reg[5]/NET0131  & \P2_addr_reg[5]/NET0131  ;
  assign n11579 = ~\P1_addr_reg[4]/NET0131  & ~\P2_addr_reg[4]/NET0131  ;
  assign n11580 = \P1_addr_reg[4]/NET0131  & \P2_addr_reg[4]/NET0131  ;
  assign n11581 = ~\P1_addr_reg[3]/NET0131  & ~\P2_addr_reg[3]/NET0131  ;
  assign n11582 = \P1_addr_reg[3]/NET0131  & \P2_addr_reg[3]/NET0131  ;
  assign n11583 = ~\P1_addr_reg[2]/NET0131  & ~\P2_addr_reg[2]/NET0131  ;
  assign n11584 = \P1_addr_reg[2]/NET0131  & \P2_addr_reg[2]/NET0131  ;
  assign n11585 = ~\P1_addr_reg[1]/NET0131  & ~\P2_addr_reg[1]/NET0131  ;
  assign n11586 = \P1_addr_reg[1]/NET0131  & \P2_addr_reg[1]/NET0131  ;
  assign n11587 = ~n11563 & ~n11586 ;
  assign n11588 = ~n11585 & ~n11587 ;
  assign n11589 = ~n11584 & ~n11588 ;
  assign n11590 = ~n11583 & ~n11589 ;
  assign n11591 = ~n11582 & ~n11590 ;
  assign n11592 = ~n11581 & ~n11591 ;
  assign n11593 = ~n11580 & ~n11592 ;
  assign n11594 = ~n11579 & ~n11593 ;
  assign n11595 = ~n11578 & ~n11594 ;
  assign n11596 = ~n11577 & ~n11595 ;
  assign n11597 = ~n11576 & ~n11596 ;
  assign n11598 = ~n11575 & ~n11597 ;
  assign n11599 = ~n11574 & ~n11598 ;
  assign n11600 = ~n11573 & ~n11599 ;
  assign n11601 = ~n11572 & ~n11600 ;
  assign n11602 = ~n11571 & ~n11601 ;
  assign n11603 = ~n11570 & ~n11602 ;
  assign n11604 = ~n11569 & ~n11603 ;
  assign n11605 = ~n11568 & n11604 ;
  assign n11606 = n11568 & ~n11604 ;
  assign n11607 = ~n11605 & ~n11606 ;
  assign n11608 = \P1_addr_reg[11]/NET0131  & \P2_addr_reg[11]/NET0131  ;
  assign n11609 = ~\P1_addr_reg[11]/NET0131  & ~\P2_addr_reg[11]/NET0131  ;
  assign n11610 = ~n11608 & ~n11609 ;
  assign n11611 = ~n11566 & ~n11604 ;
  assign n11612 = ~n11567 & ~n11611 ;
  assign n11613 = ~n11610 & n11612 ;
  assign n11614 = n11610 & ~n11612 ;
  assign n11615 = ~n11613 & ~n11614 ;
  assign n11616 = \P1_addr_reg[12]/NET0131  & \P2_addr_reg[12]/NET0131  ;
  assign n11617 = ~\P1_addr_reg[12]/NET0131  & ~\P2_addr_reg[12]/NET0131  ;
  assign n11618 = ~n11616 & ~n11617 ;
  assign n11619 = ~n11608 & ~n11612 ;
  assign n11620 = ~n11609 & ~n11619 ;
  assign n11621 = ~n11618 & n11620 ;
  assign n11622 = n11618 & ~n11620 ;
  assign n11623 = ~n11621 & ~n11622 ;
  assign n11624 = \P1_addr_reg[13]/NET0131  & \P2_addr_reg[13]/NET0131  ;
  assign n11625 = ~\P1_addr_reg[13]/NET0131  & ~\P2_addr_reg[13]/NET0131  ;
  assign n11626 = ~n11624 & ~n11625 ;
  assign n11627 = ~n11616 & ~n11620 ;
  assign n11628 = ~n11617 & ~n11627 ;
  assign n11629 = ~n11626 & n11628 ;
  assign n11630 = n11626 & ~n11628 ;
  assign n11631 = ~n11629 & ~n11630 ;
  assign n11632 = \P1_addr_reg[14]/NET0131  & \P2_addr_reg[14]/NET0131  ;
  assign n11633 = ~\P1_addr_reg[14]/NET0131  & ~\P2_addr_reg[14]/NET0131  ;
  assign n11634 = ~n11632 & ~n11633 ;
  assign n11635 = ~n11624 & ~n11628 ;
  assign n11636 = ~n11625 & ~n11635 ;
  assign n11637 = ~n11634 & n11636 ;
  assign n11638 = n11634 & ~n11636 ;
  assign n11639 = ~n11637 & ~n11638 ;
  assign n11640 = \P1_addr_reg[15]/NET0131  & \P2_addr_reg[15]/NET0131  ;
  assign n11641 = ~\P1_addr_reg[15]/NET0131  & ~\P2_addr_reg[15]/NET0131  ;
  assign n11642 = ~n11640 & ~n11641 ;
  assign n11643 = ~n11632 & ~n11636 ;
  assign n11644 = ~n11633 & ~n11643 ;
  assign n11645 = ~n11642 & n11644 ;
  assign n11646 = n11642 & ~n11644 ;
  assign n11647 = ~n11645 & ~n11646 ;
  assign n11648 = \P1_addr_reg[16]/NET0131  & \P2_addr_reg[16]/NET0131  ;
  assign n11649 = ~\P1_addr_reg[16]/NET0131  & ~\P2_addr_reg[16]/NET0131  ;
  assign n11650 = ~n11648 & ~n11649 ;
  assign n11651 = ~n11640 & ~n11644 ;
  assign n11652 = ~n11641 & ~n11651 ;
  assign n11653 = ~n11650 & n11652 ;
  assign n11654 = n11650 & ~n11652 ;
  assign n11655 = ~n11653 & ~n11654 ;
  assign n11656 = \P1_addr_reg[17]/NET0131  & \P2_addr_reg[17]/NET0131  ;
  assign n11657 = ~\P1_addr_reg[17]/NET0131  & ~\P2_addr_reg[17]/NET0131  ;
  assign n11658 = ~n11656 & ~n11657 ;
  assign n11659 = ~n11648 & ~n11652 ;
  assign n11660 = ~n11649 & ~n11659 ;
  assign n11661 = ~n11658 & n11660 ;
  assign n11662 = n11658 & ~n11660 ;
  assign n11663 = ~n11661 & ~n11662 ;
  assign n11664 = \P1_addr_reg[18]/NET0131  & \P2_addr_reg[18]/NET0131  ;
  assign n11665 = ~\P1_addr_reg[18]/NET0131  & ~\P2_addr_reg[18]/NET0131  ;
  assign n11666 = ~n11664 & ~n11665 ;
  assign n11667 = ~n11656 & ~n11660 ;
  assign n11668 = ~n11657 & ~n11667 ;
  assign n11669 = ~n11666 & n11668 ;
  assign n11670 = n11666 & ~n11668 ;
  assign n11671 = ~n11669 & ~n11670 ;
  assign n11672 = ~n538 & ~n540 ;
  assign n11673 = ~n11664 & ~n11668 ;
  assign n11674 = ~n11665 & ~n11673 ;
  assign n11675 = n11672 & ~n11674 ;
  assign n11676 = ~n11672 & n11674 ;
  assign n11677 = ~n11675 & ~n11676 ;
  assign n11678 = ~n11585 & ~n11586 ;
  assign n11679 = n11563 & ~n11678 ;
  assign n11680 = ~n11563 & n11678 ;
  assign n11681 = ~n11679 & ~n11680 ;
  assign n11682 = ~n11583 & ~n11584 ;
  assign n11683 = n11588 & ~n11682 ;
  assign n11684 = ~n11588 & n11682 ;
  assign n11685 = ~n11683 & ~n11684 ;
  assign n11686 = ~n11581 & ~n11582 ;
  assign n11687 = n11590 & ~n11686 ;
  assign n11688 = ~n11590 & n11686 ;
  assign n11689 = ~n11687 & ~n11688 ;
  assign n11690 = ~n11579 & ~n11580 ;
  assign n11691 = n11592 & ~n11690 ;
  assign n11692 = ~n11592 & n11690 ;
  assign n11693 = ~n11691 & ~n11692 ;
  assign n11694 = ~n11577 & ~n11578 ;
  assign n11695 = n11594 & ~n11694 ;
  assign n11696 = ~n11594 & n11694 ;
  assign n11697 = ~n11695 & ~n11696 ;
  assign n11698 = ~n11575 & ~n11576 ;
  assign n11699 = n11596 & ~n11698 ;
  assign n11700 = ~n11596 & n11698 ;
  assign n11701 = ~n11699 & ~n11700 ;
  assign n11702 = ~n11573 & ~n11574 ;
  assign n11703 = n11598 & ~n11702 ;
  assign n11704 = ~n11598 & n11702 ;
  assign n11705 = ~n11703 & ~n11704 ;
  assign n11706 = ~n11571 & ~n11572 ;
  assign n11707 = n11600 & ~n11706 ;
  assign n11708 = ~n11600 & n11706 ;
  assign n11709 = ~n11707 & ~n11708 ;
  assign n11710 = ~n11569 & ~n11570 ;
  assign n11711 = n11602 & ~n11710 ;
  assign n11712 = ~n11602 & n11710 ;
  assign n11713 = ~n11711 & ~n11712 ;
  assign n11714 = ~\P1_wr_reg/NET0131  & ~\P2_wr_reg/NET0131  ;
  assign n11715 = \P1_wr_reg/NET0131  & \P2_wr_reg/NET0131  ;
  assign n11716 = ~n11714 & ~n11715 ;
  assign \P1_state_reg[0]/NET0131_syn_2  = ~\P1_state_reg[0]/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g70791/_0_  = ~n1957 ;
  assign \g70792/_0_  = ~n3436 ;
  assign \g70793/_0_  = ~n3671 ;
  assign \g70794/_0_  = ~n3705 ;
  assign \g70795/_0_  = ~n3897 ;
  assign \g70796/_0_  = ~n3927 ;
  assign \g70813/_0_  = ~n4233 ;
  assign \g70814/_0_  = ~n4262 ;
  assign \g70848/_0_  = ~n4280 ;
  assign \g70849/_0_  = ~n4342 ;
  assign \g70850/_0_  = ~n4448 ;
  assign \g70851/_0_  = ~n4548 ;
  assign \g70852/_0_  = ~n4609 ;
  assign \g70856/_0_  = ~n4633 ;
  assign \g70857/_0_  = ~n4662 ;
  assign \g70858/_0_  = ~n4691 ;
  assign \g70859/_0_  = ~n4715 ;
  assign \g70860/_0_  = ~n4741 ;
  assign \g70861/_0_  = ~n4769 ;
  assign \g70862/_0_  = ~n4787 ;
  assign \g70896/_0_  = ~n4831 ;
  assign \g70902/_0_  = ~n4865 ;
  assign \g70903/_0_  = ~n4921 ;
  assign \g70904/_0_  = ~n4950 ;
  assign \g70906/_0_  = ~n4976 ;
  assign \g70907/_0_  = ~n5076 ;
  assign \g70908/_0_  = ~n5107 ;
  assign \g70909/_0_  = ~n5227 ;
  assign \g70910/_0_  = ~n5247 ;
  assign \g70911/_0_  = ~n5270 ;
  assign \g70912/_0_  = ~n5357 ;
  assign \g70913/_0_  = ~n5384 ;
  assign \g70914/_0_  = ~n5392 ;
  assign \g70915/_0_  = ~n5439 ;
  assign \g70916/_0_  = ~n5462 ;
  assign \g70917/_0_  = ~n5491 ;
  assign \g70918/_0_  = ~n5546 ;
  assign \g70919/_0_  = ~n5564 ;
  assign \g70920/_0_  = ~n5578 ;
  assign \g70921/_0_  = ~n5604 ;
  assign \g70922/_0_  = ~n5611 ;
  assign \g70923/_0_  = ~n5639 ;
  assign \g70924/_0_  = ~n5655 ;
  assign \g70925/_0_  = ~n5681 ;
  assign \g70926/_0_  = ~n5707 ;
  assign \g70927/_0_  = ~n5733 ;
  assign \g70987/_0_  = ~n5772 ;
  assign \g70988/_0_  = ~n5817 ;
  assign \g70989/_0_  = ~n5865 ;
  assign \g70990/_0_  = ~n5907 ;
  assign \g70991/_0_  = ~n5948 ;
  assign \g71006/_0_  = ~n5992 ;
  assign \g71007/_0_  = ~n6018 ;
  assign \g71009/_0_  = ~n6068 ;
  assign \g71010/_0_  = ~n6084 ;
  assign \g71011/_0_  = ~n6102 ;
  assign \g71012/_0_  = ~n6124 ;
  assign \g71013/_0_  = ~n6144 ;
  assign \g71014/_0_  = ~n6164 ;
  assign \g71015/_0_  = ~n6173 ;
  assign \g71016/_0_  = ~n6208 ;
  assign \g71017/_0_  = ~n6234 ;
  assign \g71018/_0_  = ~n6240 ;
  assign \g71019/_0_  = ~n6248 ;
  assign \g71020/_0_  = ~n6265 ;
  assign \g71021/_0_  = ~n6283 ;
  assign \g71022/_0_  = ~n6309 ;
  assign \g71023/_0_  = ~n6313 ;
  assign \g71090/_0_  = ~n6339 ;
  assign \g71091/_0_  = ~n6382 ;
  assign \g71092/_0_  = ~n6424 ;
  assign \g71093/_0_  = ~n6470 ;
  assign \g71094/_0_  = ~n6511 ;
  assign \g71125/_0_  = ~n6541 ;
  assign \g71130/_0_  = ~n6557 ;
  assign \g71131/_0_  = ~n6603 ;
  assign \g71132/_0_  = ~n6629 ;
  assign \g71133/_0_  = ~n6637 ;
  assign \g71134/_0_  = ~n6663 ;
  assign \g71135/_0_  = ~n6680 ;
  assign \g71136/_0_  = ~n6704 ;
  assign \g71137/_0_  = ~n6724 ;
  assign \g71138/_0_  = ~n6746 ;
  assign \g71139/_0_  = ~n6756 ;
  assign \g71140/_0_  = ~n6774 ;
  assign \g71141/_0_  = ~n6777 ;
  assign \g71142/_0_  = ~n6792 ;
  assign \g71143/_0_  = ~n6803 ;
  assign \g71144/_0_  = ~n6812 ;
  assign \g71145/_0_  = ~n6854 ;
  assign \g71150/_0_  = ~n6866 ;
  assign \g71151/_0_  = ~n6879 ;
  assign \g71152/_0_  = ~n6882 ;
  assign \g71153/_0_  = ~n6885 ;
  assign \g71154/_0_  = ~n6898 ;
  assign \g71155/_0_  = ~n6906 ;
  assign \g71156/_0_  = ~n6924 ;
  assign \g71157/_0_  = ~n6927 ;
  assign \g71158/_0_  = ~n6930 ;
  assign \g71230/_0_  = ~n6972 ;
  assign \g71231/_0_  = ~n7014 ;
  assign \g71232/_0_  = ~n7053 ;
  assign \g71233/_0_  = ~n7096 ;
  assign \g71234/_0_  = ~n7140 ;
  assign \g71235/_0_  = ~n7183 ;
  assign \g71236/_0_  = ~n7225 ;
  assign \g71238/_0_  = ~n7267 ;
  assign \g71239/_0_  = ~n7308 ;
  assign \g71270/_0_  = ~n7331 ;
  assign \g71275/_0_  = ~n7379 ;
  assign \g71276/_0_  = ~n7420 ;
  assign \g71277/_0_  = ~n7466 ;
  assign \g71278/_0_  = ~n7491 ;
  assign \g71279/_0_  = ~n7498 ;
  assign \g71280/_0_  = ~n7520 ;
  assign \g71281/_0_  = ~n7536 ;
  assign \g71282/_0_  = ~n7565 ;
  assign \g71283/_0_  = ~n7588 ;
  assign \g71284/_0_  = ~n7612 ;
  assign \g71285/_0_  = ~n7630 ;
  assign \g71286/_0_  = ~n7633 ;
  assign \g71287/_0_  = ~n7655 ;
  assign \g71288/_0_  = ~n7660 ;
  assign \g71289/_0_  = ~n7681 ;
  assign \g71290/_0_  = ~n7692 ;
  assign \g71291/_0_  = ~n7701 ;
  assign \g71292/_0_  = ~n7725 ;
  assign \g71293/_0_  = ~n7751 ;
  assign \g71294/_0_  = ~n7763 ;
  assign \g71295/_0_  = ~n7785 ;
  assign \g71296/_0_  = ~n7808 ;
  assign \g71297/_0_  = ~n7819 ;
  assign \g71298/_0_  = ~n7837 ;
  assign \g71299/_0_  = ~n7840 ;
  assign \g71300/_0_  = ~n7858 ;
  assign \g71301/_0_  = ~n7880 ;
  assign \g71302/_0_  = ~n7902 ;
  assign \g71303/_0_  = ~n7913 ;
  assign \g71304/_0_  = ~n7932 ;
  assign \g71305/_0_  = ~n7961 ;
  assign \g71306/_0_  = ~n7981 ;
  assign \g71307/_0_  = ~n7985 ;
  assign \g71382/_0_  = ~n8021 ;
  assign \g71384/_0_  = ~n8061 ;
  assign \g71385/_0_  = ~n8102 ;
  assign \g71387/_0_  = ~n8142 ;
  assign \g71388/_0_  = ~n8183 ;
  assign \g71389/_0_  = ~n8221 ;
  assign \g71439/_0_  = ~n8243 ;
  assign \g71440/_0_  = ~n8267 ;
  assign \g71441/_0_  = ~n8293 ;
  assign \g71442/_0_  = ~n8303 ;
  assign \g71443/_0_  = ~n8318 ;
  assign \g71444/_0_  = ~n8347 ;
  assign \g71445/_0_  = ~n8369 ;
  assign \g71446/_0_  = ~n8393 ;
  assign \g71447/_0_  = ~n8415 ;
  assign \g71448/_0_  = ~n8437 ;
  assign \g71449/_0_  = ~n8459 ;
  assign \g71450/_0_  = ~n8481 ;
  assign \g71451/_0_  = ~n8505 ;
  assign \g71452/_0_  = ~n8529 ;
  assign \g71453/_0_  = ~n8553 ;
  assign \g71454/_0_  = ~n8582 ;
  assign \g71455/_0_  = ~n8606 ;
  assign \g71456/_0_  = ~n8632 ;
  assign \g71457/_0_  = ~n8658 ;
  assign \g71458/_0_  = ~n8680 ;
  assign \g71459/_0_  = ~n8702 ;
  assign \g71460/_0_  = ~n8720 ;
  assign \g71461/_0_  = ~n8724 ;
  assign \g71536/_0_  = ~n8762 ;
  assign \g71537/_0_  = ~n8799 ;
  assign \g71538/_0_  = ~n8840 ;
  assign \g71540/_0_  = ~n8880 ;
  assign \g71541/_0_  = ~n8919 ;
  assign \g71542/_0_  = ~n8955 ;
  assign \g71602/_0_  = ~n8970 ;
  assign \g71604/_0_  = ~n8979 ;
  assign \g71610/_0_  = n8994 ;
  assign \g71611/_0_  = ~n9020 ;
  assign \g71618/_0_  = ~n9023 ;
  assign \g71619/_0_  = ~n9045 ;
  assign \g71620/_0_  = ~n9056 ;
  assign \g71621/_0_  = ~n9078 ;
  assign \g71622/_0_  = ~n9100 ;
  assign \g71623/_0_  = n9113 ;
  assign \g71624/_0_  = ~n9119 ;
  assign \g71625/_0_  = ~n9145 ;
  assign \g71626/_0_  = ~n9163 ;
  assign \g71627/_0_  = ~n9172 ;
  assign \g71629/_0_  = ~n9176 ;
  assign \g71630/_0_  = ~n9179 ;
  assign \g71631/_0_  = ~n9182 ;
  assign \g71632/_0_  = ~n9204 ;
  assign \g71633/_0_  = ~n9222 ;
  assign \g71634/_0_  = ~n9231 ;
  assign \g71635/_0_  = ~n9239 ;
  assign \g71636/_0_  = ~n9243 ;
  assign \g71710/_0_  = ~n9284 ;
  assign \g71711/_0_  = ~n9324 ;
  assign \g71782/_0_  = ~n9349 ;
  assign \g71785/_0_  = ~n9357 ;
  assign \g71786/_0_  = ~n9375 ;
  assign \g71787/_0_  = ~n9397 ;
  assign \g71788/_0_  = ~n9419 ;
  assign \g71789/_0_  = ~n9437 ;
  assign \g71790/_0_  = ~n9454 ;
  assign \g71791/_0_  = ~n9472 ;
  assign \g71792/_0_  = n9485 ;
  assign \g71793/_0_  = ~n9491 ;
  assign \g71794/_0_  = ~n9508 ;
  assign \g71795/_0_  = ~n9538 ;
  assign \g71796/_0_  = ~n9541 ;
  assign \g71797/_0_  = ~n9544 ;
  assign \g71798/_0_  = ~n9566 ;
  assign \g71799/_0_  = ~n9574 ;
  assign \g71883/_0_  = ~n9606 ;
  assign \g72000/_0_  = ~n9613 ;
  assign \g72001/_0_  = ~n9635 ;
  assign \g72002/_0_  = ~n9653 ;
  assign \g72003/_0_  = ~n9683 ;
  assign \g72004/_0_  = ~n9707 ;
  assign \g72005/_0_  = ~n9710 ;
  assign \g72236/_0_  = ~n9728 ;
  assign \g72237/_0_  = n9741 ;
  assign \g72238/_0_  = ~n9759 ;
  assign \g72239/_0_  = ~n9762 ;
  assign \g72240/_0_  = ~n9765 ;
  assign \g72372/_0_  = ~n9793 ;
  assign \g72376/_0_  = n9826 ;
  assign \g72383/_0_  = n9857 ;
  assign \g72561/_0_  = ~n9864 ;
  assign \g72562/_0_  = ~n9873 ;
  assign \g72563/_0_  = ~n9885 ;
  assign \g72564/_0_  = ~n9894 ;
  assign \g72970/_0_  = ~n9917 ;
  assign \g72980/_0_  = ~n9927 ;
  assign \g72981/_0_  = ~n9937 ;
  assign \g72982/_0_  = n9951 ;
  assign \g72983/_0_  = ~n9961 ;
  assign \g74234/_0_  = ~n9978 ;
  assign \g74260/_0_  = ~n9995 ;
  assign \g75086/_0_  = ~n10005 ;
  assign \g75087/_0_  = ~n10008 ;
  assign \g75088/_0_  = ~n10011 ;
  assign \g75089/_0_  = ~n10020 ;
  assign \g75091/_0_  = ~n10023 ;
  assign \g75092/_0_  = ~n10027 ;
  assign \g80304/_3_  = n10030 ;
  assign \g80305/_3_  = ~n10033 ;
  assign \g80306/_3_  = ~n10036 ;
  assign \g80307/_3_  = ~n10039 ;
  assign \g80308/_0_  = ~n10042 ;
  assign \g80309/_0_  = ~n10045 ;
  assign \g80815/_0_  = ~n10048 ;
  assign \g80816/_0_  = n10051 ;
  assign \g80817/_0_  = n10054 ;
  assign \g80818/_0_  = n10057 ;
  assign \g80819/_0_  = ~n10060 ;
  assign \g80820/_0_  = ~n10063 ;
  assign \g80821/_0_  = n10066 ;
  assign \g80822/_0_  = n10069 ;
  assign \g80823/_0_  = ~n10072 ;
  assign \g80824/_0_  = n10075 ;
  assign \g80825/_0_  = ~n10078 ;
  assign \g80826/_3_  = ~n10081 ;
  assign \g80827/_0_  = n10084 ;
  assign \g80828/_0_  = n10087 ;
  assign \g80829/_0_  = n10090 ;
  assign \g80830/_0_  = ~n10092 ;
  assign \g80831/_0_  = ~n10095 ;
  assign \g80832/_0_  = n10098 ;
  assign \g80833/_0_  = ~n10101 ;
  assign \g80834/_0_  = ~n10104 ;
  assign \g80835/_0_  = ~n10107 ;
  assign \g80836/_0_  = ~n10110 ;
  assign \g80837/_0_  = ~n10113 ;
  assign \g80838/_3_  = n10116 ;
  assign \g80839/_0_  = n10119 ;
  assign \g80840/_3_  = ~n10122 ;
  assign \g80841/_0_  = n10125 ;
  assign \g80859/_3_  = ~n10128 ;
  assign \g80860/_3_  = ~n10131 ;
  assign \g80861/_3_  = ~n10134 ;
  assign \g80862/_3_  = ~n10137 ;
  assign \g80863/_3_  = ~n10140 ;
  assign \g80864/_3_  = ~n10143 ;
  assign \g80865/_3_  = ~n10146 ;
  assign \g80866/_3_  = ~n10149 ;
  assign \g80867/_3_  = ~n10152 ;
  assign \g80868/_3_  = ~n10155 ;
  assign \g80869/_3_  = ~n10158 ;
  assign \g80870/_3_  = n10161 ;
  assign \g80871/_3_  = n10164 ;
  assign \g80872/_3_  = n10167 ;
  assign \g80873/_3_  = ~n10169 ;
  assign \g80874/_3_  = n10172 ;
  assign \g80875/_3_  = ~n10175 ;
  assign \g80876/_3_  = ~n10178 ;
  assign \g80877/_3_  = ~n10181 ;
  assign \g80878/_3_  = ~n10184 ;
  assign \g80879/_0_  = ~n10191 ;
  assign \g80880/_3_  = ~n10194 ;
  assign \g80881/_3_  = ~n10197 ;
  assign \g80882/_3_  = ~n10200 ;
  assign \g80883/_3_  = ~n10203 ;
  assign \g80884/_3_  = ~n10206 ;
  assign \g80885/_3_  = ~n10209 ;
  assign \g80886/_3_  = ~n10212 ;
  assign \g80888/_0_  = ~n10219 ;
  assign \g81262/_0_  = n2827 ;
  assign \g81278/_0_  = n1394 ;
  assign \g81884/_0_  = ~n10292 ;
  assign \g81893/_0_  = ~n10370 ;
  assign \g81896/_0_  = ~n10392 ;
  assign \g81897/_0_  = ~n10424 ;
  assign \g81898/_0_  = ~n10448 ;
  assign \g81899/_0_  = ~n10476 ;
  assign \g81900/_0_  = ~n10510 ;
  assign \g81901/_0_  = ~n10544 ;
  assign \g81902/_0_  = ~n10579 ;
  assign \g81903/_0_  = ~n10613 ;
  assign \g81904/_0_  = ~n10637 ;
  assign \g81905/_0_  = ~n10661 ;
  assign \g81906/_0_  = ~n10688 ;
  assign \g81907/_0_  = ~n10713 ;
  assign \g81908/_0_  = ~n10735 ;
  assign \g81909/_0_  = ~n10759 ;
  assign \g81910/_0_  = ~n10781 ;
  assign \g81911/_0_  = ~n10803 ;
  assign \g81923/_0_  = ~n10837 ;
  assign \g81924/_0_  = ~n10871 ;
  assign \g81925/_0_  = n10923 ;
  assign \g81926/_0_  = n10962 ;
  assign \g82414/_0_  = ~n10963 ;
  assign \g82532/_0_  = ~n10965 ;
  assign \g83134/_0_  = ~n11018 ;
  assign \g83135/_0_  = ~n11037 ;
  assign \g83141/_0_  = ~n11059 ;
  assign \g83142/_0_  = ~n11080 ;
  assign \g83145/_0_  = ~n11090 ;
  assign \g83146/_0_  = ~n11126 ;
  assign \g83147/_0_  = ~n11163 ;
  assign \g83148/_0_  = ~n11195 ;
  assign \g83152/_0_  = ~n11229 ;
  assign \g83153/_0_  = ~n11261 ;
  assign \g83154/_0_  = ~n11299 ;
  assign \g83155/_0_  = ~n11340 ;
  assign \g83156/_0_  = ~n11376 ;
  assign \g83157/_0_  = ~n11410 ;
  assign \g83158/_0_  = ~n11430 ;
  assign \g83159/_0_  = ~n11451 ;
  assign \g83164/_0_  = ~n11470 ;
  assign \g83165/_0_  = ~n11492 ;
  assign \g83177/_0_  = ~n2027 ;
  assign \g83178/_0_  = ~n3445 ;
  assign \g83409/_0_  = ~n2032 ;
  assign \g83411/_0_  = ~n3449 ;
  assign \g83807/u3_syn_4  = n11493 ;
  assign \g84138/u3_syn_4  = n11494 ;
  assign \g85062/_0_  = ~n3363 ;
  assign \g85079/_2_  = ~n2385 ;
  assign \g85113/_0_  = ~n2241 ;
  assign \g85121/_0_  = ~n3329 ;
  assign \g85594/_0_  = ~n3046 ;
  assign \g85663/_0_  = ~n1677 ;
  assign \g85669/_0_  = ~n1618 ;
  assign \g85749/_0_  = ~n2800 ;
  assign \g85784/_0_  = ~n2755 ;
  assign \g85809/_0_  = ~n2937 ;
  assign \g85817/_0_  = ~n3105 ;
  assign \g85828/_0_  = ~n3056 ;
  assign \g85845/_0_  = ~n2640 ;
  assign \g85851/_0_  = ~n2666 ;
  assign \g85858/_0_  = ~n2613 ;
  assign \g85871/_0_  = ~n2328 ;
  assign \g85882_dup/_0_  = ~n2588 ;
  assign \g85891/_0_  = ~n2551 ;
  assign \g85900/_0_  = ~n2531 ;
  assign \g85905/_0_  = ~n2507 ;
  assign \g85917/_0_  = ~n2433 ;
  assign \g85934/_0_  = ~n2678 ;
  assign \g85949/_0_  = ~n2911 ;
  assign \g85971/_0_  = ~n1702 ;
  assign \g85997/_0_  = ~n2823 ;
  assign \g86044/_0_  = ~n692 ;
  assign \g86053/_0_  = ~n1542 ;
  assign \g86063/_0_  = ~n1344 ;
  assign \g86082/_0_  = ~n1646 ;
  assign \g86088/_0_  = ~n921 ;
  assign \g86098/_0_  = ~n838 ;
  assign \g86105/_0_  = ~n1026 ;
  assign \g86179/_0_  = ~n999 ;
  assign \g86256_dup/_0_  = ~n1075 ;
  assign \g86264/_0_  = ~n1051 ;
  assign \g86273/_0_  = ~n1274 ;
  assign \g86281/_0_  = ~n887 ;
  assign \g86288/_0_  = ~n1115 ;
  assign \g86297/_0_  = ~n1138 ;
  assign \g86304/_0_  = ~n1189 ;
  assign \g86310/_0_  = ~n1162 ;
  assign \g86320/_0_  = ~n949 ;
  assign \g86328/_0_  = ~n973 ;
  assign \g86339/_0_  = ~n796 ;
  assign \g86353/_0_  = ~n1222 ;
  assign \g86360/_0_  = ~n1248 ;
  assign \g86368/_0_  = ~n752 ;
  assign \g86373/_0_  = ~n1298 ;
  assign \g86385/_0_  = ~n1322 ;
  assign \g86392/_0_  = ~n1390 ;
  assign \g86399/_0_  = ~n1367 ;
  assign \g86421/_0_  = ~n1570 ;
  assign \g86432/_0_  = ~n1510 ;
  assign \g87592/_1__syn_2  = n3434 ;
  assign \g87632/_1_  = n3703 ;
  assign \g92847/_0_  = ~n3082 ;
  assign \g92957/_0_  = ~n11517 ;
  assign \g93056/_0_  = ~n1478 ;
  assign \g93289/_0_  = ~n11540 ;
  assign \g93538_dup95061/_0_  = ~n2965 ;
  assign \g93856/_0_  = ~n11559 ;
  assign \g93870/_0_  = ~n2730 ;
  assign \g94004/_0_  = ~n2484 ;
  assign \g94128/_0_  = ~n2702 ;
  assign \g94173/_0_  = ~n2990 ;
  assign \g94187/_0_  = ~n2866 ;
  assign \g94191/_0_  = ~n2858 ;
  assign \g94318/_0_  = ~n2461 ;
  assign \g94505/_0_  = ~n2777 ;
  assign rd_pad = ~n11562 ;
  assign \so[0]_pad  = n11565 ;
  assign \so[10]_pad  = ~n11607 ;
  assign \so[11]_pad  = ~n11615 ;
  assign \so[12]_pad  = ~n11623 ;
  assign \so[13]_pad  = ~n11631 ;
  assign \so[14]_pad  = ~n11639 ;
  assign \so[15]_pad  = ~n11647 ;
  assign \so[16]_pad  = ~n11655 ;
  assign \so[17]_pad  = ~n11663 ;
  assign \so[18]_pad  = ~n11671 ;
  assign \so[19]_pad  = ~n11677 ;
  assign \so[1]_pad  = ~n11681 ;
  assign \so[2]_pad  = ~n11685 ;
  assign \so[3]_pad  = ~n11689 ;
  assign \so[4]_pad  = ~n11693 ;
  assign \so[5]_pad  = ~n11697 ;
  assign \so[6]_pad  = ~n11701 ;
  assign \so[7]_pad  = ~n11705 ;
  assign \so[8]_pad  = ~n11709 ;
  assign \so[9]_pad  = ~n11713 ;
  assign wr_pad = ~n11716 ;
endmodule
