module top( \ACVQN0_reg/NET0131  , \ACVQN1_reg/NET0131  , \ACVQN2_reg/NET0131  , \ACVQN3_reg/NET0131  , \AX0_reg/NET0131  , \AX1_reg/NET0131  , \AX2_reg/NET0131  , \AX3_reg/NET0131  , \B0_pad  , \B1_pad  , \B2_pad  , \B3_pad  , \CT0_reg/NET0131  , \CT1_reg/NET0131  , \CT2_reg/NET0131  , \MRVQN0_reg/NET0131  , \MRVQN1_reg/NET0131  , \MRVQN2_reg/NET0131  , \MRVQN3_reg/NET0131  , START_pad , \ACVQN0_reg/P0001  , \ACVQN1_reg/P0001  , \ACVQN2_reg/P0001  , \ACVQN3_reg/P0001  , \CNTVCON2_pad  , \MRVQN0_reg/P0001  , \P1_pad  , \P2_pad  , \P3_pad  , \_al_n0  , \_al_n1  , \g12/_2_  , \g25/_0_  , \g29/_0_  , \g614/_0_  , \g621/_0_  , \g623/_3_  , \g624/_3_  , \g625/_3_  , \g631/_0_  , \g635/_0_  , \g658/_1_  , \g765/_0_  , \g775/_2_  , \g782/_0_  );
  input \ACVQN0_reg/NET0131  ;
  input \ACVQN1_reg/NET0131  ;
  input \ACVQN2_reg/NET0131  ;
  input \ACVQN3_reg/NET0131  ;
  input \AX0_reg/NET0131  ;
  input \AX1_reg/NET0131  ;
  input \AX2_reg/NET0131  ;
  input \AX3_reg/NET0131  ;
  input \B0_pad  ;
  input \B1_pad  ;
  input \B2_pad  ;
  input \B3_pad  ;
  input \CT0_reg/NET0131  ;
  input \CT1_reg/NET0131  ;
  input \CT2_reg/NET0131  ;
  input \MRVQN0_reg/NET0131  ;
  input \MRVQN1_reg/NET0131  ;
  input \MRVQN2_reg/NET0131  ;
  input \MRVQN3_reg/NET0131  ;
  input START_pad ;
  output \ACVQN0_reg/P0001  ;
  output \ACVQN1_reg/P0001  ;
  output \ACVQN2_reg/P0001  ;
  output \ACVQN3_reg/P0001  ;
  output \CNTVCON2_pad  ;
  output \MRVQN0_reg/P0001  ;
  output \P1_pad  ;
  output \P2_pad  ;
  output \P3_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g12/_2_  ;
  output \g25/_0_  ;
  output \g29/_0_  ;
  output \g614/_0_  ;
  output \g621/_0_  ;
  output \g623/_3_  ;
  output \g624/_3_  ;
  output \g625/_3_  ;
  output \g631/_0_  ;
  output \g635/_0_  ;
  output \g658/_1_  ;
  output \g765/_0_  ;
  output \g775/_2_  ;
  output \g782/_0_  ;
  wire n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 ;
  assign n21 = \CT0_reg/NET0131  & \CT1_reg/NET0131  ;
  assign n22 = \CT2_reg/NET0131  & n21 ;
  assign n23 = \CT0_reg/NET0131  & ~\CT1_reg/NET0131  ;
  assign n24 = \CT2_reg/NET0131  & n23 ;
  assign n25 = ~\ACVQN0_reg/NET0131  & \AX0_reg/NET0131  ;
  assign n26 = ~\MRVQN0_reg/NET0131  & n25 ;
  assign n27 = \ACVQN1_reg/NET0131  & ~n26 ;
  assign n28 = ~\ACVQN1_reg/NET0131  & n26 ;
  assign n29 = \AX1_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n30 = ~n28 & ~n29 ;
  assign n31 = ~n27 & ~n30 ;
  assign n32 = ~\ACVQN2_reg/NET0131  & \AX2_reg/NET0131  ;
  assign n33 = ~\MRVQN0_reg/NET0131  & n32 ;
  assign n34 = ~n31 & ~n33 ;
  assign n35 = \AX2_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n36 = \ACVQN2_reg/NET0131  & ~n35 ;
  assign n37 = ~n34 & ~n36 ;
  assign n38 = \AX3_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n39 = \ACVQN3_reg/NET0131  & ~n38 ;
  assign n40 = ~n37 & n39 ;
  assign n42 = ~\ACVQN2_reg/NET0131  & ~\ACVQN3_reg/NET0131  ;
  assign n43 = \MRVQN0_reg/NET0131  & ~n42 ;
  assign n41 = \ACVQN2_reg/NET0131  & ~\AX2_reg/NET0131  ;
  assign n44 = \ACVQN3_reg/NET0131  & ~\AX3_reg/NET0131  ;
  assign n45 = ~n41 & ~n44 ;
  assign n46 = ~n43 & n45 ;
  assign n47 = ~n34 & n46 ;
  assign n48 = ~\ACVQN3_reg/NET0131  & n38 ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = ~n40 & n49 ;
  assign n51 = n37 & n48 ;
  assign n52 = ~\CT0_reg/NET0131  & ~\CT1_reg/NET0131  ;
  assign n53 = ~\CT2_reg/NET0131  & n52 ;
  assign n54 = ~n24 & ~n53 ;
  assign n55 = ~n51 & n54 ;
  assign n56 = ~n50 & n55 ;
  assign n57 = \ACVQN2_reg/NET0131  & ~n54 ;
  assign n58 = ~START_pad & ~n57 ;
  assign n59 = ~n56 & n58 ;
  assign n62 = n27 & ~n29 ;
  assign n63 = ~n31 & ~n62 ;
  assign n61 = \AX1_reg/NET0131  & n28 ;
  assign n64 = n54 & ~n61 ;
  assign n65 = ~n63 & n64 ;
  assign n60 = \ACVQN0_reg/NET0131  & ~n54 ;
  assign n66 = ~START_pad & ~n60 ;
  assign n67 = ~n65 & n66 ;
  assign n68 = \CT0_reg/NET0131  & ~n24 ;
  assign n69 = ~\CT1_reg/NET0131  & ~n68 ;
  assign n70 = ~START_pad & ~n21 ;
  assign n71 = ~n69 & n70 ;
  assign n72 = \AX0_reg/NET0131  & ~\MRVQN0_reg/NET0131  ;
  assign n73 = \ACVQN0_reg/NET0131  & ~n72 ;
  assign n74 = ~n26 & ~n73 ;
  assign n75 = n54 & ~n74 ;
  assign n77 = \B3_pad  & ~n24 ;
  assign n76 = ~\MRVQN3_reg/NET0131  & n24 ;
  assign n78 = ~n54 & ~n76 ;
  assign n79 = ~n77 & n78 ;
  assign n80 = ~n75 & ~n79 ;
  assign n81 = ~\B2_pad  & ~n24 ;
  assign n82 = \MRVQN2_reg/NET0131  & n24 ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = ~n54 & ~n83 ;
  assign n85 = \MRVQN3_reg/NET0131  & n54 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = ~\B0_pad  & ~n24 ;
  assign n88 = \MRVQN0_reg/NET0131  & n24 ;
  assign n89 = ~n87 & ~n88 ;
  assign n90 = ~n54 & ~n89 ;
  assign n91 = \MRVQN1_reg/NET0131  & n54 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = ~\B1_pad  & ~n24 ;
  assign n94 = \MRVQN1_reg/NET0131  & n24 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = ~n54 & ~n95 ;
  assign n97 = \MRVQN2_reg/NET0131  & n54 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = ~\CT2_reg/NET0131  & ~n21 ;
  assign n100 = ~START_pad & ~n22 ;
  assign n101 = ~n99 & n100 ;
  assign n102 = ~START_pad & ~n68 ;
  assign n105 = ~n31 & n36 ;
  assign n106 = ~n37 & ~n105 ;
  assign n104 = n31 & n33 ;
  assign n107 = n54 & ~n104 ;
  assign n108 = ~n106 & n107 ;
  assign n103 = \ACVQN1_reg/NET0131  & ~n54 ;
  assign n109 = ~START_pad & ~n103 ;
  assign n110 = ~n108 & n109 ;
  assign n112 = n49 & n54 ;
  assign n111 = \ACVQN3_reg/NET0131  & ~n54 ;
  assign n113 = ~START_pad & ~n111 ;
  assign n114 = ~n112 & n113 ;
  assign \ACVQN0_reg/P0001  = ~\ACVQN0_reg/NET0131  ;
  assign \ACVQN1_reg/P0001  = ~\ACVQN1_reg/NET0131  ;
  assign \ACVQN2_reg/P0001  = ~\ACVQN2_reg/NET0131  ;
  assign \ACVQN3_reg/P0001  = ~\ACVQN3_reg/NET0131  ;
  assign \CNTVCON2_pad  = ~n22 ;
  assign \MRVQN0_reg/P0001  = ~\MRVQN0_reg/NET0131  ;
  assign \P1_pad  = ~\MRVQN1_reg/NET0131  ;
  assign \P2_pad  = ~\MRVQN2_reg/NET0131  ;
  assign \P3_pad  = ~\MRVQN3_reg/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g12/_2_  = n24 ;
  assign \g25/_0_  = ~n59 ;
  assign \g29/_0_  = ~n67 ;
  assign \g614/_0_  = n71 ;
  assign \g621/_0_  = ~n80 ;
  assign \g623/_3_  = ~n86 ;
  assign \g624/_3_  = ~n92 ;
  assign \g625/_3_  = ~n98 ;
  assign \g631/_0_  = n101 ;
  assign \g635/_0_  = n102 ;
  assign \g658/_1_  = n22 ;
  assign \g765/_0_  = ~n110 ;
  assign \g775/_2_  = n53 ;
  assign \g782/_0_  = ~n114 ;
endmodule
