module top (\ccyc_addr_in[0]_pad , \ccyc_addr_in[11]_pad , \ccyc_addr_in[12]_pad , \ccyc_addr_in[13]_pad , \ccyc_addr_in[14]_pad , \ccyc_addr_in[15]_pad , \ccyc_addr_in[16]_pad , \ccyc_addr_in[17]_pad , \ccyc_addr_in[18]_pad , \ccyc_addr_in[19]_pad , \ccyc_addr_in[20]_pad , \ccyc_addr_in[21]_pad , \ccyc_addr_in[22]_pad , \ccyc_addr_in[23]_pad , \ccyc_addr_in[24]_pad , \ccyc_addr_in[25]_pad , \ccyc_addr_in[26]_pad , \ccyc_addr_in[27]_pad , \ccyc_addr_in[28]_pad , \ccyc_addr_in[29]_pad , \ccyc_addr_in[30]_pad , \ccyc_addr_in[31]_pad , \ccyc_addr_out[11]_pad , \ccyc_addr_out[12]_pad , \ccyc_addr_out[13]_pad , \ccyc_addr_out[14]_pad , \ccyc_addr_out[15]_pad , \ccyc_addr_out[16]_pad , \ccyc_addr_out[17]_pad , \ccyc_addr_out[18]_pad , \ccyc_addr_out[19]_pad , \ccyc_addr_out[20]_pad , \ccyc_addr_out[21]_pad , \ccyc_addr_out[22]_pad , \ccyc_addr_out[23]_pad , \ccyc_addr_out[24]_pad , \ccyc_addr_out[25]_pad , \ccyc_addr_out[26]_pad , \ccyc_addr_out[27]_pad , \ccyc_addr_out[28]_pad , \ccyc_addr_out[29]_pad , \ccyc_addr_out[30]_pad , \ccyc_addr_out[31]_pad );
	input \ccyc_addr_in[0]_pad  ;
	input \ccyc_addr_in[11]_pad  ;
	input \ccyc_addr_in[12]_pad  ;
	input \ccyc_addr_in[13]_pad  ;
	input \ccyc_addr_in[14]_pad  ;
	input \ccyc_addr_in[15]_pad  ;
	input \ccyc_addr_in[16]_pad  ;
	input \ccyc_addr_in[17]_pad  ;
	input \ccyc_addr_in[18]_pad  ;
	input \ccyc_addr_in[19]_pad  ;
	input \ccyc_addr_in[20]_pad  ;
	input \ccyc_addr_in[21]_pad  ;
	input \ccyc_addr_in[22]_pad  ;
	input \ccyc_addr_in[23]_pad  ;
	input \ccyc_addr_in[24]_pad  ;
	input \ccyc_addr_in[25]_pad  ;
	input \ccyc_addr_in[26]_pad  ;
	input \ccyc_addr_in[27]_pad  ;
	input \ccyc_addr_in[28]_pad  ;
	input \ccyc_addr_in[29]_pad  ;
	input \ccyc_addr_in[30]_pad  ;
	input \ccyc_addr_in[31]_pad  ;
	output \ccyc_addr_out[11]_pad  ;
	output \ccyc_addr_out[12]_pad  ;
	output \ccyc_addr_out[13]_pad  ;
	output \ccyc_addr_out[14]_pad  ;
	output \ccyc_addr_out[15]_pad  ;
	output \ccyc_addr_out[16]_pad  ;
	output \ccyc_addr_out[17]_pad  ;
	output \ccyc_addr_out[18]_pad  ;
	output \ccyc_addr_out[19]_pad  ;
	output \ccyc_addr_out[20]_pad  ;
	output \ccyc_addr_out[21]_pad  ;
	output \ccyc_addr_out[22]_pad  ;
	output \ccyc_addr_out[23]_pad  ;
	output \ccyc_addr_out[24]_pad  ;
	output \ccyc_addr_out[25]_pad  ;
	output \ccyc_addr_out[26]_pad  ;
	output \ccyc_addr_out[27]_pad  ;
	output \ccyc_addr_out[28]_pad  ;
	output \ccyc_addr_out[29]_pad  ;
	output \ccyc_addr_out[30]_pad  ;
	output \ccyc_addr_out[31]_pad  ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	LUT4 #(
		.INIT('h0001)
	) name0 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w24_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		_w25_
	);
	LUT3 #(
		.INIT('h98)
	) name2 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		_w24_,
		_w26_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		_w27_
	);
	LUT3 #(
		.INIT('h0b)
	) name4 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		\ccyc_addr_in[12]_pad ,
		_w28_
	);
	LUT3 #(
		.INIT('h0e)
	) name5 (
		\ccyc_addr_in[0]_pad ,
		_w24_,
		_w28_,
		_w29_
	);
	LUT4 #(
		.INIT('h0002)
	) name6 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[13]_pad ,
		_w31_
	);
	LUT3 #(
		.INIT('hf8)
	) name8 (
		_w25_,
		_w30_,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[14]_pad ,
		_w33_
	);
	LUT3 #(
		.INIT('hf8)
	) name10 (
		_w27_,
		_w30_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w35_
	);
	LUT4 #(
		.INIT('h0004)
	) name12 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w36_
	);
	LUT3 #(
		.INIT('hec)
	) name13 (
		_w25_,
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[16]_pad ,
		_w38_
	);
	LUT3 #(
		.INIT('hf8)
	) name15 (
		_w27_,
		_w36_,
		_w38_,
		_w39_
	);
	LUT4 #(
		.INIT('h0008)
	) name16 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[17]_pad ,
		_w41_
	);
	LUT3 #(
		.INIT('hf8)
	) name18 (
		_w25_,
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[18]_pad ,
		_w43_
	);
	LUT3 #(
		.INIT('hf8)
	) name20 (
		_w27_,
		_w40_,
		_w43_,
		_w44_
	);
	LUT4 #(
		.INIT('h0010)
	) name21 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[19]_pad ,
		_w46_
	);
	LUT3 #(
		.INIT('hf8)
	) name23 (
		_w25_,
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[20]_pad ,
		_w48_
	);
	LUT3 #(
		.INIT('hf8)
	) name25 (
		_w27_,
		_w45_,
		_w48_,
		_w49_
	);
	LUT4 #(
		.INIT('h0020)
	) name26 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[21]_pad ,
		_w51_
	);
	LUT3 #(
		.INIT('hf8)
	) name28 (
		_w25_,
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[22]_pad ,
		_w53_
	);
	LUT3 #(
		.INIT('hf8)
	) name30 (
		_w27_,
		_w50_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[23]_pad ,
		_w55_
	);
	LUT4 #(
		.INIT('h0040)
	) name32 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w56_
	);
	LUT3 #(
		.INIT('hec)
	) name33 (
		_w25_,
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[24]_pad ,
		_w58_
	);
	LUT3 #(
		.INIT('hf8)
	) name35 (
		_w27_,
		_w56_,
		_w58_,
		_w59_
	);
	LUT4 #(
		.INIT('h0080)
	) name36 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[25]_pad ,
		_w61_
	);
	LUT3 #(
		.INIT('hf8)
	) name38 (
		_w25_,
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[26]_pad ,
		_w63_
	);
	LUT3 #(
		.INIT('hf8)
	) name40 (
		_w27_,
		_w60_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w65_
	);
	LUT4 #(
		.INIT('h0100)
	) name42 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[27]_pad ,
		_w67_
	);
	LUT3 #(
		.INIT('hf8)
	) name44 (
		_w25_,
		_w66_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[28]_pad ,
		_w69_
	);
	LUT3 #(
		.INIT('hf8)
	) name46 (
		_w27_,
		_w66_,
		_w69_,
		_w70_
	);
	LUT4 #(
		.INIT('h0200)
	) name47 (
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		\ccyc_addr_in[14]_pad ,
		\ccyc_addr_in[15]_pad ,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[29]_pad ,
		_w72_
	);
	LUT3 #(
		.INIT('hf8)
	) name49 (
		_w25_,
		_w71_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[30]_pad ,
		_w74_
	);
	LUT3 #(
		.INIT('hf8)
	) name51 (
		_w27_,
		_w71_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[31]_pad ,
		_w76_
	);
	LUT4 #(
		.INIT('h0100)
	) name53 (
		\ccyc_addr_in[0]_pad ,
		\ccyc_addr_in[11]_pad ,
		\ccyc_addr_in[12]_pad ,
		\ccyc_addr_in[13]_pad ,
		_w77_
	);
	LUT3 #(
		.INIT('hec)
	) name54 (
		_w65_,
		_w76_,
		_w77_,
		_w78_
	);
	assign \ccyc_addr_out[11]_pad  = _w26_ ;
	assign \ccyc_addr_out[12]_pad  = _w29_ ;
	assign \ccyc_addr_out[13]_pad  = _w32_ ;
	assign \ccyc_addr_out[14]_pad  = _w34_ ;
	assign \ccyc_addr_out[15]_pad  = _w37_ ;
	assign \ccyc_addr_out[16]_pad  = _w39_ ;
	assign \ccyc_addr_out[17]_pad  = _w42_ ;
	assign \ccyc_addr_out[18]_pad  = _w44_ ;
	assign \ccyc_addr_out[19]_pad  = _w47_ ;
	assign \ccyc_addr_out[20]_pad  = _w49_ ;
	assign \ccyc_addr_out[21]_pad  = _w52_ ;
	assign \ccyc_addr_out[22]_pad  = _w54_ ;
	assign \ccyc_addr_out[23]_pad  = _w57_ ;
	assign \ccyc_addr_out[24]_pad  = _w59_ ;
	assign \ccyc_addr_out[25]_pad  = _w62_ ;
	assign \ccyc_addr_out[26]_pad  = _w64_ ;
	assign \ccyc_addr_out[27]_pad  = _w68_ ;
	assign \ccyc_addr_out[28]_pad  = _w70_ ;
	assign \ccyc_addr_out[29]_pad  = _w73_ ;
	assign \ccyc_addr_out[30]_pad  = _w75_ ;
	assign \ccyc_addr_out[31]_pad  = _w78_ ;
endmodule;