module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	output f_pad ;
	output g_pad ;
	output h_pad ;
	output i_pad ;
	output j_pad ;
	output k_pad ;
	output l_pad ;
	output m_pad ;
	output n_pad ;
	output o_pad ;
	output p_pad ;
	output q_pad ;
	output r_pad ;
	output s_pad ;
	output t_pad ;
	output u_pad ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w7_ ;
	wire _w8_ ;
	wire _w9_ ;
	wire _w10_ ;
	wire _w11_ ;
	wire _w12_ ;
	wire _w13_ ;
	wire _w14_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		a_pad,
		e_pad,
		_w7_
	);
	LUT3 #(
		.INIT('h80)
	) name1 (
		b_pad,
		c_pad,
		d_pad,
		_w8_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w7_,
		_w8_,
		_w9_
	);
	LUT3 #(
		.INIT('h08)
	) name3 (
		b_pad,
		c_pad,
		d_pad,
		_w10_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		_w7_,
		_w10_,
		_w11_
	);
	LUT3 #(
		.INIT('h20)
	) name5 (
		b_pad,
		c_pad,
		d_pad,
		_w12_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w7_,
		_w12_,
		_w13_
	);
	LUT3 #(
		.INIT('h02)
	) name7 (
		b_pad,
		c_pad,
		d_pad,
		_w14_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w7_,
		_w14_,
		_w15_
	);
	LUT3 #(
		.INIT('h40)
	) name9 (
		b_pad,
		c_pad,
		d_pad,
		_w16_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w7_,
		_w16_,
		_w17_
	);
	LUT3 #(
		.INIT('h04)
	) name11 (
		b_pad,
		c_pad,
		d_pad,
		_w18_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w7_,
		_w18_,
		_w19_
	);
	LUT3 #(
		.INIT('h10)
	) name13 (
		b_pad,
		c_pad,
		d_pad,
		_w20_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w7_,
		_w20_,
		_w21_
	);
	LUT3 #(
		.INIT('h01)
	) name15 (
		b_pad,
		c_pad,
		d_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w7_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		a_pad,
		e_pad,
		_w24_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w8_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w10_,
		_w24_,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w12_,
		_w24_,
		_w27_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w14_,
		_w24_,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w16_,
		_w24_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w18_,
		_w24_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w20_,
		_w24_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w22_,
		_w24_,
		_w32_
	);
	assign f_pad = _w9_ ;
	assign g_pad = _w11_ ;
	assign h_pad = _w13_ ;
	assign i_pad = _w15_ ;
	assign j_pad = _w17_ ;
	assign k_pad = _w19_ ;
	assign l_pad = _w21_ ;
	assign m_pad = _w23_ ;
	assign n_pad = _w25_ ;
	assign o_pad = _w26_ ;
	assign p_pad = _w27_ ;
	assign q_pad = _w28_ ;
	assign r_pad = _w29_ ;
	assign s_pad = _w30_ ;
	assign t_pad = _w31_ ;
	assign u_pad = _w32_ ;
endmodule;