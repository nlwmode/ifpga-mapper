module top (\a0_pad , a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \b0_pad , \c0_pad , \d0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad );
	input \a0_pad  ;
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \d0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		i_pad,
		j_pad,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		k_pad,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		t_pad,
		u_pad,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		v_pad,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		w_pad,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		x_pad,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		y_pad,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		z_pad,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\a0_pad ,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w29_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		a_pad,
		i_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		b_pad,
		i_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		c_pad,
		i_pad,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		d_pad,
		i_pad,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		e_pad,
		i_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		f_pad,
		i_pad,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		g_pad,
		i_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		h_pad,
		i_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		l_pad,
		_w37_,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		t_pad,
		_w29_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w38_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w46_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		t_pad,
		u_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w30_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		m_pad,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w37_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w29_,
		_w51_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w39_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w53_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		v_pad,
		_w30_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w31_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		n_pad,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w37_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w29_,
		_w58_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w40_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w60_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		w_pad,
		_w31_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w32_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		o_pad,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w37_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w29_,
		_w65_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w41_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w67_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		x_pad,
		_w32_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w33_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		p_pad,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w37_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w29_,
		_w72_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w42_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w74_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		y_pad,
		_w33_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w34_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		q_pad,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w37_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w29_,
		_w79_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w43_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w81_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		r_pad,
		_w37_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		z_pad,
		_w34_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w29_,
		_w35_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w44_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w85_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		s_pad,
		_w36_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\a0_pad ,
		_w35_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		_w29_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w91_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w45_,
		_w94_,
		_w95_
	);
	assign \b0_pad  = _w37_ ;
	assign \c0_pad  = _w38_ ;
	assign \d0_pad  = _w39_ ;
	assign \e0_pad  = _w40_ ;
	assign \f0_pad  = _w41_ ;
	assign \g0_pad  = _w42_ ;
	assign \h0_pad  = _w43_ ;
	assign \i0_pad  = _w44_ ;
	assign \j0_pad  = _w45_ ;
	assign \k0_pad  = _w49_ ;
	assign \l0_pad  = _w56_ ;
	assign \m0_pad  = _w63_ ;
	assign \n0_pad  = _w70_ ;
	assign \o0_pad  = _w77_ ;
	assign \p0_pad  = _w84_ ;
	assign \q0_pad  = _w90_ ;
	assign \r0_pad  = _w95_ ;
endmodule;