module top (\B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] , \B[8] , \B[9] , \B[10] , \M[0] , \M[1] , \M[2] , \M[3] , \E[0] , \E[1] , \E[2] );
	input \B[0]  ;
	input \B[1]  ;
	input \B[2]  ;
	input \B[3]  ;
	input \B[4]  ;
	input \B[5]  ;
	input \B[6]  ;
	input \B[7]  ;
	input \B[8]  ;
	input \B[9]  ;
	input \B[10]  ;
	output \M[0]  ;
	output \M[1]  ;
	output \M[2]  ;
	output \M[3]  ;
	output \E[0]  ;
	output \E[1]  ;
	output \E[2]  ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w14_ ;
	wire _w13_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\B[6] ,
		\B[7] ,
		_w13_
	);
	LUT3 #(
		.INIT('hea)
	) name1 (
		\B[6] ,
		\B[7] ,
		\B[10] ,
		_w14_
	);
	LUT3 #(
		.INIT('h10)
	) name2 (
		\B[6] ,
		\B[7] ,
		\B[10] ,
		_w15_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\B[7] ,
		\B[10] ,
		_w16_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\B[2] ,
		\B[3] ,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\B[2] ,
		\B[3] ,
		_w18_
	);
	LUT2 #(
		.INIT('h6)
	) name6 (
		\B[2] ,
		\B[3] ,
		_w19_
	);
	LUT3 #(
		.INIT('h01)
	) name7 (
		\B[7] ,
		\B[8] ,
		\B[9] ,
		_w20_
	);
	LUT3 #(
		.INIT('h15)
	) name8 (
		_w16_,
		_w19_,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\B[6] ,
		\B[7] ,
		_w22_
	);
	LUT3 #(
		.INIT('h40)
	) name10 (
		\B[6] ,
		\B[7] ,
		\B[10] ,
		_w23_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\B[8] ,
		\B[10] ,
		_w24_
	);
	LUT3 #(
		.INIT('h80)
	) name12 (
		\B[8] ,
		\B[9] ,
		\B[10] ,
		_w25_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w23_,
		_w25_,
		_w26_
	);
	LUT3 #(
		.INIT('h02)
	) name14 (
		\B[10] ,
		_w22_,
		_w25_,
		_w27_
	);
	LUT3 #(
		.INIT('h15)
	) name15 (
		_w15_,
		_w21_,
		_w27_,
		_w28_
	);
	LUT4 #(
		.INIT('h0040)
	) name16 (
		\B[3] ,
		\B[4] ,
		\B[7] ,
		\B[8] ,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\B[9] ,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\B[4] ,
		\B[7] ,
		_w31_
	);
	LUT4 #(
		.INIT('h0020)
	) name19 (
		\B[1] ,
		\B[2] ,
		\B[5] ,
		\B[7] ,
		_w32_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\B[3] ,
		\B[8] ,
		_w33_
	);
	LUT3 #(
		.INIT('h02)
	) name21 (
		\B[3] ,
		\B[8] ,
		\B[9] ,
		_w34_
	);
	LUT3 #(
		.INIT('he0)
	) name22 (
		_w31_,
		_w32_,
		_w34_,
		_w35_
	);
	LUT4 #(
		.INIT('h8a80)
	) name23 (
		\B[0] ,
		\B[1] ,
		\B[4] ,
		\B[8] ,
		_w36_
	);
	LUT3 #(
		.INIT('h15)
	) name24 (
		\B[0] ,
		\B[1] ,
		\B[4] ,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\B[4] ,
		\B[8] ,
		_w38_
	);
	LUT3 #(
		.INIT('h13)
	) name26 (
		\B[4] ,
		\B[5] ,
		\B[8] ,
		_w39_
	);
	LUT4 #(
		.INIT('hfd00)
	) name27 (
		_w13_,
		_w36_,
		_w37_,
		_w39_,
		_w40_
	);
	LUT4 #(
		.INIT('h0073)
	) name28 (
		\B[4] ,
		\B[5] ,
		\B[8] ,
		\B[9] ,
		_w41_
	);
	LUT4 #(
		.INIT('h1011)
	) name29 (
		_w30_,
		_w35_,
		_w40_,
		_w41_,
		_w42_
	);
	LUT3 #(
		.INIT('h2a)
	) name30 (
		_w14_,
		_w21_,
		_w26_,
		_w43_
	);
	LUT3 #(
		.INIT('h40)
	) name31 (
		\B[5] ,
		\B[6] ,
		\B[9] ,
		_w44_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\B[5] ,
		\B[6] ,
		_w45_
	);
	LUT4 #(
		.INIT('h2022)
	) name33 (
		\B[1] ,
		\B[2] ,
		\B[4] ,
		\B[7] ,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\B[3] ,
		\B[4] ,
		_w47_
	);
	LUT3 #(
		.INIT('h37)
	) name35 (
		\B[3] ,
		\B[4] ,
		\B[8] ,
		_w48_
	);
	LUT4 #(
		.INIT('h0004)
	) name36 (
		\B[1] ,
		\B[2] ,
		\B[7] ,
		\B[8] ,
		_w49_
	);
	LUT4 #(
		.INIT('h0015)
	) name37 (
		\B[9] ,
		_w46_,
		_w48_,
		_w49_,
		_w50_
	);
	LUT3 #(
		.INIT('h51)
	) name38 (
		_w44_,
		_w45_,
		_w50_,
		_w51_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name39 (
		_w28_,
		_w42_,
		_w43_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\B[7] ,
		\B[10] ,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\B[6] ,
		\B[9] ,
		_w54_
	);
	LUT3 #(
		.INIT('h80)
	) name42 (
		\B[2] ,
		\B[3] ,
		\B[4] ,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT3 #(
		.INIT('h04)
	) name44 (
		\B[4] ,
		\B[6] ,
		\B[9] ,
		_w57_
	);
	LUT3 #(
		.INIT('h04)
	) name45 (
		\B[3] ,
		\B[5] ,
		\B[6] ,
		_w58_
	);
	LUT3 #(
		.INIT('h54)
	) name46 (
		\B[2] ,
		_w57_,
		_w58_,
		_w59_
	);
	LUT3 #(
		.INIT('h04)
	) name47 (
		\B[1] ,
		\B[5] ,
		\B[6] ,
		_w60_
	);
	LUT4 #(
		.INIT('h2223)
	) name48 (
		\B[3] ,
		\B[10] ,
		_w57_,
		_w60_,
		_w61_
	);
	LUT4 #(
		.INIT('h5455)
	) name49 (
		_w53_,
		_w56_,
		_w59_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\B[6] ,
		\B[7] ,
		_w63_
	);
	LUT3 #(
		.INIT('h07)
	) name51 (
		\B[6] ,
		\B[7] ,
		\B[8] ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w62_,
		_w64_,
		_w65_
	);
	LUT3 #(
		.INIT('h08)
	) name53 (
		\B[6] ,
		\B[7] ,
		\B[9] ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w24_,
		_w66_,
		_w67_
	);
	LUT3 #(
		.INIT('h4c)
	) name55 (
		\B[8] ,
		\B[10] ,
		_w66_,
		_w68_
	);
	LUT3 #(
		.INIT('h10)
	) name56 (
		\B[5] ,
		\B[7] ,
		\B[9] ,
		_w69_
	);
	LUT3 #(
		.INIT('h70)
	) name57 (
		\B[3] ,
		\B[4] ,
		\B[7] ,
		_w70_
	);
	LUT3 #(
		.INIT('h01)
	) name58 (
		\B[5] ,
		\B[8] ,
		\B[9] ,
		_w71_
	);
	LUT3 #(
		.INIT('h15)
	) name59 (
		_w69_,
		_w70_,
		_w71_,
		_w72_
	);
	LUT3 #(
		.INIT('h2a)
	) name60 (
		\B[0] ,
		\B[1] ,
		\B[2] ,
		_w73_
	);
	LUT4 #(
		.INIT('h00b0)
	) name61 (
		\B[0] ,
		\B[2] ,
		\B[4] ,
		\B[7] ,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\B[8] ,
		\B[9] ,
		_w76_
	);
	LUT4 #(
		.INIT('hfac8)
	) name64 (
		\B[2] ,
		\B[4] ,
		\B[7] ,
		\B[9] ,
		_w77_
	);
	LUT3 #(
		.INIT('h32)
	) name65 (
		\B[1] ,
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\B[5] ,
		\B[6] ,
		_w79_
	);
	LUT4 #(
		.INIT('h20aa)
	) name67 (
		_w72_,
		_w75_,
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\B[4] ,
		\B[6] ,
		_w81_
	);
	LUT4 #(
		.INIT('h0010)
	) name69 (
		\B[4] ,
		\B[6] ,
		\B[8] ,
		\B[9] ,
		_w82_
	);
	LUT3 #(
		.INIT('h10)
	) name70 (
		\B[6] ,
		\B[7] ,
		\B[9] ,
		_w83_
	);
	LUT3 #(
		.INIT('h01)
	) name71 (
		\B[5] ,
		_w82_,
		_w83_,
		_w84_
	);
	LUT4 #(
		.INIT('h888a)
	) name72 (
		\B[3] ,
		\B[4] ,
		\B[6] ,
		\B[7] ,
		_w85_
	);
	LUT3 #(
		.INIT('ha8)
	) name73 (
		\B[4] ,
		\B[8] ,
		\B[9] ,
		_w86_
	);
	LUT3 #(
		.INIT('h07)
	) name74 (
		\B[1] ,
		\B[2] ,
		\B[7] ,
		_w87_
	);
	LUT3 #(
		.INIT('h02)
	) name75 (
		_w85_,
		_w86_,
		_w87_,
		_w88_
	);
	LUT3 #(
		.INIT('ha8)
	) name76 (
		\B[6] ,
		\B[8] ,
		\B[9] ,
		_w89_
	);
	LUT3 #(
		.INIT('hca)
	) name77 (
		\B[4] ,
		\B[7] ,
		\B[9] ,
		_w90_
	);
	LUT4 #(
		.INIT('h0111)
	) name78 (
		_w82_,
		_w83_,
		_w89_,
		_w90_,
		_w91_
	);
	LUT4 #(
		.INIT('h4544)
	) name79 (
		_w67_,
		_w84_,
		_w88_,
		_w91_,
		_w92_
	);
	LUT3 #(
		.INIT('h15)
	) name80 (
		_w68_,
		_w80_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w65_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\B[4] ,
		\B[5] ,
		_w95_
	);
	LUT4 #(
		.INIT('h0777)
	) name83 (
		\B[4] ,
		\B[5] ,
		\B[6] ,
		\B[7] ,
		_w96_
	);
	LUT4 #(
		.INIT('h0c50)
	) name84 (
		\B[2] ,
		\B[3] ,
		\B[6] ,
		\B[7] ,
		_w97_
	);
	LUT4 #(
		.INIT('hfd5d)
	) name85 (
		\B[8] ,
		_w63_,
		_w95_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\B[9] ,
		\B[10] ,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\B[5] ,
		\B[6] ,
		_w100_
	);
	LUT4 #(
		.INIT('h0080)
	) name88 (
		\B[4] ,
		\B[5] ,
		\B[6] ,
		\B[7] ,
		_w101_
	);
	LUT4 #(
		.INIT('hf07f)
	) name89 (
		\B[4] ,
		\B[5] ,
		\B[6] ,
		\B[7] ,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		\B[8] ,
		\B[10] ,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w102_,
		_w103_,
		_w104_
	);
	LUT3 #(
		.INIT('h07)
	) name92 (
		_w98_,
		_w99_,
		_w104_,
		_w105_
	);
	LUT3 #(
		.INIT('h40)
	) name93 (
		\B[3] ,
		\B[4] ,
		\B[5] ,
		_w106_
	);
	LUT4 #(
		.INIT('h0040)
	) name94 (
		\B[2] ,
		\B[3] ,
		\B[4] ,
		\B[6] ,
		_w107_
	);
	LUT3 #(
		.INIT('h54)
	) name95 (
		\B[7] ,
		_w106_,
		_w107_,
		_w108_
	);
	LUT4 #(
		.INIT('h0020)
	) name96 (
		\B[0] ,
		\B[3] ,
		\B[4] ,
		\B[6] ,
		_w109_
	);
	LUT3 #(
		.INIT('h20)
	) name97 (
		\B[3] ,
		\B[4] ,
		\B[5] ,
		_w110_
	);
	LUT3 #(
		.INIT('ha8)
	) name98 (
		\B[1] ,
		_w109_,
		_w110_,
		_w111_
	);
	LUT4 #(
		.INIT('h7000)
	) name99 (
		\B[0] ,
		\B[1] ,
		\B[3] ,
		\B[4] ,
		_w112_
	);
	LUT3 #(
		.INIT('h54)
	) name100 (
		\B[5] ,
		_w81_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\B[2] ,
		\B[7] ,
		_w114_
	);
	LUT4 #(
		.INIT('h0155)
	) name102 (
		_w108_,
		_w111_,
		_w113_,
		_w114_,
		_w115_
	);
	LUT3 #(
		.INIT('h31)
	) name103 (
		_w95_,
		_w96_,
		_w97_,
		_w116_
	);
	LUT4 #(
		.INIT('h7000)
	) name104 (
		\B[3] ,
		\B[4] ,
		\B[5] ,
		\B[6] ,
		_w117_
	);
	LUT4 #(
		.INIT('hf3af)
	) name105 (
		\B[1] ,
		\B[2] ,
		\B[5] ,
		\B[6] ,
		_w118_
	);
	LUT3 #(
		.INIT('h31)
	) name106 (
		_w47_,
		_w117_,
		_w118_,
		_w119_
	);
	LUT3 #(
		.INIT('h10)
	) name107 (
		_w104_,
		_w116_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\B[9] ,
		\B[10] ,
		_w121_
	);
	LUT4 #(
		.INIT('h7000)
	) name109 (
		\B[5] ,
		\B[7] ,
		\B[8] ,
		\B[9] ,
		_w122_
	);
	LUT4 #(
		.INIT('h13df)
	) name110 (
		\B[5] ,
		\B[8] ,
		\B[9] ,
		\B[10] ,
		_w123_
	);
	LUT4 #(
		.INIT('h0301)
	) name111 (
		_w63_,
		_w121_,
		_w122_,
		_w123_,
		_w124_
	);
	LUT4 #(
		.INIT('h15ff)
	) name112 (
		_w105_,
		_w115_,
		_w120_,
		_w124_,
		_w125_
	);
	LUT3 #(
		.INIT('h01)
	) name113 (
		\B[5] ,
		\B[7] ,
		\B[8] ,
		_w126_
	);
	LUT4 #(
		.INIT('h4000)
	) name114 (
		\B[2] ,
		\B[5] ,
		\B[6] ,
		\B[7] ,
		_w127_
	);
	LUT4 #(
		.INIT('h153f)
	) name115 (
		_w38_,
		_w81_,
		_w126_,
		_w127_,
		_w128_
	);
	LUT3 #(
		.INIT('h01)
	) name116 (
		\B[3] ,
		\B[9] ,
		\B[10] ,
		_w129_
	);
	LUT2 #(
		.INIT('hb)
	) name117 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT4 #(
		.INIT('h8000)
	) name118 (
		\B[5] ,
		\B[6] ,
		\B[7] ,
		\B[8] ,
		_w131_
	);
	LUT3 #(
		.INIT('h02)
	) name119 (
		\B[9] ,
		\B[10] ,
		_w131_,
		_w132_
	);
	LUT4 #(
		.INIT('he000)
	) name120 (
		\B[2] ,
		\B[3] ,
		\B[4] ,
		\B[5] ,
		_w133_
	);
	LUT4 #(
		.INIT('h0008)
	) name121 (
		\B[6] ,
		\B[7] ,
		\B[9] ,
		\B[10] ,
		_w134_
	);
	LUT3 #(
		.INIT('h40)
	) name122 (
		_w33_,
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w132_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\B[8] ,
		\B[10] ,
		_w137_
	);
	LUT4 #(
		.INIT('h0073)
	) name125 (
		\B[3] ,
		\B[4] ,
		\B[5] ,
		\B[6] ,
		_w138_
	);
	LUT4 #(
		.INIT('h0008)
	) name126 (
		\B[0] ,
		\B[1] ,
		\B[5] ,
		\B[6] ,
		_w139_
	);
	LUT3 #(
		.INIT('ha8)
	) name127 (
		_w18_,
		_w101_,
		_w139_,
		_w140_
	);
	LUT4 #(
		.INIT('h008f)
	) name128 (
		\B[1] ,
		\B[2] ,
		\B[5] ,
		\B[7] ,
		_w141_
	);
	LUT3 #(
		.INIT('h0b)
	) name129 (
		_w70_,
		_w100_,
		_w141_,
		_w142_
	);
	LUT4 #(
		.INIT('haaa8)
	) name130 (
		_w137_,
		_w138_,
		_w140_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w136_,
		_w143_,
		_w144_
	);
	LUT4 #(
		.INIT('h8000)
	) name132 (
		\B[0] ,
		\B[1] ,
		\B[2] ,
		\B[3] ,
		_w145_
	);
	LUT4 #(
		.INIT('h23af)
	) name133 (
		_w17_,
		_w126_,
		_w131_,
		_w145_,
		_w146_
	);
	LUT4 #(
		.INIT('h000e)
	) name134 (
		\B[5] ,
		\B[6] ,
		\B[7] ,
		\B[8] ,
		_w147_
	);
	LUT4 #(
		.INIT('h7f33)
	) name135 (
		_w55_,
		_w99_,
		_w100_,
		_w147_,
		_w148_
	);
	LUT3 #(
		.INIT('hf2)
	) name136 (
		\B[4] ,
		_w146_,
		_w148_,
		_w149_
	);
	LUT4 #(
		.INIT('h0001)
	) name137 (
		\B[7] ,
		\B[8] ,
		\B[9] ,
		\B[10] ,
		_w150_
	);
	LUT3 #(
		.INIT('h8f)
	) name138 (
		_w55_,
		_w100_,
		_w150_,
		_w151_
	);
	assign \M[0]  = _w52_ ;
	assign \M[1]  = _w94_ ;
	assign \M[2]  = _w125_ ;
	assign \M[3]  = _w130_ ;
	assign \E[0]  = _w144_ ;
	assign \E[1]  = _w149_ ;
	assign \E[2]  = _w151_ ;
endmodule;