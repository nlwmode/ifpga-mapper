module top( \v0_pad  , \v10_reg/NET0131  , \v11_reg/NET0131  , \v12_reg/NET0131  , \v1_pad  , \v2_pad  , \v3_pad  , \v4_pad  , \v5_pad  , \v6_pad  , \v7_reg/NET0131  , \v8_reg/NET0131  , \v9_reg/NET0131  , \_al_n0  , \_al_n1  , \g528/_2_  , \g534/_0_  , \g535/_0_  , \g537/_0_  , \g560/_3_  , \g722/_0_  , \g754/_0_  , \v13_D_10_pad  , \v13_D_11_pad  , \v13_D_12_pad  , \v13_D_6_pad  , \v13_D_7_pad  , \v13_D_9_pad  );
  input \v0_pad  ;
  input \v10_reg/NET0131  ;
  input \v11_reg/NET0131  ;
  input \v12_reg/NET0131  ;
  input \v1_pad  ;
  input \v2_pad  ;
  input \v3_pad  ;
  input \v4_pad  ;
  input \v5_pad  ;
  input \v6_pad  ;
  input \v7_reg/NET0131  ;
  input \v8_reg/NET0131  ;
  input \v9_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g528/_2_  ;
  output \g534/_0_  ;
  output \g535/_0_  ;
  output \g537/_0_  ;
  output \g560/_3_  ;
  output \g722/_0_  ;
  output \g754/_0_  ;
  output \v13_D_10_pad  ;
  output \v13_D_11_pad  ;
  output \v13_D_12_pad  ;
  output \v13_D_6_pad  ;
  output \v13_D_7_pad  ;
  output \v13_D_9_pad  ;
  wire n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 ;
  assign n14 = ~\v11_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n15 = ~\v5_pad  & \v9_reg/NET0131  ;
  assign n16 = n14 & n15 ;
  assign n17 = \v10_reg/NET0131  & ~n16 ;
  assign n18 = ~\v7_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n19 = ~\v0_pad  & n18 ;
  assign n20 = ~n17 & n19 ;
  assign n21 = \v1_pad  & n18 ;
  assign n22 = ~\v10_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n23 = \v0_pad  & ~\v11_reg/NET0131  ;
  assign n24 = ~\v12_reg/NET0131  & n23 ;
  assign n25 = ~n22 & ~n24 ;
  assign n26 = n21 & ~n25 ;
  assign n27 = ~\v12_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n28 = ~\v0_pad  & ~\v10_reg/NET0131  ;
  assign n29 = n27 & n28 ;
  assign n30 = ~\v12_reg/NET0131  & \v1_pad  ;
  assign n31 = n22 & n30 ;
  assign n32 = ~n29 & ~n31 ;
  assign n33 = ~n26 & n32 ;
  assign n34 = ~n20 & n33 ;
  assign n35 = \v10_reg/NET0131  & n18 ;
  assign n36 = ~\v11_reg/NET0131  & ~\v5_pad  ;
  assign n37 = n30 & n36 ;
  assign n38 = n35 & n37 ;
  assign n39 = ~n31 & ~n38 ;
  assign n40 = \v10_reg/NET0131  & ~n14 ;
  assign n41 = \v1_pad  & ~\v9_reg/NET0131  ;
  assign n42 = \v0_pad  & ~n41 ;
  assign n43 = n18 & ~n42 ;
  assign n44 = ~n40 & n43 ;
  assign n45 = ~n29 & ~n44 ;
  assign n46 = n39 & n45 ;
  assign n47 = \v11_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n48 = \v12_reg/NET0131  & n47 ;
  assign n49 = ~\v7_reg/NET0131  & n48 ;
  assign n50 = \v2_pad  & n14 ;
  assign n51 = \v3_pad  & \v8_reg/NET0131  ;
  assign n52 = ~\v7_reg/NET0131  & n51 ;
  assign n53 = n50 & n52 ;
  assign n54 = ~n49 & ~n53 ;
  assign n55 = \v11_reg/NET0131  & \v7_reg/NET0131  ;
  assign n56 = ~\v12_reg/NET0131  & \v8_reg/NET0131  ;
  assign n57 = n55 & n56 ;
  assign n58 = n54 & ~n57 ;
  assign n59 = ~\v10_reg/NET0131  & ~\v1_pad  ;
  assign n60 = \v0_pad  & ~\v9_reg/NET0131  ;
  assign n61 = n59 & n60 ;
  assign n62 = ~n58 & n61 ;
  assign n63 = ~\v12_reg/NET0131  & n61 ;
  assign n64 = ~\v11_reg/NET0131  & ~\v3_pad  ;
  assign n65 = ~\v4_pad  & \v8_reg/NET0131  ;
  assign n66 = n64 & n65 ;
  assign n67 = \v7_reg/NET0131  & \v8_reg/NET0131  ;
  assign n68 = \v11_reg/NET0131  & ~n67 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = n63 & ~n69 ;
  assign n71 = ~\v11_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n72 = ~\v12_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n73 = n71 & n72 ;
  assign n74 = \v10_reg/NET0131  & ~\v6_pad  ;
  assign n75 = n60 & n74 ;
  assign n76 = n73 & n75 ;
  assign n77 = \v3_pad  & n67 ;
  assign n78 = ~\v11_reg/NET0131  & n77 ;
  assign n79 = \v2_pad  & ~\v8_reg/NET0131  ;
  assign n80 = ~\v7_reg/NET0131  & ~n79 ;
  assign n81 = ~\v11_reg/NET0131  & \v4_pad  ;
  assign n82 = ~n80 & n81 ;
  assign n83 = ~n78 & ~n82 ;
  assign n84 = ~\v7_reg/NET0131  & ~n14 ;
  assign n85 = ~n47 & n84 ;
  assign n86 = \v5_pad  & \v7_reg/NET0131  ;
  assign n87 = n47 & n86 ;
  assign n88 = ~\v2_pad  & ~\v7_reg/NET0131  ;
  assign n89 = n51 & n88 ;
  assign n90 = ~n87 & ~n89 ;
  assign n91 = ~n85 & n90 ;
  assign n92 = n83 & n91 ;
  assign n93 = ~\v8_reg/NET0131  & n71 ;
  assign n94 = \v12_reg/NET0131  & ~n93 ;
  assign n95 = n61 & ~n94 ;
  assign n96 = ~n92 & n95 ;
  assign n97 = ~\v7_reg/NET0131  & ~n66 ;
  assign n98 = ~\v12_reg/NET0131  & ~n97 ;
  assign n99 = n14 & n79 ;
  assign n100 = \v12_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n101 = n47 & n100 ;
  assign n102 = ~\v5_pad  & n101 ;
  assign n103 = ~n99 & ~n102 ;
  assign n104 = ~n98 & n103 ;
  assign n105 = n61 & ~n104 ;
  assign n106 = \v0_pad  & \v5_pad  ;
  assign n107 = \v10_reg/NET0131  & ~n106 ;
  assign n108 = \v9_reg/NET0131  & n14 ;
  assign n109 = n21 & n108 ;
  assign n110 = ~n107 & n109 ;
  assign n111 = ~n18 & ~n27 ;
  assign n112 = n28 & ~n111 ;
  assign n113 = \v9_reg/NET0131  & ~n112 ;
  assign n114 = \v12_reg/NET0131  & ~n18 ;
  assign n115 = \v1_pad  & ~n114 ;
  assign n116 = ~\v10_reg/NET0131  & n115 ;
  assign n117 = ~\v4_pad  & n64 ;
  assign n118 = ~n55 & ~n117 ;
  assign n119 = ~\v10_reg/NET0131  & n56 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = ~n116 & ~n120 ;
  assign n122 = n24 & n35 ;
  assign n123 = ~n112 & ~n122 ;
  assign n124 = n121 & n123 ;
  assign n125 = ~n113 & ~n124 ;
  assign n126 = ~\v0_pad  & \v10_reg/NET0131  ;
  assign n127 = \v5_pad  & \v9_reg/NET0131  ;
  assign n128 = n126 & n127 ;
  assign n129 = n73 & n128 ;
  assign n130 = \v5_pad  & n101 ;
  assign n131 = n61 & n130 ;
  assign n132 = ~\v3_pad  & \v8_reg/NET0131  ;
  assign n133 = ~n88 & ~n132 ;
  assign n134 = \v4_pad  & \v7_reg/NET0131  ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = n14 & n61 ;
  assign n137 = ~n135 & n136 ;
  assign n138 = ~n131 & ~n137 ;
  assign n139 = \v7_reg/NET0131  & n47 ;
  assign n140 = ~n66 & ~n139 ;
  assign n141 = n63 & ~n140 ;
  assign n142 = \v0_pad  & \v10_reg/NET0131  ;
  assign n143 = ~\v8_reg/NET0131  & n142 ;
  assign n144 = \v4_pad  & n59 ;
  assign n145 = n132 & n144 ;
  assign n146 = ~n143 & ~n145 ;
  assign n147 = n27 & n71 ;
  assign n148 = ~n146 & n147 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g528/_2_  = ~n34 ;
  assign \g534/_0_  = ~n46 ;
  assign \g535/_0_  = n62 ;
  assign \g537/_0_  = n70 ;
  assign \g560/_3_  = n76 ;
  assign \g722/_0_  = n96 ;
  assign \g754/_0_  = n105 ;
  assign \v13_D_10_pad  = n110 ;
  assign \v13_D_11_pad  = n125 ;
  assign \v13_D_12_pad  = n129 ;
  assign \v13_D_6_pad  = ~n138 ;
  assign \v13_D_7_pad  = n141 ;
  assign \v13_D_9_pad  = n148 ;
endmodule
