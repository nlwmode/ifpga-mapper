module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	output e_pad ;
	output f_pad ;
	output g_pad ;
	output h_pad ;
	output i_pad ;
	output j_pad ;
	output k_pad ;
	output l_pad ;
	output m_pad ;
	output n_pad ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w5_ ;
	wire _w6_ ;
	wire _w7_ ;
	wire _w8_ ;
	wire _w9_ ;
	wire _w10_ ;
	wire _w11_ ;
	wire _w12_ ;
	wire _w13_ ;
	wire _w14_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		c_pad,
		d_pad,
		_w5_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		a_pad,
		b_pad,
		_w6_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w5_,
		_w6_,
		_w7_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		a_pad,
		b_pad,
		_w8_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		_w5_,
		_w8_,
		_w9_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		a_pad,
		b_pad,
		_w10_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w5_,
		_w10_,
		_w11_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		a_pad,
		b_pad,
		_w12_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w5_,
		_w12_,
		_w13_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		c_pad,
		d_pad,
		_w14_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w6_,
		_w14_,
		_w15_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w8_,
		_w14_,
		_w16_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w10_,
		_w14_,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w12_,
		_w14_,
		_w18_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		b_pad,
		c_pad,
		_w19_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		d_pad,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		a_pad,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		a_pad,
		_w20_,
		_w22_
	);
	assign e_pad = _w7_ ;
	assign f_pad = _w9_ ;
	assign g_pad = _w11_ ;
	assign h_pad = _w13_ ;
	assign i_pad = _w15_ ;
	assign j_pad = _w16_ ;
	assign k_pad = _w17_ ;
	assign l_pad = _w18_ ;
	assign m_pad = _w21_ ;
	assign n_pad = _w22_ ;
endmodule;